module AND_X1 (A, B, Y);
input A, B;
output Y;
assign Y = (A & B);
endmodule 
