`include "large_mux.v"
`include "memory_cntrl.v"
`include "register.v"
`include "full_adder.v"
`include "d_latch.v"
`include "shift_reg.v"
`include "mod_n_counter.v"
`include "decoder.v"
`include "parity_generator.v"

module design188_100_80_top #(parameter WIDTH=32,CHANNEL=100) (clk, rst, in, out);

	localparam OUT_BUS=CHANNEL*WIDTH;
	input clk,rst;
	input [WIDTH-1:0] in;
	output [WIDTH-1:0] out;

	reg [WIDTH-1:0] d_in0;
	reg [WIDTH-1:0] d_in1;
	reg [WIDTH-1:0] d_in2;
	reg [WIDTH-1:0] d_in3;
	reg [WIDTH-1:0] d_in4;
	reg [WIDTH-1:0] d_in5;
	reg [WIDTH-1:0] d_in6;
	reg [WIDTH-1:0] d_in7;
	reg [WIDTH-1:0] d_in8;
	reg [WIDTH-1:0] d_in9;
	reg [WIDTH-1:0] d_in10;
	reg [WIDTH-1:0] d_in11;
	reg [WIDTH-1:0] d_in12;
	reg [WIDTH-1:0] d_in13;
	reg [WIDTH-1:0] d_in14;
	reg [WIDTH-1:0] d_in15;
	reg [WIDTH-1:0] d_in16;
	reg [WIDTH-1:0] d_in17;
	reg [WIDTH-1:0] d_in18;
	reg [WIDTH-1:0] d_in19;
	reg [WIDTH-1:0] d_in20;
	reg [WIDTH-1:0] d_in21;
	reg [WIDTH-1:0] d_in22;
	reg [WIDTH-1:0] d_in23;
	reg [WIDTH-1:0] d_in24;
	reg [WIDTH-1:0] d_in25;
	reg [WIDTH-1:0] d_in26;
	reg [WIDTH-1:0] d_in27;
	reg [WIDTH-1:0] d_in28;
	reg [WIDTH-1:0] d_in29;
	reg [WIDTH-1:0] d_in30;
	reg [WIDTH-1:0] d_in31;
	reg [WIDTH-1:0] d_in32;
	reg [WIDTH-1:0] d_in33;
	reg [WIDTH-1:0] d_in34;
	reg [WIDTH-1:0] d_in35;
	reg [WIDTH-1:0] d_in36;
	reg [WIDTH-1:0] d_in37;
	reg [WIDTH-1:0] d_in38;
	reg [WIDTH-1:0] d_in39;
	reg [WIDTH-1:0] d_in40;
	reg [WIDTH-1:0] d_in41;
	reg [WIDTH-1:0] d_in42;
	reg [WIDTH-1:0] d_in43;
	reg [WIDTH-1:0] d_in44;
	reg [WIDTH-1:0] d_in45;
	reg [WIDTH-1:0] d_in46;
	reg [WIDTH-1:0] d_in47;
	reg [WIDTH-1:0] d_in48;
	reg [WIDTH-1:0] d_in49;
	reg [WIDTH-1:0] d_in50;
	reg [WIDTH-1:0] d_in51;
	reg [WIDTH-1:0] d_in52;
	reg [WIDTH-1:0] d_in53;
	reg [WIDTH-1:0] d_in54;
	reg [WIDTH-1:0] d_in55;
	reg [WIDTH-1:0] d_in56;
	reg [WIDTH-1:0] d_in57;
	reg [WIDTH-1:0] d_in58;
	reg [WIDTH-1:0] d_in59;
	reg [WIDTH-1:0] d_in60;
	reg [WIDTH-1:0] d_in61;
	reg [WIDTH-1:0] d_in62;
	reg [WIDTH-1:0] d_in63;
	reg [WIDTH-1:0] d_in64;
	reg [WIDTH-1:0] d_in65;
	reg [WIDTH-1:0] d_in66;
	reg [WIDTH-1:0] d_in67;
	reg [WIDTH-1:0] d_in68;
	reg [WIDTH-1:0] d_in69;
	reg [WIDTH-1:0] d_in70;
	reg [WIDTH-1:0] d_in71;
	reg [WIDTH-1:0] d_in72;
	reg [WIDTH-1:0] d_in73;
	reg [WIDTH-1:0] d_in74;
	reg [WIDTH-1:0] d_in75;
	reg [WIDTH-1:0] d_in76;
	reg [WIDTH-1:0] d_in77;
	reg [WIDTH-1:0] d_in78;
	reg [WIDTH-1:0] d_in79;
	reg [WIDTH-1:0] d_in80;
	reg [WIDTH-1:0] d_in81;
	reg [WIDTH-1:0] d_in82;
	reg [WIDTH-1:0] d_in83;
	reg [WIDTH-1:0] d_in84;
	reg [WIDTH-1:0] d_in85;
	reg [WIDTH-1:0] d_in86;
	reg [WIDTH-1:0] d_in87;
	reg [WIDTH-1:0] d_in88;
	reg [WIDTH-1:0] d_in89;
	reg [WIDTH-1:0] d_in90;
	reg [WIDTH-1:0] d_in91;
	reg [WIDTH-1:0] d_in92;
	reg [WIDTH-1:0] d_in93;
	reg [WIDTH-1:0] d_in94;
	reg [WIDTH-1:0] d_in95;
	reg [WIDTH-1:0] d_in96;
	reg [WIDTH-1:0] d_in97;
	reg [WIDTH-1:0] d_in98;
	reg [WIDTH-1:0] d_in99;
	wire [WIDTH-1:0] d_out0;
	wire [WIDTH-1:0] d_out1;
	wire [WIDTH-1:0] d_out2;
	wire [WIDTH-1:0] d_out3;
	wire [WIDTH-1:0] d_out4;
	wire [WIDTH-1:0] d_out5;
	wire [WIDTH-1:0] d_out6;
	wire [WIDTH-1:0] d_out7;
	wire [WIDTH-1:0] d_out8;
	wire [WIDTH-1:0] d_out9;
	wire [WIDTH-1:0] d_out10;
	wire [WIDTH-1:0] d_out11;
	wire [WIDTH-1:0] d_out12;
	wire [WIDTH-1:0] d_out13;
	wire [WIDTH-1:0] d_out14;
	wire [WIDTH-1:0] d_out15;
	wire [WIDTH-1:0] d_out16;
	wire [WIDTH-1:0] d_out17;
	wire [WIDTH-1:0] d_out18;
	wire [WIDTH-1:0] d_out19;
	wire [WIDTH-1:0] d_out20;
	wire [WIDTH-1:0] d_out21;
	wire [WIDTH-1:0] d_out22;
	wire [WIDTH-1:0] d_out23;
	wire [WIDTH-1:0] d_out24;
	wire [WIDTH-1:0] d_out25;
	wire [WIDTH-1:0] d_out26;
	wire [WIDTH-1:0] d_out27;
	wire [WIDTH-1:0] d_out28;
	wire [WIDTH-1:0] d_out29;
	wire [WIDTH-1:0] d_out30;
	wire [WIDTH-1:0] d_out31;
	wire [WIDTH-1:0] d_out32;
	wire [WIDTH-1:0] d_out33;
	wire [WIDTH-1:0] d_out34;
	wire [WIDTH-1:0] d_out35;
	wire [WIDTH-1:0] d_out36;
	wire [WIDTH-1:0] d_out37;
	wire [WIDTH-1:0] d_out38;
	wire [WIDTH-1:0] d_out39;
	wire [WIDTH-1:0] d_out40;
	wire [WIDTH-1:0] d_out41;
	wire [WIDTH-1:0] d_out42;
	wire [WIDTH-1:0] d_out43;
	wire [WIDTH-1:0] d_out44;
	wire [WIDTH-1:0] d_out45;
	wire [WIDTH-1:0] d_out46;
	wire [WIDTH-1:0] d_out47;
	wire [WIDTH-1:0] d_out48;
	wire [WIDTH-1:0] d_out49;
	wire [WIDTH-1:0] d_out50;
	wire [WIDTH-1:0] d_out51;
	wire [WIDTH-1:0] d_out52;
	wire [WIDTH-1:0] d_out53;
	wire [WIDTH-1:0] d_out54;
	wire [WIDTH-1:0] d_out55;
	wire [WIDTH-1:0] d_out56;
	wire [WIDTH-1:0] d_out57;
	wire [WIDTH-1:0] d_out58;
	wire [WIDTH-1:0] d_out59;
	wire [WIDTH-1:0] d_out60;
	wire [WIDTH-1:0] d_out61;
	wire [WIDTH-1:0] d_out62;
	wire [WIDTH-1:0] d_out63;
	wire [WIDTH-1:0] d_out64;
	wire [WIDTH-1:0] d_out65;
	wire [WIDTH-1:0] d_out66;
	wire [WIDTH-1:0] d_out67;
	wire [WIDTH-1:0] d_out68;
	wire [WIDTH-1:0] d_out69;
	wire [WIDTH-1:0] d_out70;
	wire [WIDTH-1:0] d_out71;
	wire [WIDTH-1:0] d_out72;
	wire [WIDTH-1:0] d_out73;
	wire [WIDTH-1:0] d_out74;
	wire [WIDTH-1:0] d_out75;
	wire [WIDTH-1:0] d_out76;
	wire [WIDTH-1:0] d_out77;
	wire [WIDTH-1:0] d_out78;
	wire [WIDTH-1:0] d_out79;
	wire [WIDTH-1:0] d_out80;
	wire [WIDTH-1:0] d_out81;
	wire [WIDTH-1:0] d_out82;
	wire [WIDTH-1:0] d_out83;
	wire [WIDTH-1:0] d_out84;
	wire [WIDTH-1:0] d_out85;
	wire [WIDTH-1:0] d_out86;
	wire [WIDTH-1:0] d_out87;
	wire [WIDTH-1:0] d_out88;
	wire [WIDTH-1:0] d_out89;
	wire [WIDTH-1:0] d_out90;
	wire [WIDTH-1:0] d_out91;
	wire [WIDTH-1:0] d_out92;
	wire [WIDTH-1:0] d_out93;
	wire [WIDTH-1:0] d_out94;
	wire [WIDTH-1:0] d_out95;
	wire [WIDTH-1:0] d_out96;
	wire [WIDTH-1:0] d_out97;
	wire [WIDTH-1:0] d_out98;
	wire [WIDTH-1:0] d_out99;

	reg [OUT_BUS-1:0] tmp;

	always @ (posedge clk or posedge rst) begin
		if (rst)
			tmp <= 0;
		else
			tmp <= {tmp[OUT_BUS-(WIDTH-1):0],in};
	end

	always @ (posedge clk) begin
		d_in0 <= tmp[WIDTH-1:0];
		d_in1 <= tmp[(WIDTH*2)-1:WIDTH*1];
		d_in2 <= tmp[(WIDTH*3)-1:WIDTH*2];
		d_in3 <= tmp[(WIDTH*4)-1:WIDTH*3];
		d_in4 <= tmp[(WIDTH*5)-1:WIDTH*4];
		d_in5 <= tmp[(WIDTH*6)-1:WIDTH*5];
		d_in6 <= tmp[(WIDTH*7)-1:WIDTH*6];
		d_in7 <= tmp[(WIDTH*8)-1:WIDTH*7];
		d_in8 <= tmp[(WIDTH*9)-1:WIDTH*8];
		d_in9 <= tmp[(WIDTH*10)-1:WIDTH*9];
		d_in10 <= tmp[(WIDTH*11)-1:WIDTH*10];
		d_in11 <= tmp[(WIDTH*12)-1:WIDTH*11];
		d_in12 <= tmp[(WIDTH*13)-1:WIDTH*12];
		d_in13 <= tmp[(WIDTH*14)-1:WIDTH*13];
		d_in14 <= tmp[(WIDTH*15)-1:WIDTH*14];
		d_in15 <= tmp[(WIDTH*16)-1:WIDTH*15];
		d_in16 <= tmp[(WIDTH*17)-1:WIDTH*16];
		d_in17 <= tmp[(WIDTH*18)-1:WIDTH*17];
		d_in18 <= tmp[(WIDTH*19)-1:WIDTH*18];
		d_in19 <= tmp[(WIDTH*20)-1:WIDTH*19];
		d_in20 <= tmp[(WIDTH*21)-1:WIDTH*20];
		d_in21 <= tmp[(WIDTH*22)-1:WIDTH*21];
		d_in22 <= tmp[(WIDTH*23)-1:WIDTH*22];
		d_in23 <= tmp[(WIDTH*24)-1:WIDTH*23];
		d_in24 <= tmp[(WIDTH*25)-1:WIDTH*24];
		d_in25 <= tmp[(WIDTH*26)-1:WIDTH*25];
		d_in26 <= tmp[(WIDTH*27)-1:WIDTH*26];
		d_in27 <= tmp[(WIDTH*28)-1:WIDTH*27];
		d_in28 <= tmp[(WIDTH*29)-1:WIDTH*28];
		d_in29 <= tmp[(WIDTH*30)-1:WIDTH*29];
		d_in30 <= tmp[(WIDTH*31)-1:WIDTH*30];
		d_in31 <= tmp[(WIDTH*32)-1:WIDTH*31];
		d_in32 <= tmp[(WIDTH*33)-1:WIDTH*32];
		d_in33 <= tmp[(WIDTH*34)-1:WIDTH*33];
		d_in34 <= tmp[(WIDTH*35)-1:WIDTH*34];
		d_in35 <= tmp[(WIDTH*36)-1:WIDTH*35];
		d_in36 <= tmp[(WIDTH*37)-1:WIDTH*36];
		d_in37 <= tmp[(WIDTH*38)-1:WIDTH*37];
		d_in38 <= tmp[(WIDTH*39)-1:WIDTH*38];
		d_in39 <= tmp[(WIDTH*40)-1:WIDTH*39];
		d_in40 <= tmp[(WIDTH*41)-1:WIDTH*40];
		d_in41 <= tmp[(WIDTH*42)-1:WIDTH*41];
		d_in42 <= tmp[(WIDTH*43)-1:WIDTH*42];
		d_in43 <= tmp[(WIDTH*44)-1:WIDTH*43];
		d_in44 <= tmp[(WIDTH*45)-1:WIDTH*44];
		d_in45 <= tmp[(WIDTH*46)-1:WIDTH*45];
		d_in46 <= tmp[(WIDTH*47)-1:WIDTH*46];
		d_in47 <= tmp[(WIDTH*48)-1:WIDTH*47];
		d_in48 <= tmp[(WIDTH*49)-1:WIDTH*48];
		d_in49 <= tmp[(WIDTH*50)-1:WIDTH*49];
		d_in50 <= tmp[(WIDTH*51)-1:WIDTH*50];
		d_in51 <= tmp[(WIDTH*52)-1:WIDTH*51];
		d_in52 <= tmp[(WIDTH*53)-1:WIDTH*52];
		d_in53 <= tmp[(WIDTH*54)-1:WIDTH*53];
		d_in54 <= tmp[(WIDTH*55)-1:WIDTH*54];
		d_in55 <= tmp[(WIDTH*56)-1:WIDTH*55];
		d_in56 <= tmp[(WIDTH*57)-1:WIDTH*56];
		d_in57 <= tmp[(WIDTH*58)-1:WIDTH*57];
		d_in58 <= tmp[(WIDTH*59)-1:WIDTH*58];
		d_in59 <= tmp[(WIDTH*60)-1:WIDTH*59];
		d_in60 <= tmp[(WIDTH*61)-1:WIDTH*60];
		d_in61 <= tmp[(WIDTH*62)-1:WIDTH*61];
		d_in62 <= tmp[(WIDTH*63)-1:WIDTH*62];
		d_in63 <= tmp[(WIDTH*64)-1:WIDTH*63];
		d_in64 <= tmp[(WIDTH*65)-1:WIDTH*64];
		d_in65 <= tmp[(WIDTH*66)-1:WIDTH*65];
		d_in66 <= tmp[(WIDTH*67)-1:WIDTH*66];
		d_in67 <= tmp[(WIDTH*68)-1:WIDTH*67];
		d_in68 <= tmp[(WIDTH*69)-1:WIDTH*68];
		d_in69 <= tmp[(WIDTH*70)-1:WIDTH*69];
		d_in70 <= tmp[(WIDTH*71)-1:WIDTH*70];
		d_in71 <= tmp[(WIDTH*72)-1:WIDTH*71];
		d_in72 <= tmp[(WIDTH*73)-1:WIDTH*72];
		d_in73 <= tmp[(WIDTH*74)-1:WIDTH*73];
		d_in74 <= tmp[(WIDTH*75)-1:WIDTH*74];
		d_in75 <= tmp[(WIDTH*76)-1:WIDTH*75];
		d_in76 <= tmp[(WIDTH*77)-1:WIDTH*76];
		d_in77 <= tmp[(WIDTH*78)-1:WIDTH*77];
		d_in78 <= tmp[(WIDTH*79)-1:WIDTH*78];
		d_in79 <= tmp[(WIDTH*80)-1:WIDTH*79];
		d_in80 <= tmp[(WIDTH*81)-1:WIDTH*80];
		d_in81 <= tmp[(WIDTH*82)-1:WIDTH*81];
		d_in82 <= tmp[(WIDTH*83)-1:WIDTH*82];
		d_in83 <= tmp[(WIDTH*84)-1:WIDTH*83];
		d_in84 <= tmp[(WIDTH*85)-1:WIDTH*84];
		d_in85 <= tmp[(WIDTH*86)-1:WIDTH*85];
		d_in86 <= tmp[(WIDTH*87)-1:WIDTH*86];
		d_in87 <= tmp[(WIDTH*88)-1:WIDTH*87];
		d_in88 <= tmp[(WIDTH*89)-1:WIDTH*88];
		d_in89 <= tmp[(WIDTH*90)-1:WIDTH*89];
		d_in90 <= tmp[(WIDTH*91)-1:WIDTH*90];
		d_in91 <= tmp[(WIDTH*92)-1:WIDTH*91];
		d_in92 <= tmp[(WIDTH*93)-1:WIDTH*92];
		d_in93 <= tmp[(WIDTH*94)-1:WIDTH*93];
		d_in94 <= tmp[(WIDTH*95)-1:WIDTH*94];
		d_in95 <= tmp[(WIDTH*96)-1:WIDTH*95];
		d_in96 <= tmp[(WIDTH*97)-1:WIDTH*96];
		d_in97 <= tmp[(WIDTH*98)-1:WIDTH*97];
		d_in98 <= tmp[(WIDTH*99)-1:WIDTH*98];
		d_in99 <= tmp[(WIDTH*100)-1:WIDTH*99];
	end

	design188_100_80 #(.WIDTH(WIDTH)) design188_100_80_inst(.d_in0(d_in0),.d_in1(d_in1),.d_in2(d_in2),.d_in3(d_in3),.d_in4(d_in4),.d_in5(d_in5),.d_in6(d_in6),.d_in7(d_in7),.d_in8(d_in8),.d_in9(d_in9),.d_in10(d_in10),.d_in11(d_in11),.d_in12(d_in12),.d_in13(d_in13),.d_in14(d_in14),.d_in15(d_in15),.d_in16(d_in16),.d_in17(d_in17),.d_in18(d_in18),.d_in19(d_in19),.d_in20(d_in20),.d_in21(d_in21),.d_in22(d_in22),.d_in23(d_in23),.d_in24(d_in24),.d_in25(d_in25),.d_in26(d_in26),.d_in27(d_in27),.d_in28(d_in28),.d_in29(d_in29),.d_in30(d_in30),.d_in31(d_in31),.d_in32(d_in32),.d_in33(d_in33),.d_in34(d_in34),.d_in35(d_in35),.d_in36(d_in36),.d_in37(d_in37),.d_in38(d_in38),.d_in39(d_in39),.d_in40(d_in40),.d_in41(d_in41),.d_in42(d_in42),.d_in43(d_in43),.d_in44(d_in44),.d_in45(d_in45),.d_in46(d_in46),.d_in47(d_in47),.d_in48(d_in48),.d_in49(d_in49),.d_in50(d_in50),.d_in51(d_in51),.d_in52(d_in52),.d_in53(d_in53),.d_in54(d_in54),.d_in55(d_in55),.d_in56(d_in56),.d_in57(d_in57),.d_in58(d_in58),.d_in59(d_in59),.d_in60(d_in60),.d_in61(d_in61),.d_in62(d_in62),.d_in63(d_in63),.d_in64(d_in64),.d_in65(d_in65),.d_in66(d_in66),.d_in67(d_in67),.d_in68(d_in68),.d_in69(d_in69),.d_in70(d_in70),.d_in71(d_in71),.d_in72(d_in72),.d_in73(d_in73),.d_in74(d_in74),.d_in75(d_in75),.d_in76(d_in76),.d_in77(d_in77),.d_in78(d_in78),.d_in79(d_in79),.d_in80(d_in80),.d_in81(d_in81),.d_in82(d_in82),.d_in83(d_in83),.d_in84(d_in84),.d_in85(d_in85),.d_in86(d_in86),.d_in87(d_in87),.d_in88(d_in88),.d_in89(d_in89),.d_in90(d_in90),.d_in91(d_in91),.d_in92(d_in92),.d_in93(d_in93),.d_in94(d_in94),.d_in95(d_in95),.d_in96(d_in96),.d_in97(d_in97),.d_in98(d_in98),.d_in99(d_in99),.d_out0(d_out0),.d_out1(d_out1),.d_out2(d_out2),.d_out3(d_out3),.d_out4(d_out4),.d_out5(d_out5),.d_out6(d_out6),.d_out7(d_out7),.d_out8(d_out8),.d_out9(d_out9),.d_out10(d_out10),.d_out11(d_out11),.d_out12(d_out12),.d_out13(d_out13),.d_out14(d_out14),.d_out15(d_out15),.d_out16(d_out16),.d_out17(d_out17),.d_out18(d_out18),.d_out19(d_out19),.d_out20(d_out20),.d_out21(d_out21),.d_out22(d_out22),.d_out23(d_out23),.d_out24(d_out24),.d_out25(d_out25),.d_out26(d_out26),.d_out27(d_out27),.d_out28(d_out28),.d_out29(d_out29),.d_out30(d_out30),.d_out31(d_out31),.d_out32(d_out32),.d_out33(d_out33),.d_out34(d_out34),.d_out35(d_out35),.d_out36(d_out36),.d_out37(d_out37),.d_out38(d_out38),.d_out39(d_out39),.d_out40(d_out40),.d_out41(d_out41),.d_out42(d_out42),.d_out43(d_out43),.d_out44(d_out44),.d_out45(d_out45),.d_out46(d_out46),.d_out47(d_out47),.d_out48(d_out48),.d_out49(d_out49),.d_out50(d_out50),.d_out51(d_out51),.d_out52(d_out52),.d_out53(d_out53),.d_out54(d_out54),.d_out55(d_out55),.d_out56(d_out56),.d_out57(d_out57),.d_out58(d_out58),.d_out59(d_out59),.d_out60(d_out60),.d_out61(d_out61),.d_out62(d_out62),.d_out63(d_out63),.d_out64(d_out64),.d_out65(d_out65),.d_out66(d_out66),.d_out67(d_out67),.d_out68(d_out68),.d_out69(d_out69),.d_out70(d_out70),.d_out71(d_out71),.d_out72(d_out72),.d_out73(d_out73),.d_out74(d_out74),.d_out75(d_out75),.d_out76(d_out76),.d_out77(d_out77),.d_out78(d_out78),.d_out79(d_out79),.d_out80(d_out80),.d_out81(d_out81),.d_out82(d_out82),.d_out83(d_out83),.d_out84(d_out84),.d_out85(d_out85),.d_out86(d_out86),.d_out87(d_out87),.d_out88(d_out88),.d_out89(d_out89),.d_out90(d_out90),.d_out91(d_out91),.d_out92(d_out92),.d_out93(d_out93),.d_out94(d_out94),.d_out95(d_out95),.d_out96(d_out96),.d_out97(d_out97),.d_out98(d_out98),.d_out99(d_out99),.clk(clk),.rst(rst));

	assign out = d_out0^d_out1^d_out2^d_out3^d_out4^d_out5^d_out6^d_out7^d_out8^d_out9^d_out10^d_out11^d_out12^d_out13^d_out14^d_out15^d_out16^d_out17^d_out18^d_out19^d_out20^d_out21^d_out22^d_out23^d_out24^d_out25^d_out26^d_out27^d_out28^d_out29^d_out30^d_out31^d_out32^d_out33^d_out34^d_out35^d_out36^d_out37^d_out38^d_out39^d_out40^d_out41^d_out42^d_out43^d_out44^d_out45^d_out46^d_out47^d_out48^d_out49^d_out50^d_out51^d_out52^d_out53^d_out54^d_out55^d_out56^d_out57^d_out58^d_out59^d_out60^d_out61^d_out62^d_out63^d_out64^d_out65^d_out66^d_out67^d_out68^d_out69^d_out70^d_out71^d_out72^d_out73^d_out74^d_out75^d_out76^d_out77^d_out78^d_out79^d_out80^d_out81^d_out82^d_out83^d_out84^d_out85^d_out86^d_out87^d_out88^d_out89^d_out90^d_out91^d_out92^d_out93^d_out94^d_out95^d_out96^d_out97^d_out98^d_out99;

endmodule

module design188_100_80 #(parameter WIDTH=32) (d_in0, d_in1, d_in2, d_in3, d_in4, d_in5, d_in6, d_in7, d_in8, d_in9, d_in10, d_in11, d_in12, d_in13, d_in14, d_in15, d_in16, d_in17, d_in18, d_in19, d_in20, d_in21, d_in22, d_in23, d_in24, d_in25, d_in26, d_in27, d_in28, d_in29, d_in30, d_in31, d_in32, d_in33, d_in34, d_in35, d_in36, d_in37, d_in38, d_in39, d_in40, d_in41, d_in42, d_in43, d_in44, d_in45, d_in46, d_in47, d_in48, d_in49, d_in50, d_in51, d_in52, d_in53, d_in54, d_in55, d_in56, d_in57, d_in58, d_in59, d_in60, d_in61, d_in62, d_in63, d_in64, d_in65, d_in66, d_in67, d_in68, d_in69, d_in70, d_in71, d_in72, d_in73, d_in74, d_in75, d_in76, d_in77, d_in78, d_in79, d_in80, d_in81, d_in82, d_in83, d_in84, d_in85, d_in86, d_in87, d_in88, d_in89, d_in90, d_in91, d_in92, d_in93, d_in94, d_in95, d_in96, d_in97, d_in98, d_in99, d_out0, d_out1, d_out2, d_out3, d_out4, d_out5, d_out6, d_out7, d_out8, d_out9, d_out10, d_out11, d_out12, d_out13, d_out14, d_out15, d_out16, d_out17, d_out18, d_out19, d_out20, d_out21, d_out22, d_out23, d_out24, d_out25, d_out26, d_out27, d_out28, d_out29, d_out30, d_out31, d_out32, d_out33, d_out34, d_out35, d_out36, d_out37, d_out38, d_out39, d_out40, d_out41, d_out42, d_out43, d_out44, d_out45, d_out46, d_out47, d_out48, d_out49, d_out50, d_out51, d_out52, d_out53, d_out54, d_out55, d_out56, d_out57, d_out58, d_out59, d_out60, d_out61, d_out62, d_out63, d_out64, d_out65, d_out66, d_out67, d_out68, d_out69, d_out70, d_out71, d_out72, d_out73, d_out74, d_out75, d_out76, d_out77, d_out78, d_out79, d_out80, d_out81, d_out82, d_out83, d_out84, d_out85, d_out86, d_out87, d_out88, d_out89, d_out90, d_out91, d_out92, d_out93, d_out94, d_out95, d_out96, d_out97, d_out98, d_out99, clk, rst);
	input clk;
	input rst;
	input [WIDTH-1:0] d_in0; 
	input [WIDTH-1:0] d_in1; 
	input [WIDTH-1:0] d_in2; 
	input [WIDTH-1:0] d_in3; 
	input [WIDTH-1:0] d_in4; 
	input [WIDTH-1:0] d_in5; 
	input [WIDTH-1:0] d_in6; 
	input [WIDTH-1:0] d_in7; 
	input [WIDTH-1:0] d_in8; 
	input [WIDTH-1:0] d_in9; 
	input [WIDTH-1:0] d_in10; 
	input [WIDTH-1:0] d_in11; 
	input [WIDTH-1:0] d_in12; 
	input [WIDTH-1:0] d_in13; 
	input [WIDTH-1:0] d_in14; 
	input [WIDTH-1:0] d_in15; 
	input [WIDTH-1:0] d_in16; 
	input [WIDTH-1:0] d_in17; 
	input [WIDTH-1:0] d_in18; 
	input [WIDTH-1:0] d_in19; 
	input [WIDTH-1:0] d_in20; 
	input [WIDTH-1:0] d_in21; 
	input [WIDTH-1:0] d_in22; 
	input [WIDTH-1:0] d_in23; 
	input [WIDTH-1:0] d_in24; 
	input [WIDTH-1:0] d_in25; 
	input [WIDTH-1:0] d_in26; 
	input [WIDTH-1:0] d_in27; 
	input [WIDTH-1:0] d_in28; 
	input [WIDTH-1:0] d_in29; 
	input [WIDTH-1:0] d_in30; 
	input [WIDTH-1:0] d_in31; 
	input [WIDTH-1:0] d_in32; 
	input [WIDTH-1:0] d_in33; 
	input [WIDTH-1:0] d_in34; 
	input [WIDTH-1:0] d_in35; 
	input [WIDTH-1:0] d_in36; 
	input [WIDTH-1:0] d_in37; 
	input [WIDTH-1:0] d_in38; 
	input [WIDTH-1:0] d_in39; 
	input [WIDTH-1:0] d_in40; 
	input [WIDTH-1:0] d_in41; 
	input [WIDTH-1:0] d_in42; 
	input [WIDTH-1:0] d_in43; 
	input [WIDTH-1:0] d_in44; 
	input [WIDTH-1:0] d_in45; 
	input [WIDTH-1:0] d_in46; 
	input [WIDTH-1:0] d_in47; 
	input [WIDTH-1:0] d_in48; 
	input [WIDTH-1:0] d_in49; 
	input [WIDTH-1:0] d_in50; 
	input [WIDTH-1:0] d_in51; 
	input [WIDTH-1:0] d_in52; 
	input [WIDTH-1:0] d_in53; 
	input [WIDTH-1:0] d_in54; 
	input [WIDTH-1:0] d_in55; 
	input [WIDTH-1:0] d_in56; 
	input [WIDTH-1:0] d_in57; 
	input [WIDTH-1:0] d_in58; 
	input [WIDTH-1:0] d_in59; 
	input [WIDTH-1:0] d_in60; 
	input [WIDTH-1:0] d_in61; 
	input [WIDTH-1:0] d_in62; 
	input [WIDTH-1:0] d_in63; 
	input [WIDTH-1:0] d_in64; 
	input [WIDTH-1:0] d_in65; 
	input [WIDTH-1:0] d_in66; 
	input [WIDTH-1:0] d_in67; 
	input [WIDTH-1:0] d_in68; 
	input [WIDTH-1:0] d_in69; 
	input [WIDTH-1:0] d_in70; 
	input [WIDTH-1:0] d_in71; 
	input [WIDTH-1:0] d_in72; 
	input [WIDTH-1:0] d_in73; 
	input [WIDTH-1:0] d_in74; 
	input [WIDTH-1:0] d_in75; 
	input [WIDTH-1:0] d_in76; 
	input [WIDTH-1:0] d_in77; 
	input [WIDTH-1:0] d_in78; 
	input [WIDTH-1:0] d_in79; 
	input [WIDTH-1:0] d_in80; 
	input [WIDTH-1:0] d_in81; 
	input [WIDTH-1:0] d_in82; 
	input [WIDTH-1:0] d_in83; 
	input [WIDTH-1:0] d_in84; 
	input [WIDTH-1:0] d_in85; 
	input [WIDTH-1:0] d_in86; 
	input [WIDTH-1:0] d_in87; 
	input [WIDTH-1:0] d_in88; 
	input [WIDTH-1:0] d_in89; 
	input [WIDTH-1:0] d_in90; 
	input [WIDTH-1:0] d_in91; 
	input [WIDTH-1:0] d_in92; 
	input [WIDTH-1:0] d_in93; 
	input [WIDTH-1:0] d_in94; 
	input [WIDTH-1:0] d_in95; 
	input [WIDTH-1:0] d_in96; 
	input [WIDTH-1:0] d_in97; 
	input [WIDTH-1:0] d_in98; 
	input [WIDTH-1:0] d_in99; 
	output [WIDTH-1:0] d_out0; 
	output [WIDTH-1:0] d_out1; 
	output [WIDTH-1:0] d_out2; 
	output [WIDTH-1:0] d_out3; 
	output [WIDTH-1:0] d_out4; 
	output [WIDTH-1:0] d_out5; 
	output [WIDTH-1:0] d_out6; 
	output [WIDTH-1:0] d_out7; 
	output [WIDTH-1:0] d_out8; 
	output [WIDTH-1:0] d_out9; 
	output [WIDTH-1:0] d_out10; 
	output [WIDTH-1:0] d_out11; 
	output [WIDTH-1:0] d_out12; 
	output [WIDTH-1:0] d_out13; 
	output [WIDTH-1:0] d_out14; 
	output [WIDTH-1:0] d_out15; 
	output [WIDTH-1:0] d_out16; 
	output [WIDTH-1:0] d_out17; 
	output [WIDTH-1:0] d_out18; 
	output [WIDTH-1:0] d_out19; 
	output [WIDTH-1:0] d_out20; 
	output [WIDTH-1:0] d_out21; 
	output [WIDTH-1:0] d_out22; 
	output [WIDTH-1:0] d_out23; 
	output [WIDTH-1:0] d_out24; 
	output [WIDTH-1:0] d_out25; 
	output [WIDTH-1:0] d_out26; 
	output [WIDTH-1:0] d_out27; 
	output [WIDTH-1:0] d_out28; 
	output [WIDTH-1:0] d_out29; 
	output [WIDTH-1:0] d_out30; 
	output [WIDTH-1:0] d_out31; 
	output [WIDTH-1:0] d_out32; 
	output [WIDTH-1:0] d_out33; 
	output [WIDTH-1:0] d_out34; 
	output [WIDTH-1:0] d_out35; 
	output [WIDTH-1:0] d_out36; 
	output [WIDTH-1:0] d_out37; 
	output [WIDTH-1:0] d_out38; 
	output [WIDTH-1:0] d_out39; 
	output [WIDTH-1:0] d_out40; 
	output [WIDTH-1:0] d_out41; 
	output [WIDTH-1:0] d_out42; 
	output [WIDTH-1:0] d_out43; 
	output [WIDTH-1:0] d_out44; 
	output [WIDTH-1:0] d_out45; 
	output [WIDTH-1:0] d_out46; 
	output [WIDTH-1:0] d_out47; 
	output [WIDTH-1:0] d_out48; 
	output [WIDTH-1:0] d_out49; 
	output [WIDTH-1:0] d_out50; 
	output [WIDTH-1:0] d_out51; 
	output [WIDTH-1:0] d_out52; 
	output [WIDTH-1:0] d_out53; 
	output [WIDTH-1:0] d_out54; 
	output [WIDTH-1:0] d_out55; 
	output [WIDTH-1:0] d_out56; 
	output [WIDTH-1:0] d_out57; 
	output [WIDTH-1:0] d_out58; 
	output [WIDTH-1:0] d_out59; 
	output [WIDTH-1:0] d_out60; 
	output [WIDTH-1:0] d_out61; 
	output [WIDTH-1:0] d_out62; 
	output [WIDTH-1:0] d_out63; 
	output [WIDTH-1:0] d_out64; 
	output [WIDTH-1:0] d_out65; 
	output [WIDTH-1:0] d_out66; 
	output [WIDTH-1:0] d_out67; 
	output [WIDTH-1:0] d_out68; 
	output [WIDTH-1:0] d_out69; 
	output [WIDTH-1:0] d_out70; 
	output [WIDTH-1:0] d_out71; 
	output [WIDTH-1:0] d_out72; 
	output [WIDTH-1:0] d_out73; 
	output [WIDTH-1:0] d_out74; 
	output [WIDTH-1:0] d_out75; 
	output [WIDTH-1:0] d_out76; 
	output [WIDTH-1:0] d_out77; 
	output [WIDTH-1:0] d_out78; 
	output [WIDTH-1:0] d_out79; 
	output [WIDTH-1:0] d_out80; 
	output [WIDTH-1:0] d_out81; 
	output [WIDTH-1:0] d_out82; 
	output [WIDTH-1:0] d_out83; 
	output [WIDTH-1:0] d_out84; 
	output [WIDTH-1:0] d_out85; 
	output [WIDTH-1:0] d_out86; 
	output [WIDTH-1:0] d_out87; 
	output [WIDTH-1:0] d_out88; 
	output [WIDTH-1:0] d_out89; 
	output [WIDTH-1:0] d_out90; 
	output [WIDTH-1:0] d_out91; 
	output [WIDTH-1:0] d_out92; 
	output [WIDTH-1:0] d_out93; 
	output [WIDTH-1:0] d_out94; 
	output [WIDTH-1:0] d_out95; 
	output [WIDTH-1:0] d_out96; 
	output [WIDTH-1:0] d_out97; 
	output [WIDTH-1:0] d_out98; 
	output [WIDTH-1:0] d_out99; 

	wire [WIDTH-1:0] wire_d0_0;
	wire [WIDTH-1:0] wire_d0_1;
	wire [WIDTH-1:0] wire_d0_2;
	wire [WIDTH-1:0] wire_d0_3;
	wire [WIDTH-1:0] wire_d0_4;
	wire [WIDTH-1:0] wire_d0_5;
	wire [WIDTH-1:0] wire_d0_6;
	wire [WIDTH-1:0] wire_d0_7;
	wire [WIDTH-1:0] wire_d0_8;
	wire [WIDTH-1:0] wire_d0_9;
	wire [WIDTH-1:0] wire_d0_10;
	wire [WIDTH-1:0] wire_d0_11;
	wire [WIDTH-1:0] wire_d0_12;
	wire [WIDTH-1:0] wire_d0_13;
	wire [WIDTH-1:0] wire_d0_14;
	wire [WIDTH-1:0] wire_d0_15;
	wire [WIDTH-1:0] wire_d0_16;
	wire [WIDTH-1:0] wire_d0_17;
	wire [WIDTH-1:0] wire_d0_18;
	wire [WIDTH-1:0] wire_d0_19;
	wire [WIDTH-1:0] wire_d0_20;
	wire [WIDTH-1:0] wire_d0_21;
	wire [WIDTH-1:0] wire_d0_22;
	wire [WIDTH-1:0] wire_d0_23;
	wire [WIDTH-1:0] wire_d0_24;
	wire [WIDTH-1:0] wire_d0_25;
	wire [WIDTH-1:0] wire_d0_26;
	wire [WIDTH-1:0] wire_d0_27;
	wire [WIDTH-1:0] wire_d0_28;
	wire [WIDTH-1:0] wire_d0_29;
	wire [WIDTH-1:0] wire_d0_30;
	wire [WIDTH-1:0] wire_d0_31;
	wire [WIDTH-1:0] wire_d0_32;
	wire [WIDTH-1:0] wire_d0_33;
	wire [WIDTH-1:0] wire_d0_34;
	wire [WIDTH-1:0] wire_d0_35;
	wire [WIDTH-1:0] wire_d0_36;
	wire [WIDTH-1:0] wire_d0_37;
	wire [WIDTH-1:0] wire_d0_38;
	wire [WIDTH-1:0] wire_d0_39;
	wire [WIDTH-1:0] wire_d0_40;
	wire [WIDTH-1:0] wire_d0_41;
	wire [WIDTH-1:0] wire_d0_42;
	wire [WIDTH-1:0] wire_d0_43;
	wire [WIDTH-1:0] wire_d0_44;
	wire [WIDTH-1:0] wire_d0_45;
	wire [WIDTH-1:0] wire_d0_46;
	wire [WIDTH-1:0] wire_d0_47;
	wire [WIDTH-1:0] wire_d0_48;
	wire [WIDTH-1:0] wire_d0_49;
	wire [WIDTH-1:0] wire_d0_50;
	wire [WIDTH-1:0] wire_d0_51;
	wire [WIDTH-1:0] wire_d0_52;
	wire [WIDTH-1:0] wire_d0_53;
	wire [WIDTH-1:0] wire_d0_54;
	wire [WIDTH-1:0] wire_d0_55;
	wire [WIDTH-1:0] wire_d0_56;
	wire [WIDTH-1:0] wire_d0_57;
	wire [WIDTH-1:0] wire_d0_58;
	wire [WIDTH-1:0] wire_d0_59;
	wire [WIDTH-1:0] wire_d0_60;
	wire [WIDTH-1:0] wire_d0_61;
	wire [WIDTH-1:0] wire_d0_62;
	wire [WIDTH-1:0] wire_d0_63;
	wire [WIDTH-1:0] wire_d0_64;
	wire [WIDTH-1:0] wire_d0_65;
	wire [WIDTH-1:0] wire_d0_66;
	wire [WIDTH-1:0] wire_d0_67;
	wire [WIDTH-1:0] wire_d0_68;
	wire [WIDTH-1:0] wire_d0_69;
	wire [WIDTH-1:0] wire_d0_70;
	wire [WIDTH-1:0] wire_d0_71;
	wire [WIDTH-1:0] wire_d0_72;
	wire [WIDTH-1:0] wire_d0_73;
	wire [WIDTH-1:0] wire_d0_74;
	wire [WIDTH-1:0] wire_d0_75;
	wire [WIDTH-1:0] wire_d0_76;
	wire [WIDTH-1:0] wire_d0_77;
	wire [WIDTH-1:0] wire_d0_78;
	wire [WIDTH-1:0] wire_d1_0;
	wire [WIDTH-1:0] wire_d1_1;
	wire [WIDTH-1:0] wire_d1_2;
	wire [WIDTH-1:0] wire_d1_3;
	wire [WIDTH-1:0] wire_d1_4;
	wire [WIDTH-1:0] wire_d1_5;
	wire [WIDTH-1:0] wire_d1_6;
	wire [WIDTH-1:0] wire_d1_7;
	wire [WIDTH-1:0] wire_d1_8;
	wire [WIDTH-1:0] wire_d1_9;
	wire [WIDTH-1:0] wire_d1_10;
	wire [WIDTH-1:0] wire_d1_11;
	wire [WIDTH-1:0] wire_d1_12;
	wire [WIDTH-1:0] wire_d1_13;
	wire [WIDTH-1:0] wire_d1_14;
	wire [WIDTH-1:0] wire_d1_15;
	wire [WIDTH-1:0] wire_d1_16;
	wire [WIDTH-1:0] wire_d1_17;
	wire [WIDTH-1:0] wire_d1_18;
	wire [WIDTH-1:0] wire_d1_19;
	wire [WIDTH-1:0] wire_d1_20;
	wire [WIDTH-1:0] wire_d1_21;
	wire [WIDTH-1:0] wire_d1_22;
	wire [WIDTH-1:0] wire_d1_23;
	wire [WIDTH-1:0] wire_d1_24;
	wire [WIDTH-1:0] wire_d1_25;
	wire [WIDTH-1:0] wire_d1_26;
	wire [WIDTH-1:0] wire_d1_27;
	wire [WIDTH-1:0] wire_d1_28;
	wire [WIDTH-1:0] wire_d1_29;
	wire [WIDTH-1:0] wire_d1_30;
	wire [WIDTH-1:0] wire_d1_31;
	wire [WIDTH-1:0] wire_d1_32;
	wire [WIDTH-1:0] wire_d1_33;
	wire [WIDTH-1:0] wire_d1_34;
	wire [WIDTH-1:0] wire_d1_35;
	wire [WIDTH-1:0] wire_d1_36;
	wire [WIDTH-1:0] wire_d1_37;
	wire [WIDTH-1:0] wire_d1_38;
	wire [WIDTH-1:0] wire_d1_39;
	wire [WIDTH-1:0] wire_d1_40;
	wire [WIDTH-1:0] wire_d1_41;
	wire [WIDTH-1:0] wire_d1_42;
	wire [WIDTH-1:0] wire_d1_43;
	wire [WIDTH-1:0] wire_d1_44;
	wire [WIDTH-1:0] wire_d1_45;
	wire [WIDTH-1:0] wire_d1_46;
	wire [WIDTH-1:0] wire_d1_47;
	wire [WIDTH-1:0] wire_d1_48;
	wire [WIDTH-1:0] wire_d1_49;
	wire [WIDTH-1:0] wire_d1_50;
	wire [WIDTH-1:0] wire_d1_51;
	wire [WIDTH-1:0] wire_d1_52;
	wire [WIDTH-1:0] wire_d1_53;
	wire [WIDTH-1:0] wire_d1_54;
	wire [WIDTH-1:0] wire_d1_55;
	wire [WIDTH-1:0] wire_d1_56;
	wire [WIDTH-1:0] wire_d1_57;
	wire [WIDTH-1:0] wire_d1_58;
	wire [WIDTH-1:0] wire_d1_59;
	wire [WIDTH-1:0] wire_d1_60;
	wire [WIDTH-1:0] wire_d1_61;
	wire [WIDTH-1:0] wire_d1_62;
	wire [WIDTH-1:0] wire_d1_63;
	wire [WIDTH-1:0] wire_d1_64;
	wire [WIDTH-1:0] wire_d1_65;
	wire [WIDTH-1:0] wire_d1_66;
	wire [WIDTH-1:0] wire_d1_67;
	wire [WIDTH-1:0] wire_d1_68;
	wire [WIDTH-1:0] wire_d1_69;
	wire [WIDTH-1:0] wire_d1_70;
	wire [WIDTH-1:0] wire_d1_71;
	wire [WIDTH-1:0] wire_d1_72;
	wire [WIDTH-1:0] wire_d1_73;
	wire [WIDTH-1:0] wire_d1_74;
	wire [WIDTH-1:0] wire_d1_75;
	wire [WIDTH-1:0] wire_d1_76;
	wire [WIDTH-1:0] wire_d1_77;
	wire [WIDTH-1:0] wire_d1_78;
	wire [WIDTH-1:0] wire_d2_0;
	wire [WIDTH-1:0] wire_d2_1;
	wire [WIDTH-1:0] wire_d2_2;
	wire [WIDTH-1:0] wire_d2_3;
	wire [WIDTH-1:0] wire_d2_4;
	wire [WIDTH-1:0] wire_d2_5;
	wire [WIDTH-1:0] wire_d2_6;
	wire [WIDTH-1:0] wire_d2_7;
	wire [WIDTH-1:0] wire_d2_8;
	wire [WIDTH-1:0] wire_d2_9;
	wire [WIDTH-1:0] wire_d2_10;
	wire [WIDTH-1:0] wire_d2_11;
	wire [WIDTH-1:0] wire_d2_12;
	wire [WIDTH-1:0] wire_d2_13;
	wire [WIDTH-1:0] wire_d2_14;
	wire [WIDTH-1:0] wire_d2_15;
	wire [WIDTH-1:0] wire_d2_16;
	wire [WIDTH-1:0] wire_d2_17;
	wire [WIDTH-1:0] wire_d2_18;
	wire [WIDTH-1:0] wire_d2_19;
	wire [WIDTH-1:0] wire_d2_20;
	wire [WIDTH-1:0] wire_d2_21;
	wire [WIDTH-1:0] wire_d2_22;
	wire [WIDTH-1:0] wire_d2_23;
	wire [WIDTH-1:0] wire_d2_24;
	wire [WIDTH-1:0] wire_d2_25;
	wire [WIDTH-1:0] wire_d2_26;
	wire [WIDTH-1:0] wire_d2_27;
	wire [WIDTH-1:0] wire_d2_28;
	wire [WIDTH-1:0] wire_d2_29;
	wire [WIDTH-1:0] wire_d2_30;
	wire [WIDTH-1:0] wire_d2_31;
	wire [WIDTH-1:0] wire_d2_32;
	wire [WIDTH-1:0] wire_d2_33;
	wire [WIDTH-1:0] wire_d2_34;
	wire [WIDTH-1:0] wire_d2_35;
	wire [WIDTH-1:0] wire_d2_36;
	wire [WIDTH-1:0] wire_d2_37;
	wire [WIDTH-1:0] wire_d2_38;
	wire [WIDTH-1:0] wire_d2_39;
	wire [WIDTH-1:0] wire_d2_40;
	wire [WIDTH-1:0] wire_d2_41;
	wire [WIDTH-1:0] wire_d2_42;
	wire [WIDTH-1:0] wire_d2_43;
	wire [WIDTH-1:0] wire_d2_44;
	wire [WIDTH-1:0] wire_d2_45;
	wire [WIDTH-1:0] wire_d2_46;
	wire [WIDTH-1:0] wire_d2_47;
	wire [WIDTH-1:0] wire_d2_48;
	wire [WIDTH-1:0] wire_d2_49;
	wire [WIDTH-1:0] wire_d2_50;
	wire [WIDTH-1:0] wire_d2_51;
	wire [WIDTH-1:0] wire_d2_52;
	wire [WIDTH-1:0] wire_d2_53;
	wire [WIDTH-1:0] wire_d2_54;
	wire [WIDTH-1:0] wire_d2_55;
	wire [WIDTH-1:0] wire_d2_56;
	wire [WIDTH-1:0] wire_d2_57;
	wire [WIDTH-1:0] wire_d2_58;
	wire [WIDTH-1:0] wire_d2_59;
	wire [WIDTH-1:0] wire_d2_60;
	wire [WIDTH-1:0] wire_d2_61;
	wire [WIDTH-1:0] wire_d2_62;
	wire [WIDTH-1:0] wire_d2_63;
	wire [WIDTH-1:0] wire_d2_64;
	wire [WIDTH-1:0] wire_d2_65;
	wire [WIDTH-1:0] wire_d2_66;
	wire [WIDTH-1:0] wire_d2_67;
	wire [WIDTH-1:0] wire_d2_68;
	wire [WIDTH-1:0] wire_d2_69;
	wire [WIDTH-1:0] wire_d2_70;
	wire [WIDTH-1:0] wire_d2_71;
	wire [WIDTH-1:0] wire_d2_72;
	wire [WIDTH-1:0] wire_d2_73;
	wire [WIDTH-1:0] wire_d2_74;
	wire [WIDTH-1:0] wire_d2_75;
	wire [WIDTH-1:0] wire_d2_76;
	wire [WIDTH-1:0] wire_d2_77;
	wire [WIDTH-1:0] wire_d2_78;
	wire [WIDTH-1:0] wire_d3_0;
	wire [WIDTH-1:0] wire_d3_1;
	wire [WIDTH-1:0] wire_d3_2;
	wire [WIDTH-1:0] wire_d3_3;
	wire [WIDTH-1:0] wire_d3_4;
	wire [WIDTH-1:0] wire_d3_5;
	wire [WIDTH-1:0] wire_d3_6;
	wire [WIDTH-1:0] wire_d3_7;
	wire [WIDTH-1:0] wire_d3_8;
	wire [WIDTH-1:0] wire_d3_9;
	wire [WIDTH-1:0] wire_d3_10;
	wire [WIDTH-1:0] wire_d3_11;
	wire [WIDTH-1:0] wire_d3_12;
	wire [WIDTH-1:0] wire_d3_13;
	wire [WIDTH-1:0] wire_d3_14;
	wire [WIDTH-1:0] wire_d3_15;
	wire [WIDTH-1:0] wire_d3_16;
	wire [WIDTH-1:0] wire_d3_17;
	wire [WIDTH-1:0] wire_d3_18;
	wire [WIDTH-1:0] wire_d3_19;
	wire [WIDTH-1:0] wire_d3_20;
	wire [WIDTH-1:0] wire_d3_21;
	wire [WIDTH-1:0] wire_d3_22;
	wire [WIDTH-1:0] wire_d3_23;
	wire [WIDTH-1:0] wire_d3_24;
	wire [WIDTH-1:0] wire_d3_25;
	wire [WIDTH-1:0] wire_d3_26;
	wire [WIDTH-1:0] wire_d3_27;
	wire [WIDTH-1:0] wire_d3_28;
	wire [WIDTH-1:0] wire_d3_29;
	wire [WIDTH-1:0] wire_d3_30;
	wire [WIDTH-1:0] wire_d3_31;
	wire [WIDTH-1:0] wire_d3_32;
	wire [WIDTH-1:0] wire_d3_33;
	wire [WIDTH-1:0] wire_d3_34;
	wire [WIDTH-1:0] wire_d3_35;
	wire [WIDTH-1:0] wire_d3_36;
	wire [WIDTH-1:0] wire_d3_37;
	wire [WIDTH-1:0] wire_d3_38;
	wire [WIDTH-1:0] wire_d3_39;
	wire [WIDTH-1:0] wire_d3_40;
	wire [WIDTH-1:0] wire_d3_41;
	wire [WIDTH-1:0] wire_d3_42;
	wire [WIDTH-1:0] wire_d3_43;
	wire [WIDTH-1:0] wire_d3_44;
	wire [WIDTH-1:0] wire_d3_45;
	wire [WIDTH-1:0] wire_d3_46;
	wire [WIDTH-1:0] wire_d3_47;
	wire [WIDTH-1:0] wire_d3_48;
	wire [WIDTH-1:0] wire_d3_49;
	wire [WIDTH-1:0] wire_d3_50;
	wire [WIDTH-1:0] wire_d3_51;
	wire [WIDTH-1:0] wire_d3_52;
	wire [WIDTH-1:0] wire_d3_53;
	wire [WIDTH-1:0] wire_d3_54;
	wire [WIDTH-1:0] wire_d3_55;
	wire [WIDTH-1:0] wire_d3_56;
	wire [WIDTH-1:0] wire_d3_57;
	wire [WIDTH-1:0] wire_d3_58;
	wire [WIDTH-1:0] wire_d3_59;
	wire [WIDTH-1:0] wire_d3_60;
	wire [WIDTH-1:0] wire_d3_61;
	wire [WIDTH-1:0] wire_d3_62;
	wire [WIDTH-1:0] wire_d3_63;
	wire [WIDTH-1:0] wire_d3_64;
	wire [WIDTH-1:0] wire_d3_65;
	wire [WIDTH-1:0] wire_d3_66;
	wire [WIDTH-1:0] wire_d3_67;
	wire [WIDTH-1:0] wire_d3_68;
	wire [WIDTH-1:0] wire_d3_69;
	wire [WIDTH-1:0] wire_d3_70;
	wire [WIDTH-1:0] wire_d3_71;
	wire [WIDTH-1:0] wire_d3_72;
	wire [WIDTH-1:0] wire_d3_73;
	wire [WIDTH-1:0] wire_d3_74;
	wire [WIDTH-1:0] wire_d3_75;
	wire [WIDTH-1:0] wire_d3_76;
	wire [WIDTH-1:0] wire_d3_77;
	wire [WIDTH-1:0] wire_d3_78;
	wire [WIDTH-1:0] wire_d4_0;
	wire [WIDTH-1:0] wire_d4_1;
	wire [WIDTH-1:0] wire_d4_2;
	wire [WIDTH-1:0] wire_d4_3;
	wire [WIDTH-1:0] wire_d4_4;
	wire [WIDTH-1:0] wire_d4_5;
	wire [WIDTH-1:0] wire_d4_6;
	wire [WIDTH-1:0] wire_d4_7;
	wire [WIDTH-1:0] wire_d4_8;
	wire [WIDTH-1:0] wire_d4_9;
	wire [WIDTH-1:0] wire_d4_10;
	wire [WIDTH-1:0] wire_d4_11;
	wire [WIDTH-1:0] wire_d4_12;
	wire [WIDTH-1:0] wire_d4_13;
	wire [WIDTH-1:0] wire_d4_14;
	wire [WIDTH-1:0] wire_d4_15;
	wire [WIDTH-1:0] wire_d4_16;
	wire [WIDTH-1:0] wire_d4_17;
	wire [WIDTH-1:0] wire_d4_18;
	wire [WIDTH-1:0] wire_d4_19;
	wire [WIDTH-1:0] wire_d4_20;
	wire [WIDTH-1:0] wire_d4_21;
	wire [WIDTH-1:0] wire_d4_22;
	wire [WIDTH-1:0] wire_d4_23;
	wire [WIDTH-1:0] wire_d4_24;
	wire [WIDTH-1:0] wire_d4_25;
	wire [WIDTH-1:0] wire_d4_26;
	wire [WIDTH-1:0] wire_d4_27;
	wire [WIDTH-1:0] wire_d4_28;
	wire [WIDTH-1:0] wire_d4_29;
	wire [WIDTH-1:0] wire_d4_30;
	wire [WIDTH-1:0] wire_d4_31;
	wire [WIDTH-1:0] wire_d4_32;
	wire [WIDTH-1:0] wire_d4_33;
	wire [WIDTH-1:0] wire_d4_34;
	wire [WIDTH-1:0] wire_d4_35;
	wire [WIDTH-1:0] wire_d4_36;
	wire [WIDTH-1:0] wire_d4_37;
	wire [WIDTH-1:0] wire_d4_38;
	wire [WIDTH-1:0] wire_d4_39;
	wire [WIDTH-1:0] wire_d4_40;
	wire [WIDTH-1:0] wire_d4_41;
	wire [WIDTH-1:0] wire_d4_42;
	wire [WIDTH-1:0] wire_d4_43;
	wire [WIDTH-1:0] wire_d4_44;
	wire [WIDTH-1:0] wire_d4_45;
	wire [WIDTH-1:0] wire_d4_46;
	wire [WIDTH-1:0] wire_d4_47;
	wire [WIDTH-1:0] wire_d4_48;
	wire [WIDTH-1:0] wire_d4_49;
	wire [WIDTH-1:0] wire_d4_50;
	wire [WIDTH-1:0] wire_d4_51;
	wire [WIDTH-1:0] wire_d4_52;
	wire [WIDTH-1:0] wire_d4_53;
	wire [WIDTH-1:0] wire_d4_54;
	wire [WIDTH-1:0] wire_d4_55;
	wire [WIDTH-1:0] wire_d4_56;
	wire [WIDTH-1:0] wire_d4_57;
	wire [WIDTH-1:0] wire_d4_58;
	wire [WIDTH-1:0] wire_d4_59;
	wire [WIDTH-1:0] wire_d4_60;
	wire [WIDTH-1:0] wire_d4_61;
	wire [WIDTH-1:0] wire_d4_62;
	wire [WIDTH-1:0] wire_d4_63;
	wire [WIDTH-1:0] wire_d4_64;
	wire [WIDTH-1:0] wire_d4_65;
	wire [WIDTH-1:0] wire_d4_66;
	wire [WIDTH-1:0] wire_d4_67;
	wire [WIDTH-1:0] wire_d4_68;
	wire [WIDTH-1:0] wire_d4_69;
	wire [WIDTH-1:0] wire_d4_70;
	wire [WIDTH-1:0] wire_d4_71;
	wire [WIDTH-1:0] wire_d4_72;
	wire [WIDTH-1:0] wire_d4_73;
	wire [WIDTH-1:0] wire_d4_74;
	wire [WIDTH-1:0] wire_d4_75;
	wire [WIDTH-1:0] wire_d4_76;
	wire [WIDTH-1:0] wire_d4_77;
	wire [WIDTH-1:0] wire_d4_78;
	wire [WIDTH-1:0] wire_d5_0;
	wire [WIDTH-1:0] wire_d5_1;
	wire [WIDTH-1:0] wire_d5_2;
	wire [WIDTH-1:0] wire_d5_3;
	wire [WIDTH-1:0] wire_d5_4;
	wire [WIDTH-1:0] wire_d5_5;
	wire [WIDTH-1:0] wire_d5_6;
	wire [WIDTH-1:0] wire_d5_7;
	wire [WIDTH-1:0] wire_d5_8;
	wire [WIDTH-1:0] wire_d5_9;
	wire [WIDTH-1:0] wire_d5_10;
	wire [WIDTH-1:0] wire_d5_11;
	wire [WIDTH-1:0] wire_d5_12;
	wire [WIDTH-1:0] wire_d5_13;
	wire [WIDTH-1:0] wire_d5_14;
	wire [WIDTH-1:0] wire_d5_15;
	wire [WIDTH-1:0] wire_d5_16;
	wire [WIDTH-1:0] wire_d5_17;
	wire [WIDTH-1:0] wire_d5_18;
	wire [WIDTH-1:0] wire_d5_19;
	wire [WIDTH-1:0] wire_d5_20;
	wire [WIDTH-1:0] wire_d5_21;
	wire [WIDTH-1:0] wire_d5_22;
	wire [WIDTH-1:0] wire_d5_23;
	wire [WIDTH-1:0] wire_d5_24;
	wire [WIDTH-1:0] wire_d5_25;
	wire [WIDTH-1:0] wire_d5_26;
	wire [WIDTH-1:0] wire_d5_27;
	wire [WIDTH-1:0] wire_d5_28;
	wire [WIDTH-1:0] wire_d5_29;
	wire [WIDTH-1:0] wire_d5_30;
	wire [WIDTH-1:0] wire_d5_31;
	wire [WIDTH-1:0] wire_d5_32;
	wire [WIDTH-1:0] wire_d5_33;
	wire [WIDTH-1:0] wire_d5_34;
	wire [WIDTH-1:0] wire_d5_35;
	wire [WIDTH-1:0] wire_d5_36;
	wire [WIDTH-1:0] wire_d5_37;
	wire [WIDTH-1:0] wire_d5_38;
	wire [WIDTH-1:0] wire_d5_39;
	wire [WIDTH-1:0] wire_d5_40;
	wire [WIDTH-1:0] wire_d5_41;
	wire [WIDTH-1:0] wire_d5_42;
	wire [WIDTH-1:0] wire_d5_43;
	wire [WIDTH-1:0] wire_d5_44;
	wire [WIDTH-1:0] wire_d5_45;
	wire [WIDTH-1:0] wire_d5_46;
	wire [WIDTH-1:0] wire_d5_47;
	wire [WIDTH-1:0] wire_d5_48;
	wire [WIDTH-1:0] wire_d5_49;
	wire [WIDTH-1:0] wire_d5_50;
	wire [WIDTH-1:0] wire_d5_51;
	wire [WIDTH-1:0] wire_d5_52;
	wire [WIDTH-1:0] wire_d5_53;
	wire [WIDTH-1:0] wire_d5_54;
	wire [WIDTH-1:0] wire_d5_55;
	wire [WIDTH-1:0] wire_d5_56;
	wire [WIDTH-1:0] wire_d5_57;
	wire [WIDTH-1:0] wire_d5_58;
	wire [WIDTH-1:0] wire_d5_59;
	wire [WIDTH-1:0] wire_d5_60;
	wire [WIDTH-1:0] wire_d5_61;
	wire [WIDTH-1:0] wire_d5_62;
	wire [WIDTH-1:0] wire_d5_63;
	wire [WIDTH-1:0] wire_d5_64;
	wire [WIDTH-1:0] wire_d5_65;
	wire [WIDTH-1:0] wire_d5_66;
	wire [WIDTH-1:0] wire_d5_67;
	wire [WIDTH-1:0] wire_d5_68;
	wire [WIDTH-1:0] wire_d5_69;
	wire [WIDTH-1:0] wire_d5_70;
	wire [WIDTH-1:0] wire_d5_71;
	wire [WIDTH-1:0] wire_d5_72;
	wire [WIDTH-1:0] wire_d5_73;
	wire [WIDTH-1:0] wire_d5_74;
	wire [WIDTH-1:0] wire_d5_75;
	wire [WIDTH-1:0] wire_d5_76;
	wire [WIDTH-1:0] wire_d5_77;
	wire [WIDTH-1:0] wire_d5_78;
	wire [WIDTH-1:0] wire_d6_0;
	wire [WIDTH-1:0] wire_d6_1;
	wire [WIDTH-1:0] wire_d6_2;
	wire [WIDTH-1:0] wire_d6_3;
	wire [WIDTH-1:0] wire_d6_4;
	wire [WIDTH-1:0] wire_d6_5;
	wire [WIDTH-1:0] wire_d6_6;
	wire [WIDTH-1:0] wire_d6_7;
	wire [WIDTH-1:0] wire_d6_8;
	wire [WIDTH-1:0] wire_d6_9;
	wire [WIDTH-1:0] wire_d6_10;
	wire [WIDTH-1:0] wire_d6_11;
	wire [WIDTH-1:0] wire_d6_12;
	wire [WIDTH-1:0] wire_d6_13;
	wire [WIDTH-1:0] wire_d6_14;
	wire [WIDTH-1:0] wire_d6_15;
	wire [WIDTH-1:0] wire_d6_16;
	wire [WIDTH-1:0] wire_d6_17;
	wire [WIDTH-1:0] wire_d6_18;
	wire [WIDTH-1:0] wire_d6_19;
	wire [WIDTH-1:0] wire_d6_20;
	wire [WIDTH-1:0] wire_d6_21;
	wire [WIDTH-1:0] wire_d6_22;
	wire [WIDTH-1:0] wire_d6_23;
	wire [WIDTH-1:0] wire_d6_24;
	wire [WIDTH-1:0] wire_d6_25;
	wire [WIDTH-1:0] wire_d6_26;
	wire [WIDTH-1:0] wire_d6_27;
	wire [WIDTH-1:0] wire_d6_28;
	wire [WIDTH-1:0] wire_d6_29;
	wire [WIDTH-1:0] wire_d6_30;
	wire [WIDTH-1:0] wire_d6_31;
	wire [WIDTH-1:0] wire_d6_32;
	wire [WIDTH-1:0] wire_d6_33;
	wire [WIDTH-1:0] wire_d6_34;
	wire [WIDTH-1:0] wire_d6_35;
	wire [WIDTH-1:0] wire_d6_36;
	wire [WIDTH-1:0] wire_d6_37;
	wire [WIDTH-1:0] wire_d6_38;
	wire [WIDTH-1:0] wire_d6_39;
	wire [WIDTH-1:0] wire_d6_40;
	wire [WIDTH-1:0] wire_d6_41;
	wire [WIDTH-1:0] wire_d6_42;
	wire [WIDTH-1:0] wire_d6_43;
	wire [WIDTH-1:0] wire_d6_44;
	wire [WIDTH-1:0] wire_d6_45;
	wire [WIDTH-1:0] wire_d6_46;
	wire [WIDTH-1:0] wire_d6_47;
	wire [WIDTH-1:0] wire_d6_48;
	wire [WIDTH-1:0] wire_d6_49;
	wire [WIDTH-1:0] wire_d6_50;
	wire [WIDTH-1:0] wire_d6_51;
	wire [WIDTH-1:0] wire_d6_52;
	wire [WIDTH-1:0] wire_d6_53;
	wire [WIDTH-1:0] wire_d6_54;
	wire [WIDTH-1:0] wire_d6_55;
	wire [WIDTH-1:0] wire_d6_56;
	wire [WIDTH-1:0] wire_d6_57;
	wire [WIDTH-1:0] wire_d6_58;
	wire [WIDTH-1:0] wire_d6_59;
	wire [WIDTH-1:0] wire_d6_60;
	wire [WIDTH-1:0] wire_d6_61;
	wire [WIDTH-1:0] wire_d6_62;
	wire [WIDTH-1:0] wire_d6_63;
	wire [WIDTH-1:0] wire_d6_64;
	wire [WIDTH-1:0] wire_d6_65;
	wire [WIDTH-1:0] wire_d6_66;
	wire [WIDTH-1:0] wire_d6_67;
	wire [WIDTH-1:0] wire_d6_68;
	wire [WIDTH-1:0] wire_d6_69;
	wire [WIDTH-1:0] wire_d6_70;
	wire [WIDTH-1:0] wire_d6_71;
	wire [WIDTH-1:0] wire_d6_72;
	wire [WIDTH-1:0] wire_d6_73;
	wire [WIDTH-1:0] wire_d6_74;
	wire [WIDTH-1:0] wire_d6_75;
	wire [WIDTH-1:0] wire_d6_76;
	wire [WIDTH-1:0] wire_d6_77;
	wire [WIDTH-1:0] wire_d6_78;
	wire [WIDTH-1:0] wire_d7_0;
	wire [WIDTH-1:0] wire_d7_1;
	wire [WIDTH-1:0] wire_d7_2;
	wire [WIDTH-1:0] wire_d7_3;
	wire [WIDTH-1:0] wire_d7_4;
	wire [WIDTH-1:0] wire_d7_5;
	wire [WIDTH-1:0] wire_d7_6;
	wire [WIDTH-1:0] wire_d7_7;
	wire [WIDTH-1:0] wire_d7_8;
	wire [WIDTH-1:0] wire_d7_9;
	wire [WIDTH-1:0] wire_d7_10;
	wire [WIDTH-1:0] wire_d7_11;
	wire [WIDTH-1:0] wire_d7_12;
	wire [WIDTH-1:0] wire_d7_13;
	wire [WIDTH-1:0] wire_d7_14;
	wire [WIDTH-1:0] wire_d7_15;
	wire [WIDTH-1:0] wire_d7_16;
	wire [WIDTH-1:0] wire_d7_17;
	wire [WIDTH-1:0] wire_d7_18;
	wire [WIDTH-1:0] wire_d7_19;
	wire [WIDTH-1:0] wire_d7_20;
	wire [WIDTH-1:0] wire_d7_21;
	wire [WIDTH-1:0] wire_d7_22;
	wire [WIDTH-1:0] wire_d7_23;
	wire [WIDTH-1:0] wire_d7_24;
	wire [WIDTH-1:0] wire_d7_25;
	wire [WIDTH-1:0] wire_d7_26;
	wire [WIDTH-1:0] wire_d7_27;
	wire [WIDTH-1:0] wire_d7_28;
	wire [WIDTH-1:0] wire_d7_29;
	wire [WIDTH-1:0] wire_d7_30;
	wire [WIDTH-1:0] wire_d7_31;
	wire [WIDTH-1:0] wire_d7_32;
	wire [WIDTH-1:0] wire_d7_33;
	wire [WIDTH-1:0] wire_d7_34;
	wire [WIDTH-1:0] wire_d7_35;
	wire [WIDTH-1:0] wire_d7_36;
	wire [WIDTH-1:0] wire_d7_37;
	wire [WIDTH-1:0] wire_d7_38;
	wire [WIDTH-1:0] wire_d7_39;
	wire [WIDTH-1:0] wire_d7_40;
	wire [WIDTH-1:0] wire_d7_41;
	wire [WIDTH-1:0] wire_d7_42;
	wire [WIDTH-1:0] wire_d7_43;
	wire [WIDTH-1:0] wire_d7_44;
	wire [WIDTH-1:0] wire_d7_45;
	wire [WIDTH-1:0] wire_d7_46;
	wire [WIDTH-1:0] wire_d7_47;
	wire [WIDTH-1:0] wire_d7_48;
	wire [WIDTH-1:0] wire_d7_49;
	wire [WIDTH-1:0] wire_d7_50;
	wire [WIDTH-1:0] wire_d7_51;
	wire [WIDTH-1:0] wire_d7_52;
	wire [WIDTH-1:0] wire_d7_53;
	wire [WIDTH-1:0] wire_d7_54;
	wire [WIDTH-1:0] wire_d7_55;
	wire [WIDTH-1:0] wire_d7_56;
	wire [WIDTH-1:0] wire_d7_57;
	wire [WIDTH-1:0] wire_d7_58;
	wire [WIDTH-1:0] wire_d7_59;
	wire [WIDTH-1:0] wire_d7_60;
	wire [WIDTH-1:0] wire_d7_61;
	wire [WIDTH-1:0] wire_d7_62;
	wire [WIDTH-1:0] wire_d7_63;
	wire [WIDTH-1:0] wire_d7_64;
	wire [WIDTH-1:0] wire_d7_65;
	wire [WIDTH-1:0] wire_d7_66;
	wire [WIDTH-1:0] wire_d7_67;
	wire [WIDTH-1:0] wire_d7_68;
	wire [WIDTH-1:0] wire_d7_69;
	wire [WIDTH-1:0] wire_d7_70;
	wire [WIDTH-1:0] wire_d7_71;
	wire [WIDTH-1:0] wire_d7_72;
	wire [WIDTH-1:0] wire_d7_73;
	wire [WIDTH-1:0] wire_d7_74;
	wire [WIDTH-1:0] wire_d7_75;
	wire [WIDTH-1:0] wire_d7_76;
	wire [WIDTH-1:0] wire_d7_77;
	wire [WIDTH-1:0] wire_d7_78;
	wire [WIDTH-1:0] wire_d8_0;
	wire [WIDTH-1:0] wire_d8_1;
	wire [WIDTH-1:0] wire_d8_2;
	wire [WIDTH-1:0] wire_d8_3;
	wire [WIDTH-1:0] wire_d8_4;
	wire [WIDTH-1:0] wire_d8_5;
	wire [WIDTH-1:0] wire_d8_6;
	wire [WIDTH-1:0] wire_d8_7;
	wire [WIDTH-1:0] wire_d8_8;
	wire [WIDTH-1:0] wire_d8_9;
	wire [WIDTH-1:0] wire_d8_10;
	wire [WIDTH-1:0] wire_d8_11;
	wire [WIDTH-1:0] wire_d8_12;
	wire [WIDTH-1:0] wire_d8_13;
	wire [WIDTH-1:0] wire_d8_14;
	wire [WIDTH-1:0] wire_d8_15;
	wire [WIDTH-1:0] wire_d8_16;
	wire [WIDTH-1:0] wire_d8_17;
	wire [WIDTH-1:0] wire_d8_18;
	wire [WIDTH-1:0] wire_d8_19;
	wire [WIDTH-1:0] wire_d8_20;
	wire [WIDTH-1:0] wire_d8_21;
	wire [WIDTH-1:0] wire_d8_22;
	wire [WIDTH-1:0] wire_d8_23;
	wire [WIDTH-1:0] wire_d8_24;
	wire [WIDTH-1:0] wire_d8_25;
	wire [WIDTH-1:0] wire_d8_26;
	wire [WIDTH-1:0] wire_d8_27;
	wire [WIDTH-1:0] wire_d8_28;
	wire [WIDTH-1:0] wire_d8_29;
	wire [WIDTH-1:0] wire_d8_30;
	wire [WIDTH-1:0] wire_d8_31;
	wire [WIDTH-1:0] wire_d8_32;
	wire [WIDTH-1:0] wire_d8_33;
	wire [WIDTH-1:0] wire_d8_34;
	wire [WIDTH-1:0] wire_d8_35;
	wire [WIDTH-1:0] wire_d8_36;
	wire [WIDTH-1:0] wire_d8_37;
	wire [WIDTH-1:0] wire_d8_38;
	wire [WIDTH-1:0] wire_d8_39;
	wire [WIDTH-1:0] wire_d8_40;
	wire [WIDTH-1:0] wire_d8_41;
	wire [WIDTH-1:0] wire_d8_42;
	wire [WIDTH-1:0] wire_d8_43;
	wire [WIDTH-1:0] wire_d8_44;
	wire [WIDTH-1:0] wire_d8_45;
	wire [WIDTH-1:0] wire_d8_46;
	wire [WIDTH-1:0] wire_d8_47;
	wire [WIDTH-1:0] wire_d8_48;
	wire [WIDTH-1:0] wire_d8_49;
	wire [WIDTH-1:0] wire_d8_50;
	wire [WIDTH-1:0] wire_d8_51;
	wire [WIDTH-1:0] wire_d8_52;
	wire [WIDTH-1:0] wire_d8_53;
	wire [WIDTH-1:0] wire_d8_54;
	wire [WIDTH-1:0] wire_d8_55;
	wire [WIDTH-1:0] wire_d8_56;
	wire [WIDTH-1:0] wire_d8_57;
	wire [WIDTH-1:0] wire_d8_58;
	wire [WIDTH-1:0] wire_d8_59;
	wire [WIDTH-1:0] wire_d8_60;
	wire [WIDTH-1:0] wire_d8_61;
	wire [WIDTH-1:0] wire_d8_62;
	wire [WIDTH-1:0] wire_d8_63;
	wire [WIDTH-1:0] wire_d8_64;
	wire [WIDTH-1:0] wire_d8_65;
	wire [WIDTH-1:0] wire_d8_66;
	wire [WIDTH-1:0] wire_d8_67;
	wire [WIDTH-1:0] wire_d8_68;
	wire [WIDTH-1:0] wire_d8_69;
	wire [WIDTH-1:0] wire_d8_70;
	wire [WIDTH-1:0] wire_d8_71;
	wire [WIDTH-1:0] wire_d8_72;
	wire [WIDTH-1:0] wire_d8_73;
	wire [WIDTH-1:0] wire_d8_74;
	wire [WIDTH-1:0] wire_d8_75;
	wire [WIDTH-1:0] wire_d8_76;
	wire [WIDTH-1:0] wire_d8_77;
	wire [WIDTH-1:0] wire_d8_78;
	wire [WIDTH-1:0] wire_d9_0;
	wire [WIDTH-1:0] wire_d9_1;
	wire [WIDTH-1:0] wire_d9_2;
	wire [WIDTH-1:0] wire_d9_3;
	wire [WIDTH-1:0] wire_d9_4;
	wire [WIDTH-1:0] wire_d9_5;
	wire [WIDTH-1:0] wire_d9_6;
	wire [WIDTH-1:0] wire_d9_7;
	wire [WIDTH-1:0] wire_d9_8;
	wire [WIDTH-1:0] wire_d9_9;
	wire [WIDTH-1:0] wire_d9_10;
	wire [WIDTH-1:0] wire_d9_11;
	wire [WIDTH-1:0] wire_d9_12;
	wire [WIDTH-1:0] wire_d9_13;
	wire [WIDTH-1:0] wire_d9_14;
	wire [WIDTH-1:0] wire_d9_15;
	wire [WIDTH-1:0] wire_d9_16;
	wire [WIDTH-1:0] wire_d9_17;
	wire [WIDTH-1:0] wire_d9_18;
	wire [WIDTH-1:0] wire_d9_19;
	wire [WIDTH-1:0] wire_d9_20;
	wire [WIDTH-1:0] wire_d9_21;
	wire [WIDTH-1:0] wire_d9_22;
	wire [WIDTH-1:0] wire_d9_23;
	wire [WIDTH-1:0] wire_d9_24;
	wire [WIDTH-1:0] wire_d9_25;
	wire [WIDTH-1:0] wire_d9_26;
	wire [WIDTH-1:0] wire_d9_27;
	wire [WIDTH-1:0] wire_d9_28;
	wire [WIDTH-1:0] wire_d9_29;
	wire [WIDTH-1:0] wire_d9_30;
	wire [WIDTH-1:0] wire_d9_31;
	wire [WIDTH-1:0] wire_d9_32;
	wire [WIDTH-1:0] wire_d9_33;
	wire [WIDTH-1:0] wire_d9_34;
	wire [WIDTH-1:0] wire_d9_35;
	wire [WIDTH-1:0] wire_d9_36;
	wire [WIDTH-1:0] wire_d9_37;
	wire [WIDTH-1:0] wire_d9_38;
	wire [WIDTH-1:0] wire_d9_39;
	wire [WIDTH-1:0] wire_d9_40;
	wire [WIDTH-1:0] wire_d9_41;
	wire [WIDTH-1:0] wire_d9_42;
	wire [WIDTH-1:0] wire_d9_43;
	wire [WIDTH-1:0] wire_d9_44;
	wire [WIDTH-1:0] wire_d9_45;
	wire [WIDTH-1:0] wire_d9_46;
	wire [WIDTH-1:0] wire_d9_47;
	wire [WIDTH-1:0] wire_d9_48;
	wire [WIDTH-1:0] wire_d9_49;
	wire [WIDTH-1:0] wire_d9_50;
	wire [WIDTH-1:0] wire_d9_51;
	wire [WIDTH-1:0] wire_d9_52;
	wire [WIDTH-1:0] wire_d9_53;
	wire [WIDTH-1:0] wire_d9_54;
	wire [WIDTH-1:0] wire_d9_55;
	wire [WIDTH-1:0] wire_d9_56;
	wire [WIDTH-1:0] wire_d9_57;
	wire [WIDTH-1:0] wire_d9_58;
	wire [WIDTH-1:0] wire_d9_59;
	wire [WIDTH-1:0] wire_d9_60;
	wire [WIDTH-1:0] wire_d9_61;
	wire [WIDTH-1:0] wire_d9_62;
	wire [WIDTH-1:0] wire_d9_63;
	wire [WIDTH-1:0] wire_d9_64;
	wire [WIDTH-1:0] wire_d9_65;
	wire [WIDTH-1:0] wire_d9_66;
	wire [WIDTH-1:0] wire_d9_67;
	wire [WIDTH-1:0] wire_d9_68;
	wire [WIDTH-1:0] wire_d9_69;
	wire [WIDTH-1:0] wire_d9_70;
	wire [WIDTH-1:0] wire_d9_71;
	wire [WIDTH-1:0] wire_d9_72;
	wire [WIDTH-1:0] wire_d9_73;
	wire [WIDTH-1:0] wire_d9_74;
	wire [WIDTH-1:0] wire_d9_75;
	wire [WIDTH-1:0] wire_d9_76;
	wire [WIDTH-1:0] wire_d9_77;
	wire [WIDTH-1:0] wire_d9_78;
	wire [WIDTH-1:0] wire_d10_0;
	wire [WIDTH-1:0] wire_d10_1;
	wire [WIDTH-1:0] wire_d10_2;
	wire [WIDTH-1:0] wire_d10_3;
	wire [WIDTH-1:0] wire_d10_4;
	wire [WIDTH-1:0] wire_d10_5;
	wire [WIDTH-1:0] wire_d10_6;
	wire [WIDTH-1:0] wire_d10_7;
	wire [WIDTH-1:0] wire_d10_8;
	wire [WIDTH-1:0] wire_d10_9;
	wire [WIDTH-1:0] wire_d10_10;
	wire [WIDTH-1:0] wire_d10_11;
	wire [WIDTH-1:0] wire_d10_12;
	wire [WIDTH-1:0] wire_d10_13;
	wire [WIDTH-1:0] wire_d10_14;
	wire [WIDTH-1:0] wire_d10_15;
	wire [WIDTH-1:0] wire_d10_16;
	wire [WIDTH-1:0] wire_d10_17;
	wire [WIDTH-1:0] wire_d10_18;
	wire [WIDTH-1:0] wire_d10_19;
	wire [WIDTH-1:0] wire_d10_20;
	wire [WIDTH-1:0] wire_d10_21;
	wire [WIDTH-1:0] wire_d10_22;
	wire [WIDTH-1:0] wire_d10_23;
	wire [WIDTH-1:0] wire_d10_24;
	wire [WIDTH-1:0] wire_d10_25;
	wire [WIDTH-1:0] wire_d10_26;
	wire [WIDTH-1:0] wire_d10_27;
	wire [WIDTH-1:0] wire_d10_28;
	wire [WIDTH-1:0] wire_d10_29;
	wire [WIDTH-1:0] wire_d10_30;
	wire [WIDTH-1:0] wire_d10_31;
	wire [WIDTH-1:0] wire_d10_32;
	wire [WIDTH-1:0] wire_d10_33;
	wire [WIDTH-1:0] wire_d10_34;
	wire [WIDTH-1:0] wire_d10_35;
	wire [WIDTH-1:0] wire_d10_36;
	wire [WIDTH-1:0] wire_d10_37;
	wire [WIDTH-1:0] wire_d10_38;
	wire [WIDTH-1:0] wire_d10_39;
	wire [WIDTH-1:0] wire_d10_40;
	wire [WIDTH-1:0] wire_d10_41;
	wire [WIDTH-1:0] wire_d10_42;
	wire [WIDTH-1:0] wire_d10_43;
	wire [WIDTH-1:0] wire_d10_44;
	wire [WIDTH-1:0] wire_d10_45;
	wire [WIDTH-1:0] wire_d10_46;
	wire [WIDTH-1:0] wire_d10_47;
	wire [WIDTH-1:0] wire_d10_48;
	wire [WIDTH-1:0] wire_d10_49;
	wire [WIDTH-1:0] wire_d10_50;
	wire [WIDTH-1:0] wire_d10_51;
	wire [WIDTH-1:0] wire_d10_52;
	wire [WIDTH-1:0] wire_d10_53;
	wire [WIDTH-1:0] wire_d10_54;
	wire [WIDTH-1:0] wire_d10_55;
	wire [WIDTH-1:0] wire_d10_56;
	wire [WIDTH-1:0] wire_d10_57;
	wire [WIDTH-1:0] wire_d10_58;
	wire [WIDTH-1:0] wire_d10_59;
	wire [WIDTH-1:0] wire_d10_60;
	wire [WIDTH-1:0] wire_d10_61;
	wire [WIDTH-1:0] wire_d10_62;
	wire [WIDTH-1:0] wire_d10_63;
	wire [WIDTH-1:0] wire_d10_64;
	wire [WIDTH-1:0] wire_d10_65;
	wire [WIDTH-1:0] wire_d10_66;
	wire [WIDTH-1:0] wire_d10_67;
	wire [WIDTH-1:0] wire_d10_68;
	wire [WIDTH-1:0] wire_d10_69;
	wire [WIDTH-1:0] wire_d10_70;
	wire [WIDTH-1:0] wire_d10_71;
	wire [WIDTH-1:0] wire_d10_72;
	wire [WIDTH-1:0] wire_d10_73;
	wire [WIDTH-1:0] wire_d10_74;
	wire [WIDTH-1:0] wire_d10_75;
	wire [WIDTH-1:0] wire_d10_76;
	wire [WIDTH-1:0] wire_d10_77;
	wire [WIDTH-1:0] wire_d10_78;
	wire [WIDTH-1:0] wire_d11_0;
	wire [WIDTH-1:0] wire_d11_1;
	wire [WIDTH-1:0] wire_d11_2;
	wire [WIDTH-1:0] wire_d11_3;
	wire [WIDTH-1:0] wire_d11_4;
	wire [WIDTH-1:0] wire_d11_5;
	wire [WIDTH-1:0] wire_d11_6;
	wire [WIDTH-1:0] wire_d11_7;
	wire [WIDTH-1:0] wire_d11_8;
	wire [WIDTH-1:0] wire_d11_9;
	wire [WIDTH-1:0] wire_d11_10;
	wire [WIDTH-1:0] wire_d11_11;
	wire [WIDTH-1:0] wire_d11_12;
	wire [WIDTH-1:0] wire_d11_13;
	wire [WIDTH-1:0] wire_d11_14;
	wire [WIDTH-1:0] wire_d11_15;
	wire [WIDTH-1:0] wire_d11_16;
	wire [WIDTH-1:0] wire_d11_17;
	wire [WIDTH-1:0] wire_d11_18;
	wire [WIDTH-1:0] wire_d11_19;
	wire [WIDTH-1:0] wire_d11_20;
	wire [WIDTH-1:0] wire_d11_21;
	wire [WIDTH-1:0] wire_d11_22;
	wire [WIDTH-1:0] wire_d11_23;
	wire [WIDTH-1:0] wire_d11_24;
	wire [WIDTH-1:0] wire_d11_25;
	wire [WIDTH-1:0] wire_d11_26;
	wire [WIDTH-1:0] wire_d11_27;
	wire [WIDTH-1:0] wire_d11_28;
	wire [WIDTH-1:0] wire_d11_29;
	wire [WIDTH-1:0] wire_d11_30;
	wire [WIDTH-1:0] wire_d11_31;
	wire [WIDTH-1:0] wire_d11_32;
	wire [WIDTH-1:0] wire_d11_33;
	wire [WIDTH-1:0] wire_d11_34;
	wire [WIDTH-1:0] wire_d11_35;
	wire [WIDTH-1:0] wire_d11_36;
	wire [WIDTH-1:0] wire_d11_37;
	wire [WIDTH-1:0] wire_d11_38;
	wire [WIDTH-1:0] wire_d11_39;
	wire [WIDTH-1:0] wire_d11_40;
	wire [WIDTH-1:0] wire_d11_41;
	wire [WIDTH-1:0] wire_d11_42;
	wire [WIDTH-1:0] wire_d11_43;
	wire [WIDTH-1:0] wire_d11_44;
	wire [WIDTH-1:0] wire_d11_45;
	wire [WIDTH-1:0] wire_d11_46;
	wire [WIDTH-1:0] wire_d11_47;
	wire [WIDTH-1:0] wire_d11_48;
	wire [WIDTH-1:0] wire_d11_49;
	wire [WIDTH-1:0] wire_d11_50;
	wire [WIDTH-1:0] wire_d11_51;
	wire [WIDTH-1:0] wire_d11_52;
	wire [WIDTH-1:0] wire_d11_53;
	wire [WIDTH-1:0] wire_d11_54;
	wire [WIDTH-1:0] wire_d11_55;
	wire [WIDTH-1:0] wire_d11_56;
	wire [WIDTH-1:0] wire_d11_57;
	wire [WIDTH-1:0] wire_d11_58;
	wire [WIDTH-1:0] wire_d11_59;
	wire [WIDTH-1:0] wire_d11_60;
	wire [WIDTH-1:0] wire_d11_61;
	wire [WIDTH-1:0] wire_d11_62;
	wire [WIDTH-1:0] wire_d11_63;
	wire [WIDTH-1:0] wire_d11_64;
	wire [WIDTH-1:0] wire_d11_65;
	wire [WIDTH-1:0] wire_d11_66;
	wire [WIDTH-1:0] wire_d11_67;
	wire [WIDTH-1:0] wire_d11_68;
	wire [WIDTH-1:0] wire_d11_69;
	wire [WIDTH-1:0] wire_d11_70;
	wire [WIDTH-1:0] wire_d11_71;
	wire [WIDTH-1:0] wire_d11_72;
	wire [WIDTH-1:0] wire_d11_73;
	wire [WIDTH-1:0] wire_d11_74;
	wire [WIDTH-1:0] wire_d11_75;
	wire [WIDTH-1:0] wire_d11_76;
	wire [WIDTH-1:0] wire_d11_77;
	wire [WIDTH-1:0] wire_d11_78;
	wire [WIDTH-1:0] wire_d12_0;
	wire [WIDTH-1:0] wire_d12_1;
	wire [WIDTH-1:0] wire_d12_2;
	wire [WIDTH-1:0] wire_d12_3;
	wire [WIDTH-1:0] wire_d12_4;
	wire [WIDTH-1:0] wire_d12_5;
	wire [WIDTH-1:0] wire_d12_6;
	wire [WIDTH-1:0] wire_d12_7;
	wire [WIDTH-1:0] wire_d12_8;
	wire [WIDTH-1:0] wire_d12_9;
	wire [WIDTH-1:0] wire_d12_10;
	wire [WIDTH-1:0] wire_d12_11;
	wire [WIDTH-1:0] wire_d12_12;
	wire [WIDTH-1:0] wire_d12_13;
	wire [WIDTH-1:0] wire_d12_14;
	wire [WIDTH-1:0] wire_d12_15;
	wire [WIDTH-1:0] wire_d12_16;
	wire [WIDTH-1:0] wire_d12_17;
	wire [WIDTH-1:0] wire_d12_18;
	wire [WIDTH-1:0] wire_d12_19;
	wire [WIDTH-1:0] wire_d12_20;
	wire [WIDTH-1:0] wire_d12_21;
	wire [WIDTH-1:0] wire_d12_22;
	wire [WIDTH-1:0] wire_d12_23;
	wire [WIDTH-1:0] wire_d12_24;
	wire [WIDTH-1:0] wire_d12_25;
	wire [WIDTH-1:0] wire_d12_26;
	wire [WIDTH-1:0] wire_d12_27;
	wire [WIDTH-1:0] wire_d12_28;
	wire [WIDTH-1:0] wire_d12_29;
	wire [WIDTH-1:0] wire_d12_30;
	wire [WIDTH-1:0] wire_d12_31;
	wire [WIDTH-1:0] wire_d12_32;
	wire [WIDTH-1:0] wire_d12_33;
	wire [WIDTH-1:0] wire_d12_34;
	wire [WIDTH-1:0] wire_d12_35;
	wire [WIDTH-1:0] wire_d12_36;
	wire [WIDTH-1:0] wire_d12_37;
	wire [WIDTH-1:0] wire_d12_38;
	wire [WIDTH-1:0] wire_d12_39;
	wire [WIDTH-1:0] wire_d12_40;
	wire [WIDTH-1:0] wire_d12_41;
	wire [WIDTH-1:0] wire_d12_42;
	wire [WIDTH-1:0] wire_d12_43;
	wire [WIDTH-1:0] wire_d12_44;
	wire [WIDTH-1:0] wire_d12_45;
	wire [WIDTH-1:0] wire_d12_46;
	wire [WIDTH-1:0] wire_d12_47;
	wire [WIDTH-1:0] wire_d12_48;
	wire [WIDTH-1:0] wire_d12_49;
	wire [WIDTH-1:0] wire_d12_50;
	wire [WIDTH-1:0] wire_d12_51;
	wire [WIDTH-1:0] wire_d12_52;
	wire [WIDTH-1:0] wire_d12_53;
	wire [WIDTH-1:0] wire_d12_54;
	wire [WIDTH-1:0] wire_d12_55;
	wire [WIDTH-1:0] wire_d12_56;
	wire [WIDTH-1:0] wire_d12_57;
	wire [WIDTH-1:0] wire_d12_58;
	wire [WIDTH-1:0] wire_d12_59;
	wire [WIDTH-1:0] wire_d12_60;
	wire [WIDTH-1:0] wire_d12_61;
	wire [WIDTH-1:0] wire_d12_62;
	wire [WIDTH-1:0] wire_d12_63;
	wire [WIDTH-1:0] wire_d12_64;
	wire [WIDTH-1:0] wire_d12_65;
	wire [WIDTH-1:0] wire_d12_66;
	wire [WIDTH-1:0] wire_d12_67;
	wire [WIDTH-1:0] wire_d12_68;
	wire [WIDTH-1:0] wire_d12_69;
	wire [WIDTH-1:0] wire_d12_70;
	wire [WIDTH-1:0] wire_d12_71;
	wire [WIDTH-1:0] wire_d12_72;
	wire [WIDTH-1:0] wire_d12_73;
	wire [WIDTH-1:0] wire_d12_74;
	wire [WIDTH-1:0] wire_d12_75;
	wire [WIDTH-1:0] wire_d12_76;
	wire [WIDTH-1:0] wire_d12_77;
	wire [WIDTH-1:0] wire_d12_78;
	wire [WIDTH-1:0] wire_d13_0;
	wire [WIDTH-1:0] wire_d13_1;
	wire [WIDTH-1:0] wire_d13_2;
	wire [WIDTH-1:0] wire_d13_3;
	wire [WIDTH-1:0] wire_d13_4;
	wire [WIDTH-1:0] wire_d13_5;
	wire [WIDTH-1:0] wire_d13_6;
	wire [WIDTH-1:0] wire_d13_7;
	wire [WIDTH-1:0] wire_d13_8;
	wire [WIDTH-1:0] wire_d13_9;
	wire [WIDTH-1:0] wire_d13_10;
	wire [WIDTH-1:0] wire_d13_11;
	wire [WIDTH-1:0] wire_d13_12;
	wire [WIDTH-1:0] wire_d13_13;
	wire [WIDTH-1:0] wire_d13_14;
	wire [WIDTH-1:0] wire_d13_15;
	wire [WIDTH-1:0] wire_d13_16;
	wire [WIDTH-1:0] wire_d13_17;
	wire [WIDTH-1:0] wire_d13_18;
	wire [WIDTH-1:0] wire_d13_19;
	wire [WIDTH-1:0] wire_d13_20;
	wire [WIDTH-1:0] wire_d13_21;
	wire [WIDTH-1:0] wire_d13_22;
	wire [WIDTH-1:0] wire_d13_23;
	wire [WIDTH-1:0] wire_d13_24;
	wire [WIDTH-1:0] wire_d13_25;
	wire [WIDTH-1:0] wire_d13_26;
	wire [WIDTH-1:0] wire_d13_27;
	wire [WIDTH-1:0] wire_d13_28;
	wire [WIDTH-1:0] wire_d13_29;
	wire [WIDTH-1:0] wire_d13_30;
	wire [WIDTH-1:0] wire_d13_31;
	wire [WIDTH-1:0] wire_d13_32;
	wire [WIDTH-1:0] wire_d13_33;
	wire [WIDTH-1:0] wire_d13_34;
	wire [WIDTH-1:0] wire_d13_35;
	wire [WIDTH-1:0] wire_d13_36;
	wire [WIDTH-1:0] wire_d13_37;
	wire [WIDTH-1:0] wire_d13_38;
	wire [WIDTH-1:0] wire_d13_39;
	wire [WIDTH-1:0] wire_d13_40;
	wire [WIDTH-1:0] wire_d13_41;
	wire [WIDTH-1:0] wire_d13_42;
	wire [WIDTH-1:0] wire_d13_43;
	wire [WIDTH-1:0] wire_d13_44;
	wire [WIDTH-1:0] wire_d13_45;
	wire [WIDTH-1:0] wire_d13_46;
	wire [WIDTH-1:0] wire_d13_47;
	wire [WIDTH-1:0] wire_d13_48;
	wire [WIDTH-1:0] wire_d13_49;
	wire [WIDTH-1:0] wire_d13_50;
	wire [WIDTH-1:0] wire_d13_51;
	wire [WIDTH-1:0] wire_d13_52;
	wire [WIDTH-1:0] wire_d13_53;
	wire [WIDTH-1:0] wire_d13_54;
	wire [WIDTH-1:0] wire_d13_55;
	wire [WIDTH-1:0] wire_d13_56;
	wire [WIDTH-1:0] wire_d13_57;
	wire [WIDTH-1:0] wire_d13_58;
	wire [WIDTH-1:0] wire_d13_59;
	wire [WIDTH-1:0] wire_d13_60;
	wire [WIDTH-1:0] wire_d13_61;
	wire [WIDTH-1:0] wire_d13_62;
	wire [WIDTH-1:0] wire_d13_63;
	wire [WIDTH-1:0] wire_d13_64;
	wire [WIDTH-1:0] wire_d13_65;
	wire [WIDTH-1:0] wire_d13_66;
	wire [WIDTH-1:0] wire_d13_67;
	wire [WIDTH-1:0] wire_d13_68;
	wire [WIDTH-1:0] wire_d13_69;
	wire [WIDTH-1:0] wire_d13_70;
	wire [WIDTH-1:0] wire_d13_71;
	wire [WIDTH-1:0] wire_d13_72;
	wire [WIDTH-1:0] wire_d13_73;
	wire [WIDTH-1:0] wire_d13_74;
	wire [WIDTH-1:0] wire_d13_75;
	wire [WIDTH-1:0] wire_d13_76;
	wire [WIDTH-1:0] wire_d13_77;
	wire [WIDTH-1:0] wire_d13_78;
	wire [WIDTH-1:0] wire_d14_0;
	wire [WIDTH-1:0] wire_d14_1;
	wire [WIDTH-1:0] wire_d14_2;
	wire [WIDTH-1:0] wire_d14_3;
	wire [WIDTH-1:0] wire_d14_4;
	wire [WIDTH-1:0] wire_d14_5;
	wire [WIDTH-1:0] wire_d14_6;
	wire [WIDTH-1:0] wire_d14_7;
	wire [WIDTH-1:0] wire_d14_8;
	wire [WIDTH-1:0] wire_d14_9;
	wire [WIDTH-1:0] wire_d14_10;
	wire [WIDTH-1:0] wire_d14_11;
	wire [WIDTH-1:0] wire_d14_12;
	wire [WIDTH-1:0] wire_d14_13;
	wire [WIDTH-1:0] wire_d14_14;
	wire [WIDTH-1:0] wire_d14_15;
	wire [WIDTH-1:0] wire_d14_16;
	wire [WIDTH-1:0] wire_d14_17;
	wire [WIDTH-1:0] wire_d14_18;
	wire [WIDTH-1:0] wire_d14_19;
	wire [WIDTH-1:0] wire_d14_20;
	wire [WIDTH-1:0] wire_d14_21;
	wire [WIDTH-1:0] wire_d14_22;
	wire [WIDTH-1:0] wire_d14_23;
	wire [WIDTH-1:0] wire_d14_24;
	wire [WIDTH-1:0] wire_d14_25;
	wire [WIDTH-1:0] wire_d14_26;
	wire [WIDTH-1:0] wire_d14_27;
	wire [WIDTH-1:0] wire_d14_28;
	wire [WIDTH-1:0] wire_d14_29;
	wire [WIDTH-1:0] wire_d14_30;
	wire [WIDTH-1:0] wire_d14_31;
	wire [WIDTH-1:0] wire_d14_32;
	wire [WIDTH-1:0] wire_d14_33;
	wire [WIDTH-1:0] wire_d14_34;
	wire [WIDTH-1:0] wire_d14_35;
	wire [WIDTH-1:0] wire_d14_36;
	wire [WIDTH-1:0] wire_d14_37;
	wire [WIDTH-1:0] wire_d14_38;
	wire [WIDTH-1:0] wire_d14_39;
	wire [WIDTH-1:0] wire_d14_40;
	wire [WIDTH-1:0] wire_d14_41;
	wire [WIDTH-1:0] wire_d14_42;
	wire [WIDTH-1:0] wire_d14_43;
	wire [WIDTH-1:0] wire_d14_44;
	wire [WIDTH-1:0] wire_d14_45;
	wire [WIDTH-1:0] wire_d14_46;
	wire [WIDTH-1:0] wire_d14_47;
	wire [WIDTH-1:0] wire_d14_48;
	wire [WIDTH-1:0] wire_d14_49;
	wire [WIDTH-1:0] wire_d14_50;
	wire [WIDTH-1:0] wire_d14_51;
	wire [WIDTH-1:0] wire_d14_52;
	wire [WIDTH-1:0] wire_d14_53;
	wire [WIDTH-1:0] wire_d14_54;
	wire [WIDTH-1:0] wire_d14_55;
	wire [WIDTH-1:0] wire_d14_56;
	wire [WIDTH-1:0] wire_d14_57;
	wire [WIDTH-1:0] wire_d14_58;
	wire [WIDTH-1:0] wire_d14_59;
	wire [WIDTH-1:0] wire_d14_60;
	wire [WIDTH-1:0] wire_d14_61;
	wire [WIDTH-1:0] wire_d14_62;
	wire [WIDTH-1:0] wire_d14_63;
	wire [WIDTH-1:0] wire_d14_64;
	wire [WIDTH-1:0] wire_d14_65;
	wire [WIDTH-1:0] wire_d14_66;
	wire [WIDTH-1:0] wire_d14_67;
	wire [WIDTH-1:0] wire_d14_68;
	wire [WIDTH-1:0] wire_d14_69;
	wire [WIDTH-1:0] wire_d14_70;
	wire [WIDTH-1:0] wire_d14_71;
	wire [WIDTH-1:0] wire_d14_72;
	wire [WIDTH-1:0] wire_d14_73;
	wire [WIDTH-1:0] wire_d14_74;
	wire [WIDTH-1:0] wire_d14_75;
	wire [WIDTH-1:0] wire_d14_76;
	wire [WIDTH-1:0] wire_d14_77;
	wire [WIDTH-1:0] wire_d14_78;
	wire [WIDTH-1:0] wire_d15_0;
	wire [WIDTH-1:0] wire_d15_1;
	wire [WIDTH-1:0] wire_d15_2;
	wire [WIDTH-1:0] wire_d15_3;
	wire [WIDTH-1:0] wire_d15_4;
	wire [WIDTH-1:0] wire_d15_5;
	wire [WIDTH-1:0] wire_d15_6;
	wire [WIDTH-1:0] wire_d15_7;
	wire [WIDTH-1:0] wire_d15_8;
	wire [WIDTH-1:0] wire_d15_9;
	wire [WIDTH-1:0] wire_d15_10;
	wire [WIDTH-1:0] wire_d15_11;
	wire [WIDTH-1:0] wire_d15_12;
	wire [WIDTH-1:0] wire_d15_13;
	wire [WIDTH-1:0] wire_d15_14;
	wire [WIDTH-1:0] wire_d15_15;
	wire [WIDTH-1:0] wire_d15_16;
	wire [WIDTH-1:0] wire_d15_17;
	wire [WIDTH-1:0] wire_d15_18;
	wire [WIDTH-1:0] wire_d15_19;
	wire [WIDTH-1:0] wire_d15_20;
	wire [WIDTH-1:0] wire_d15_21;
	wire [WIDTH-1:0] wire_d15_22;
	wire [WIDTH-1:0] wire_d15_23;
	wire [WIDTH-1:0] wire_d15_24;
	wire [WIDTH-1:0] wire_d15_25;
	wire [WIDTH-1:0] wire_d15_26;
	wire [WIDTH-1:0] wire_d15_27;
	wire [WIDTH-1:0] wire_d15_28;
	wire [WIDTH-1:0] wire_d15_29;
	wire [WIDTH-1:0] wire_d15_30;
	wire [WIDTH-1:0] wire_d15_31;
	wire [WIDTH-1:0] wire_d15_32;
	wire [WIDTH-1:0] wire_d15_33;
	wire [WIDTH-1:0] wire_d15_34;
	wire [WIDTH-1:0] wire_d15_35;
	wire [WIDTH-1:0] wire_d15_36;
	wire [WIDTH-1:0] wire_d15_37;
	wire [WIDTH-1:0] wire_d15_38;
	wire [WIDTH-1:0] wire_d15_39;
	wire [WIDTH-1:0] wire_d15_40;
	wire [WIDTH-1:0] wire_d15_41;
	wire [WIDTH-1:0] wire_d15_42;
	wire [WIDTH-1:0] wire_d15_43;
	wire [WIDTH-1:0] wire_d15_44;
	wire [WIDTH-1:0] wire_d15_45;
	wire [WIDTH-1:0] wire_d15_46;
	wire [WIDTH-1:0] wire_d15_47;
	wire [WIDTH-1:0] wire_d15_48;
	wire [WIDTH-1:0] wire_d15_49;
	wire [WIDTH-1:0] wire_d15_50;
	wire [WIDTH-1:0] wire_d15_51;
	wire [WIDTH-1:0] wire_d15_52;
	wire [WIDTH-1:0] wire_d15_53;
	wire [WIDTH-1:0] wire_d15_54;
	wire [WIDTH-1:0] wire_d15_55;
	wire [WIDTH-1:0] wire_d15_56;
	wire [WIDTH-1:0] wire_d15_57;
	wire [WIDTH-1:0] wire_d15_58;
	wire [WIDTH-1:0] wire_d15_59;
	wire [WIDTH-1:0] wire_d15_60;
	wire [WIDTH-1:0] wire_d15_61;
	wire [WIDTH-1:0] wire_d15_62;
	wire [WIDTH-1:0] wire_d15_63;
	wire [WIDTH-1:0] wire_d15_64;
	wire [WIDTH-1:0] wire_d15_65;
	wire [WIDTH-1:0] wire_d15_66;
	wire [WIDTH-1:0] wire_d15_67;
	wire [WIDTH-1:0] wire_d15_68;
	wire [WIDTH-1:0] wire_d15_69;
	wire [WIDTH-1:0] wire_d15_70;
	wire [WIDTH-1:0] wire_d15_71;
	wire [WIDTH-1:0] wire_d15_72;
	wire [WIDTH-1:0] wire_d15_73;
	wire [WIDTH-1:0] wire_d15_74;
	wire [WIDTH-1:0] wire_d15_75;
	wire [WIDTH-1:0] wire_d15_76;
	wire [WIDTH-1:0] wire_d15_77;
	wire [WIDTH-1:0] wire_d15_78;
	wire [WIDTH-1:0] wire_d16_0;
	wire [WIDTH-1:0] wire_d16_1;
	wire [WIDTH-1:0] wire_d16_2;
	wire [WIDTH-1:0] wire_d16_3;
	wire [WIDTH-1:0] wire_d16_4;
	wire [WIDTH-1:0] wire_d16_5;
	wire [WIDTH-1:0] wire_d16_6;
	wire [WIDTH-1:0] wire_d16_7;
	wire [WIDTH-1:0] wire_d16_8;
	wire [WIDTH-1:0] wire_d16_9;
	wire [WIDTH-1:0] wire_d16_10;
	wire [WIDTH-1:0] wire_d16_11;
	wire [WIDTH-1:0] wire_d16_12;
	wire [WIDTH-1:0] wire_d16_13;
	wire [WIDTH-1:0] wire_d16_14;
	wire [WIDTH-1:0] wire_d16_15;
	wire [WIDTH-1:0] wire_d16_16;
	wire [WIDTH-1:0] wire_d16_17;
	wire [WIDTH-1:0] wire_d16_18;
	wire [WIDTH-1:0] wire_d16_19;
	wire [WIDTH-1:0] wire_d16_20;
	wire [WIDTH-1:0] wire_d16_21;
	wire [WIDTH-1:0] wire_d16_22;
	wire [WIDTH-1:0] wire_d16_23;
	wire [WIDTH-1:0] wire_d16_24;
	wire [WIDTH-1:0] wire_d16_25;
	wire [WIDTH-1:0] wire_d16_26;
	wire [WIDTH-1:0] wire_d16_27;
	wire [WIDTH-1:0] wire_d16_28;
	wire [WIDTH-1:0] wire_d16_29;
	wire [WIDTH-1:0] wire_d16_30;
	wire [WIDTH-1:0] wire_d16_31;
	wire [WIDTH-1:0] wire_d16_32;
	wire [WIDTH-1:0] wire_d16_33;
	wire [WIDTH-1:0] wire_d16_34;
	wire [WIDTH-1:0] wire_d16_35;
	wire [WIDTH-1:0] wire_d16_36;
	wire [WIDTH-1:0] wire_d16_37;
	wire [WIDTH-1:0] wire_d16_38;
	wire [WIDTH-1:0] wire_d16_39;
	wire [WIDTH-1:0] wire_d16_40;
	wire [WIDTH-1:0] wire_d16_41;
	wire [WIDTH-1:0] wire_d16_42;
	wire [WIDTH-1:0] wire_d16_43;
	wire [WIDTH-1:0] wire_d16_44;
	wire [WIDTH-1:0] wire_d16_45;
	wire [WIDTH-1:0] wire_d16_46;
	wire [WIDTH-1:0] wire_d16_47;
	wire [WIDTH-1:0] wire_d16_48;
	wire [WIDTH-1:0] wire_d16_49;
	wire [WIDTH-1:0] wire_d16_50;
	wire [WIDTH-1:0] wire_d16_51;
	wire [WIDTH-1:0] wire_d16_52;
	wire [WIDTH-1:0] wire_d16_53;
	wire [WIDTH-1:0] wire_d16_54;
	wire [WIDTH-1:0] wire_d16_55;
	wire [WIDTH-1:0] wire_d16_56;
	wire [WIDTH-1:0] wire_d16_57;
	wire [WIDTH-1:0] wire_d16_58;
	wire [WIDTH-1:0] wire_d16_59;
	wire [WIDTH-1:0] wire_d16_60;
	wire [WIDTH-1:0] wire_d16_61;
	wire [WIDTH-1:0] wire_d16_62;
	wire [WIDTH-1:0] wire_d16_63;
	wire [WIDTH-1:0] wire_d16_64;
	wire [WIDTH-1:0] wire_d16_65;
	wire [WIDTH-1:0] wire_d16_66;
	wire [WIDTH-1:0] wire_d16_67;
	wire [WIDTH-1:0] wire_d16_68;
	wire [WIDTH-1:0] wire_d16_69;
	wire [WIDTH-1:0] wire_d16_70;
	wire [WIDTH-1:0] wire_d16_71;
	wire [WIDTH-1:0] wire_d16_72;
	wire [WIDTH-1:0] wire_d16_73;
	wire [WIDTH-1:0] wire_d16_74;
	wire [WIDTH-1:0] wire_d16_75;
	wire [WIDTH-1:0] wire_d16_76;
	wire [WIDTH-1:0] wire_d16_77;
	wire [WIDTH-1:0] wire_d16_78;
	wire [WIDTH-1:0] wire_d17_0;
	wire [WIDTH-1:0] wire_d17_1;
	wire [WIDTH-1:0] wire_d17_2;
	wire [WIDTH-1:0] wire_d17_3;
	wire [WIDTH-1:0] wire_d17_4;
	wire [WIDTH-1:0] wire_d17_5;
	wire [WIDTH-1:0] wire_d17_6;
	wire [WIDTH-1:0] wire_d17_7;
	wire [WIDTH-1:0] wire_d17_8;
	wire [WIDTH-1:0] wire_d17_9;
	wire [WIDTH-1:0] wire_d17_10;
	wire [WIDTH-1:0] wire_d17_11;
	wire [WIDTH-1:0] wire_d17_12;
	wire [WIDTH-1:0] wire_d17_13;
	wire [WIDTH-1:0] wire_d17_14;
	wire [WIDTH-1:0] wire_d17_15;
	wire [WIDTH-1:0] wire_d17_16;
	wire [WIDTH-1:0] wire_d17_17;
	wire [WIDTH-1:0] wire_d17_18;
	wire [WIDTH-1:0] wire_d17_19;
	wire [WIDTH-1:0] wire_d17_20;
	wire [WIDTH-1:0] wire_d17_21;
	wire [WIDTH-1:0] wire_d17_22;
	wire [WIDTH-1:0] wire_d17_23;
	wire [WIDTH-1:0] wire_d17_24;
	wire [WIDTH-1:0] wire_d17_25;
	wire [WIDTH-1:0] wire_d17_26;
	wire [WIDTH-1:0] wire_d17_27;
	wire [WIDTH-1:0] wire_d17_28;
	wire [WIDTH-1:0] wire_d17_29;
	wire [WIDTH-1:0] wire_d17_30;
	wire [WIDTH-1:0] wire_d17_31;
	wire [WIDTH-1:0] wire_d17_32;
	wire [WIDTH-1:0] wire_d17_33;
	wire [WIDTH-1:0] wire_d17_34;
	wire [WIDTH-1:0] wire_d17_35;
	wire [WIDTH-1:0] wire_d17_36;
	wire [WIDTH-1:0] wire_d17_37;
	wire [WIDTH-1:0] wire_d17_38;
	wire [WIDTH-1:0] wire_d17_39;
	wire [WIDTH-1:0] wire_d17_40;
	wire [WIDTH-1:0] wire_d17_41;
	wire [WIDTH-1:0] wire_d17_42;
	wire [WIDTH-1:0] wire_d17_43;
	wire [WIDTH-1:0] wire_d17_44;
	wire [WIDTH-1:0] wire_d17_45;
	wire [WIDTH-1:0] wire_d17_46;
	wire [WIDTH-1:0] wire_d17_47;
	wire [WIDTH-1:0] wire_d17_48;
	wire [WIDTH-1:0] wire_d17_49;
	wire [WIDTH-1:0] wire_d17_50;
	wire [WIDTH-1:0] wire_d17_51;
	wire [WIDTH-1:0] wire_d17_52;
	wire [WIDTH-1:0] wire_d17_53;
	wire [WIDTH-1:0] wire_d17_54;
	wire [WIDTH-1:0] wire_d17_55;
	wire [WIDTH-1:0] wire_d17_56;
	wire [WIDTH-1:0] wire_d17_57;
	wire [WIDTH-1:0] wire_d17_58;
	wire [WIDTH-1:0] wire_d17_59;
	wire [WIDTH-1:0] wire_d17_60;
	wire [WIDTH-1:0] wire_d17_61;
	wire [WIDTH-1:0] wire_d17_62;
	wire [WIDTH-1:0] wire_d17_63;
	wire [WIDTH-1:0] wire_d17_64;
	wire [WIDTH-1:0] wire_d17_65;
	wire [WIDTH-1:0] wire_d17_66;
	wire [WIDTH-1:0] wire_d17_67;
	wire [WIDTH-1:0] wire_d17_68;
	wire [WIDTH-1:0] wire_d17_69;
	wire [WIDTH-1:0] wire_d17_70;
	wire [WIDTH-1:0] wire_d17_71;
	wire [WIDTH-1:0] wire_d17_72;
	wire [WIDTH-1:0] wire_d17_73;
	wire [WIDTH-1:0] wire_d17_74;
	wire [WIDTH-1:0] wire_d17_75;
	wire [WIDTH-1:0] wire_d17_76;
	wire [WIDTH-1:0] wire_d17_77;
	wire [WIDTH-1:0] wire_d17_78;
	wire [WIDTH-1:0] wire_d18_0;
	wire [WIDTH-1:0] wire_d18_1;
	wire [WIDTH-1:0] wire_d18_2;
	wire [WIDTH-1:0] wire_d18_3;
	wire [WIDTH-1:0] wire_d18_4;
	wire [WIDTH-1:0] wire_d18_5;
	wire [WIDTH-1:0] wire_d18_6;
	wire [WIDTH-1:0] wire_d18_7;
	wire [WIDTH-1:0] wire_d18_8;
	wire [WIDTH-1:0] wire_d18_9;
	wire [WIDTH-1:0] wire_d18_10;
	wire [WIDTH-1:0] wire_d18_11;
	wire [WIDTH-1:0] wire_d18_12;
	wire [WIDTH-1:0] wire_d18_13;
	wire [WIDTH-1:0] wire_d18_14;
	wire [WIDTH-1:0] wire_d18_15;
	wire [WIDTH-1:0] wire_d18_16;
	wire [WIDTH-1:0] wire_d18_17;
	wire [WIDTH-1:0] wire_d18_18;
	wire [WIDTH-1:0] wire_d18_19;
	wire [WIDTH-1:0] wire_d18_20;
	wire [WIDTH-1:0] wire_d18_21;
	wire [WIDTH-1:0] wire_d18_22;
	wire [WIDTH-1:0] wire_d18_23;
	wire [WIDTH-1:0] wire_d18_24;
	wire [WIDTH-1:0] wire_d18_25;
	wire [WIDTH-1:0] wire_d18_26;
	wire [WIDTH-1:0] wire_d18_27;
	wire [WIDTH-1:0] wire_d18_28;
	wire [WIDTH-1:0] wire_d18_29;
	wire [WIDTH-1:0] wire_d18_30;
	wire [WIDTH-1:0] wire_d18_31;
	wire [WIDTH-1:0] wire_d18_32;
	wire [WIDTH-1:0] wire_d18_33;
	wire [WIDTH-1:0] wire_d18_34;
	wire [WIDTH-1:0] wire_d18_35;
	wire [WIDTH-1:0] wire_d18_36;
	wire [WIDTH-1:0] wire_d18_37;
	wire [WIDTH-1:0] wire_d18_38;
	wire [WIDTH-1:0] wire_d18_39;
	wire [WIDTH-1:0] wire_d18_40;
	wire [WIDTH-1:0] wire_d18_41;
	wire [WIDTH-1:0] wire_d18_42;
	wire [WIDTH-1:0] wire_d18_43;
	wire [WIDTH-1:0] wire_d18_44;
	wire [WIDTH-1:0] wire_d18_45;
	wire [WIDTH-1:0] wire_d18_46;
	wire [WIDTH-1:0] wire_d18_47;
	wire [WIDTH-1:0] wire_d18_48;
	wire [WIDTH-1:0] wire_d18_49;
	wire [WIDTH-1:0] wire_d18_50;
	wire [WIDTH-1:0] wire_d18_51;
	wire [WIDTH-1:0] wire_d18_52;
	wire [WIDTH-1:0] wire_d18_53;
	wire [WIDTH-1:0] wire_d18_54;
	wire [WIDTH-1:0] wire_d18_55;
	wire [WIDTH-1:0] wire_d18_56;
	wire [WIDTH-1:0] wire_d18_57;
	wire [WIDTH-1:0] wire_d18_58;
	wire [WIDTH-1:0] wire_d18_59;
	wire [WIDTH-1:0] wire_d18_60;
	wire [WIDTH-1:0] wire_d18_61;
	wire [WIDTH-1:0] wire_d18_62;
	wire [WIDTH-1:0] wire_d18_63;
	wire [WIDTH-1:0] wire_d18_64;
	wire [WIDTH-1:0] wire_d18_65;
	wire [WIDTH-1:0] wire_d18_66;
	wire [WIDTH-1:0] wire_d18_67;
	wire [WIDTH-1:0] wire_d18_68;
	wire [WIDTH-1:0] wire_d18_69;
	wire [WIDTH-1:0] wire_d18_70;
	wire [WIDTH-1:0] wire_d18_71;
	wire [WIDTH-1:0] wire_d18_72;
	wire [WIDTH-1:0] wire_d18_73;
	wire [WIDTH-1:0] wire_d18_74;
	wire [WIDTH-1:0] wire_d18_75;
	wire [WIDTH-1:0] wire_d18_76;
	wire [WIDTH-1:0] wire_d18_77;
	wire [WIDTH-1:0] wire_d18_78;
	wire [WIDTH-1:0] wire_d19_0;
	wire [WIDTH-1:0] wire_d19_1;
	wire [WIDTH-1:0] wire_d19_2;
	wire [WIDTH-1:0] wire_d19_3;
	wire [WIDTH-1:0] wire_d19_4;
	wire [WIDTH-1:0] wire_d19_5;
	wire [WIDTH-1:0] wire_d19_6;
	wire [WIDTH-1:0] wire_d19_7;
	wire [WIDTH-1:0] wire_d19_8;
	wire [WIDTH-1:0] wire_d19_9;
	wire [WIDTH-1:0] wire_d19_10;
	wire [WIDTH-1:0] wire_d19_11;
	wire [WIDTH-1:0] wire_d19_12;
	wire [WIDTH-1:0] wire_d19_13;
	wire [WIDTH-1:0] wire_d19_14;
	wire [WIDTH-1:0] wire_d19_15;
	wire [WIDTH-1:0] wire_d19_16;
	wire [WIDTH-1:0] wire_d19_17;
	wire [WIDTH-1:0] wire_d19_18;
	wire [WIDTH-1:0] wire_d19_19;
	wire [WIDTH-1:0] wire_d19_20;
	wire [WIDTH-1:0] wire_d19_21;
	wire [WIDTH-1:0] wire_d19_22;
	wire [WIDTH-1:0] wire_d19_23;
	wire [WIDTH-1:0] wire_d19_24;
	wire [WIDTH-1:0] wire_d19_25;
	wire [WIDTH-1:0] wire_d19_26;
	wire [WIDTH-1:0] wire_d19_27;
	wire [WIDTH-1:0] wire_d19_28;
	wire [WIDTH-1:0] wire_d19_29;
	wire [WIDTH-1:0] wire_d19_30;
	wire [WIDTH-1:0] wire_d19_31;
	wire [WIDTH-1:0] wire_d19_32;
	wire [WIDTH-1:0] wire_d19_33;
	wire [WIDTH-1:0] wire_d19_34;
	wire [WIDTH-1:0] wire_d19_35;
	wire [WIDTH-1:0] wire_d19_36;
	wire [WIDTH-1:0] wire_d19_37;
	wire [WIDTH-1:0] wire_d19_38;
	wire [WIDTH-1:0] wire_d19_39;
	wire [WIDTH-1:0] wire_d19_40;
	wire [WIDTH-1:0] wire_d19_41;
	wire [WIDTH-1:0] wire_d19_42;
	wire [WIDTH-1:0] wire_d19_43;
	wire [WIDTH-1:0] wire_d19_44;
	wire [WIDTH-1:0] wire_d19_45;
	wire [WIDTH-1:0] wire_d19_46;
	wire [WIDTH-1:0] wire_d19_47;
	wire [WIDTH-1:0] wire_d19_48;
	wire [WIDTH-1:0] wire_d19_49;
	wire [WIDTH-1:0] wire_d19_50;
	wire [WIDTH-1:0] wire_d19_51;
	wire [WIDTH-1:0] wire_d19_52;
	wire [WIDTH-1:0] wire_d19_53;
	wire [WIDTH-1:0] wire_d19_54;
	wire [WIDTH-1:0] wire_d19_55;
	wire [WIDTH-1:0] wire_d19_56;
	wire [WIDTH-1:0] wire_d19_57;
	wire [WIDTH-1:0] wire_d19_58;
	wire [WIDTH-1:0] wire_d19_59;
	wire [WIDTH-1:0] wire_d19_60;
	wire [WIDTH-1:0] wire_d19_61;
	wire [WIDTH-1:0] wire_d19_62;
	wire [WIDTH-1:0] wire_d19_63;
	wire [WIDTH-1:0] wire_d19_64;
	wire [WIDTH-1:0] wire_d19_65;
	wire [WIDTH-1:0] wire_d19_66;
	wire [WIDTH-1:0] wire_d19_67;
	wire [WIDTH-1:0] wire_d19_68;
	wire [WIDTH-1:0] wire_d19_69;
	wire [WIDTH-1:0] wire_d19_70;
	wire [WIDTH-1:0] wire_d19_71;
	wire [WIDTH-1:0] wire_d19_72;
	wire [WIDTH-1:0] wire_d19_73;
	wire [WIDTH-1:0] wire_d19_74;
	wire [WIDTH-1:0] wire_d19_75;
	wire [WIDTH-1:0] wire_d19_76;
	wire [WIDTH-1:0] wire_d19_77;
	wire [WIDTH-1:0] wire_d19_78;
	wire [WIDTH-1:0] wire_d20_0;
	wire [WIDTH-1:0] wire_d20_1;
	wire [WIDTH-1:0] wire_d20_2;
	wire [WIDTH-1:0] wire_d20_3;
	wire [WIDTH-1:0] wire_d20_4;
	wire [WIDTH-1:0] wire_d20_5;
	wire [WIDTH-1:0] wire_d20_6;
	wire [WIDTH-1:0] wire_d20_7;
	wire [WIDTH-1:0] wire_d20_8;
	wire [WIDTH-1:0] wire_d20_9;
	wire [WIDTH-1:0] wire_d20_10;
	wire [WIDTH-1:0] wire_d20_11;
	wire [WIDTH-1:0] wire_d20_12;
	wire [WIDTH-1:0] wire_d20_13;
	wire [WIDTH-1:0] wire_d20_14;
	wire [WIDTH-1:0] wire_d20_15;
	wire [WIDTH-1:0] wire_d20_16;
	wire [WIDTH-1:0] wire_d20_17;
	wire [WIDTH-1:0] wire_d20_18;
	wire [WIDTH-1:0] wire_d20_19;
	wire [WIDTH-1:0] wire_d20_20;
	wire [WIDTH-1:0] wire_d20_21;
	wire [WIDTH-1:0] wire_d20_22;
	wire [WIDTH-1:0] wire_d20_23;
	wire [WIDTH-1:0] wire_d20_24;
	wire [WIDTH-1:0] wire_d20_25;
	wire [WIDTH-1:0] wire_d20_26;
	wire [WIDTH-1:0] wire_d20_27;
	wire [WIDTH-1:0] wire_d20_28;
	wire [WIDTH-1:0] wire_d20_29;
	wire [WIDTH-1:0] wire_d20_30;
	wire [WIDTH-1:0] wire_d20_31;
	wire [WIDTH-1:0] wire_d20_32;
	wire [WIDTH-1:0] wire_d20_33;
	wire [WIDTH-1:0] wire_d20_34;
	wire [WIDTH-1:0] wire_d20_35;
	wire [WIDTH-1:0] wire_d20_36;
	wire [WIDTH-1:0] wire_d20_37;
	wire [WIDTH-1:0] wire_d20_38;
	wire [WIDTH-1:0] wire_d20_39;
	wire [WIDTH-1:0] wire_d20_40;
	wire [WIDTH-1:0] wire_d20_41;
	wire [WIDTH-1:0] wire_d20_42;
	wire [WIDTH-1:0] wire_d20_43;
	wire [WIDTH-1:0] wire_d20_44;
	wire [WIDTH-1:0] wire_d20_45;
	wire [WIDTH-1:0] wire_d20_46;
	wire [WIDTH-1:0] wire_d20_47;
	wire [WIDTH-1:0] wire_d20_48;
	wire [WIDTH-1:0] wire_d20_49;
	wire [WIDTH-1:0] wire_d20_50;
	wire [WIDTH-1:0] wire_d20_51;
	wire [WIDTH-1:0] wire_d20_52;
	wire [WIDTH-1:0] wire_d20_53;
	wire [WIDTH-1:0] wire_d20_54;
	wire [WIDTH-1:0] wire_d20_55;
	wire [WIDTH-1:0] wire_d20_56;
	wire [WIDTH-1:0] wire_d20_57;
	wire [WIDTH-1:0] wire_d20_58;
	wire [WIDTH-1:0] wire_d20_59;
	wire [WIDTH-1:0] wire_d20_60;
	wire [WIDTH-1:0] wire_d20_61;
	wire [WIDTH-1:0] wire_d20_62;
	wire [WIDTH-1:0] wire_d20_63;
	wire [WIDTH-1:0] wire_d20_64;
	wire [WIDTH-1:0] wire_d20_65;
	wire [WIDTH-1:0] wire_d20_66;
	wire [WIDTH-1:0] wire_d20_67;
	wire [WIDTH-1:0] wire_d20_68;
	wire [WIDTH-1:0] wire_d20_69;
	wire [WIDTH-1:0] wire_d20_70;
	wire [WIDTH-1:0] wire_d20_71;
	wire [WIDTH-1:0] wire_d20_72;
	wire [WIDTH-1:0] wire_d20_73;
	wire [WIDTH-1:0] wire_d20_74;
	wire [WIDTH-1:0] wire_d20_75;
	wire [WIDTH-1:0] wire_d20_76;
	wire [WIDTH-1:0] wire_d20_77;
	wire [WIDTH-1:0] wire_d20_78;
	wire [WIDTH-1:0] wire_d21_0;
	wire [WIDTH-1:0] wire_d21_1;
	wire [WIDTH-1:0] wire_d21_2;
	wire [WIDTH-1:0] wire_d21_3;
	wire [WIDTH-1:0] wire_d21_4;
	wire [WIDTH-1:0] wire_d21_5;
	wire [WIDTH-1:0] wire_d21_6;
	wire [WIDTH-1:0] wire_d21_7;
	wire [WIDTH-1:0] wire_d21_8;
	wire [WIDTH-1:0] wire_d21_9;
	wire [WIDTH-1:0] wire_d21_10;
	wire [WIDTH-1:0] wire_d21_11;
	wire [WIDTH-1:0] wire_d21_12;
	wire [WIDTH-1:0] wire_d21_13;
	wire [WIDTH-1:0] wire_d21_14;
	wire [WIDTH-1:0] wire_d21_15;
	wire [WIDTH-1:0] wire_d21_16;
	wire [WIDTH-1:0] wire_d21_17;
	wire [WIDTH-1:0] wire_d21_18;
	wire [WIDTH-1:0] wire_d21_19;
	wire [WIDTH-1:0] wire_d21_20;
	wire [WIDTH-1:0] wire_d21_21;
	wire [WIDTH-1:0] wire_d21_22;
	wire [WIDTH-1:0] wire_d21_23;
	wire [WIDTH-1:0] wire_d21_24;
	wire [WIDTH-1:0] wire_d21_25;
	wire [WIDTH-1:0] wire_d21_26;
	wire [WIDTH-1:0] wire_d21_27;
	wire [WIDTH-1:0] wire_d21_28;
	wire [WIDTH-1:0] wire_d21_29;
	wire [WIDTH-1:0] wire_d21_30;
	wire [WIDTH-1:0] wire_d21_31;
	wire [WIDTH-1:0] wire_d21_32;
	wire [WIDTH-1:0] wire_d21_33;
	wire [WIDTH-1:0] wire_d21_34;
	wire [WIDTH-1:0] wire_d21_35;
	wire [WIDTH-1:0] wire_d21_36;
	wire [WIDTH-1:0] wire_d21_37;
	wire [WIDTH-1:0] wire_d21_38;
	wire [WIDTH-1:0] wire_d21_39;
	wire [WIDTH-1:0] wire_d21_40;
	wire [WIDTH-1:0] wire_d21_41;
	wire [WIDTH-1:0] wire_d21_42;
	wire [WIDTH-1:0] wire_d21_43;
	wire [WIDTH-1:0] wire_d21_44;
	wire [WIDTH-1:0] wire_d21_45;
	wire [WIDTH-1:0] wire_d21_46;
	wire [WIDTH-1:0] wire_d21_47;
	wire [WIDTH-1:0] wire_d21_48;
	wire [WIDTH-1:0] wire_d21_49;
	wire [WIDTH-1:0] wire_d21_50;
	wire [WIDTH-1:0] wire_d21_51;
	wire [WIDTH-1:0] wire_d21_52;
	wire [WIDTH-1:0] wire_d21_53;
	wire [WIDTH-1:0] wire_d21_54;
	wire [WIDTH-1:0] wire_d21_55;
	wire [WIDTH-1:0] wire_d21_56;
	wire [WIDTH-1:0] wire_d21_57;
	wire [WIDTH-1:0] wire_d21_58;
	wire [WIDTH-1:0] wire_d21_59;
	wire [WIDTH-1:0] wire_d21_60;
	wire [WIDTH-1:0] wire_d21_61;
	wire [WIDTH-1:0] wire_d21_62;
	wire [WIDTH-1:0] wire_d21_63;
	wire [WIDTH-1:0] wire_d21_64;
	wire [WIDTH-1:0] wire_d21_65;
	wire [WIDTH-1:0] wire_d21_66;
	wire [WIDTH-1:0] wire_d21_67;
	wire [WIDTH-1:0] wire_d21_68;
	wire [WIDTH-1:0] wire_d21_69;
	wire [WIDTH-1:0] wire_d21_70;
	wire [WIDTH-1:0] wire_d21_71;
	wire [WIDTH-1:0] wire_d21_72;
	wire [WIDTH-1:0] wire_d21_73;
	wire [WIDTH-1:0] wire_d21_74;
	wire [WIDTH-1:0] wire_d21_75;
	wire [WIDTH-1:0] wire_d21_76;
	wire [WIDTH-1:0] wire_d21_77;
	wire [WIDTH-1:0] wire_d21_78;
	wire [WIDTH-1:0] wire_d22_0;
	wire [WIDTH-1:0] wire_d22_1;
	wire [WIDTH-1:0] wire_d22_2;
	wire [WIDTH-1:0] wire_d22_3;
	wire [WIDTH-1:0] wire_d22_4;
	wire [WIDTH-1:0] wire_d22_5;
	wire [WIDTH-1:0] wire_d22_6;
	wire [WIDTH-1:0] wire_d22_7;
	wire [WIDTH-1:0] wire_d22_8;
	wire [WIDTH-1:0] wire_d22_9;
	wire [WIDTH-1:0] wire_d22_10;
	wire [WIDTH-1:0] wire_d22_11;
	wire [WIDTH-1:0] wire_d22_12;
	wire [WIDTH-1:0] wire_d22_13;
	wire [WIDTH-1:0] wire_d22_14;
	wire [WIDTH-1:0] wire_d22_15;
	wire [WIDTH-1:0] wire_d22_16;
	wire [WIDTH-1:0] wire_d22_17;
	wire [WIDTH-1:0] wire_d22_18;
	wire [WIDTH-1:0] wire_d22_19;
	wire [WIDTH-1:0] wire_d22_20;
	wire [WIDTH-1:0] wire_d22_21;
	wire [WIDTH-1:0] wire_d22_22;
	wire [WIDTH-1:0] wire_d22_23;
	wire [WIDTH-1:0] wire_d22_24;
	wire [WIDTH-1:0] wire_d22_25;
	wire [WIDTH-1:0] wire_d22_26;
	wire [WIDTH-1:0] wire_d22_27;
	wire [WIDTH-1:0] wire_d22_28;
	wire [WIDTH-1:0] wire_d22_29;
	wire [WIDTH-1:0] wire_d22_30;
	wire [WIDTH-1:0] wire_d22_31;
	wire [WIDTH-1:0] wire_d22_32;
	wire [WIDTH-1:0] wire_d22_33;
	wire [WIDTH-1:0] wire_d22_34;
	wire [WIDTH-1:0] wire_d22_35;
	wire [WIDTH-1:0] wire_d22_36;
	wire [WIDTH-1:0] wire_d22_37;
	wire [WIDTH-1:0] wire_d22_38;
	wire [WIDTH-1:0] wire_d22_39;
	wire [WIDTH-1:0] wire_d22_40;
	wire [WIDTH-1:0] wire_d22_41;
	wire [WIDTH-1:0] wire_d22_42;
	wire [WIDTH-1:0] wire_d22_43;
	wire [WIDTH-1:0] wire_d22_44;
	wire [WIDTH-1:0] wire_d22_45;
	wire [WIDTH-1:0] wire_d22_46;
	wire [WIDTH-1:0] wire_d22_47;
	wire [WIDTH-1:0] wire_d22_48;
	wire [WIDTH-1:0] wire_d22_49;
	wire [WIDTH-1:0] wire_d22_50;
	wire [WIDTH-1:0] wire_d22_51;
	wire [WIDTH-1:0] wire_d22_52;
	wire [WIDTH-1:0] wire_d22_53;
	wire [WIDTH-1:0] wire_d22_54;
	wire [WIDTH-1:0] wire_d22_55;
	wire [WIDTH-1:0] wire_d22_56;
	wire [WIDTH-1:0] wire_d22_57;
	wire [WIDTH-1:0] wire_d22_58;
	wire [WIDTH-1:0] wire_d22_59;
	wire [WIDTH-1:0] wire_d22_60;
	wire [WIDTH-1:0] wire_d22_61;
	wire [WIDTH-1:0] wire_d22_62;
	wire [WIDTH-1:0] wire_d22_63;
	wire [WIDTH-1:0] wire_d22_64;
	wire [WIDTH-1:0] wire_d22_65;
	wire [WIDTH-1:0] wire_d22_66;
	wire [WIDTH-1:0] wire_d22_67;
	wire [WIDTH-1:0] wire_d22_68;
	wire [WIDTH-1:0] wire_d22_69;
	wire [WIDTH-1:0] wire_d22_70;
	wire [WIDTH-1:0] wire_d22_71;
	wire [WIDTH-1:0] wire_d22_72;
	wire [WIDTH-1:0] wire_d22_73;
	wire [WIDTH-1:0] wire_d22_74;
	wire [WIDTH-1:0] wire_d22_75;
	wire [WIDTH-1:0] wire_d22_76;
	wire [WIDTH-1:0] wire_d22_77;
	wire [WIDTH-1:0] wire_d22_78;
	wire [WIDTH-1:0] wire_d23_0;
	wire [WIDTH-1:0] wire_d23_1;
	wire [WIDTH-1:0] wire_d23_2;
	wire [WIDTH-1:0] wire_d23_3;
	wire [WIDTH-1:0] wire_d23_4;
	wire [WIDTH-1:0] wire_d23_5;
	wire [WIDTH-1:0] wire_d23_6;
	wire [WIDTH-1:0] wire_d23_7;
	wire [WIDTH-1:0] wire_d23_8;
	wire [WIDTH-1:0] wire_d23_9;
	wire [WIDTH-1:0] wire_d23_10;
	wire [WIDTH-1:0] wire_d23_11;
	wire [WIDTH-1:0] wire_d23_12;
	wire [WIDTH-1:0] wire_d23_13;
	wire [WIDTH-1:0] wire_d23_14;
	wire [WIDTH-1:0] wire_d23_15;
	wire [WIDTH-1:0] wire_d23_16;
	wire [WIDTH-1:0] wire_d23_17;
	wire [WIDTH-1:0] wire_d23_18;
	wire [WIDTH-1:0] wire_d23_19;
	wire [WIDTH-1:0] wire_d23_20;
	wire [WIDTH-1:0] wire_d23_21;
	wire [WIDTH-1:0] wire_d23_22;
	wire [WIDTH-1:0] wire_d23_23;
	wire [WIDTH-1:0] wire_d23_24;
	wire [WIDTH-1:0] wire_d23_25;
	wire [WIDTH-1:0] wire_d23_26;
	wire [WIDTH-1:0] wire_d23_27;
	wire [WIDTH-1:0] wire_d23_28;
	wire [WIDTH-1:0] wire_d23_29;
	wire [WIDTH-1:0] wire_d23_30;
	wire [WIDTH-1:0] wire_d23_31;
	wire [WIDTH-1:0] wire_d23_32;
	wire [WIDTH-1:0] wire_d23_33;
	wire [WIDTH-1:0] wire_d23_34;
	wire [WIDTH-1:0] wire_d23_35;
	wire [WIDTH-1:0] wire_d23_36;
	wire [WIDTH-1:0] wire_d23_37;
	wire [WIDTH-1:0] wire_d23_38;
	wire [WIDTH-1:0] wire_d23_39;
	wire [WIDTH-1:0] wire_d23_40;
	wire [WIDTH-1:0] wire_d23_41;
	wire [WIDTH-1:0] wire_d23_42;
	wire [WIDTH-1:0] wire_d23_43;
	wire [WIDTH-1:0] wire_d23_44;
	wire [WIDTH-1:0] wire_d23_45;
	wire [WIDTH-1:0] wire_d23_46;
	wire [WIDTH-1:0] wire_d23_47;
	wire [WIDTH-1:0] wire_d23_48;
	wire [WIDTH-1:0] wire_d23_49;
	wire [WIDTH-1:0] wire_d23_50;
	wire [WIDTH-1:0] wire_d23_51;
	wire [WIDTH-1:0] wire_d23_52;
	wire [WIDTH-1:0] wire_d23_53;
	wire [WIDTH-1:0] wire_d23_54;
	wire [WIDTH-1:0] wire_d23_55;
	wire [WIDTH-1:0] wire_d23_56;
	wire [WIDTH-1:0] wire_d23_57;
	wire [WIDTH-1:0] wire_d23_58;
	wire [WIDTH-1:0] wire_d23_59;
	wire [WIDTH-1:0] wire_d23_60;
	wire [WIDTH-1:0] wire_d23_61;
	wire [WIDTH-1:0] wire_d23_62;
	wire [WIDTH-1:0] wire_d23_63;
	wire [WIDTH-1:0] wire_d23_64;
	wire [WIDTH-1:0] wire_d23_65;
	wire [WIDTH-1:0] wire_d23_66;
	wire [WIDTH-1:0] wire_d23_67;
	wire [WIDTH-1:0] wire_d23_68;
	wire [WIDTH-1:0] wire_d23_69;
	wire [WIDTH-1:0] wire_d23_70;
	wire [WIDTH-1:0] wire_d23_71;
	wire [WIDTH-1:0] wire_d23_72;
	wire [WIDTH-1:0] wire_d23_73;
	wire [WIDTH-1:0] wire_d23_74;
	wire [WIDTH-1:0] wire_d23_75;
	wire [WIDTH-1:0] wire_d23_76;
	wire [WIDTH-1:0] wire_d23_77;
	wire [WIDTH-1:0] wire_d23_78;
	wire [WIDTH-1:0] wire_d24_0;
	wire [WIDTH-1:0] wire_d24_1;
	wire [WIDTH-1:0] wire_d24_2;
	wire [WIDTH-1:0] wire_d24_3;
	wire [WIDTH-1:0] wire_d24_4;
	wire [WIDTH-1:0] wire_d24_5;
	wire [WIDTH-1:0] wire_d24_6;
	wire [WIDTH-1:0] wire_d24_7;
	wire [WIDTH-1:0] wire_d24_8;
	wire [WIDTH-1:0] wire_d24_9;
	wire [WIDTH-1:0] wire_d24_10;
	wire [WIDTH-1:0] wire_d24_11;
	wire [WIDTH-1:0] wire_d24_12;
	wire [WIDTH-1:0] wire_d24_13;
	wire [WIDTH-1:0] wire_d24_14;
	wire [WIDTH-1:0] wire_d24_15;
	wire [WIDTH-1:0] wire_d24_16;
	wire [WIDTH-1:0] wire_d24_17;
	wire [WIDTH-1:0] wire_d24_18;
	wire [WIDTH-1:0] wire_d24_19;
	wire [WIDTH-1:0] wire_d24_20;
	wire [WIDTH-1:0] wire_d24_21;
	wire [WIDTH-1:0] wire_d24_22;
	wire [WIDTH-1:0] wire_d24_23;
	wire [WIDTH-1:0] wire_d24_24;
	wire [WIDTH-1:0] wire_d24_25;
	wire [WIDTH-1:0] wire_d24_26;
	wire [WIDTH-1:0] wire_d24_27;
	wire [WIDTH-1:0] wire_d24_28;
	wire [WIDTH-1:0] wire_d24_29;
	wire [WIDTH-1:0] wire_d24_30;
	wire [WIDTH-1:0] wire_d24_31;
	wire [WIDTH-1:0] wire_d24_32;
	wire [WIDTH-1:0] wire_d24_33;
	wire [WIDTH-1:0] wire_d24_34;
	wire [WIDTH-1:0] wire_d24_35;
	wire [WIDTH-1:0] wire_d24_36;
	wire [WIDTH-1:0] wire_d24_37;
	wire [WIDTH-1:0] wire_d24_38;
	wire [WIDTH-1:0] wire_d24_39;
	wire [WIDTH-1:0] wire_d24_40;
	wire [WIDTH-1:0] wire_d24_41;
	wire [WIDTH-1:0] wire_d24_42;
	wire [WIDTH-1:0] wire_d24_43;
	wire [WIDTH-1:0] wire_d24_44;
	wire [WIDTH-1:0] wire_d24_45;
	wire [WIDTH-1:0] wire_d24_46;
	wire [WIDTH-1:0] wire_d24_47;
	wire [WIDTH-1:0] wire_d24_48;
	wire [WIDTH-1:0] wire_d24_49;
	wire [WIDTH-1:0] wire_d24_50;
	wire [WIDTH-1:0] wire_d24_51;
	wire [WIDTH-1:0] wire_d24_52;
	wire [WIDTH-1:0] wire_d24_53;
	wire [WIDTH-1:0] wire_d24_54;
	wire [WIDTH-1:0] wire_d24_55;
	wire [WIDTH-1:0] wire_d24_56;
	wire [WIDTH-1:0] wire_d24_57;
	wire [WIDTH-1:0] wire_d24_58;
	wire [WIDTH-1:0] wire_d24_59;
	wire [WIDTH-1:0] wire_d24_60;
	wire [WIDTH-1:0] wire_d24_61;
	wire [WIDTH-1:0] wire_d24_62;
	wire [WIDTH-1:0] wire_d24_63;
	wire [WIDTH-1:0] wire_d24_64;
	wire [WIDTH-1:0] wire_d24_65;
	wire [WIDTH-1:0] wire_d24_66;
	wire [WIDTH-1:0] wire_d24_67;
	wire [WIDTH-1:0] wire_d24_68;
	wire [WIDTH-1:0] wire_d24_69;
	wire [WIDTH-1:0] wire_d24_70;
	wire [WIDTH-1:0] wire_d24_71;
	wire [WIDTH-1:0] wire_d24_72;
	wire [WIDTH-1:0] wire_d24_73;
	wire [WIDTH-1:0] wire_d24_74;
	wire [WIDTH-1:0] wire_d24_75;
	wire [WIDTH-1:0] wire_d24_76;
	wire [WIDTH-1:0] wire_d24_77;
	wire [WIDTH-1:0] wire_d24_78;
	wire [WIDTH-1:0] wire_d25_0;
	wire [WIDTH-1:0] wire_d25_1;
	wire [WIDTH-1:0] wire_d25_2;
	wire [WIDTH-1:0] wire_d25_3;
	wire [WIDTH-1:0] wire_d25_4;
	wire [WIDTH-1:0] wire_d25_5;
	wire [WIDTH-1:0] wire_d25_6;
	wire [WIDTH-1:0] wire_d25_7;
	wire [WIDTH-1:0] wire_d25_8;
	wire [WIDTH-1:0] wire_d25_9;
	wire [WIDTH-1:0] wire_d25_10;
	wire [WIDTH-1:0] wire_d25_11;
	wire [WIDTH-1:0] wire_d25_12;
	wire [WIDTH-1:0] wire_d25_13;
	wire [WIDTH-1:0] wire_d25_14;
	wire [WIDTH-1:0] wire_d25_15;
	wire [WIDTH-1:0] wire_d25_16;
	wire [WIDTH-1:0] wire_d25_17;
	wire [WIDTH-1:0] wire_d25_18;
	wire [WIDTH-1:0] wire_d25_19;
	wire [WIDTH-1:0] wire_d25_20;
	wire [WIDTH-1:0] wire_d25_21;
	wire [WIDTH-1:0] wire_d25_22;
	wire [WIDTH-1:0] wire_d25_23;
	wire [WIDTH-1:0] wire_d25_24;
	wire [WIDTH-1:0] wire_d25_25;
	wire [WIDTH-1:0] wire_d25_26;
	wire [WIDTH-1:0] wire_d25_27;
	wire [WIDTH-1:0] wire_d25_28;
	wire [WIDTH-1:0] wire_d25_29;
	wire [WIDTH-1:0] wire_d25_30;
	wire [WIDTH-1:0] wire_d25_31;
	wire [WIDTH-1:0] wire_d25_32;
	wire [WIDTH-1:0] wire_d25_33;
	wire [WIDTH-1:0] wire_d25_34;
	wire [WIDTH-1:0] wire_d25_35;
	wire [WIDTH-1:0] wire_d25_36;
	wire [WIDTH-1:0] wire_d25_37;
	wire [WIDTH-1:0] wire_d25_38;
	wire [WIDTH-1:0] wire_d25_39;
	wire [WIDTH-1:0] wire_d25_40;
	wire [WIDTH-1:0] wire_d25_41;
	wire [WIDTH-1:0] wire_d25_42;
	wire [WIDTH-1:0] wire_d25_43;
	wire [WIDTH-1:0] wire_d25_44;
	wire [WIDTH-1:0] wire_d25_45;
	wire [WIDTH-1:0] wire_d25_46;
	wire [WIDTH-1:0] wire_d25_47;
	wire [WIDTH-1:0] wire_d25_48;
	wire [WIDTH-1:0] wire_d25_49;
	wire [WIDTH-1:0] wire_d25_50;
	wire [WIDTH-1:0] wire_d25_51;
	wire [WIDTH-1:0] wire_d25_52;
	wire [WIDTH-1:0] wire_d25_53;
	wire [WIDTH-1:0] wire_d25_54;
	wire [WIDTH-1:0] wire_d25_55;
	wire [WIDTH-1:0] wire_d25_56;
	wire [WIDTH-1:0] wire_d25_57;
	wire [WIDTH-1:0] wire_d25_58;
	wire [WIDTH-1:0] wire_d25_59;
	wire [WIDTH-1:0] wire_d25_60;
	wire [WIDTH-1:0] wire_d25_61;
	wire [WIDTH-1:0] wire_d25_62;
	wire [WIDTH-1:0] wire_d25_63;
	wire [WIDTH-1:0] wire_d25_64;
	wire [WIDTH-1:0] wire_d25_65;
	wire [WIDTH-1:0] wire_d25_66;
	wire [WIDTH-1:0] wire_d25_67;
	wire [WIDTH-1:0] wire_d25_68;
	wire [WIDTH-1:0] wire_d25_69;
	wire [WIDTH-1:0] wire_d25_70;
	wire [WIDTH-1:0] wire_d25_71;
	wire [WIDTH-1:0] wire_d25_72;
	wire [WIDTH-1:0] wire_d25_73;
	wire [WIDTH-1:0] wire_d25_74;
	wire [WIDTH-1:0] wire_d25_75;
	wire [WIDTH-1:0] wire_d25_76;
	wire [WIDTH-1:0] wire_d25_77;
	wire [WIDTH-1:0] wire_d25_78;
	wire [WIDTH-1:0] wire_d26_0;
	wire [WIDTH-1:0] wire_d26_1;
	wire [WIDTH-1:0] wire_d26_2;
	wire [WIDTH-1:0] wire_d26_3;
	wire [WIDTH-1:0] wire_d26_4;
	wire [WIDTH-1:0] wire_d26_5;
	wire [WIDTH-1:0] wire_d26_6;
	wire [WIDTH-1:0] wire_d26_7;
	wire [WIDTH-1:0] wire_d26_8;
	wire [WIDTH-1:0] wire_d26_9;
	wire [WIDTH-1:0] wire_d26_10;
	wire [WIDTH-1:0] wire_d26_11;
	wire [WIDTH-1:0] wire_d26_12;
	wire [WIDTH-1:0] wire_d26_13;
	wire [WIDTH-1:0] wire_d26_14;
	wire [WIDTH-1:0] wire_d26_15;
	wire [WIDTH-1:0] wire_d26_16;
	wire [WIDTH-1:0] wire_d26_17;
	wire [WIDTH-1:0] wire_d26_18;
	wire [WIDTH-1:0] wire_d26_19;
	wire [WIDTH-1:0] wire_d26_20;
	wire [WIDTH-1:0] wire_d26_21;
	wire [WIDTH-1:0] wire_d26_22;
	wire [WIDTH-1:0] wire_d26_23;
	wire [WIDTH-1:0] wire_d26_24;
	wire [WIDTH-1:0] wire_d26_25;
	wire [WIDTH-1:0] wire_d26_26;
	wire [WIDTH-1:0] wire_d26_27;
	wire [WIDTH-1:0] wire_d26_28;
	wire [WIDTH-1:0] wire_d26_29;
	wire [WIDTH-1:0] wire_d26_30;
	wire [WIDTH-1:0] wire_d26_31;
	wire [WIDTH-1:0] wire_d26_32;
	wire [WIDTH-1:0] wire_d26_33;
	wire [WIDTH-1:0] wire_d26_34;
	wire [WIDTH-1:0] wire_d26_35;
	wire [WIDTH-1:0] wire_d26_36;
	wire [WIDTH-1:0] wire_d26_37;
	wire [WIDTH-1:0] wire_d26_38;
	wire [WIDTH-1:0] wire_d26_39;
	wire [WIDTH-1:0] wire_d26_40;
	wire [WIDTH-1:0] wire_d26_41;
	wire [WIDTH-1:0] wire_d26_42;
	wire [WIDTH-1:0] wire_d26_43;
	wire [WIDTH-1:0] wire_d26_44;
	wire [WIDTH-1:0] wire_d26_45;
	wire [WIDTH-1:0] wire_d26_46;
	wire [WIDTH-1:0] wire_d26_47;
	wire [WIDTH-1:0] wire_d26_48;
	wire [WIDTH-1:0] wire_d26_49;
	wire [WIDTH-1:0] wire_d26_50;
	wire [WIDTH-1:0] wire_d26_51;
	wire [WIDTH-1:0] wire_d26_52;
	wire [WIDTH-1:0] wire_d26_53;
	wire [WIDTH-1:0] wire_d26_54;
	wire [WIDTH-1:0] wire_d26_55;
	wire [WIDTH-1:0] wire_d26_56;
	wire [WIDTH-1:0] wire_d26_57;
	wire [WIDTH-1:0] wire_d26_58;
	wire [WIDTH-1:0] wire_d26_59;
	wire [WIDTH-1:0] wire_d26_60;
	wire [WIDTH-1:0] wire_d26_61;
	wire [WIDTH-1:0] wire_d26_62;
	wire [WIDTH-1:0] wire_d26_63;
	wire [WIDTH-1:0] wire_d26_64;
	wire [WIDTH-1:0] wire_d26_65;
	wire [WIDTH-1:0] wire_d26_66;
	wire [WIDTH-1:0] wire_d26_67;
	wire [WIDTH-1:0] wire_d26_68;
	wire [WIDTH-1:0] wire_d26_69;
	wire [WIDTH-1:0] wire_d26_70;
	wire [WIDTH-1:0] wire_d26_71;
	wire [WIDTH-1:0] wire_d26_72;
	wire [WIDTH-1:0] wire_d26_73;
	wire [WIDTH-1:0] wire_d26_74;
	wire [WIDTH-1:0] wire_d26_75;
	wire [WIDTH-1:0] wire_d26_76;
	wire [WIDTH-1:0] wire_d26_77;
	wire [WIDTH-1:0] wire_d26_78;
	wire [WIDTH-1:0] wire_d27_0;
	wire [WIDTH-1:0] wire_d27_1;
	wire [WIDTH-1:0] wire_d27_2;
	wire [WIDTH-1:0] wire_d27_3;
	wire [WIDTH-1:0] wire_d27_4;
	wire [WIDTH-1:0] wire_d27_5;
	wire [WIDTH-1:0] wire_d27_6;
	wire [WIDTH-1:0] wire_d27_7;
	wire [WIDTH-1:0] wire_d27_8;
	wire [WIDTH-1:0] wire_d27_9;
	wire [WIDTH-1:0] wire_d27_10;
	wire [WIDTH-1:0] wire_d27_11;
	wire [WIDTH-1:0] wire_d27_12;
	wire [WIDTH-1:0] wire_d27_13;
	wire [WIDTH-1:0] wire_d27_14;
	wire [WIDTH-1:0] wire_d27_15;
	wire [WIDTH-1:0] wire_d27_16;
	wire [WIDTH-1:0] wire_d27_17;
	wire [WIDTH-1:0] wire_d27_18;
	wire [WIDTH-1:0] wire_d27_19;
	wire [WIDTH-1:0] wire_d27_20;
	wire [WIDTH-1:0] wire_d27_21;
	wire [WIDTH-1:0] wire_d27_22;
	wire [WIDTH-1:0] wire_d27_23;
	wire [WIDTH-1:0] wire_d27_24;
	wire [WIDTH-1:0] wire_d27_25;
	wire [WIDTH-1:0] wire_d27_26;
	wire [WIDTH-1:0] wire_d27_27;
	wire [WIDTH-1:0] wire_d27_28;
	wire [WIDTH-1:0] wire_d27_29;
	wire [WIDTH-1:0] wire_d27_30;
	wire [WIDTH-1:0] wire_d27_31;
	wire [WIDTH-1:0] wire_d27_32;
	wire [WIDTH-1:0] wire_d27_33;
	wire [WIDTH-1:0] wire_d27_34;
	wire [WIDTH-1:0] wire_d27_35;
	wire [WIDTH-1:0] wire_d27_36;
	wire [WIDTH-1:0] wire_d27_37;
	wire [WIDTH-1:0] wire_d27_38;
	wire [WIDTH-1:0] wire_d27_39;
	wire [WIDTH-1:0] wire_d27_40;
	wire [WIDTH-1:0] wire_d27_41;
	wire [WIDTH-1:0] wire_d27_42;
	wire [WIDTH-1:0] wire_d27_43;
	wire [WIDTH-1:0] wire_d27_44;
	wire [WIDTH-1:0] wire_d27_45;
	wire [WIDTH-1:0] wire_d27_46;
	wire [WIDTH-1:0] wire_d27_47;
	wire [WIDTH-1:0] wire_d27_48;
	wire [WIDTH-1:0] wire_d27_49;
	wire [WIDTH-1:0] wire_d27_50;
	wire [WIDTH-1:0] wire_d27_51;
	wire [WIDTH-1:0] wire_d27_52;
	wire [WIDTH-1:0] wire_d27_53;
	wire [WIDTH-1:0] wire_d27_54;
	wire [WIDTH-1:0] wire_d27_55;
	wire [WIDTH-1:0] wire_d27_56;
	wire [WIDTH-1:0] wire_d27_57;
	wire [WIDTH-1:0] wire_d27_58;
	wire [WIDTH-1:0] wire_d27_59;
	wire [WIDTH-1:0] wire_d27_60;
	wire [WIDTH-1:0] wire_d27_61;
	wire [WIDTH-1:0] wire_d27_62;
	wire [WIDTH-1:0] wire_d27_63;
	wire [WIDTH-1:0] wire_d27_64;
	wire [WIDTH-1:0] wire_d27_65;
	wire [WIDTH-1:0] wire_d27_66;
	wire [WIDTH-1:0] wire_d27_67;
	wire [WIDTH-1:0] wire_d27_68;
	wire [WIDTH-1:0] wire_d27_69;
	wire [WIDTH-1:0] wire_d27_70;
	wire [WIDTH-1:0] wire_d27_71;
	wire [WIDTH-1:0] wire_d27_72;
	wire [WIDTH-1:0] wire_d27_73;
	wire [WIDTH-1:0] wire_d27_74;
	wire [WIDTH-1:0] wire_d27_75;
	wire [WIDTH-1:0] wire_d27_76;
	wire [WIDTH-1:0] wire_d27_77;
	wire [WIDTH-1:0] wire_d27_78;
	wire [WIDTH-1:0] wire_d28_0;
	wire [WIDTH-1:0] wire_d28_1;
	wire [WIDTH-1:0] wire_d28_2;
	wire [WIDTH-1:0] wire_d28_3;
	wire [WIDTH-1:0] wire_d28_4;
	wire [WIDTH-1:0] wire_d28_5;
	wire [WIDTH-1:0] wire_d28_6;
	wire [WIDTH-1:0] wire_d28_7;
	wire [WIDTH-1:0] wire_d28_8;
	wire [WIDTH-1:0] wire_d28_9;
	wire [WIDTH-1:0] wire_d28_10;
	wire [WIDTH-1:0] wire_d28_11;
	wire [WIDTH-1:0] wire_d28_12;
	wire [WIDTH-1:0] wire_d28_13;
	wire [WIDTH-1:0] wire_d28_14;
	wire [WIDTH-1:0] wire_d28_15;
	wire [WIDTH-1:0] wire_d28_16;
	wire [WIDTH-1:0] wire_d28_17;
	wire [WIDTH-1:0] wire_d28_18;
	wire [WIDTH-1:0] wire_d28_19;
	wire [WIDTH-1:0] wire_d28_20;
	wire [WIDTH-1:0] wire_d28_21;
	wire [WIDTH-1:0] wire_d28_22;
	wire [WIDTH-1:0] wire_d28_23;
	wire [WIDTH-1:0] wire_d28_24;
	wire [WIDTH-1:0] wire_d28_25;
	wire [WIDTH-1:0] wire_d28_26;
	wire [WIDTH-1:0] wire_d28_27;
	wire [WIDTH-1:0] wire_d28_28;
	wire [WIDTH-1:0] wire_d28_29;
	wire [WIDTH-1:0] wire_d28_30;
	wire [WIDTH-1:0] wire_d28_31;
	wire [WIDTH-1:0] wire_d28_32;
	wire [WIDTH-1:0] wire_d28_33;
	wire [WIDTH-1:0] wire_d28_34;
	wire [WIDTH-1:0] wire_d28_35;
	wire [WIDTH-1:0] wire_d28_36;
	wire [WIDTH-1:0] wire_d28_37;
	wire [WIDTH-1:0] wire_d28_38;
	wire [WIDTH-1:0] wire_d28_39;
	wire [WIDTH-1:0] wire_d28_40;
	wire [WIDTH-1:0] wire_d28_41;
	wire [WIDTH-1:0] wire_d28_42;
	wire [WIDTH-1:0] wire_d28_43;
	wire [WIDTH-1:0] wire_d28_44;
	wire [WIDTH-1:0] wire_d28_45;
	wire [WIDTH-1:0] wire_d28_46;
	wire [WIDTH-1:0] wire_d28_47;
	wire [WIDTH-1:0] wire_d28_48;
	wire [WIDTH-1:0] wire_d28_49;
	wire [WIDTH-1:0] wire_d28_50;
	wire [WIDTH-1:0] wire_d28_51;
	wire [WIDTH-1:0] wire_d28_52;
	wire [WIDTH-1:0] wire_d28_53;
	wire [WIDTH-1:0] wire_d28_54;
	wire [WIDTH-1:0] wire_d28_55;
	wire [WIDTH-1:0] wire_d28_56;
	wire [WIDTH-1:0] wire_d28_57;
	wire [WIDTH-1:0] wire_d28_58;
	wire [WIDTH-1:0] wire_d28_59;
	wire [WIDTH-1:0] wire_d28_60;
	wire [WIDTH-1:0] wire_d28_61;
	wire [WIDTH-1:0] wire_d28_62;
	wire [WIDTH-1:0] wire_d28_63;
	wire [WIDTH-1:0] wire_d28_64;
	wire [WIDTH-1:0] wire_d28_65;
	wire [WIDTH-1:0] wire_d28_66;
	wire [WIDTH-1:0] wire_d28_67;
	wire [WIDTH-1:0] wire_d28_68;
	wire [WIDTH-1:0] wire_d28_69;
	wire [WIDTH-1:0] wire_d28_70;
	wire [WIDTH-1:0] wire_d28_71;
	wire [WIDTH-1:0] wire_d28_72;
	wire [WIDTH-1:0] wire_d28_73;
	wire [WIDTH-1:0] wire_d28_74;
	wire [WIDTH-1:0] wire_d28_75;
	wire [WIDTH-1:0] wire_d28_76;
	wire [WIDTH-1:0] wire_d28_77;
	wire [WIDTH-1:0] wire_d28_78;
	wire [WIDTH-1:0] wire_d29_0;
	wire [WIDTH-1:0] wire_d29_1;
	wire [WIDTH-1:0] wire_d29_2;
	wire [WIDTH-1:0] wire_d29_3;
	wire [WIDTH-1:0] wire_d29_4;
	wire [WIDTH-1:0] wire_d29_5;
	wire [WIDTH-1:0] wire_d29_6;
	wire [WIDTH-1:0] wire_d29_7;
	wire [WIDTH-1:0] wire_d29_8;
	wire [WIDTH-1:0] wire_d29_9;
	wire [WIDTH-1:0] wire_d29_10;
	wire [WIDTH-1:0] wire_d29_11;
	wire [WIDTH-1:0] wire_d29_12;
	wire [WIDTH-1:0] wire_d29_13;
	wire [WIDTH-1:0] wire_d29_14;
	wire [WIDTH-1:0] wire_d29_15;
	wire [WIDTH-1:0] wire_d29_16;
	wire [WIDTH-1:0] wire_d29_17;
	wire [WIDTH-1:0] wire_d29_18;
	wire [WIDTH-1:0] wire_d29_19;
	wire [WIDTH-1:0] wire_d29_20;
	wire [WIDTH-1:0] wire_d29_21;
	wire [WIDTH-1:0] wire_d29_22;
	wire [WIDTH-1:0] wire_d29_23;
	wire [WIDTH-1:0] wire_d29_24;
	wire [WIDTH-1:0] wire_d29_25;
	wire [WIDTH-1:0] wire_d29_26;
	wire [WIDTH-1:0] wire_d29_27;
	wire [WIDTH-1:0] wire_d29_28;
	wire [WIDTH-1:0] wire_d29_29;
	wire [WIDTH-1:0] wire_d29_30;
	wire [WIDTH-1:0] wire_d29_31;
	wire [WIDTH-1:0] wire_d29_32;
	wire [WIDTH-1:0] wire_d29_33;
	wire [WIDTH-1:0] wire_d29_34;
	wire [WIDTH-1:0] wire_d29_35;
	wire [WIDTH-1:0] wire_d29_36;
	wire [WIDTH-1:0] wire_d29_37;
	wire [WIDTH-1:0] wire_d29_38;
	wire [WIDTH-1:0] wire_d29_39;
	wire [WIDTH-1:0] wire_d29_40;
	wire [WIDTH-1:0] wire_d29_41;
	wire [WIDTH-1:0] wire_d29_42;
	wire [WIDTH-1:0] wire_d29_43;
	wire [WIDTH-1:0] wire_d29_44;
	wire [WIDTH-1:0] wire_d29_45;
	wire [WIDTH-1:0] wire_d29_46;
	wire [WIDTH-1:0] wire_d29_47;
	wire [WIDTH-1:0] wire_d29_48;
	wire [WIDTH-1:0] wire_d29_49;
	wire [WIDTH-1:0] wire_d29_50;
	wire [WIDTH-1:0] wire_d29_51;
	wire [WIDTH-1:0] wire_d29_52;
	wire [WIDTH-1:0] wire_d29_53;
	wire [WIDTH-1:0] wire_d29_54;
	wire [WIDTH-1:0] wire_d29_55;
	wire [WIDTH-1:0] wire_d29_56;
	wire [WIDTH-1:0] wire_d29_57;
	wire [WIDTH-1:0] wire_d29_58;
	wire [WIDTH-1:0] wire_d29_59;
	wire [WIDTH-1:0] wire_d29_60;
	wire [WIDTH-1:0] wire_d29_61;
	wire [WIDTH-1:0] wire_d29_62;
	wire [WIDTH-1:0] wire_d29_63;
	wire [WIDTH-1:0] wire_d29_64;
	wire [WIDTH-1:0] wire_d29_65;
	wire [WIDTH-1:0] wire_d29_66;
	wire [WIDTH-1:0] wire_d29_67;
	wire [WIDTH-1:0] wire_d29_68;
	wire [WIDTH-1:0] wire_d29_69;
	wire [WIDTH-1:0] wire_d29_70;
	wire [WIDTH-1:0] wire_d29_71;
	wire [WIDTH-1:0] wire_d29_72;
	wire [WIDTH-1:0] wire_d29_73;
	wire [WIDTH-1:0] wire_d29_74;
	wire [WIDTH-1:0] wire_d29_75;
	wire [WIDTH-1:0] wire_d29_76;
	wire [WIDTH-1:0] wire_d29_77;
	wire [WIDTH-1:0] wire_d29_78;
	wire [WIDTH-1:0] wire_d30_0;
	wire [WIDTH-1:0] wire_d30_1;
	wire [WIDTH-1:0] wire_d30_2;
	wire [WIDTH-1:0] wire_d30_3;
	wire [WIDTH-1:0] wire_d30_4;
	wire [WIDTH-1:0] wire_d30_5;
	wire [WIDTH-1:0] wire_d30_6;
	wire [WIDTH-1:0] wire_d30_7;
	wire [WIDTH-1:0] wire_d30_8;
	wire [WIDTH-1:0] wire_d30_9;
	wire [WIDTH-1:0] wire_d30_10;
	wire [WIDTH-1:0] wire_d30_11;
	wire [WIDTH-1:0] wire_d30_12;
	wire [WIDTH-1:0] wire_d30_13;
	wire [WIDTH-1:0] wire_d30_14;
	wire [WIDTH-1:0] wire_d30_15;
	wire [WIDTH-1:0] wire_d30_16;
	wire [WIDTH-1:0] wire_d30_17;
	wire [WIDTH-1:0] wire_d30_18;
	wire [WIDTH-1:0] wire_d30_19;
	wire [WIDTH-1:0] wire_d30_20;
	wire [WIDTH-1:0] wire_d30_21;
	wire [WIDTH-1:0] wire_d30_22;
	wire [WIDTH-1:0] wire_d30_23;
	wire [WIDTH-1:0] wire_d30_24;
	wire [WIDTH-1:0] wire_d30_25;
	wire [WIDTH-1:0] wire_d30_26;
	wire [WIDTH-1:0] wire_d30_27;
	wire [WIDTH-1:0] wire_d30_28;
	wire [WIDTH-1:0] wire_d30_29;
	wire [WIDTH-1:0] wire_d30_30;
	wire [WIDTH-1:0] wire_d30_31;
	wire [WIDTH-1:0] wire_d30_32;
	wire [WIDTH-1:0] wire_d30_33;
	wire [WIDTH-1:0] wire_d30_34;
	wire [WIDTH-1:0] wire_d30_35;
	wire [WIDTH-1:0] wire_d30_36;
	wire [WIDTH-1:0] wire_d30_37;
	wire [WIDTH-1:0] wire_d30_38;
	wire [WIDTH-1:0] wire_d30_39;
	wire [WIDTH-1:0] wire_d30_40;
	wire [WIDTH-1:0] wire_d30_41;
	wire [WIDTH-1:0] wire_d30_42;
	wire [WIDTH-1:0] wire_d30_43;
	wire [WIDTH-1:0] wire_d30_44;
	wire [WIDTH-1:0] wire_d30_45;
	wire [WIDTH-1:0] wire_d30_46;
	wire [WIDTH-1:0] wire_d30_47;
	wire [WIDTH-1:0] wire_d30_48;
	wire [WIDTH-1:0] wire_d30_49;
	wire [WIDTH-1:0] wire_d30_50;
	wire [WIDTH-1:0] wire_d30_51;
	wire [WIDTH-1:0] wire_d30_52;
	wire [WIDTH-1:0] wire_d30_53;
	wire [WIDTH-1:0] wire_d30_54;
	wire [WIDTH-1:0] wire_d30_55;
	wire [WIDTH-1:0] wire_d30_56;
	wire [WIDTH-1:0] wire_d30_57;
	wire [WIDTH-1:0] wire_d30_58;
	wire [WIDTH-1:0] wire_d30_59;
	wire [WIDTH-1:0] wire_d30_60;
	wire [WIDTH-1:0] wire_d30_61;
	wire [WIDTH-1:0] wire_d30_62;
	wire [WIDTH-1:0] wire_d30_63;
	wire [WIDTH-1:0] wire_d30_64;
	wire [WIDTH-1:0] wire_d30_65;
	wire [WIDTH-1:0] wire_d30_66;
	wire [WIDTH-1:0] wire_d30_67;
	wire [WIDTH-1:0] wire_d30_68;
	wire [WIDTH-1:0] wire_d30_69;
	wire [WIDTH-1:0] wire_d30_70;
	wire [WIDTH-1:0] wire_d30_71;
	wire [WIDTH-1:0] wire_d30_72;
	wire [WIDTH-1:0] wire_d30_73;
	wire [WIDTH-1:0] wire_d30_74;
	wire [WIDTH-1:0] wire_d30_75;
	wire [WIDTH-1:0] wire_d30_76;
	wire [WIDTH-1:0] wire_d30_77;
	wire [WIDTH-1:0] wire_d30_78;
	wire [WIDTH-1:0] wire_d31_0;
	wire [WIDTH-1:0] wire_d31_1;
	wire [WIDTH-1:0] wire_d31_2;
	wire [WIDTH-1:0] wire_d31_3;
	wire [WIDTH-1:0] wire_d31_4;
	wire [WIDTH-1:0] wire_d31_5;
	wire [WIDTH-1:0] wire_d31_6;
	wire [WIDTH-1:0] wire_d31_7;
	wire [WIDTH-1:0] wire_d31_8;
	wire [WIDTH-1:0] wire_d31_9;
	wire [WIDTH-1:0] wire_d31_10;
	wire [WIDTH-1:0] wire_d31_11;
	wire [WIDTH-1:0] wire_d31_12;
	wire [WIDTH-1:0] wire_d31_13;
	wire [WIDTH-1:0] wire_d31_14;
	wire [WIDTH-1:0] wire_d31_15;
	wire [WIDTH-1:0] wire_d31_16;
	wire [WIDTH-1:0] wire_d31_17;
	wire [WIDTH-1:0] wire_d31_18;
	wire [WIDTH-1:0] wire_d31_19;
	wire [WIDTH-1:0] wire_d31_20;
	wire [WIDTH-1:0] wire_d31_21;
	wire [WIDTH-1:0] wire_d31_22;
	wire [WIDTH-1:0] wire_d31_23;
	wire [WIDTH-1:0] wire_d31_24;
	wire [WIDTH-1:0] wire_d31_25;
	wire [WIDTH-1:0] wire_d31_26;
	wire [WIDTH-1:0] wire_d31_27;
	wire [WIDTH-1:0] wire_d31_28;
	wire [WIDTH-1:0] wire_d31_29;
	wire [WIDTH-1:0] wire_d31_30;
	wire [WIDTH-1:0] wire_d31_31;
	wire [WIDTH-1:0] wire_d31_32;
	wire [WIDTH-1:0] wire_d31_33;
	wire [WIDTH-1:0] wire_d31_34;
	wire [WIDTH-1:0] wire_d31_35;
	wire [WIDTH-1:0] wire_d31_36;
	wire [WIDTH-1:0] wire_d31_37;
	wire [WIDTH-1:0] wire_d31_38;
	wire [WIDTH-1:0] wire_d31_39;
	wire [WIDTH-1:0] wire_d31_40;
	wire [WIDTH-1:0] wire_d31_41;
	wire [WIDTH-1:0] wire_d31_42;
	wire [WIDTH-1:0] wire_d31_43;
	wire [WIDTH-1:0] wire_d31_44;
	wire [WIDTH-1:0] wire_d31_45;
	wire [WIDTH-1:0] wire_d31_46;
	wire [WIDTH-1:0] wire_d31_47;
	wire [WIDTH-1:0] wire_d31_48;
	wire [WIDTH-1:0] wire_d31_49;
	wire [WIDTH-1:0] wire_d31_50;
	wire [WIDTH-1:0] wire_d31_51;
	wire [WIDTH-1:0] wire_d31_52;
	wire [WIDTH-1:0] wire_d31_53;
	wire [WIDTH-1:0] wire_d31_54;
	wire [WIDTH-1:0] wire_d31_55;
	wire [WIDTH-1:0] wire_d31_56;
	wire [WIDTH-1:0] wire_d31_57;
	wire [WIDTH-1:0] wire_d31_58;
	wire [WIDTH-1:0] wire_d31_59;
	wire [WIDTH-1:0] wire_d31_60;
	wire [WIDTH-1:0] wire_d31_61;
	wire [WIDTH-1:0] wire_d31_62;
	wire [WIDTH-1:0] wire_d31_63;
	wire [WIDTH-1:0] wire_d31_64;
	wire [WIDTH-1:0] wire_d31_65;
	wire [WIDTH-1:0] wire_d31_66;
	wire [WIDTH-1:0] wire_d31_67;
	wire [WIDTH-1:0] wire_d31_68;
	wire [WIDTH-1:0] wire_d31_69;
	wire [WIDTH-1:0] wire_d31_70;
	wire [WIDTH-1:0] wire_d31_71;
	wire [WIDTH-1:0] wire_d31_72;
	wire [WIDTH-1:0] wire_d31_73;
	wire [WIDTH-1:0] wire_d31_74;
	wire [WIDTH-1:0] wire_d31_75;
	wire [WIDTH-1:0] wire_d31_76;
	wire [WIDTH-1:0] wire_d31_77;
	wire [WIDTH-1:0] wire_d31_78;
	wire [WIDTH-1:0] wire_d32_0;
	wire [WIDTH-1:0] wire_d32_1;
	wire [WIDTH-1:0] wire_d32_2;
	wire [WIDTH-1:0] wire_d32_3;
	wire [WIDTH-1:0] wire_d32_4;
	wire [WIDTH-1:0] wire_d32_5;
	wire [WIDTH-1:0] wire_d32_6;
	wire [WIDTH-1:0] wire_d32_7;
	wire [WIDTH-1:0] wire_d32_8;
	wire [WIDTH-1:0] wire_d32_9;
	wire [WIDTH-1:0] wire_d32_10;
	wire [WIDTH-1:0] wire_d32_11;
	wire [WIDTH-1:0] wire_d32_12;
	wire [WIDTH-1:0] wire_d32_13;
	wire [WIDTH-1:0] wire_d32_14;
	wire [WIDTH-1:0] wire_d32_15;
	wire [WIDTH-1:0] wire_d32_16;
	wire [WIDTH-1:0] wire_d32_17;
	wire [WIDTH-1:0] wire_d32_18;
	wire [WIDTH-1:0] wire_d32_19;
	wire [WIDTH-1:0] wire_d32_20;
	wire [WIDTH-1:0] wire_d32_21;
	wire [WIDTH-1:0] wire_d32_22;
	wire [WIDTH-1:0] wire_d32_23;
	wire [WIDTH-1:0] wire_d32_24;
	wire [WIDTH-1:0] wire_d32_25;
	wire [WIDTH-1:0] wire_d32_26;
	wire [WIDTH-1:0] wire_d32_27;
	wire [WIDTH-1:0] wire_d32_28;
	wire [WIDTH-1:0] wire_d32_29;
	wire [WIDTH-1:0] wire_d32_30;
	wire [WIDTH-1:0] wire_d32_31;
	wire [WIDTH-1:0] wire_d32_32;
	wire [WIDTH-1:0] wire_d32_33;
	wire [WIDTH-1:0] wire_d32_34;
	wire [WIDTH-1:0] wire_d32_35;
	wire [WIDTH-1:0] wire_d32_36;
	wire [WIDTH-1:0] wire_d32_37;
	wire [WIDTH-1:0] wire_d32_38;
	wire [WIDTH-1:0] wire_d32_39;
	wire [WIDTH-1:0] wire_d32_40;
	wire [WIDTH-1:0] wire_d32_41;
	wire [WIDTH-1:0] wire_d32_42;
	wire [WIDTH-1:0] wire_d32_43;
	wire [WIDTH-1:0] wire_d32_44;
	wire [WIDTH-1:0] wire_d32_45;
	wire [WIDTH-1:0] wire_d32_46;
	wire [WIDTH-1:0] wire_d32_47;
	wire [WIDTH-1:0] wire_d32_48;
	wire [WIDTH-1:0] wire_d32_49;
	wire [WIDTH-1:0] wire_d32_50;
	wire [WIDTH-1:0] wire_d32_51;
	wire [WIDTH-1:0] wire_d32_52;
	wire [WIDTH-1:0] wire_d32_53;
	wire [WIDTH-1:0] wire_d32_54;
	wire [WIDTH-1:0] wire_d32_55;
	wire [WIDTH-1:0] wire_d32_56;
	wire [WIDTH-1:0] wire_d32_57;
	wire [WIDTH-1:0] wire_d32_58;
	wire [WIDTH-1:0] wire_d32_59;
	wire [WIDTH-1:0] wire_d32_60;
	wire [WIDTH-1:0] wire_d32_61;
	wire [WIDTH-1:0] wire_d32_62;
	wire [WIDTH-1:0] wire_d32_63;
	wire [WIDTH-1:0] wire_d32_64;
	wire [WIDTH-1:0] wire_d32_65;
	wire [WIDTH-1:0] wire_d32_66;
	wire [WIDTH-1:0] wire_d32_67;
	wire [WIDTH-1:0] wire_d32_68;
	wire [WIDTH-1:0] wire_d32_69;
	wire [WIDTH-1:0] wire_d32_70;
	wire [WIDTH-1:0] wire_d32_71;
	wire [WIDTH-1:0] wire_d32_72;
	wire [WIDTH-1:0] wire_d32_73;
	wire [WIDTH-1:0] wire_d32_74;
	wire [WIDTH-1:0] wire_d32_75;
	wire [WIDTH-1:0] wire_d32_76;
	wire [WIDTH-1:0] wire_d32_77;
	wire [WIDTH-1:0] wire_d32_78;
	wire [WIDTH-1:0] wire_d33_0;
	wire [WIDTH-1:0] wire_d33_1;
	wire [WIDTH-1:0] wire_d33_2;
	wire [WIDTH-1:0] wire_d33_3;
	wire [WIDTH-1:0] wire_d33_4;
	wire [WIDTH-1:0] wire_d33_5;
	wire [WIDTH-1:0] wire_d33_6;
	wire [WIDTH-1:0] wire_d33_7;
	wire [WIDTH-1:0] wire_d33_8;
	wire [WIDTH-1:0] wire_d33_9;
	wire [WIDTH-1:0] wire_d33_10;
	wire [WIDTH-1:0] wire_d33_11;
	wire [WIDTH-1:0] wire_d33_12;
	wire [WIDTH-1:0] wire_d33_13;
	wire [WIDTH-1:0] wire_d33_14;
	wire [WIDTH-1:0] wire_d33_15;
	wire [WIDTH-1:0] wire_d33_16;
	wire [WIDTH-1:0] wire_d33_17;
	wire [WIDTH-1:0] wire_d33_18;
	wire [WIDTH-1:0] wire_d33_19;
	wire [WIDTH-1:0] wire_d33_20;
	wire [WIDTH-1:0] wire_d33_21;
	wire [WIDTH-1:0] wire_d33_22;
	wire [WIDTH-1:0] wire_d33_23;
	wire [WIDTH-1:0] wire_d33_24;
	wire [WIDTH-1:0] wire_d33_25;
	wire [WIDTH-1:0] wire_d33_26;
	wire [WIDTH-1:0] wire_d33_27;
	wire [WIDTH-1:0] wire_d33_28;
	wire [WIDTH-1:0] wire_d33_29;
	wire [WIDTH-1:0] wire_d33_30;
	wire [WIDTH-1:0] wire_d33_31;
	wire [WIDTH-1:0] wire_d33_32;
	wire [WIDTH-1:0] wire_d33_33;
	wire [WIDTH-1:0] wire_d33_34;
	wire [WIDTH-1:0] wire_d33_35;
	wire [WIDTH-1:0] wire_d33_36;
	wire [WIDTH-1:0] wire_d33_37;
	wire [WIDTH-1:0] wire_d33_38;
	wire [WIDTH-1:0] wire_d33_39;
	wire [WIDTH-1:0] wire_d33_40;
	wire [WIDTH-1:0] wire_d33_41;
	wire [WIDTH-1:0] wire_d33_42;
	wire [WIDTH-1:0] wire_d33_43;
	wire [WIDTH-1:0] wire_d33_44;
	wire [WIDTH-1:0] wire_d33_45;
	wire [WIDTH-1:0] wire_d33_46;
	wire [WIDTH-1:0] wire_d33_47;
	wire [WIDTH-1:0] wire_d33_48;
	wire [WIDTH-1:0] wire_d33_49;
	wire [WIDTH-1:0] wire_d33_50;
	wire [WIDTH-1:0] wire_d33_51;
	wire [WIDTH-1:0] wire_d33_52;
	wire [WIDTH-1:0] wire_d33_53;
	wire [WIDTH-1:0] wire_d33_54;
	wire [WIDTH-1:0] wire_d33_55;
	wire [WIDTH-1:0] wire_d33_56;
	wire [WIDTH-1:0] wire_d33_57;
	wire [WIDTH-1:0] wire_d33_58;
	wire [WIDTH-1:0] wire_d33_59;
	wire [WIDTH-1:0] wire_d33_60;
	wire [WIDTH-1:0] wire_d33_61;
	wire [WIDTH-1:0] wire_d33_62;
	wire [WIDTH-1:0] wire_d33_63;
	wire [WIDTH-1:0] wire_d33_64;
	wire [WIDTH-1:0] wire_d33_65;
	wire [WIDTH-1:0] wire_d33_66;
	wire [WIDTH-1:0] wire_d33_67;
	wire [WIDTH-1:0] wire_d33_68;
	wire [WIDTH-1:0] wire_d33_69;
	wire [WIDTH-1:0] wire_d33_70;
	wire [WIDTH-1:0] wire_d33_71;
	wire [WIDTH-1:0] wire_d33_72;
	wire [WIDTH-1:0] wire_d33_73;
	wire [WIDTH-1:0] wire_d33_74;
	wire [WIDTH-1:0] wire_d33_75;
	wire [WIDTH-1:0] wire_d33_76;
	wire [WIDTH-1:0] wire_d33_77;
	wire [WIDTH-1:0] wire_d33_78;
	wire [WIDTH-1:0] wire_d34_0;
	wire [WIDTH-1:0] wire_d34_1;
	wire [WIDTH-1:0] wire_d34_2;
	wire [WIDTH-1:0] wire_d34_3;
	wire [WIDTH-1:0] wire_d34_4;
	wire [WIDTH-1:0] wire_d34_5;
	wire [WIDTH-1:0] wire_d34_6;
	wire [WIDTH-1:0] wire_d34_7;
	wire [WIDTH-1:0] wire_d34_8;
	wire [WIDTH-1:0] wire_d34_9;
	wire [WIDTH-1:0] wire_d34_10;
	wire [WIDTH-1:0] wire_d34_11;
	wire [WIDTH-1:0] wire_d34_12;
	wire [WIDTH-1:0] wire_d34_13;
	wire [WIDTH-1:0] wire_d34_14;
	wire [WIDTH-1:0] wire_d34_15;
	wire [WIDTH-1:0] wire_d34_16;
	wire [WIDTH-1:0] wire_d34_17;
	wire [WIDTH-1:0] wire_d34_18;
	wire [WIDTH-1:0] wire_d34_19;
	wire [WIDTH-1:0] wire_d34_20;
	wire [WIDTH-1:0] wire_d34_21;
	wire [WIDTH-1:0] wire_d34_22;
	wire [WIDTH-1:0] wire_d34_23;
	wire [WIDTH-1:0] wire_d34_24;
	wire [WIDTH-1:0] wire_d34_25;
	wire [WIDTH-1:0] wire_d34_26;
	wire [WIDTH-1:0] wire_d34_27;
	wire [WIDTH-1:0] wire_d34_28;
	wire [WIDTH-1:0] wire_d34_29;
	wire [WIDTH-1:0] wire_d34_30;
	wire [WIDTH-1:0] wire_d34_31;
	wire [WIDTH-1:0] wire_d34_32;
	wire [WIDTH-1:0] wire_d34_33;
	wire [WIDTH-1:0] wire_d34_34;
	wire [WIDTH-1:0] wire_d34_35;
	wire [WIDTH-1:0] wire_d34_36;
	wire [WIDTH-1:0] wire_d34_37;
	wire [WIDTH-1:0] wire_d34_38;
	wire [WIDTH-1:0] wire_d34_39;
	wire [WIDTH-1:0] wire_d34_40;
	wire [WIDTH-1:0] wire_d34_41;
	wire [WIDTH-1:0] wire_d34_42;
	wire [WIDTH-1:0] wire_d34_43;
	wire [WIDTH-1:0] wire_d34_44;
	wire [WIDTH-1:0] wire_d34_45;
	wire [WIDTH-1:0] wire_d34_46;
	wire [WIDTH-1:0] wire_d34_47;
	wire [WIDTH-1:0] wire_d34_48;
	wire [WIDTH-1:0] wire_d34_49;
	wire [WIDTH-1:0] wire_d34_50;
	wire [WIDTH-1:0] wire_d34_51;
	wire [WIDTH-1:0] wire_d34_52;
	wire [WIDTH-1:0] wire_d34_53;
	wire [WIDTH-1:0] wire_d34_54;
	wire [WIDTH-1:0] wire_d34_55;
	wire [WIDTH-1:0] wire_d34_56;
	wire [WIDTH-1:0] wire_d34_57;
	wire [WIDTH-1:0] wire_d34_58;
	wire [WIDTH-1:0] wire_d34_59;
	wire [WIDTH-1:0] wire_d34_60;
	wire [WIDTH-1:0] wire_d34_61;
	wire [WIDTH-1:0] wire_d34_62;
	wire [WIDTH-1:0] wire_d34_63;
	wire [WIDTH-1:0] wire_d34_64;
	wire [WIDTH-1:0] wire_d34_65;
	wire [WIDTH-1:0] wire_d34_66;
	wire [WIDTH-1:0] wire_d34_67;
	wire [WIDTH-1:0] wire_d34_68;
	wire [WIDTH-1:0] wire_d34_69;
	wire [WIDTH-1:0] wire_d34_70;
	wire [WIDTH-1:0] wire_d34_71;
	wire [WIDTH-1:0] wire_d34_72;
	wire [WIDTH-1:0] wire_d34_73;
	wire [WIDTH-1:0] wire_d34_74;
	wire [WIDTH-1:0] wire_d34_75;
	wire [WIDTH-1:0] wire_d34_76;
	wire [WIDTH-1:0] wire_d34_77;
	wire [WIDTH-1:0] wire_d34_78;
	wire [WIDTH-1:0] wire_d35_0;
	wire [WIDTH-1:0] wire_d35_1;
	wire [WIDTH-1:0] wire_d35_2;
	wire [WIDTH-1:0] wire_d35_3;
	wire [WIDTH-1:0] wire_d35_4;
	wire [WIDTH-1:0] wire_d35_5;
	wire [WIDTH-1:0] wire_d35_6;
	wire [WIDTH-1:0] wire_d35_7;
	wire [WIDTH-1:0] wire_d35_8;
	wire [WIDTH-1:0] wire_d35_9;
	wire [WIDTH-1:0] wire_d35_10;
	wire [WIDTH-1:0] wire_d35_11;
	wire [WIDTH-1:0] wire_d35_12;
	wire [WIDTH-1:0] wire_d35_13;
	wire [WIDTH-1:0] wire_d35_14;
	wire [WIDTH-1:0] wire_d35_15;
	wire [WIDTH-1:0] wire_d35_16;
	wire [WIDTH-1:0] wire_d35_17;
	wire [WIDTH-1:0] wire_d35_18;
	wire [WIDTH-1:0] wire_d35_19;
	wire [WIDTH-1:0] wire_d35_20;
	wire [WIDTH-1:0] wire_d35_21;
	wire [WIDTH-1:0] wire_d35_22;
	wire [WIDTH-1:0] wire_d35_23;
	wire [WIDTH-1:0] wire_d35_24;
	wire [WIDTH-1:0] wire_d35_25;
	wire [WIDTH-1:0] wire_d35_26;
	wire [WIDTH-1:0] wire_d35_27;
	wire [WIDTH-1:0] wire_d35_28;
	wire [WIDTH-1:0] wire_d35_29;
	wire [WIDTH-1:0] wire_d35_30;
	wire [WIDTH-1:0] wire_d35_31;
	wire [WIDTH-1:0] wire_d35_32;
	wire [WIDTH-1:0] wire_d35_33;
	wire [WIDTH-1:0] wire_d35_34;
	wire [WIDTH-1:0] wire_d35_35;
	wire [WIDTH-1:0] wire_d35_36;
	wire [WIDTH-1:0] wire_d35_37;
	wire [WIDTH-1:0] wire_d35_38;
	wire [WIDTH-1:0] wire_d35_39;
	wire [WIDTH-1:0] wire_d35_40;
	wire [WIDTH-1:0] wire_d35_41;
	wire [WIDTH-1:0] wire_d35_42;
	wire [WIDTH-1:0] wire_d35_43;
	wire [WIDTH-1:0] wire_d35_44;
	wire [WIDTH-1:0] wire_d35_45;
	wire [WIDTH-1:0] wire_d35_46;
	wire [WIDTH-1:0] wire_d35_47;
	wire [WIDTH-1:0] wire_d35_48;
	wire [WIDTH-1:0] wire_d35_49;
	wire [WIDTH-1:0] wire_d35_50;
	wire [WIDTH-1:0] wire_d35_51;
	wire [WIDTH-1:0] wire_d35_52;
	wire [WIDTH-1:0] wire_d35_53;
	wire [WIDTH-1:0] wire_d35_54;
	wire [WIDTH-1:0] wire_d35_55;
	wire [WIDTH-1:0] wire_d35_56;
	wire [WIDTH-1:0] wire_d35_57;
	wire [WIDTH-1:0] wire_d35_58;
	wire [WIDTH-1:0] wire_d35_59;
	wire [WIDTH-1:0] wire_d35_60;
	wire [WIDTH-1:0] wire_d35_61;
	wire [WIDTH-1:0] wire_d35_62;
	wire [WIDTH-1:0] wire_d35_63;
	wire [WIDTH-1:0] wire_d35_64;
	wire [WIDTH-1:0] wire_d35_65;
	wire [WIDTH-1:0] wire_d35_66;
	wire [WIDTH-1:0] wire_d35_67;
	wire [WIDTH-1:0] wire_d35_68;
	wire [WIDTH-1:0] wire_d35_69;
	wire [WIDTH-1:0] wire_d35_70;
	wire [WIDTH-1:0] wire_d35_71;
	wire [WIDTH-1:0] wire_d35_72;
	wire [WIDTH-1:0] wire_d35_73;
	wire [WIDTH-1:0] wire_d35_74;
	wire [WIDTH-1:0] wire_d35_75;
	wire [WIDTH-1:0] wire_d35_76;
	wire [WIDTH-1:0] wire_d35_77;
	wire [WIDTH-1:0] wire_d35_78;
	wire [WIDTH-1:0] wire_d36_0;
	wire [WIDTH-1:0] wire_d36_1;
	wire [WIDTH-1:0] wire_d36_2;
	wire [WIDTH-1:0] wire_d36_3;
	wire [WIDTH-1:0] wire_d36_4;
	wire [WIDTH-1:0] wire_d36_5;
	wire [WIDTH-1:0] wire_d36_6;
	wire [WIDTH-1:0] wire_d36_7;
	wire [WIDTH-1:0] wire_d36_8;
	wire [WIDTH-1:0] wire_d36_9;
	wire [WIDTH-1:0] wire_d36_10;
	wire [WIDTH-1:0] wire_d36_11;
	wire [WIDTH-1:0] wire_d36_12;
	wire [WIDTH-1:0] wire_d36_13;
	wire [WIDTH-1:0] wire_d36_14;
	wire [WIDTH-1:0] wire_d36_15;
	wire [WIDTH-1:0] wire_d36_16;
	wire [WIDTH-1:0] wire_d36_17;
	wire [WIDTH-1:0] wire_d36_18;
	wire [WIDTH-1:0] wire_d36_19;
	wire [WIDTH-1:0] wire_d36_20;
	wire [WIDTH-1:0] wire_d36_21;
	wire [WIDTH-1:0] wire_d36_22;
	wire [WIDTH-1:0] wire_d36_23;
	wire [WIDTH-1:0] wire_d36_24;
	wire [WIDTH-1:0] wire_d36_25;
	wire [WIDTH-1:0] wire_d36_26;
	wire [WIDTH-1:0] wire_d36_27;
	wire [WIDTH-1:0] wire_d36_28;
	wire [WIDTH-1:0] wire_d36_29;
	wire [WIDTH-1:0] wire_d36_30;
	wire [WIDTH-1:0] wire_d36_31;
	wire [WIDTH-1:0] wire_d36_32;
	wire [WIDTH-1:0] wire_d36_33;
	wire [WIDTH-1:0] wire_d36_34;
	wire [WIDTH-1:0] wire_d36_35;
	wire [WIDTH-1:0] wire_d36_36;
	wire [WIDTH-1:0] wire_d36_37;
	wire [WIDTH-1:0] wire_d36_38;
	wire [WIDTH-1:0] wire_d36_39;
	wire [WIDTH-1:0] wire_d36_40;
	wire [WIDTH-1:0] wire_d36_41;
	wire [WIDTH-1:0] wire_d36_42;
	wire [WIDTH-1:0] wire_d36_43;
	wire [WIDTH-1:0] wire_d36_44;
	wire [WIDTH-1:0] wire_d36_45;
	wire [WIDTH-1:0] wire_d36_46;
	wire [WIDTH-1:0] wire_d36_47;
	wire [WIDTH-1:0] wire_d36_48;
	wire [WIDTH-1:0] wire_d36_49;
	wire [WIDTH-1:0] wire_d36_50;
	wire [WIDTH-1:0] wire_d36_51;
	wire [WIDTH-1:0] wire_d36_52;
	wire [WIDTH-1:0] wire_d36_53;
	wire [WIDTH-1:0] wire_d36_54;
	wire [WIDTH-1:0] wire_d36_55;
	wire [WIDTH-1:0] wire_d36_56;
	wire [WIDTH-1:0] wire_d36_57;
	wire [WIDTH-1:0] wire_d36_58;
	wire [WIDTH-1:0] wire_d36_59;
	wire [WIDTH-1:0] wire_d36_60;
	wire [WIDTH-1:0] wire_d36_61;
	wire [WIDTH-1:0] wire_d36_62;
	wire [WIDTH-1:0] wire_d36_63;
	wire [WIDTH-1:0] wire_d36_64;
	wire [WIDTH-1:0] wire_d36_65;
	wire [WIDTH-1:0] wire_d36_66;
	wire [WIDTH-1:0] wire_d36_67;
	wire [WIDTH-1:0] wire_d36_68;
	wire [WIDTH-1:0] wire_d36_69;
	wire [WIDTH-1:0] wire_d36_70;
	wire [WIDTH-1:0] wire_d36_71;
	wire [WIDTH-1:0] wire_d36_72;
	wire [WIDTH-1:0] wire_d36_73;
	wire [WIDTH-1:0] wire_d36_74;
	wire [WIDTH-1:0] wire_d36_75;
	wire [WIDTH-1:0] wire_d36_76;
	wire [WIDTH-1:0] wire_d36_77;
	wire [WIDTH-1:0] wire_d36_78;
	wire [WIDTH-1:0] wire_d37_0;
	wire [WIDTH-1:0] wire_d37_1;
	wire [WIDTH-1:0] wire_d37_2;
	wire [WIDTH-1:0] wire_d37_3;
	wire [WIDTH-1:0] wire_d37_4;
	wire [WIDTH-1:0] wire_d37_5;
	wire [WIDTH-1:0] wire_d37_6;
	wire [WIDTH-1:0] wire_d37_7;
	wire [WIDTH-1:0] wire_d37_8;
	wire [WIDTH-1:0] wire_d37_9;
	wire [WIDTH-1:0] wire_d37_10;
	wire [WIDTH-1:0] wire_d37_11;
	wire [WIDTH-1:0] wire_d37_12;
	wire [WIDTH-1:0] wire_d37_13;
	wire [WIDTH-1:0] wire_d37_14;
	wire [WIDTH-1:0] wire_d37_15;
	wire [WIDTH-1:0] wire_d37_16;
	wire [WIDTH-1:0] wire_d37_17;
	wire [WIDTH-1:0] wire_d37_18;
	wire [WIDTH-1:0] wire_d37_19;
	wire [WIDTH-1:0] wire_d37_20;
	wire [WIDTH-1:0] wire_d37_21;
	wire [WIDTH-1:0] wire_d37_22;
	wire [WIDTH-1:0] wire_d37_23;
	wire [WIDTH-1:0] wire_d37_24;
	wire [WIDTH-1:0] wire_d37_25;
	wire [WIDTH-1:0] wire_d37_26;
	wire [WIDTH-1:0] wire_d37_27;
	wire [WIDTH-1:0] wire_d37_28;
	wire [WIDTH-1:0] wire_d37_29;
	wire [WIDTH-1:0] wire_d37_30;
	wire [WIDTH-1:0] wire_d37_31;
	wire [WIDTH-1:0] wire_d37_32;
	wire [WIDTH-1:0] wire_d37_33;
	wire [WIDTH-1:0] wire_d37_34;
	wire [WIDTH-1:0] wire_d37_35;
	wire [WIDTH-1:0] wire_d37_36;
	wire [WIDTH-1:0] wire_d37_37;
	wire [WIDTH-1:0] wire_d37_38;
	wire [WIDTH-1:0] wire_d37_39;
	wire [WIDTH-1:0] wire_d37_40;
	wire [WIDTH-1:0] wire_d37_41;
	wire [WIDTH-1:0] wire_d37_42;
	wire [WIDTH-1:0] wire_d37_43;
	wire [WIDTH-1:0] wire_d37_44;
	wire [WIDTH-1:0] wire_d37_45;
	wire [WIDTH-1:0] wire_d37_46;
	wire [WIDTH-1:0] wire_d37_47;
	wire [WIDTH-1:0] wire_d37_48;
	wire [WIDTH-1:0] wire_d37_49;
	wire [WIDTH-1:0] wire_d37_50;
	wire [WIDTH-1:0] wire_d37_51;
	wire [WIDTH-1:0] wire_d37_52;
	wire [WIDTH-1:0] wire_d37_53;
	wire [WIDTH-1:0] wire_d37_54;
	wire [WIDTH-1:0] wire_d37_55;
	wire [WIDTH-1:0] wire_d37_56;
	wire [WIDTH-1:0] wire_d37_57;
	wire [WIDTH-1:0] wire_d37_58;
	wire [WIDTH-1:0] wire_d37_59;
	wire [WIDTH-1:0] wire_d37_60;
	wire [WIDTH-1:0] wire_d37_61;
	wire [WIDTH-1:0] wire_d37_62;
	wire [WIDTH-1:0] wire_d37_63;
	wire [WIDTH-1:0] wire_d37_64;
	wire [WIDTH-1:0] wire_d37_65;
	wire [WIDTH-1:0] wire_d37_66;
	wire [WIDTH-1:0] wire_d37_67;
	wire [WIDTH-1:0] wire_d37_68;
	wire [WIDTH-1:0] wire_d37_69;
	wire [WIDTH-1:0] wire_d37_70;
	wire [WIDTH-1:0] wire_d37_71;
	wire [WIDTH-1:0] wire_d37_72;
	wire [WIDTH-1:0] wire_d37_73;
	wire [WIDTH-1:0] wire_d37_74;
	wire [WIDTH-1:0] wire_d37_75;
	wire [WIDTH-1:0] wire_d37_76;
	wire [WIDTH-1:0] wire_d37_77;
	wire [WIDTH-1:0] wire_d37_78;
	wire [WIDTH-1:0] wire_d38_0;
	wire [WIDTH-1:0] wire_d38_1;
	wire [WIDTH-1:0] wire_d38_2;
	wire [WIDTH-1:0] wire_d38_3;
	wire [WIDTH-1:0] wire_d38_4;
	wire [WIDTH-1:0] wire_d38_5;
	wire [WIDTH-1:0] wire_d38_6;
	wire [WIDTH-1:0] wire_d38_7;
	wire [WIDTH-1:0] wire_d38_8;
	wire [WIDTH-1:0] wire_d38_9;
	wire [WIDTH-1:0] wire_d38_10;
	wire [WIDTH-1:0] wire_d38_11;
	wire [WIDTH-1:0] wire_d38_12;
	wire [WIDTH-1:0] wire_d38_13;
	wire [WIDTH-1:0] wire_d38_14;
	wire [WIDTH-1:0] wire_d38_15;
	wire [WIDTH-1:0] wire_d38_16;
	wire [WIDTH-1:0] wire_d38_17;
	wire [WIDTH-1:0] wire_d38_18;
	wire [WIDTH-1:0] wire_d38_19;
	wire [WIDTH-1:0] wire_d38_20;
	wire [WIDTH-1:0] wire_d38_21;
	wire [WIDTH-1:0] wire_d38_22;
	wire [WIDTH-1:0] wire_d38_23;
	wire [WIDTH-1:0] wire_d38_24;
	wire [WIDTH-1:0] wire_d38_25;
	wire [WIDTH-1:0] wire_d38_26;
	wire [WIDTH-1:0] wire_d38_27;
	wire [WIDTH-1:0] wire_d38_28;
	wire [WIDTH-1:0] wire_d38_29;
	wire [WIDTH-1:0] wire_d38_30;
	wire [WIDTH-1:0] wire_d38_31;
	wire [WIDTH-1:0] wire_d38_32;
	wire [WIDTH-1:0] wire_d38_33;
	wire [WIDTH-1:0] wire_d38_34;
	wire [WIDTH-1:0] wire_d38_35;
	wire [WIDTH-1:0] wire_d38_36;
	wire [WIDTH-1:0] wire_d38_37;
	wire [WIDTH-1:0] wire_d38_38;
	wire [WIDTH-1:0] wire_d38_39;
	wire [WIDTH-1:0] wire_d38_40;
	wire [WIDTH-1:0] wire_d38_41;
	wire [WIDTH-1:0] wire_d38_42;
	wire [WIDTH-1:0] wire_d38_43;
	wire [WIDTH-1:0] wire_d38_44;
	wire [WIDTH-1:0] wire_d38_45;
	wire [WIDTH-1:0] wire_d38_46;
	wire [WIDTH-1:0] wire_d38_47;
	wire [WIDTH-1:0] wire_d38_48;
	wire [WIDTH-1:0] wire_d38_49;
	wire [WIDTH-1:0] wire_d38_50;
	wire [WIDTH-1:0] wire_d38_51;
	wire [WIDTH-1:0] wire_d38_52;
	wire [WIDTH-1:0] wire_d38_53;
	wire [WIDTH-1:0] wire_d38_54;
	wire [WIDTH-1:0] wire_d38_55;
	wire [WIDTH-1:0] wire_d38_56;
	wire [WIDTH-1:0] wire_d38_57;
	wire [WIDTH-1:0] wire_d38_58;
	wire [WIDTH-1:0] wire_d38_59;
	wire [WIDTH-1:0] wire_d38_60;
	wire [WIDTH-1:0] wire_d38_61;
	wire [WIDTH-1:0] wire_d38_62;
	wire [WIDTH-1:0] wire_d38_63;
	wire [WIDTH-1:0] wire_d38_64;
	wire [WIDTH-1:0] wire_d38_65;
	wire [WIDTH-1:0] wire_d38_66;
	wire [WIDTH-1:0] wire_d38_67;
	wire [WIDTH-1:0] wire_d38_68;
	wire [WIDTH-1:0] wire_d38_69;
	wire [WIDTH-1:0] wire_d38_70;
	wire [WIDTH-1:0] wire_d38_71;
	wire [WIDTH-1:0] wire_d38_72;
	wire [WIDTH-1:0] wire_d38_73;
	wire [WIDTH-1:0] wire_d38_74;
	wire [WIDTH-1:0] wire_d38_75;
	wire [WIDTH-1:0] wire_d38_76;
	wire [WIDTH-1:0] wire_d38_77;
	wire [WIDTH-1:0] wire_d38_78;
	wire [WIDTH-1:0] wire_d39_0;
	wire [WIDTH-1:0] wire_d39_1;
	wire [WIDTH-1:0] wire_d39_2;
	wire [WIDTH-1:0] wire_d39_3;
	wire [WIDTH-1:0] wire_d39_4;
	wire [WIDTH-1:0] wire_d39_5;
	wire [WIDTH-1:0] wire_d39_6;
	wire [WIDTH-1:0] wire_d39_7;
	wire [WIDTH-1:0] wire_d39_8;
	wire [WIDTH-1:0] wire_d39_9;
	wire [WIDTH-1:0] wire_d39_10;
	wire [WIDTH-1:0] wire_d39_11;
	wire [WIDTH-1:0] wire_d39_12;
	wire [WIDTH-1:0] wire_d39_13;
	wire [WIDTH-1:0] wire_d39_14;
	wire [WIDTH-1:0] wire_d39_15;
	wire [WIDTH-1:0] wire_d39_16;
	wire [WIDTH-1:0] wire_d39_17;
	wire [WIDTH-1:0] wire_d39_18;
	wire [WIDTH-1:0] wire_d39_19;
	wire [WIDTH-1:0] wire_d39_20;
	wire [WIDTH-1:0] wire_d39_21;
	wire [WIDTH-1:0] wire_d39_22;
	wire [WIDTH-1:0] wire_d39_23;
	wire [WIDTH-1:0] wire_d39_24;
	wire [WIDTH-1:0] wire_d39_25;
	wire [WIDTH-1:0] wire_d39_26;
	wire [WIDTH-1:0] wire_d39_27;
	wire [WIDTH-1:0] wire_d39_28;
	wire [WIDTH-1:0] wire_d39_29;
	wire [WIDTH-1:0] wire_d39_30;
	wire [WIDTH-1:0] wire_d39_31;
	wire [WIDTH-1:0] wire_d39_32;
	wire [WIDTH-1:0] wire_d39_33;
	wire [WIDTH-1:0] wire_d39_34;
	wire [WIDTH-1:0] wire_d39_35;
	wire [WIDTH-1:0] wire_d39_36;
	wire [WIDTH-1:0] wire_d39_37;
	wire [WIDTH-1:0] wire_d39_38;
	wire [WIDTH-1:0] wire_d39_39;
	wire [WIDTH-1:0] wire_d39_40;
	wire [WIDTH-1:0] wire_d39_41;
	wire [WIDTH-1:0] wire_d39_42;
	wire [WIDTH-1:0] wire_d39_43;
	wire [WIDTH-1:0] wire_d39_44;
	wire [WIDTH-1:0] wire_d39_45;
	wire [WIDTH-1:0] wire_d39_46;
	wire [WIDTH-1:0] wire_d39_47;
	wire [WIDTH-1:0] wire_d39_48;
	wire [WIDTH-1:0] wire_d39_49;
	wire [WIDTH-1:0] wire_d39_50;
	wire [WIDTH-1:0] wire_d39_51;
	wire [WIDTH-1:0] wire_d39_52;
	wire [WIDTH-1:0] wire_d39_53;
	wire [WIDTH-1:0] wire_d39_54;
	wire [WIDTH-1:0] wire_d39_55;
	wire [WIDTH-1:0] wire_d39_56;
	wire [WIDTH-1:0] wire_d39_57;
	wire [WIDTH-1:0] wire_d39_58;
	wire [WIDTH-1:0] wire_d39_59;
	wire [WIDTH-1:0] wire_d39_60;
	wire [WIDTH-1:0] wire_d39_61;
	wire [WIDTH-1:0] wire_d39_62;
	wire [WIDTH-1:0] wire_d39_63;
	wire [WIDTH-1:0] wire_d39_64;
	wire [WIDTH-1:0] wire_d39_65;
	wire [WIDTH-1:0] wire_d39_66;
	wire [WIDTH-1:0] wire_d39_67;
	wire [WIDTH-1:0] wire_d39_68;
	wire [WIDTH-1:0] wire_d39_69;
	wire [WIDTH-1:0] wire_d39_70;
	wire [WIDTH-1:0] wire_d39_71;
	wire [WIDTH-1:0] wire_d39_72;
	wire [WIDTH-1:0] wire_d39_73;
	wire [WIDTH-1:0] wire_d39_74;
	wire [WIDTH-1:0] wire_d39_75;
	wire [WIDTH-1:0] wire_d39_76;
	wire [WIDTH-1:0] wire_d39_77;
	wire [WIDTH-1:0] wire_d39_78;
	wire [WIDTH-1:0] wire_d40_0;
	wire [WIDTH-1:0] wire_d40_1;
	wire [WIDTH-1:0] wire_d40_2;
	wire [WIDTH-1:0] wire_d40_3;
	wire [WIDTH-1:0] wire_d40_4;
	wire [WIDTH-1:0] wire_d40_5;
	wire [WIDTH-1:0] wire_d40_6;
	wire [WIDTH-1:0] wire_d40_7;
	wire [WIDTH-1:0] wire_d40_8;
	wire [WIDTH-1:0] wire_d40_9;
	wire [WIDTH-1:0] wire_d40_10;
	wire [WIDTH-1:0] wire_d40_11;
	wire [WIDTH-1:0] wire_d40_12;
	wire [WIDTH-1:0] wire_d40_13;
	wire [WIDTH-1:0] wire_d40_14;
	wire [WIDTH-1:0] wire_d40_15;
	wire [WIDTH-1:0] wire_d40_16;
	wire [WIDTH-1:0] wire_d40_17;
	wire [WIDTH-1:0] wire_d40_18;
	wire [WIDTH-1:0] wire_d40_19;
	wire [WIDTH-1:0] wire_d40_20;
	wire [WIDTH-1:0] wire_d40_21;
	wire [WIDTH-1:0] wire_d40_22;
	wire [WIDTH-1:0] wire_d40_23;
	wire [WIDTH-1:0] wire_d40_24;
	wire [WIDTH-1:0] wire_d40_25;
	wire [WIDTH-1:0] wire_d40_26;
	wire [WIDTH-1:0] wire_d40_27;
	wire [WIDTH-1:0] wire_d40_28;
	wire [WIDTH-1:0] wire_d40_29;
	wire [WIDTH-1:0] wire_d40_30;
	wire [WIDTH-1:0] wire_d40_31;
	wire [WIDTH-1:0] wire_d40_32;
	wire [WIDTH-1:0] wire_d40_33;
	wire [WIDTH-1:0] wire_d40_34;
	wire [WIDTH-1:0] wire_d40_35;
	wire [WIDTH-1:0] wire_d40_36;
	wire [WIDTH-1:0] wire_d40_37;
	wire [WIDTH-1:0] wire_d40_38;
	wire [WIDTH-1:0] wire_d40_39;
	wire [WIDTH-1:0] wire_d40_40;
	wire [WIDTH-1:0] wire_d40_41;
	wire [WIDTH-1:0] wire_d40_42;
	wire [WIDTH-1:0] wire_d40_43;
	wire [WIDTH-1:0] wire_d40_44;
	wire [WIDTH-1:0] wire_d40_45;
	wire [WIDTH-1:0] wire_d40_46;
	wire [WIDTH-1:0] wire_d40_47;
	wire [WIDTH-1:0] wire_d40_48;
	wire [WIDTH-1:0] wire_d40_49;
	wire [WIDTH-1:0] wire_d40_50;
	wire [WIDTH-1:0] wire_d40_51;
	wire [WIDTH-1:0] wire_d40_52;
	wire [WIDTH-1:0] wire_d40_53;
	wire [WIDTH-1:0] wire_d40_54;
	wire [WIDTH-1:0] wire_d40_55;
	wire [WIDTH-1:0] wire_d40_56;
	wire [WIDTH-1:0] wire_d40_57;
	wire [WIDTH-1:0] wire_d40_58;
	wire [WIDTH-1:0] wire_d40_59;
	wire [WIDTH-1:0] wire_d40_60;
	wire [WIDTH-1:0] wire_d40_61;
	wire [WIDTH-1:0] wire_d40_62;
	wire [WIDTH-1:0] wire_d40_63;
	wire [WIDTH-1:0] wire_d40_64;
	wire [WIDTH-1:0] wire_d40_65;
	wire [WIDTH-1:0] wire_d40_66;
	wire [WIDTH-1:0] wire_d40_67;
	wire [WIDTH-1:0] wire_d40_68;
	wire [WIDTH-1:0] wire_d40_69;
	wire [WIDTH-1:0] wire_d40_70;
	wire [WIDTH-1:0] wire_d40_71;
	wire [WIDTH-1:0] wire_d40_72;
	wire [WIDTH-1:0] wire_d40_73;
	wire [WIDTH-1:0] wire_d40_74;
	wire [WIDTH-1:0] wire_d40_75;
	wire [WIDTH-1:0] wire_d40_76;
	wire [WIDTH-1:0] wire_d40_77;
	wire [WIDTH-1:0] wire_d40_78;
	wire [WIDTH-1:0] wire_d41_0;
	wire [WIDTH-1:0] wire_d41_1;
	wire [WIDTH-1:0] wire_d41_2;
	wire [WIDTH-1:0] wire_d41_3;
	wire [WIDTH-1:0] wire_d41_4;
	wire [WIDTH-1:0] wire_d41_5;
	wire [WIDTH-1:0] wire_d41_6;
	wire [WIDTH-1:0] wire_d41_7;
	wire [WIDTH-1:0] wire_d41_8;
	wire [WIDTH-1:0] wire_d41_9;
	wire [WIDTH-1:0] wire_d41_10;
	wire [WIDTH-1:0] wire_d41_11;
	wire [WIDTH-1:0] wire_d41_12;
	wire [WIDTH-1:0] wire_d41_13;
	wire [WIDTH-1:0] wire_d41_14;
	wire [WIDTH-1:0] wire_d41_15;
	wire [WIDTH-1:0] wire_d41_16;
	wire [WIDTH-1:0] wire_d41_17;
	wire [WIDTH-1:0] wire_d41_18;
	wire [WIDTH-1:0] wire_d41_19;
	wire [WIDTH-1:0] wire_d41_20;
	wire [WIDTH-1:0] wire_d41_21;
	wire [WIDTH-1:0] wire_d41_22;
	wire [WIDTH-1:0] wire_d41_23;
	wire [WIDTH-1:0] wire_d41_24;
	wire [WIDTH-1:0] wire_d41_25;
	wire [WIDTH-1:0] wire_d41_26;
	wire [WIDTH-1:0] wire_d41_27;
	wire [WIDTH-1:0] wire_d41_28;
	wire [WIDTH-1:0] wire_d41_29;
	wire [WIDTH-1:0] wire_d41_30;
	wire [WIDTH-1:0] wire_d41_31;
	wire [WIDTH-1:0] wire_d41_32;
	wire [WIDTH-1:0] wire_d41_33;
	wire [WIDTH-1:0] wire_d41_34;
	wire [WIDTH-1:0] wire_d41_35;
	wire [WIDTH-1:0] wire_d41_36;
	wire [WIDTH-1:0] wire_d41_37;
	wire [WIDTH-1:0] wire_d41_38;
	wire [WIDTH-1:0] wire_d41_39;
	wire [WIDTH-1:0] wire_d41_40;
	wire [WIDTH-1:0] wire_d41_41;
	wire [WIDTH-1:0] wire_d41_42;
	wire [WIDTH-1:0] wire_d41_43;
	wire [WIDTH-1:0] wire_d41_44;
	wire [WIDTH-1:0] wire_d41_45;
	wire [WIDTH-1:0] wire_d41_46;
	wire [WIDTH-1:0] wire_d41_47;
	wire [WIDTH-1:0] wire_d41_48;
	wire [WIDTH-1:0] wire_d41_49;
	wire [WIDTH-1:0] wire_d41_50;
	wire [WIDTH-1:0] wire_d41_51;
	wire [WIDTH-1:0] wire_d41_52;
	wire [WIDTH-1:0] wire_d41_53;
	wire [WIDTH-1:0] wire_d41_54;
	wire [WIDTH-1:0] wire_d41_55;
	wire [WIDTH-1:0] wire_d41_56;
	wire [WIDTH-1:0] wire_d41_57;
	wire [WIDTH-1:0] wire_d41_58;
	wire [WIDTH-1:0] wire_d41_59;
	wire [WIDTH-1:0] wire_d41_60;
	wire [WIDTH-1:0] wire_d41_61;
	wire [WIDTH-1:0] wire_d41_62;
	wire [WIDTH-1:0] wire_d41_63;
	wire [WIDTH-1:0] wire_d41_64;
	wire [WIDTH-1:0] wire_d41_65;
	wire [WIDTH-1:0] wire_d41_66;
	wire [WIDTH-1:0] wire_d41_67;
	wire [WIDTH-1:0] wire_d41_68;
	wire [WIDTH-1:0] wire_d41_69;
	wire [WIDTH-1:0] wire_d41_70;
	wire [WIDTH-1:0] wire_d41_71;
	wire [WIDTH-1:0] wire_d41_72;
	wire [WIDTH-1:0] wire_d41_73;
	wire [WIDTH-1:0] wire_d41_74;
	wire [WIDTH-1:0] wire_d41_75;
	wire [WIDTH-1:0] wire_d41_76;
	wire [WIDTH-1:0] wire_d41_77;
	wire [WIDTH-1:0] wire_d41_78;
	wire [WIDTH-1:0] wire_d42_0;
	wire [WIDTH-1:0] wire_d42_1;
	wire [WIDTH-1:0] wire_d42_2;
	wire [WIDTH-1:0] wire_d42_3;
	wire [WIDTH-1:0] wire_d42_4;
	wire [WIDTH-1:0] wire_d42_5;
	wire [WIDTH-1:0] wire_d42_6;
	wire [WIDTH-1:0] wire_d42_7;
	wire [WIDTH-1:0] wire_d42_8;
	wire [WIDTH-1:0] wire_d42_9;
	wire [WIDTH-1:0] wire_d42_10;
	wire [WIDTH-1:0] wire_d42_11;
	wire [WIDTH-1:0] wire_d42_12;
	wire [WIDTH-1:0] wire_d42_13;
	wire [WIDTH-1:0] wire_d42_14;
	wire [WIDTH-1:0] wire_d42_15;
	wire [WIDTH-1:0] wire_d42_16;
	wire [WIDTH-1:0] wire_d42_17;
	wire [WIDTH-1:0] wire_d42_18;
	wire [WIDTH-1:0] wire_d42_19;
	wire [WIDTH-1:0] wire_d42_20;
	wire [WIDTH-1:0] wire_d42_21;
	wire [WIDTH-1:0] wire_d42_22;
	wire [WIDTH-1:0] wire_d42_23;
	wire [WIDTH-1:0] wire_d42_24;
	wire [WIDTH-1:0] wire_d42_25;
	wire [WIDTH-1:0] wire_d42_26;
	wire [WIDTH-1:0] wire_d42_27;
	wire [WIDTH-1:0] wire_d42_28;
	wire [WIDTH-1:0] wire_d42_29;
	wire [WIDTH-1:0] wire_d42_30;
	wire [WIDTH-1:0] wire_d42_31;
	wire [WIDTH-1:0] wire_d42_32;
	wire [WIDTH-1:0] wire_d42_33;
	wire [WIDTH-1:0] wire_d42_34;
	wire [WIDTH-1:0] wire_d42_35;
	wire [WIDTH-1:0] wire_d42_36;
	wire [WIDTH-1:0] wire_d42_37;
	wire [WIDTH-1:0] wire_d42_38;
	wire [WIDTH-1:0] wire_d42_39;
	wire [WIDTH-1:0] wire_d42_40;
	wire [WIDTH-1:0] wire_d42_41;
	wire [WIDTH-1:0] wire_d42_42;
	wire [WIDTH-1:0] wire_d42_43;
	wire [WIDTH-1:0] wire_d42_44;
	wire [WIDTH-1:0] wire_d42_45;
	wire [WIDTH-1:0] wire_d42_46;
	wire [WIDTH-1:0] wire_d42_47;
	wire [WIDTH-1:0] wire_d42_48;
	wire [WIDTH-1:0] wire_d42_49;
	wire [WIDTH-1:0] wire_d42_50;
	wire [WIDTH-1:0] wire_d42_51;
	wire [WIDTH-1:0] wire_d42_52;
	wire [WIDTH-1:0] wire_d42_53;
	wire [WIDTH-1:0] wire_d42_54;
	wire [WIDTH-1:0] wire_d42_55;
	wire [WIDTH-1:0] wire_d42_56;
	wire [WIDTH-1:0] wire_d42_57;
	wire [WIDTH-1:0] wire_d42_58;
	wire [WIDTH-1:0] wire_d42_59;
	wire [WIDTH-1:0] wire_d42_60;
	wire [WIDTH-1:0] wire_d42_61;
	wire [WIDTH-1:0] wire_d42_62;
	wire [WIDTH-1:0] wire_d42_63;
	wire [WIDTH-1:0] wire_d42_64;
	wire [WIDTH-1:0] wire_d42_65;
	wire [WIDTH-1:0] wire_d42_66;
	wire [WIDTH-1:0] wire_d42_67;
	wire [WIDTH-1:0] wire_d42_68;
	wire [WIDTH-1:0] wire_d42_69;
	wire [WIDTH-1:0] wire_d42_70;
	wire [WIDTH-1:0] wire_d42_71;
	wire [WIDTH-1:0] wire_d42_72;
	wire [WIDTH-1:0] wire_d42_73;
	wire [WIDTH-1:0] wire_d42_74;
	wire [WIDTH-1:0] wire_d42_75;
	wire [WIDTH-1:0] wire_d42_76;
	wire [WIDTH-1:0] wire_d42_77;
	wire [WIDTH-1:0] wire_d42_78;
	wire [WIDTH-1:0] wire_d43_0;
	wire [WIDTH-1:0] wire_d43_1;
	wire [WIDTH-1:0] wire_d43_2;
	wire [WIDTH-1:0] wire_d43_3;
	wire [WIDTH-1:0] wire_d43_4;
	wire [WIDTH-1:0] wire_d43_5;
	wire [WIDTH-1:0] wire_d43_6;
	wire [WIDTH-1:0] wire_d43_7;
	wire [WIDTH-1:0] wire_d43_8;
	wire [WIDTH-1:0] wire_d43_9;
	wire [WIDTH-1:0] wire_d43_10;
	wire [WIDTH-1:0] wire_d43_11;
	wire [WIDTH-1:0] wire_d43_12;
	wire [WIDTH-1:0] wire_d43_13;
	wire [WIDTH-1:0] wire_d43_14;
	wire [WIDTH-1:0] wire_d43_15;
	wire [WIDTH-1:0] wire_d43_16;
	wire [WIDTH-1:0] wire_d43_17;
	wire [WIDTH-1:0] wire_d43_18;
	wire [WIDTH-1:0] wire_d43_19;
	wire [WIDTH-1:0] wire_d43_20;
	wire [WIDTH-1:0] wire_d43_21;
	wire [WIDTH-1:0] wire_d43_22;
	wire [WIDTH-1:0] wire_d43_23;
	wire [WIDTH-1:0] wire_d43_24;
	wire [WIDTH-1:0] wire_d43_25;
	wire [WIDTH-1:0] wire_d43_26;
	wire [WIDTH-1:0] wire_d43_27;
	wire [WIDTH-1:0] wire_d43_28;
	wire [WIDTH-1:0] wire_d43_29;
	wire [WIDTH-1:0] wire_d43_30;
	wire [WIDTH-1:0] wire_d43_31;
	wire [WIDTH-1:0] wire_d43_32;
	wire [WIDTH-1:0] wire_d43_33;
	wire [WIDTH-1:0] wire_d43_34;
	wire [WIDTH-1:0] wire_d43_35;
	wire [WIDTH-1:0] wire_d43_36;
	wire [WIDTH-1:0] wire_d43_37;
	wire [WIDTH-1:0] wire_d43_38;
	wire [WIDTH-1:0] wire_d43_39;
	wire [WIDTH-1:0] wire_d43_40;
	wire [WIDTH-1:0] wire_d43_41;
	wire [WIDTH-1:0] wire_d43_42;
	wire [WIDTH-1:0] wire_d43_43;
	wire [WIDTH-1:0] wire_d43_44;
	wire [WIDTH-1:0] wire_d43_45;
	wire [WIDTH-1:0] wire_d43_46;
	wire [WIDTH-1:0] wire_d43_47;
	wire [WIDTH-1:0] wire_d43_48;
	wire [WIDTH-1:0] wire_d43_49;
	wire [WIDTH-1:0] wire_d43_50;
	wire [WIDTH-1:0] wire_d43_51;
	wire [WIDTH-1:0] wire_d43_52;
	wire [WIDTH-1:0] wire_d43_53;
	wire [WIDTH-1:0] wire_d43_54;
	wire [WIDTH-1:0] wire_d43_55;
	wire [WIDTH-1:0] wire_d43_56;
	wire [WIDTH-1:0] wire_d43_57;
	wire [WIDTH-1:0] wire_d43_58;
	wire [WIDTH-1:0] wire_d43_59;
	wire [WIDTH-1:0] wire_d43_60;
	wire [WIDTH-1:0] wire_d43_61;
	wire [WIDTH-1:0] wire_d43_62;
	wire [WIDTH-1:0] wire_d43_63;
	wire [WIDTH-1:0] wire_d43_64;
	wire [WIDTH-1:0] wire_d43_65;
	wire [WIDTH-1:0] wire_d43_66;
	wire [WIDTH-1:0] wire_d43_67;
	wire [WIDTH-1:0] wire_d43_68;
	wire [WIDTH-1:0] wire_d43_69;
	wire [WIDTH-1:0] wire_d43_70;
	wire [WIDTH-1:0] wire_d43_71;
	wire [WIDTH-1:0] wire_d43_72;
	wire [WIDTH-1:0] wire_d43_73;
	wire [WIDTH-1:0] wire_d43_74;
	wire [WIDTH-1:0] wire_d43_75;
	wire [WIDTH-1:0] wire_d43_76;
	wire [WIDTH-1:0] wire_d43_77;
	wire [WIDTH-1:0] wire_d43_78;
	wire [WIDTH-1:0] wire_d44_0;
	wire [WIDTH-1:0] wire_d44_1;
	wire [WIDTH-1:0] wire_d44_2;
	wire [WIDTH-1:0] wire_d44_3;
	wire [WIDTH-1:0] wire_d44_4;
	wire [WIDTH-1:0] wire_d44_5;
	wire [WIDTH-1:0] wire_d44_6;
	wire [WIDTH-1:0] wire_d44_7;
	wire [WIDTH-1:0] wire_d44_8;
	wire [WIDTH-1:0] wire_d44_9;
	wire [WIDTH-1:0] wire_d44_10;
	wire [WIDTH-1:0] wire_d44_11;
	wire [WIDTH-1:0] wire_d44_12;
	wire [WIDTH-1:0] wire_d44_13;
	wire [WIDTH-1:0] wire_d44_14;
	wire [WIDTH-1:0] wire_d44_15;
	wire [WIDTH-1:0] wire_d44_16;
	wire [WIDTH-1:0] wire_d44_17;
	wire [WIDTH-1:0] wire_d44_18;
	wire [WIDTH-1:0] wire_d44_19;
	wire [WIDTH-1:0] wire_d44_20;
	wire [WIDTH-1:0] wire_d44_21;
	wire [WIDTH-1:0] wire_d44_22;
	wire [WIDTH-1:0] wire_d44_23;
	wire [WIDTH-1:0] wire_d44_24;
	wire [WIDTH-1:0] wire_d44_25;
	wire [WIDTH-1:0] wire_d44_26;
	wire [WIDTH-1:0] wire_d44_27;
	wire [WIDTH-1:0] wire_d44_28;
	wire [WIDTH-1:0] wire_d44_29;
	wire [WIDTH-1:0] wire_d44_30;
	wire [WIDTH-1:0] wire_d44_31;
	wire [WIDTH-1:0] wire_d44_32;
	wire [WIDTH-1:0] wire_d44_33;
	wire [WIDTH-1:0] wire_d44_34;
	wire [WIDTH-1:0] wire_d44_35;
	wire [WIDTH-1:0] wire_d44_36;
	wire [WIDTH-1:0] wire_d44_37;
	wire [WIDTH-1:0] wire_d44_38;
	wire [WIDTH-1:0] wire_d44_39;
	wire [WIDTH-1:0] wire_d44_40;
	wire [WIDTH-1:0] wire_d44_41;
	wire [WIDTH-1:0] wire_d44_42;
	wire [WIDTH-1:0] wire_d44_43;
	wire [WIDTH-1:0] wire_d44_44;
	wire [WIDTH-1:0] wire_d44_45;
	wire [WIDTH-1:0] wire_d44_46;
	wire [WIDTH-1:0] wire_d44_47;
	wire [WIDTH-1:0] wire_d44_48;
	wire [WIDTH-1:0] wire_d44_49;
	wire [WIDTH-1:0] wire_d44_50;
	wire [WIDTH-1:0] wire_d44_51;
	wire [WIDTH-1:0] wire_d44_52;
	wire [WIDTH-1:0] wire_d44_53;
	wire [WIDTH-1:0] wire_d44_54;
	wire [WIDTH-1:0] wire_d44_55;
	wire [WIDTH-1:0] wire_d44_56;
	wire [WIDTH-1:0] wire_d44_57;
	wire [WIDTH-1:0] wire_d44_58;
	wire [WIDTH-1:0] wire_d44_59;
	wire [WIDTH-1:0] wire_d44_60;
	wire [WIDTH-1:0] wire_d44_61;
	wire [WIDTH-1:0] wire_d44_62;
	wire [WIDTH-1:0] wire_d44_63;
	wire [WIDTH-1:0] wire_d44_64;
	wire [WIDTH-1:0] wire_d44_65;
	wire [WIDTH-1:0] wire_d44_66;
	wire [WIDTH-1:0] wire_d44_67;
	wire [WIDTH-1:0] wire_d44_68;
	wire [WIDTH-1:0] wire_d44_69;
	wire [WIDTH-1:0] wire_d44_70;
	wire [WIDTH-1:0] wire_d44_71;
	wire [WIDTH-1:0] wire_d44_72;
	wire [WIDTH-1:0] wire_d44_73;
	wire [WIDTH-1:0] wire_d44_74;
	wire [WIDTH-1:0] wire_d44_75;
	wire [WIDTH-1:0] wire_d44_76;
	wire [WIDTH-1:0] wire_d44_77;
	wire [WIDTH-1:0] wire_d44_78;
	wire [WIDTH-1:0] wire_d45_0;
	wire [WIDTH-1:0] wire_d45_1;
	wire [WIDTH-1:0] wire_d45_2;
	wire [WIDTH-1:0] wire_d45_3;
	wire [WIDTH-1:0] wire_d45_4;
	wire [WIDTH-1:0] wire_d45_5;
	wire [WIDTH-1:0] wire_d45_6;
	wire [WIDTH-1:0] wire_d45_7;
	wire [WIDTH-1:0] wire_d45_8;
	wire [WIDTH-1:0] wire_d45_9;
	wire [WIDTH-1:0] wire_d45_10;
	wire [WIDTH-1:0] wire_d45_11;
	wire [WIDTH-1:0] wire_d45_12;
	wire [WIDTH-1:0] wire_d45_13;
	wire [WIDTH-1:0] wire_d45_14;
	wire [WIDTH-1:0] wire_d45_15;
	wire [WIDTH-1:0] wire_d45_16;
	wire [WIDTH-1:0] wire_d45_17;
	wire [WIDTH-1:0] wire_d45_18;
	wire [WIDTH-1:0] wire_d45_19;
	wire [WIDTH-1:0] wire_d45_20;
	wire [WIDTH-1:0] wire_d45_21;
	wire [WIDTH-1:0] wire_d45_22;
	wire [WIDTH-1:0] wire_d45_23;
	wire [WIDTH-1:0] wire_d45_24;
	wire [WIDTH-1:0] wire_d45_25;
	wire [WIDTH-1:0] wire_d45_26;
	wire [WIDTH-1:0] wire_d45_27;
	wire [WIDTH-1:0] wire_d45_28;
	wire [WIDTH-1:0] wire_d45_29;
	wire [WIDTH-1:0] wire_d45_30;
	wire [WIDTH-1:0] wire_d45_31;
	wire [WIDTH-1:0] wire_d45_32;
	wire [WIDTH-1:0] wire_d45_33;
	wire [WIDTH-1:0] wire_d45_34;
	wire [WIDTH-1:0] wire_d45_35;
	wire [WIDTH-1:0] wire_d45_36;
	wire [WIDTH-1:0] wire_d45_37;
	wire [WIDTH-1:0] wire_d45_38;
	wire [WIDTH-1:0] wire_d45_39;
	wire [WIDTH-1:0] wire_d45_40;
	wire [WIDTH-1:0] wire_d45_41;
	wire [WIDTH-1:0] wire_d45_42;
	wire [WIDTH-1:0] wire_d45_43;
	wire [WIDTH-1:0] wire_d45_44;
	wire [WIDTH-1:0] wire_d45_45;
	wire [WIDTH-1:0] wire_d45_46;
	wire [WIDTH-1:0] wire_d45_47;
	wire [WIDTH-1:0] wire_d45_48;
	wire [WIDTH-1:0] wire_d45_49;
	wire [WIDTH-1:0] wire_d45_50;
	wire [WIDTH-1:0] wire_d45_51;
	wire [WIDTH-1:0] wire_d45_52;
	wire [WIDTH-1:0] wire_d45_53;
	wire [WIDTH-1:0] wire_d45_54;
	wire [WIDTH-1:0] wire_d45_55;
	wire [WIDTH-1:0] wire_d45_56;
	wire [WIDTH-1:0] wire_d45_57;
	wire [WIDTH-1:0] wire_d45_58;
	wire [WIDTH-1:0] wire_d45_59;
	wire [WIDTH-1:0] wire_d45_60;
	wire [WIDTH-1:0] wire_d45_61;
	wire [WIDTH-1:0] wire_d45_62;
	wire [WIDTH-1:0] wire_d45_63;
	wire [WIDTH-1:0] wire_d45_64;
	wire [WIDTH-1:0] wire_d45_65;
	wire [WIDTH-1:0] wire_d45_66;
	wire [WIDTH-1:0] wire_d45_67;
	wire [WIDTH-1:0] wire_d45_68;
	wire [WIDTH-1:0] wire_d45_69;
	wire [WIDTH-1:0] wire_d45_70;
	wire [WIDTH-1:0] wire_d45_71;
	wire [WIDTH-1:0] wire_d45_72;
	wire [WIDTH-1:0] wire_d45_73;
	wire [WIDTH-1:0] wire_d45_74;
	wire [WIDTH-1:0] wire_d45_75;
	wire [WIDTH-1:0] wire_d45_76;
	wire [WIDTH-1:0] wire_d45_77;
	wire [WIDTH-1:0] wire_d45_78;
	wire [WIDTH-1:0] wire_d46_0;
	wire [WIDTH-1:0] wire_d46_1;
	wire [WIDTH-1:0] wire_d46_2;
	wire [WIDTH-1:0] wire_d46_3;
	wire [WIDTH-1:0] wire_d46_4;
	wire [WIDTH-1:0] wire_d46_5;
	wire [WIDTH-1:0] wire_d46_6;
	wire [WIDTH-1:0] wire_d46_7;
	wire [WIDTH-1:0] wire_d46_8;
	wire [WIDTH-1:0] wire_d46_9;
	wire [WIDTH-1:0] wire_d46_10;
	wire [WIDTH-1:0] wire_d46_11;
	wire [WIDTH-1:0] wire_d46_12;
	wire [WIDTH-1:0] wire_d46_13;
	wire [WIDTH-1:0] wire_d46_14;
	wire [WIDTH-1:0] wire_d46_15;
	wire [WIDTH-1:0] wire_d46_16;
	wire [WIDTH-1:0] wire_d46_17;
	wire [WIDTH-1:0] wire_d46_18;
	wire [WIDTH-1:0] wire_d46_19;
	wire [WIDTH-1:0] wire_d46_20;
	wire [WIDTH-1:0] wire_d46_21;
	wire [WIDTH-1:0] wire_d46_22;
	wire [WIDTH-1:0] wire_d46_23;
	wire [WIDTH-1:0] wire_d46_24;
	wire [WIDTH-1:0] wire_d46_25;
	wire [WIDTH-1:0] wire_d46_26;
	wire [WIDTH-1:0] wire_d46_27;
	wire [WIDTH-1:0] wire_d46_28;
	wire [WIDTH-1:0] wire_d46_29;
	wire [WIDTH-1:0] wire_d46_30;
	wire [WIDTH-1:0] wire_d46_31;
	wire [WIDTH-1:0] wire_d46_32;
	wire [WIDTH-1:0] wire_d46_33;
	wire [WIDTH-1:0] wire_d46_34;
	wire [WIDTH-1:0] wire_d46_35;
	wire [WIDTH-1:0] wire_d46_36;
	wire [WIDTH-1:0] wire_d46_37;
	wire [WIDTH-1:0] wire_d46_38;
	wire [WIDTH-1:0] wire_d46_39;
	wire [WIDTH-1:0] wire_d46_40;
	wire [WIDTH-1:0] wire_d46_41;
	wire [WIDTH-1:0] wire_d46_42;
	wire [WIDTH-1:0] wire_d46_43;
	wire [WIDTH-1:0] wire_d46_44;
	wire [WIDTH-1:0] wire_d46_45;
	wire [WIDTH-1:0] wire_d46_46;
	wire [WIDTH-1:0] wire_d46_47;
	wire [WIDTH-1:0] wire_d46_48;
	wire [WIDTH-1:0] wire_d46_49;
	wire [WIDTH-1:0] wire_d46_50;
	wire [WIDTH-1:0] wire_d46_51;
	wire [WIDTH-1:0] wire_d46_52;
	wire [WIDTH-1:0] wire_d46_53;
	wire [WIDTH-1:0] wire_d46_54;
	wire [WIDTH-1:0] wire_d46_55;
	wire [WIDTH-1:0] wire_d46_56;
	wire [WIDTH-1:0] wire_d46_57;
	wire [WIDTH-1:0] wire_d46_58;
	wire [WIDTH-1:0] wire_d46_59;
	wire [WIDTH-1:0] wire_d46_60;
	wire [WIDTH-1:0] wire_d46_61;
	wire [WIDTH-1:0] wire_d46_62;
	wire [WIDTH-1:0] wire_d46_63;
	wire [WIDTH-1:0] wire_d46_64;
	wire [WIDTH-1:0] wire_d46_65;
	wire [WIDTH-1:0] wire_d46_66;
	wire [WIDTH-1:0] wire_d46_67;
	wire [WIDTH-1:0] wire_d46_68;
	wire [WIDTH-1:0] wire_d46_69;
	wire [WIDTH-1:0] wire_d46_70;
	wire [WIDTH-1:0] wire_d46_71;
	wire [WIDTH-1:0] wire_d46_72;
	wire [WIDTH-1:0] wire_d46_73;
	wire [WIDTH-1:0] wire_d46_74;
	wire [WIDTH-1:0] wire_d46_75;
	wire [WIDTH-1:0] wire_d46_76;
	wire [WIDTH-1:0] wire_d46_77;
	wire [WIDTH-1:0] wire_d46_78;
	wire [WIDTH-1:0] wire_d47_0;
	wire [WIDTH-1:0] wire_d47_1;
	wire [WIDTH-1:0] wire_d47_2;
	wire [WIDTH-1:0] wire_d47_3;
	wire [WIDTH-1:0] wire_d47_4;
	wire [WIDTH-1:0] wire_d47_5;
	wire [WIDTH-1:0] wire_d47_6;
	wire [WIDTH-1:0] wire_d47_7;
	wire [WIDTH-1:0] wire_d47_8;
	wire [WIDTH-1:0] wire_d47_9;
	wire [WIDTH-1:0] wire_d47_10;
	wire [WIDTH-1:0] wire_d47_11;
	wire [WIDTH-1:0] wire_d47_12;
	wire [WIDTH-1:0] wire_d47_13;
	wire [WIDTH-1:0] wire_d47_14;
	wire [WIDTH-1:0] wire_d47_15;
	wire [WIDTH-1:0] wire_d47_16;
	wire [WIDTH-1:0] wire_d47_17;
	wire [WIDTH-1:0] wire_d47_18;
	wire [WIDTH-1:0] wire_d47_19;
	wire [WIDTH-1:0] wire_d47_20;
	wire [WIDTH-1:0] wire_d47_21;
	wire [WIDTH-1:0] wire_d47_22;
	wire [WIDTH-1:0] wire_d47_23;
	wire [WIDTH-1:0] wire_d47_24;
	wire [WIDTH-1:0] wire_d47_25;
	wire [WIDTH-1:0] wire_d47_26;
	wire [WIDTH-1:0] wire_d47_27;
	wire [WIDTH-1:0] wire_d47_28;
	wire [WIDTH-1:0] wire_d47_29;
	wire [WIDTH-1:0] wire_d47_30;
	wire [WIDTH-1:0] wire_d47_31;
	wire [WIDTH-1:0] wire_d47_32;
	wire [WIDTH-1:0] wire_d47_33;
	wire [WIDTH-1:0] wire_d47_34;
	wire [WIDTH-1:0] wire_d47_35;
	wire [WIDTH-1:0] wire_d47_36;
	wire [WIDTH-1:0] wire_d47_37;
	wire [WIDTH-1:0] wire_d47_38;
	wire [WIDTH-1:0] wire_d47_39;
	wire [WIDTH-1:0] wire_d47_40;
	wire [WIDTH-1:0] wire_d47_41;
	wire [WIDTH-1:0] wire_d47_42;
	wire [WIDTH-1:0] wire_d47_43;
	wire [WIDTH-1:0] wire_d47_44;
	wire [WIDTH-1:0] wire_d47_45;
	wire [WIDTH-1:0] wire_d47_46;
	wire [WIDTH-1:0] wire_d47_47;
	wire [WIDTH-1:0] wire_d47_48;
	wire [WIDTH-1:0] wire_d47_49;
	wire [WIDTH-1:0] wire_d47_50;
	wire [WIDTH-1:0] wire_d47_51;
	wire [WIDTH-1:0] wire_d47_52;
	wire [WIDTH-1:0] wire_d47_53;
	wire [WIDTH-1:0] wire_d47_54;
	wire [WIDTH-1:0] wire_d47_55;
	wire [WIDTH-1:0] wire_d47_56;
	wire [WIDTH-1:0] wire_d47_57;
	wire [WIDTH-1:0] wire_d47_58;
	wire [WIDTH-1:0] wire_d47_59;
	wire [WIDTH-1:0] wire_d47_60;
	wire [WIDTH-1:0] wire_d47_61;
	wire [WIDTH-1:0] wire_d47_62;
	wire [WIDTH-1:0] wire_d47_63;
	wire [WIDTH-1:0] wire_d47_64;
	wire [WIDTH-1:0] wire_d47_65;
	wire [WIDTH-1:0] wire_d47_66;
	wire [WIDTH-1:0] wire_d47_67;
	wire [WIDTH-1:0] wire_d47_68;
	wire [WIDTH-1:0] wire_d47_69;
	wire [WIDTH-1:0] wire_d47_70;
	wire [WIDTH-1:0] wire_d47_71;
	wire [WIDTH-1:0] wire_d47_72;
	wire [WIDTH-1:0] wire_d47_73;
	wire [WIDTH-1:0] wire_d47_74;
	wire [WIDTH-1:0] wire_d47_75;
	wire [WIDTH-1:0] wire_d47_76;
	wire [WIDTH-1:0] wire_d47_77;
	wire [WIDTH-1:0] wire_d47_78;
	wire [WIDTH-1:0] wire_d48_0;
	wire [WIDTH-1:0] wire_d48_1;
	wire [WIDTH-1:0] wire_d48_2;
	wire [WIDTH-1:0] wire_d48_3;
	wire [WIDTH-1:0] wire_d48_4;
	wire [WIDTH-1:0] wire_d48_5;
	wire [WIDTH-1:0] wire_d48_6;
	wire [WIDTH-1:0] wire_d48_7;
	wire [WIDTH-1:0] wire_d48_8;
	wire [WIDTH-1:0] wire_d48_9;
	wire [WIDTH-1:0] wire_d48_10;
	wire [WIDTH-1:0] wire_d48_11;
	wire [WIDTH-1:0] wire_d48_12;
	wire [WIDTH-1:0] wire_d48_13;
	wire [WIDTH-1:0] wire_d48_14;
	wire [WIDTH-1:0] wire_d48_15;
	wire [WIDTH-1:0] wire_d48_16;
	wire [WIDTH-1:0] wire_d48_17;
	wire [WIDTH-1:0] wire_d48_18;
	wire [WIDTH-1:0] wire_d48_19;
	wire [WIDTH-1:0] wire_d48_20;
	wire [WIDTH-1:0] wire_d48_21;
	wire [WIDTH-1:0] wire_d48_22;
	wire [WIDTH-1:0] wire_d48_23;
	wire [WIDTH-1:0] wire_d48_24;
	wire [WIDTH-1:0] wire_d48_25;
	wire [WIDTH-1:0] wire_d48_26;
	wire [WIDTH-1:0] wire_d48_27;
	wire [WIDTH-1:0] wire_d48_28;
	wire [WIDTH-1:0] wire_d48_29;
	wire [WIDTH-1:0] wire_d48_30;
	wire [WIDTH-1:0] wire_d48_31;
	wire [WIDTH-1:0] wire_d48_32;
	wire [WIDTH-1:0] wire_d48_33;
	wire [WIDTH-1:0] wire_d48_34;
	wire [WIDTH-1:0] wire_d48_35;
	wire [WIDTH-1:0] wire_d48_36;
	wire [WIDTH-1:0] wire_d48_37;
	wire [WIDTH-1:0] wire_d48_38;
	wire [WIDTH-1:0] wire_d48_39;
	wire [WIDTH-1:0] wire_d48_40;
	wire [WIDTH-1:0] wire_d48_41;
	wire [WIDTH-1:0] wire_d48_42;
	wire [WIDTH-1:0] wire_d48_43;
	wire [WIDTH-1:0] wire_d48_44;
	wire [WIDTH-1:0] wire_d48_45;
	wire [WIDTH-1:0] wire_d48_46;
	wire [WIDTH-1:0] wire_d48_47;
	wire [WIDTH-1:0] wire_d48_48;
	wire [WIDTH-1:0] wire_d48_49;
	wire [WIDTH-1:0] wire_d48_50;
	wire [WIDTH-1:0] wire_d48_51;
	wire [WIDTH-1:0] wire_d48_52;
	wire [WIDTH-1:0] wire_d48_53;
	wire [WIDTH-1:0] wire_d48_54;
	wire [WIDTH-1:0] wire_d48_55;
	wire [WIDTH-1:0] wire_d48_56;
	wire [WIDTH-1:0] wire_d48_57;
	wire [WIDTH-1:0] wire_d48_58;
	wire [WIDTH-1:0] wire_d48_59;
	wire [WIDTH-1:0] wire_d48_60;
	wire [WIDTH-1:0] wire_d48_61;
	wire [WIDTH-1:0] wire_d48_62;
	wire [WIDTH-1:0] wire_d48_63;
	wire [WIDTH-1:0] wire_d48_64;
	wire [WIDTH-1:0] wire_d48_65;
	wire [WIDTH-1:0] wire_d48_66;
	wire [WIDTH-1:0] wire_d48_67;
	wire [WIDTH-1:0] wire_d48_68;
	wire [WIDTH-1:0] wire_d48_69;
	wire [WIDTH-1:0] wire_d48_70;
	wire [WIDTH-1:0] wire_d48_71;
	wire [WIDTH-1:0] wire_d48_72;
	wire [WIDTH-1:0] wire_d48_73;
	wire [WIDTH-1:0] wire_d48_74;
	wire [WIDTH-1:0] wire_d48_75;
	wire [WIDTH-1:0] wire_d48_76;
	wire [WIDTH-1:0] wire_d48_77;
	wire [WIDTH-1:0] wire_d48_78;
	wire [WIDTH-1:0] wire_d49_0;
	wire [WIDTH-1:0] wire_d49_1;
	wire [WIDTH-1:0] wire_d49_2;
	wire [WIDTH-1:0] wire_d49_3;
	wire [WIDTH-1:0] wire_d49_4;
	wire [WIDTH-1:0] wire_d49_5;
	wire [WIDTH-1:0] wire_d49_6;
	wire [WIDTH-1:0] wire_d49_7;
	wire [WIDTH-1:0] wire_d49_8;
	wire [WIDTH-1:0] wire_d49_9;
	wire [WIDTH-1:0] wire_d49_10;
	wire [WIDTH-1:0] wire_d49_11;
	wire [WIDTH-1:0] wire_d49_12;
	wire [WIDTH-1:0] wire_d49_13;
	wire [WIDTH-1:0] wire_d49_14;
	wire [WIDTH-1:0] wire_d49_15;
	wire [WIDTH-1:0] wire_d49_16;
	wire [WIDTH-1:0] wire_d49_17;
	wire [WIDTH-1:0] wire_d49_18;
	wire [WIDTH-1:0] wire_d49_19;
	wire [WIDTH-1:0] wire_d49_20;
	wire [WIDTH-1:0] wire_d49_21;
	wire [WIDTH-1:0] wire_d49_22;
	wire [WIDTH-1:0] wire_d49_23;
	wire [WIDTH-1:0] wire_d49_24;
	wire [WIDTH-1:0] wire_d49_25;
	wire [WIDTH-1:0] wire_d49_26;
	wire [WIDTH-1:0] wire_d49_27;
	wire [WIDTH-1:0] wire_d49_28;
	wire [WIDTH-1:0] wire_d49_29;
	wire [WIDTH-1:0] wire_d49_30;
	wire [WIDTH-1:0] wire_d49_31;
	wire [WIDTH-1:0] wire_d49_32;
	wire [WIDTH-1:0] wire_d49_33;
	wire [WIDTH-1:0] wire_d49_34;
	wire [WIDTH-1:0] wire_d49_35;
	wire [WIDTH-1:0] wire_d49_36;
	wire [WIDTH-1:0] wire_d49_37;
	wire [WIDTH-1:0] wire_d49_38;
	wire [WIDTH-1:0] wire_d49_39;
	wire [WIDTH-1:0] wire_d49_40;
	wire [WIDTH-1:0] wire_d49_41;
	wire [WIDTH-1:0] wire_d49_42;
	wire [WIDTH-1:0] wire_d49_43;
	wire [WIDTH-1:0] wire_d49_44;
	wire [WIDTH-1:0] wire_d49_45;
	wire [WIDTH-1:0] wire_d49_46;
	wire [WIDTH-1:0] wire_d49_47;
	wire [WIDTH-1:0] wire_d49_48;
	wire [WIDTH-1:0] wire_d49_49;
	wire [WIDTH-1:0] wire_d49_50;
	wire [WIDTH-1:0] wire_d49_51;
	wire [WIDTH-1:0] wire_d49_52;
	wire [WIDTH-1:0] wire_d49_53;
	wire [WIDTH-1:0] wire_d49_54;
	wire [WIDTH-1:0] wire_d49_55;
	wire [WIDTH-1:0] wire_d49_56;
	wire [WIDTH-1:0] wire_d49_57;
	wire [WIDTH-1:0] wire_d49_58;
	wire [WIDTH-1:0] wire_d49_59;
	wire [WIDTH-1:0] wire_d49_60;
	wire [WIDTH-1:0] wire_d49_61;
	wire [WIDTH-1:0] wire_d49_62;
	wire [WIDTH-1:0] wire_d49_63;
	wire [WIDTH-1:0] wire_d49_64;
	wire [WIDTH-1:0] wire_d49_65;
	wire [WIDTH-1:0] wire_d49_66;
	wire [WIDTH-1:0] wire_d49_67;
	wire [WIDTH-1:0] wire_d49_68;
	wire [WIDTH-1:0] wire_d49_69;
	wire [WIDTH-1:0] wire_d49_70;
	wire [WIDTH-1:0] wire_d49_71;
	wire [WIDTH-1:0] wire_d49_72;
	wire [WIDTH-1:0] wire_d49_73;
	wire [WIDTH-1:0] wire_d49_74;
	wire [WIDTH-1:0] wire_d49_75;
	wire [WIDTH-1:0] wire_d49_76;
	wire [WIDTH-1:0] wire_d49_77;
	wire [WIDTH-1:0] wire_d49_78;
	wire [WIDTH-1:0] wire_d50_0;
	wire [WIDTH-1:0] wire_d50_1;
	wire [WIDTH-1:0] wire_d50_2;
	wire [WIDTH-1:0] wire_d50_3;
	wire [WIDTH-1:0] wire_d50_4;
	wire [WIDTH-1:0] wire_d50_5;
	wire [WIDTH-1:0] wire_d50_6;
	wire [WIDTH-1:0] wire_d50_7;
	wire [WIDTH-1:0] wire_d50_8;
	wire [WIDTH-1:0] wire_d50_9;
	wire [WIDTH-1:0] wire_d50_10;
	wire [WIDTH-1:0] wire_d50_11;
	wire [WIDTH-1:0] wire_d50_12;
	wire [WIDTH-1:0] wire_d50_13;
	wire [WIDTH-1:0] wire_d50_14;
	wire [WIDTH-1:0] wire_d50_15;
	wire [WIDTH-1:0] wire_d50_16;
	wire [WIDTH-1:0] wire_d50_17;
	wire [WIDTH-1:0] wire_d50_18;
	wire [WIDTH-1:0] wire_d50_19;
	wire [WIDTH-1:0] wire_d50_20;
	wire [WIDTH-1:0] wire_d50_21;
	wire [WIDTH-1:0] wire_d50_22;
	wire [WIDTH-1:0] wire_d50_23;
	wire [WIDTH-1:0] wire_d50_24;
	wire [WIDTH-1:0] wire_d50_25;
	wire [WIDTH-1:0] wire_d50_26;
	wire [WIDTH-1:0] wire_d50_27;
	wire [WIDTH-1:0] wire_d50_28;
	wire [WIDTH-1:0] wire_d50_29;
	wire [WIDTH-1:0] wire_d50_30;
	wire [WIDTH-1:0] wire_d50_31;
	wire [WIDTH-1:0] wire_d50_32;
	wire [WIDTH-1:0] wire_d50_33;
	wire [WIDTH-1:0] wire_d50_34;
	wire [WIDTH-1:0] wire_d50_35;
	wire [WIDTH-1:0] wire_d50_36;
	wire [WIDTH-1:0] wire_d50_37;
	wire [WIDTH-1:0] wire_d50_38;
	wire [WIDTH-1:0] wire_d50_39;
	wire [WIDTH-1:0] wire_d50_40;
	wire [WIDTH-1:0] wire_d50_41;
	wire [WIDTH-1:0] wire_d50_42;
	wire [WIDTH-1:0] wire_d50_43;
	wire [WIDTH-1:0] wire_d50_44;
	wire [WIDTH-1:0] wire_d50_45;
	wire [WIDTH-1:0] wire_d50_46;
	wire [WIDTH-1:0] wire_d50_47;
	wire [WIDTH-1:0] wire_d50_48;
	wire [WIDTH-1:0] wire_d50_49;
	wire [WIDTH-1:0] wire_d50_50;
	wire [WIDTH-1:0] wire_d50_51;
	wire [WIDTH-1:0] wire_d50_52;
	wire [WIDTH-1:0] wire_d50_53;
	wire [WIDTH-1:0] wire_d50_54;
	wire [WIDTH-1:0] wire_d50_55;
	wire [WIDTH-1:0] wire_d50_56;
	wire [WIDTH-1:0] wire_d50_57;
	wire [WIDTH-1:0] wire_d50_58;
	wire [WIDTH-1:0] wire_d50_59;
	wire [WIDTH-1:0] wire_d50_60;
	wire [WIDTH-1:0] wire_d50_61;
	wire [WIDTH-1:0] wire_d50_62;
	wire [WIDTH-1:0] wire_d50_63;
	wire [WIDTH-1:0] wire_d50_64;
	wire [WIDTH-1:0] wire_d50_65;
	wire [WIDTH-1:0] wire_d50_66;
	wire [WIDTH-1:0] wire_d50_67;
	wire [WIDTH-1:0] wire_d50_68;
	wire [WIDTH-1:0] wire_d50_69;
	wire [WIDTH-1:0] wire_d50_70;
	wire [WIDTH-1:0] wire_d50_71;
	wire [WIDTH-1:0] wire_d50_72;
	wire [WIDTH-1:0] wire_d50_73;
	wire [WIDTH-1:0] wire_d50_74;
	wire [WIDTH-1:0] wire_d50_75;
	wire [WIDTH-1:0] wire_d50_76;
	wire [WIDTH-1:0] wire_d50_77;
	wire [WIDTH-1:0] wire_d50_78;
	wire [WIDTH-1:0] wire_d51_0;
	wire [WIDTH-1:0] wire_d51_1;
	wire [WIDTH-1:0] wire_d51_2;
	wire [WIDTH-1:0] wire_d51_3;
	wire [WIDTH-1:0] wire_d51_4;
	wire [WIDTH-1:0] wire_d51_5;
	wire [WIDTH-1:0] wire_d51_6;
	wire [WIDTH-1:0] wire_d51_7;
	wire [WIDTH-1:0] wire_d51_8;
	wire [WIDTH-1:0] wire_d51_9;
	wire [WIDTH-1:0] wire_d51_10;
	wire [WIDTH-1:0] wire_d51_11;
	wire [WIDTH-1:0] wire_d51_12;
	wire [WIDTH-1:0] wire_d51_13;
	wire [WIDTH-1:0] wire_d51_14;
	wire [WIDTH-1:0] wire_d51_15;
	wire [WIDTH-1:0] wire_d51_16;
	wire [WIDTH-1:0] wire_d51_17;
	wire [WIDTH-1:0] wire_d51_18;
	wire [WIDTH-1:0] wire_d51_19;
	wire [WIDTH-1:0] wire_d51_20;
	wire [WIDTH-1:0] wire_d51_21;
	wire [WIDTH-1:0] wire_d51_22;
	wire [WIDTH-1:0] wire_d51_23;
	wire [WIDTH-1:0] wire_d51_24;
	wire [WIDTH-1:0] wire_d51_25;
	wire [WIDTH-1:0] wire_d51_26;
	wire [WIDTH-1:0] wire_d51_27;
	wire [WIDTH-1:0] wire_d51_28;
	wire [WIDTH-1:0] wire_d51_29;
	wire [WIDTH-1:0] wire_d51_30;
	wire [WIDTH-1:0] wire_d51_31;
	wire [WIDTH-1:0] wire_d51_32;
	wire [WIDTH-1:0] wire_d51_33;
	wire [WIDTH-1:0] wire_d51_34;
	wire [WIDTH-1:0] wire_d51_35;
	wire [WIDTH-1:0] wire_d51_36;
	wire [WIDTH-1:0] wire_d51_37;
	wire [WIDTH-1:0] wire_d51_38;
	wire [WIDTH-1:0] wire_d51_39;
	wire [WIDTH-1:0] wire_d51_40;
	wire [WIDTH-1:0] wire_d51_41;
	wire [WIDTH-1:0] wire_d51_42;
	wire [WIDTH-1:0] wire_d51_43;
	wire [WIDTH-1:0] wire_d51_44;
	wire [WIDTH-1:0] wire_d51_45;
	wire [WIDTH-1:0] wire_d51_46;
	wire [WIDTH-1:0] wire_d51_47;
	wire [WIDTH-1:0] wire_d51_48;
	wire [WIDTH-1:0] wire_d51_49;
	wire [WIDTH-1:0] wire_d51_50;
	wire [WIDTH-1:0] wire_d51_51;
	wire [WIDTH-1:0] wire_d51_52;
	wire [WIDTH-1:0] wire_d51_53;
	wire [WIDTH-1:0] wire_d51_54;
	wire [WIDTH-1:0] wire_d51_55;
	wire [WIDTH-1:0] wire_d51_56;
	wire [WIDTH-1:0] wire_d51_57;
	wire [WIDTH-1:0] wire_d51_58;
	wire [WIDTH-1:0] wire_d51_59;
	wire [WIDTH-1:0] wire_d51_60;
	wire [WIDTH-1:0] wire_d51_61;
	wire [WIDTH-1:0] wire_d51_62;
	wire [WIDTH-1:0] wire_d51_63;
	wire [WIDTH-1:0] wire_d51_64;
	wire [WIDTH-1:0] wire_d51_65;
	wire [WIDTH-1:0] wire_d51_66;
	wire [WIDTH-1:0] wire_d51_67;
	wire [WIDTH-1:0] wire_d51_68;
	wire [WIDTH-1:0] wire_d51_69;
	wire [WIDTH-1:0] wire_d51_70;
	wire [WIDTH-1:0] wire_d51_71;
	wire [WIDTH-1:0] wire_d51_72;
	wire [WIDTH-1:0] wire_d51_73;
	wire [WIDTH-1:0] wire_d51_74;
	wire [WIDTH-1:0] wire_d51_75;
	wire [WIDTH-1:0] wire_d51_76;
	wire [WIDTH-1:0] wire_d51_77;
	wire [WIDTH-1:0] wire_d51_78;
	wire [WIDTH-1:0] wire_d52_0;
	wire [WIDTH-1:0] wire_d52_1;
	wire [WIDTH-1:0] wire_d52_2;
	wire [WIDTH-1:0] wire_d52_3;
	wire [WIDTH-1:0] wire_d52_4;
	wire [WIDTH-1:0] wire_d52_5;
	wire [WIDTH-1:0] wire_d52_6;
	wire [WIDTH-1:0] wire_d52_7;
	wire [WIDTH-1:0] wire_d52_8;
	wire [WIDTH-1:0] wire_d52_9;
	wire [WIDTH-1:0] wire_d52_10;
	wire [WIDTH-1:0] wire_d52_11;
	wire [WIDTH-1:0] wire_d52_12;
	wire [WIDTH-1:0] wire_d52_13;
	wire [WIDTH-1:0] wire_d52_14;
	wire [WIDTH-1:0] wire_d52_15;
	wire [WIDTH-1:0] wire_d52_16;
	wire [WIDTH-1:0] wire_d52_17;
	wire [WIDTH-1:0] wire_d52_18;
	wire [WIDTH-1:0] wire_d52_19;
	wire [WIDTH-1:0] wire_d52_20;
	wire [WIDTH-1:0] wire_d52_21;
	wire [WIDTH-1:0] wire_d52_22;
	wire [WIDTH-1:0] wire_d52_23;
	wire [WIDTH-1:0] wire_d52_24;
	wire [WIDTH-1:0] wire_d52_25;
	wire [WIDTH-1:0] wire_d52_26;
	wire [WIDTH-1:0] wire_d52_27;
	wire [WIDTH-1:0] wire_d52_28;
	wire [WIDTH-1:0] wire_d52_29;
	wire [WIDTH-1:0] wire_d52_30;
	wire [WIDTH-1:0] wire_d52_31;
	wire [WIDTH-1:0] wire_d52_32;
	wire [WIDTH-1:0] wire_d52_33;
	wire [WIDTH-1:0] wire_d52_34;
	wire [WIDTH-1:0] wire_d52_35;
	wire [WIDTH-1:0] wire_d52_36;
	wire [WIDTH-1:0] wire_d52_37;
	wire [WIDTH-1:0] wire_d52_38;
	wire [WIDTH-1:0] wire_d52_39;
	wire [WIDTH-1:0] wire_d52_40;
	wire [WIDTH-1:0] wire_d52_41;
	wire [WIDTH-1:0] wire_d52_42;
	wire [WIDTH-1:0] wire_d52_43;
	wire [WIDTH-1:0] wire_d52_44;
	wire [WIDTH-1:0] wire_d52_45;
	wire [WIDTH-1:0] wire_d52_46;
	wire [WIDTH-1:0] wire_d52_47;
	wire [WIDTH-1:0] wire_d52_48;
	wire [WIDTH-1:0] wire_d52_49;
	wire [WIDTH-1:0] wire_d52_50;
	wire [WIDTH-1:0] wire_d52_51;
	wire [WIDTH-1:0] wire_d52_52;
	wire [WIDTH-1:0] wire_d52_53;
	wire [WIDTH-1:0] wire_d52_54;
	wire [WIDTH-1:0] wire_d52_55;
	wire [WIDTH-1:0] wire_d52_56;
	wire [WIDTH-1:0] wire_d52_57;
	wire [WIDTH-1:0] wire_d52_58;
	wire [WIDTH-1:0] wire_d52_59;
	wire [WIDTH-1:0] wire_d52_60;
	wire [WIDTH-1:0] wire_d52_61;
	wire [WIDTH-1:0] wire_d52_62;
	wire [WIDTH-1:0] wire_d52_63;
	wire [WIDTH-1:0] wire_d52_64;
	wire [WIDTH-1:0] wire_d52_65;
	wire [WIDTH-1:0] wire_d52_66;
	wire [WIDTH-1:0] wire_d52_67;
	wire [WIDTH-1:0] wire_d52_68;
	wire [WIDTH-1:0] wire_d52_69;
	wire [WIDTH-1:0] wire_d52_70;
	wire [WIDTH-1:0] wire_d52_71;
	wire [WIDTH-1:0] wire_d52_72;
	wire [WIDTH-1:0] wire_d52_73;
	wire [WIDTH-1:0] wire_d52_74;
	wire [WIDTH-1:0] wire_d52_75;
	wire [WIDTH-1:0] wire_d52_76;
	wire [WIDTH-1:0] wire_d52_77;
	wire [WIDTH-1:0] wire_d52_78;
	wire [WIDTH-1:0] wire_d53_0;
	wire [WIDTH-1:0] wire_d53_1;
	wire [WIDTH-1:0] wire_d53_2;
	wire [WIDTH-1:0] wire_d53_3;
	wire [WIDTH-1:0] wire_d53_4;
	wire [WIDTH-1:0] wire_d53_5;
	wire [WIDTH-1:0] wire_d53_6;
	wire [WIDTH-1:0] wire_d53_7;
	wire [WIDTH-1:0] wire_d53_8;
	wire [WIDTH-1:0] wire_d53_9;
	wire [WIDTH-1:0] wire_d53_10;
	wire [WIDTH-1:0] wire_d53_11;
	wire [WIDTH-1:0] wire_d53_12;
	wire [WIDTH-1:0] wire_d53_13;
	wire [WIDTH-1:0] wire_d53_14;
	wire [WIDTH-1:0] wire_d53_15;
	wire [WIDTH-1:0] wire_d53_16;
	wire [WIDTH-1:0] wire_d53_17;
	wire [WIDTH-1:0] wire_d53_18;
	wire [WIDTH-1:0] wire_d53_19;
	wire [WIDTH-1:0] wire_d53_20;
	wire [WIDTH-1:0] wire_d53_21;
	wire [WIDTH-1:0] wire_d53_22;
	wire [WIDTH-1:0] wire_d53_23;
	wire [WIDTH-1:0] wire_d53_24;
	wire [WIDTH-1:0] wire_d53_25;
	wire [WIDTH-1:0] wire_d53_26;
	wire [WIDTH-1:0] wire_d53_27;
	wire [WIDTH-1:0] wire_d53_28;
	wire [WIDTH-1:0] wire_d53_29;
	wire [WIDTH-1:0] wire_d53_30;
	wire [WIDTH-1:0] wire_d53_31;
	wire [WIDTH-1:0] wire_d53_32;
	wire [WIDTH-1:0] wire_d53_33;
	wire [WIDTH-1:0] wire_d53_34;
	wire [WIDTH-1:0] wire_d53_35;
	wire [WIDTH-1:0] wire_d53_36;
	wire [WIDTH-1:0] wire_d53_37;
	wire [WIDTH-1:0] wire_d53_38;
	wire [WIDTH-1:0] wire_d53_39;
	wire [WIDTH-1:0] wire_d53_40;
	wire [WIDTH-1:0] wire_d53_41;
	wire [WIDTH-1:0] wire_d53_42;
	wire [WIDTH-1:0] wire_d53_43;
	wire [WIDTH-1:0] wire_d53_44;
	wire [WIDTH-1:0] wire_d53_45;
	wire [WIDTH-1:0] wire_d53_46;
	wire [WIDTH-1:0] wire_d53_47;
	wire [WIDTH-1:0] wire_d53_48;
	wire [WIDTH-1:0] wire_d53_49;
	wire [WIDTH-1:0] wire_d53_50;
	wire [WIDTH-1:0] wire_d53_51;
	wire [WIDTH-1:0] wire_d53_52;
	wire [WIDTH-1:0] wire_d53_53;
	wire [WIDTH-1:0] wire_d53_54;
	wire [WIDTH-1:0] wire_d53_55;
	wire [WIDTH-1:0] wire_d53_56;
	wire [WIDTH-1:0] wire_d53_57;
	wire [WIDTH-1:0] wire_d53_58;
	wire [WIDTH-1:0] wire_d53_59;
	wire [WIDTH-1:0] wire_d53_60;
	wire [WIDTH-1:0] wire_d53_61;
	wire [WIDTH-1:0] wire_d53_62;
	wire [WIDTH-1:0] wire_d53_63;
	wire [WIDTH-1:0] wire_d53_64;
	wire [WIDTH-1:0] wire_d53_65;
	wire [WIDTH-1:0] wire_d53_66;
	wire [WIDTH-1:0] wire_d53_67;
	wire [WIDTH-1:0] wire_d53_68;
	wire [WIDTH-1:0] wire_d53_69;
	wire [WIDTH-1:0] wire_d53_70;
	wire [WIDTH-1:0] wire_d53_71;
	wire [WIDTH-1:0] wire_d53_72;
	wire [WIDTH-1:0] wire_d53_73;
	wire [WIDTH-1:0] wire_d53_74;
	wire [WIDTH-1:0] wire_d53_75;
	wire [WIDTH-1:0] wire_d53_76;
	wire [WIDTH-1:0] wire_d53_77;
	wire [WIDTH-1:0] wire_d53_78;
	wire [WIDTH-1:0] wire_d54_0;
	wire [WIDTH-1:0] wire_d54_1;
	wire [WIDTH-1:0] wire_d54_2;
	wire [WIDTH-1:0] wire_d54_3;
	wire [WIDTH-1:0] wire_d54_4;
	wire [WIDTH-1:0] wire_d54_5;
	wire [WIDTH-1:0] wire_d54_6;
	wire [WIDTH-1:0] wire_d54_7;
	wire [WIDTH-1:0] wire_d54_8;
	wire [WIDTH-1:0] wire_d54_9;
	wire [WIDTH-1:0] wire_d54_10;
	wire [WIDTH-1:0] wire_d54_11;
	wire [WIDTH-1:0] wire_d54_12;
	wire [WIDTH-1:0] wire_d54_13;
	wire [WIDTH-1:0] wire_d54_14;
	wire [WIDTH-1:0] wire_d54_15;
	wire [WIDTH-1:0] wire_d54_16;
	wire [WIDTH-1:0] wire_d54_17;
	wire [WIDTH-1:0] wire_d54_18;
	wire [WIDTH-1:0] wire_d54_19;
	wire [WIDTH-1:0] wire_d54_20;
	wire [WIDTH-1:0] wire_d54_21;
	wire [WIDTH-1:0] wire_d54_22;
	wire [WIDTH-1:0] wire_d54_23;
	wire [WIDTH-1:0] wire_d54_24;
	wire [WIDTH-1:0] wire_d54_25;
	wire [WIDTH-1:0] wire_d54_26;
	wire [WIDTH-1:0] wire_d54_27;
	wire [WIDTH-1:0] wire_d54_28;
	wire [WIDTH-1:0] wire_d54_29;
	wire [WIDTH-1:0] wire_d54_30;
	wire [WIDTH-1:0] wire_d54_31;
	wire [WIDTH-1:0] wire_d54_32;
	wire [WIDTH-1:0] wire_d54_33;
	wire [WIDTH-1:0] wire_d54_34;
	wire [WIDTH-1:0] wire_d54_35;
	wire [WIDTH-1:0] wire_d54_36;
	wire [WIDTH-1:0] wire_d54_37;
	wire [WIDTH-1:0] wire_d54_38;
	wire [WIDTH-1:0] wire_d54_39;
	wire [WIDTH-1:0] wire_d54_40;
	wire [WIDTH-1:0] wire_d54_41;
	wire [WIDTH-1:0] wire_d54_42;
	wire [WIDTH-1:0] wire_d54_43;
	wire [WIDTH-1:0] wire_d54_44;
	wire [WIDTH-1:0] wire_d54_45;
	wire [WIDTH-1:0] wire_d54_46;
	wire [WIDTH-1:0] wire_d54_47;
	wire [WIDTH-1:0] wire_d54_48;
	wire [WIDTH-1:0] wire_d54_49;
	wire [WIDTH-1:0] wire_d54_50;
	wire [WIDTH-1:0] wire_d54_51;
	wire [WIDTH-1:0] wire_d54_52;
	wire [WIDTH-1:0] wire_d54_53;
	wire [WIDTH-1:0] wire_d54_54;
	wire [WIDTH-1:0] wire_d54_55;
	wire [WIDTH-1:0] wire_d54_56;
	wire [WIDTH-1:0] wire_d54_57;
	wire [WIDTH-1:0] wire_d54_58;
	wire [WIDTH-1:0] wire_d54_59;
	wire [WIDTH-1:0] wire_d54_60;
	wire [WIDTH-1:0] wire_d54_61;
	wire [WIDTH-1:0] wire_d54_62;
	wire [WIDTH-1:0] wire_d54_63;
	wire [WIDTH-1:0] wire_d54_64;
	wire [WIDTH-1:0] wire_d54_65;
	wire [WIDTH-1:0] wire_d54_66;
	wire [WIDTH-1:0] wire_d54_67;
	wire [WIDTH-1:0] wire_d54_68;
	wire [WIDTH-1:0] wire_d54_69;
	wire [WIDTH-1:0] wire_d54_70;
	wire [WIDTH-1:0] wire_d54_71;
	wire [WIDTH-1:0] wire_d54_72;
	wire [WIDTH-1:0] wire_d54_73;
	wire [WIDTH-1:0] wire_d54_74;
	wire [WIDTH-1:0] wire_d54_75;
	wire [WIDTH-1:0] wire_d54_76;
	wire [WIDTH-1:0] wire_d54_77;
	wire [WIDTH-1:0] wire_d54_78;
	wire [WIDTH-1:0] wire_d55_0;
	wire [WIDTH-1:0] wire_d55_1;
	wire [WIDTH-1:0] wire_d55_2;
	wire [WIDTH-1:0] wire_d55_3;
	wire [WIDTH-1:0] wire_d55_4;
	wire [WIDTH-1:0] wire_d55_5;
	wire [WIDTH-1:0] wire_d55_6;
	wire [WIDTH-1:0] wire_d55_7;
	wire [WIDTH-1:0] wire_d55_8;
	wire [WIDTH-1:0] wire_d55_9;
	wire [WIDTH-1:0] wire_d55_10;
	wire [WIDTH-1:0] wire_d55_11;
	wire [WIDTH-1:0] wire_d55_12;
	wire [WIDTH-1:0] wire_d55_13;
	wire [WIDTH-1:0] wire_d55_14;
	wire [WIDTH-1:0] wire_d55_15;
	wire [WIDTH-1:0] wire_d55_16;
	wire [WIDTH-1:0] wire_d55_17;
	wire [WIDTH-1:0] wire_d55_18;
	wire [WIDTH-1:0] wire_d55_19;
	wire [WIDTH-1:0] wire_d55_20;
	wire [WIDTH-1:0] wire_d55_21;
	wire [WIDTH-1:0] wire_d55_22;
	wire [WIDTH-1:0] wire_d55_23;
	wire [WIDTH-1:0] wire_d55_24;
	wire [WIDTH-1:0] wire_d55_25;
	wire [WIDTH-1:0] wire_d55_26;
	wire [WIDTH-1:0] wire_d55_27;
	wire [WIDTH-1:0] wire_d55_28;
	wire [WIDTH-1:0] wire_d55_29;
	wire [WIDTH-1:0] wire_d55_30;
	wire [WIDTH-1:0] wire_d55_31;
	wire [WIDTH-1:0] wire_d55_32;
	wire [WIDTH-1:0] wire_d55_33;
	wire [WIDTH-1:0] wire_d55_34;
	wire [WIDTH-1:0] wire_d55_35;
	wire [WIDTH-1:0] wire_d55_36;
	wire [WIDTH-1:0] wire_d55_37;
	wire [WIDTH-1:0] wire_d55_38;
	wire [WIDTH-1:0] wire_d55_39;
	wire [WIDTH-1:0] wire_d55_40;
	wire [WIDTH-1:0] wire_d55_41;
	wire [WIDTH-1:0] wire_d55_42;
	wire [WIDTH-1:0] wire_d55_43;
	wire [WIDTH-1:0] wire_d55_44;
	wire [WIDTH-1:0] wire_d55_45;
	wire [WIDTH-1:0] wire_d55_46;
	wire [WIDTH-1:0] wire_d55_47;
	wire [WIDTH-1:0] wire_d55_48;
	wire [WIDTH-1:0] wire_d55_49;
	wire [WIDTH-1:0] wire_d55_50;
	wire [WIDTH-1:0] wire_d55_51;
	wire [WIDTH-1:0] wire_d55_52;
	wire [WIDTH-1:0] wire_d55_53;
	wire [WIDTH-1:0] wire_d55_54;
	wire [WIDTH-1:0] wire_d55_55;
	wire [WIDTH-1:0] wire_d55_56;
	wire [WIDTH-1:0] wire_d55_57;
	wire [WIDTH-1:0] wire_d55_58;
	wire [WIDTH-1:0] wire_d55_59;
	wire [WIDTH-1:0] wire_d55_60;
	wire [WIDTH-1:0] wire_d55_61;
	wire [WIDTH-1:0] wire_d55_62;
	wire [WIDTH-1:0] wire_d55_63;
	wire [WIDTH-1:0] wire_d55_64;
	wire [WIDTH-1:0] wire_d55_65;
	wire [WIDTH-1:0] wire_d55_66;
	wire [WIDTH-1:0] wire_d55_67;
	wire [WIDTH-1:0] wire_d55_68;
	wire [WIDTH-1:0] wire_d55_69;
	wire [WIDTH-1:0] wire_d55_70;
	wire [WIDTH-1:0] wire_d55_71;
	wire [WIDTH-1:0] wire_d55_72;
	wire [WIDTH-1:0] wire_d55_73;
	wire [WIDTH-1:0] wire_d55_74;
	wire [WIDTH-1:0] wire_d55_75;
	wire [WIDTH-1:0] wire_d55_76;
	wire [WIDTH-1:0] wire_d55_77;
	wire [WIDTH-1:0] wire_d55_78;
	wire [WIDTH-1:0] wire_d56_0;
	wire [WIDTH-1:0] wire_d56_1;
	wire [WIDTH-1:0] wire_d56_2;
	wire [WIDTH-1:0] wire_d56_3;
	wire [WIDTH-1:0] wire_d56_4;
	wire [WIDTH-1:0] wire_d56_5;
	wire [WIDTH-1:0] wire_d56_6;
	wire [WIDTH-1:0] wire_d56_7;
	wire [WIDTH-1:0] wire_d56_8;
	wire [WIDTH-1:0] wire_d56_9;
	wire [WIDTH-1:0] wire_d56_10;
	wire [WIDTH-1:0] wire_d56_11;
	wire [WIDTH-1:0] wire_d56_12;
	wire [WIDTH-1:0] wire_d56_13;
	wire [WIDTH-1:0] wire_d56_14;
	wire [WIDTH-1:0] wire_d56_15;
	wire [WIDTH-1:0] wire_d56_16;
	wire [WIDTH-1:0] wire_d56_17;
	wire [WIDTH-1:0] wire_d56_18;
	wire [WIDTH-1:0] wire_d56_19;
	wire [WIDTH-1:0] wire_d56_20;
	wire [WIDTH-1:0] wire_d56_21;
	wire [WIDTH-1:0] wire_d56_22;
	wire [WIDTH-1:0] wire_d56_23;
	wire [WIDTH-1:0] wire_d56_24;
	wire [WIDTH-1:0] wire_d56_25;
	wire [WIDTH-1:0] wire_d56_26;
	wire [WIDTH-1:0] wire_d56_27;
	wire [WIDTH-1:0] wire_d56_28;
	wire [WIDTH-1:0] wire_d56_29;
	wire [WIDTH-1:0] wire_d56_30;
	wire [WIDTH-1:0] wire_d56_31;
	wire [WIDTH-1:0] wire_d56_32;
	wire [WIDTH-1:0] wire_d56_33;
	wire [WIDTH-1:0] wire_d56_34;
	wire [WIDTH-1:0] wire_d56_35;
	wire [WIDTH-1:0] wire_d56_36;
	wire [WIDTH-1:0] wire_d56_37;
	wire [WIDTH-1:0] wire_d56_38;
	wire [WIDTH-1:0] wire_d56_39;
	wire [WIDTH-1:0] wire_d56_40;
	wire [WIDTH-1:0] wire_d56_41;
	wire [WIDTH-1:0] wire_d56_42;
	wire [WIDTH-1:0] wire_d56_43;
	wire [WIDTH-1:0] wire_d56_44;
	wire [WIDTH-1:0] wire_d56_45;
	wire [WIDTH-1:0] wire_d56_46;
	wire [WIDTH-1:0] wire_d56_47;
	wire [WIDTH-1:0] wire_d56_48;
	wire [WIDTH-1:0] wire_d56_49;
	wire [WIDTH-1:0] wire_d56_50;
	wire [WIDTH-1:0] wire_d56_51;
	wire [WIDTH-1:0] wire_d56_52;
	wire [WIDTH-1:0] wire_d56_53;
	wire [WIDTH-1:0] wire_d56_54;
	wire [WIDTH-1:0] wire_d56_55;
	wire [WIDTH-1:0] wire_d56_56;
	wire [WIDTH-1:0] wire_d56_57;
	wire [WIDTH-1:0] wire_d56_58;
	wire [WIDTH-1:0] wire_d56_59;
	wire [WIDTH-1:0] wire_d56_60;
	wire [WIDTH-1:0] wire_d56_61;
	wire [WIDTH-1:0] wire_d56_62;
	wire [WIDTH-1:0] wire_d56_63;
	wire [WIDTH-1:0] wire_d56_64;
	wire [WIDTH-1:0] wire_d56_65;
	wire [WIDTH-1:0] wire_d56_66;
	wire [WIDTH-1:0] wire_d56_67;
	wire [WIDTH-1:0] wire_d56_68;
	wire [WIDTH-1:0] wire_d56_69;
	wire [WIDTH-1:0] wire_d56_70;
	wire [WIDTH-1:0] wire_d56_71;
	wire [WIDTH-1:0] wire_d56_72;
	wire [WIDTH-1:0] wire_d56_73;
	wire [WIDTH-1:0] wire_d56_74;
	wire [WIDTH-1:0] wire_d56_75;
	wire [WIDTH-1:0] wire_d56_76;
	wire [WIDTH-1:0] wire_d56_77;
	wire [WIDTH-1:0] wire_d56_78;
	wire [WIDTH-1:0] wire_d57_0;
	wire [WIDTH-1:0] wire_d57_1;
	wire [WIDTH-1:0] wire_d57_2;
	wire [WIDTH-1:0] wire_d57_3;
	wire [WIDTH-1:0] wire_d57_4;
	wire [WIDTH-1:0] wire_d57_5;
	wire [WIDTH-1:0] wire_d57_6;
	wire [WIDTH-1:0] wire_d57_7;
	wire [WIDTH-1:0] wire_d57_8;
	wire [WIDTH-1:0] wire_d57_9;
	wire [WIDTH-1:0] wire_d57_10;
	wire [WIDTH-1:0] wire_d57_11;
	wire [WIDTH-1:0] wire_d57_12;
	wire [WIDTH-1:0] wire_d57_13;
	wire [WIDTH-1:0] wire_d57_14;
	wire [WIDTH-1:0] wire_d57_15;
	wire [WIDTH-1:0] wire_d57_16;
	wire [WIDTH-1:0] wire_d57_17;
	wire [WIDTH-1:0] wire_d57_18;
	wire [WIDTH-1:0] wire_d57_19;
	wire [WIDTH-1:0] wire_d57_20;
	wire [WIDTH-1:0] wire_d57_21;
	wire [WIDTH-1:0] wire_d57_22;
	wire [WIDTH-1:0] wire_d57_23;
	wire [WIDTH-1:0] wire_d57_24;
	wire [WIDTH-1:0] wire_d57_25;
	wire [WIDTH-1:0] wire_d57_26;
	wire [WIDTH-1:0] wire_d57_27;
	wire [WIDTH-1:0] wire_d57_28;
	wire [WIDTH-1:0] wire_d57_29;
	wire [WIDTH-1:0] wire_d57_30;
	wire [WIDTH-1:0] wire_d57_31;
	wire [WIDTH-1:0] wire_d57_32;
	wire [WIDTH-1:0] wire_d57_33;
	wire [WIDTH-1:0] wire_d57_34;
	wire [WIDTH-1:0] wire_d57_35;
	wire [WIDTH-1:0] wire_d57_36;
	wire [WIDTH-1:0] wire_d57_37;
	wire [WIDTH-1:0] wire_d57_38;
	wire [WIDTH-1:0] wire_d57_39;
	wire [WIDTH-1:0] wire_d57_40;
	wire [WIDTH-1:0] wire_d57_41;
	wire [WIDTH-1:0] wire_d57_42;
	wire [WIDTH-1:0] wire_d57_43;
	wire [WIDTH-1:0] wire_d57_44;
	wire [WIDTH-1:0] wire_d57_45;
	wire [WIDTH-1:0] wire_d57_46;
	wire [WIDTH-1:0] wire_d57_47;
	wire [WIDTH-1:0] wire_d57_48;
	wire [WIDTH-1:0] wire_d57_49;
	wire [WIDTH-1:0] wire_d57_50;
	wire [WIDTH-1:0] wire_d57_51;
	wire [WIDTH-1:0] wire_d57_52;
	wire [WIDTH-1:0] wire_d57_53;
	wire [WIDTH-1:0] wire_d57_54;
	wire [WIDTH-1:0] wire_d57_55;
	wire [WIDTH-1:0] wire_d57_56;
	wire [WIDTH-1:0] wire_d57_57;
	wire [WIDTH-1:0] wire_d57_58;
	wire [WIDTH-1:0] wire_d57_59;
	wire [WIDTH-1:0] wire_d57_60;
	wire [WIDTH-1:0] wire_d57_61;
	wire [WIDTH-1:0] wire_d57_62;
	wire [WIDTH-1:0] wire_d57_63;
	wire [WIDTH-1:0] wire_d57_64;
	wire [WIDTH-1:0] wire_d57_65;
	wire [WIDTH-1:0] wire_d57_66;
	wire [WIDTH-1:0] wire_d57_67;
	wire [WIDTH-1:0] wire_d57_68;
	wire [WIDTH-1:0] wire_d57_69;
	wire [WIDTH-1:0] wire_d57_70;
	wire [WIDTH-1:0] wire_d57_71;
	wire [WIDTH-1:0] wire_d57_72;
	wire [WIDTH-1:0] wire_d57_73;
	wire [WIDTH-1:0] wire_d57_74;
	wire [WIDTH-1:0] wire_d57_75;
	wire [WIDTH-1:0] wire_d57_76;
	wire [WIDTH-1:0] wire_d57_77;
	wire [WIDTH-1:0] wire_d57_78;
	wire [WIDTH-1:0] wire_d58_0;
	wire [WIDTH-1:0] wire_d58_1;
	wire [WIDTH-1:0] wire_d58_2;
	wire [WIDTH-1:0] wire_d58_3;
	wire [WIDTH-1:0] wire_d58_4;
	wire [WIDTH-1:0] wire_d58_5;
	wire [WIDTH-1:0] wire_d58_6;
	wire [WIDTH-1:0] wire_d58_7;
	wire [WIDTH-1:0] wire_d58_8;
	wire [WIDTH-1:0] wire_d58_9;
	wire [WIDTH-1:0] wire_d58_10;
	wire [WIDTH-1:0] wire_d58_11;
	wire [WIDTH-1:0] wire_d58_12;
	wire [WIDTH-1:0] wire_d58_13;
	wire [WIDTH-1:0] wire_d58_14;
	wire [WIDTH-1:0] wire_d58_15;
	wire [WIDTH-1:0] wire_d58_16;
	wire [WIDTH-1:0] wire_d58_17;
	wire [WIDTH-1:0] wire_d58_18;
	wire [WIDTH-1:0] wire_d58_19;
	wire [WIDTH-1:0] wire_d58_20;
	wire [WIDTH-1:0] wire_d58_21;
	wire [WIDTH-1:0] wire_d58_22;
	wire [WIDTH-1:0] wire_d58_23;
	wire [WIDTH-1:0] wire_d58_24;
	wire [WIDTH-1:0] wire_d58_25;
	wire [WIDTH-1:0] wire_d58_26;
	wire [WIDTH-1:0] wire_d58_27;
	wire [WIDTH-1:0] wire_d58_28;
	wire [WIDTH-1:0] wire_d58_29;
	wire [WIDTH-1:0] wire_d58_30;
	wire [WIDTH-1:0] wire_d58_31;
	wire [WIDTH-1:0] wire_d58_32;
	wire [WIDTH-1:0] wire_d58_33;
	wire [WIDTH-1:0] wire_d58_34;
	wire [WIDTH-1:0] wire_d58_35;
	wire [WIDTH-1:0] wire_d58_36;
	wire [WIDTH-1:0] wire_d58_37;
	wire [WIDTH-1:0] wire_d58_38;
	wire [WIDTH-1:0] wire_d58_39;
	wire [WIDTH-1:0] wire_d58_40;
	wire [WIDTH-1:0] wire_d58_41;
	wire [WIDTH-1:0] wire_d58_42;
	wire [WIDTH-1:0] wire_d58_43;
	wire [WIDTH-1:0] wire_d58_44;
	wire [WIDTH-1:0] wire_d58_45;
	wire [WIDTH-1:0] wire_d58_46;
	wire [WIDTH-1:0] wire_d58_47;
	wire [WIDTH-1:0] wire_d58_48;
	wire [WIDTH-1:0] wire_d58_49;
	wire [WIDTH-1:0] wire_d58_50;
	wire [WIDTH-1:0] wire_d58_51;
	wire [WIDTH-1:0] wire_d58_52;
	wire [WIDTH-1:0] wire_d58_53;
	wire [WIDTH-1:0] wire_d58_54;
	wire [WIDTH-1:0] wire_d58_55;
	wire [WIDTH-1:0] wire_d58_56;
	wire [WIDTH-1:0] wire_d58_57;
	wire [WIDTH-1:0] wire_d58_58;
	wire [WIDTH-1:0] wire_d58_59;
	wire [WIDTH-1:0] wire_d58_60;
	wire [WIDTH-1:0] wire_d58_61;
	wire [WIDTH-1:0] wire_d58_62;
	wire [WIDTH-1:0] wire_d58_63;
	wire [WIDTH-1:0] wire_d58_64;
	wire [WIDTH-1:0] wire_d58_65;
	wire [WIDTH-1:0] wire_d58_66;
	wire [WIDTH-1:0] wire_d58_67;
	wire [WIDTH-1:0] wire_d58_68;
	wire [WIDTH-1:0] wire_d58_69;
	wire [WIDTH-1:0] wire_d58_70;
	wire [WIDTH-1:0] wire_d58_71;
	wire [WIDTH-1:0] wire_d58_72;
	wire [WIDTH-1:0] wire_d58_73;
	wire [WIDTH-1:0] wire_d58_74;
	wire [WIDTH-1:0] wire_d58_75;
	wire [WIDTH-1:0] wire_d58_76;
	wire [WIDTH-1:0] wire_d58_77;
	wire [WIDTH-1:0] wire_d58_78;
	wire [WIDTH-1:0] wire_d59_0;
	wire [WIDTH-1:0] wire_d59_1;
	wire [WIDTH-1:0] wire_d59_2;
	wire [WIDTH-1:0] wire_d59_3;
	wire [WIDTH-1:0] wire_d59_4;
	wire [WIDTH-1:0] wire_d59_5;
	wire [WIDTH-1:0] wire_d59_6;
	wire [WIDTH-1:0] wire_d59_7;
	wire [WIDTH-1:0] wire_d59_8;
	wire [WIDTH-1:0] wire_d59_9;
	wire [WIDTH-1:0] wire_d59_10;
	wire [WIDTH-1:0] wire_d59_11;
	wire [WIDTH-1:0] wire_d59_12;
	wire [WIDTH-1:0] wire_d59_13;
	wire [WIDTH-1:0] wire_d59_14;
	wire [WIDTH-1:0] wire_d59_15;
	wire [WIDTH-1:0] wire_d59_16;
	wire [WIDTH-1:0] wire_d59_17;
	wire [WIDTH-1:0] wire_d59_18;
	wire [WIDTH-1:0] wire_d59_19;
	wire [WIDTH-1:0] wire_d59_20;
	wire [WIDTH-1:0] wire_d59_21;
	wire [WIDTH-1:0] wire_d59_22;
	wire [WIDTH-1:0] wire_d59_23;
	wire [WIDTH-1:0] wire_d59_24;
	wire [WIDTH-1:0] wire_d59_25;
	wire [WIDTH-1:0] wire_d59_26;
	wire [WIDTH-1:0] wire_d59_27;
	wire [WIDTH-1:0] wire_d59_28;
	wire [WIDTH-1:0] wire_d59_29;
	wire [WIDTH-1:0] wire_d59_30;
	wire [WIDTH-1:0] wire_d59_31;
	wire [WIDTH-1:0] wire_d59_32;
	wire [WIDTH-1:0] wire_d59_33;
	wire [WIDTH-1:0] wire_d59_34;
	wire [WIDTH-1:0] wire_d59_35;
	wire [WIDTH-1:0] wire_d59_36;
	wire [WIDTH-1:0] wire_d59_37;
	wire [WIDTH-1:0] wire_d59_38;
	wire [WIDTH-1:0] wire_d59_39;
	wire [WIDTH-1:0] wire_d59_40;
	wire [WIDTH-1:0] wire_d59_41;
	wire [WIDTH-1:0] wire_d59_42;
	wire [WIDTH-1:0] wire_d59_43;
	wire [WIDTH-1:0] wire_d59_44;
	wire [WIDTH-1:0] wire_d59_45;
	wire [WIDTH-1:0] wire_d59_46;
	wire [WIDTH-1:0] wire_d59_47;
	wire [WIDTH-1:0] wire_d59_48;
	wire [WIDTH-1:0] wire_d59_49;
	wire [WIDTH-1:0] wire_d59_50;
	wire [WIDTH-1:0] wire_d59_51;
	wire [WIDTH-1:0] wire_d59_52;
	wire [WIDTH-1:0] wire_d59_53;
	wire [WIDTH-1:0] wire_d59_54;
	wire [WIDTH-1:0] wire_d59_55;
	wire [WIDTH-1:0] wire_d59_56;
	wire [WIDTH-1:0] wire_d59_57;
	wire [WIDTH-1:0] wire_d59_58;
	wire [WIDTH-1:0] wire_d59_59;
	wire [WIDTH-1:0] wire_d59_60;
	wire [WIDTH-1:0] wire_d59_61;
	wire [WIDTH-1:0] wire_d59_62;
	wire [WIDTH-1:0] wire_d59_63;
	wire [WIDTH-1:0] wire_d59_64;
	wire [WIDTH-1:0] wire_d59_65;
	wire [WIDTH-1:0] wire_d59_66;
	wire [WIDTH-1:0] wire_d59_67;
	wire [WIDTH-1:0] wire_d59_68;
	wire [WIDTH-1:0] wire_d59_69;
	wire [WIDTH-1:0] wire_d59_70;
	wire [WIDTH-1:0] wire_d59_71;
	wire [WIDTH-1:0] wire_d59_72;
	wire [WIDTH-1:0] wire_d59_73;
	wire [WIDTH-1:0] wire_d59_74;
	wire [WIDTH-1:0] wire_d59_75;
	wire [WIDTH-1:0] wire_d59_76;
	wire [WIDTH-1:0] wire_d59_77;
	wire [WIDTH-1:0] wire_d59_78;
	wire [WIDTH-1:0] wire_d60_0;
	wire [WIDTH-1:0] wire_d60_1;
	wire [WIDTH-1:0] wire_d60_2;
	wire [WIDTH-1:0] wire_d60_3;
	wire [WIDTH-1:0] wire_d60_4;
	wire [WIDTH-1:0] wire_d60_5;
	wire [WIDTH-1:0] wire_d60_6;
	wire [WIDTH-1:0] wire_d60_7;
	wire [WIDTH-1:0] wire_d60_8;
	wire [WIDTH-1:0] wire_d60_9;
	wire [WIDTH-1:0] wire_d60_10;
	wire [WIDTH-1:0] wire_d60_11;
	wire [WIDTH-1:0] wire_d60_12;
	wire [WIDTH-1:0] wire_d60_13;
	wire [WIDTH-1:0] wire_d60_14;
	wire [WIDTH-1:0] wire_d60_15;
	wire [WIDTH-1:0] wire_d60_16;
	wire [WIDTH-1:0] wire_d60_17;
	wire [WIDTH-1:0] wire_d60_18;
	wire [WIDTH-1:0] wire_d60_19;
	wire [WIDTH-1:0] wire_d60_20;
	wire [WIDTH-1:0] wire_d60_21;
	wire [WIDTH-1:0] wire_d60_22;
	wire [WIDTH-1:0] wire_d60_23;
	wire [WIDTH-1:0] wire_d60_24;
	wire [WIDTH-1:0] wire_d60_25;
	wire [WIDTH-1:0] wire_d60_26;
	wire [WIDTH-1:0] wire_d60_27;
	wire [WIDTH-1:0] wire_d60_28;
	wire [WIDTH-1:0] wire_d60_29;
	wire [WIDTH-1:0] wire_d60_30;
	wire [WIDTH-1:0] wire_d60_31;
	wire [WIDTH-1:0] wire_d60_32;
	wire [WIDTH-1:0] wire_d60_33;
	wire [WIDTH-1:0] wire_d60_34;
	wire [WIDTH-1:0] wire_d60_35;
	wire [WIDTH-1:0] wire_d60_36;
	wire [WIDTH-1:0] wire_d60_37;
	wire [WIDTH-1:0] wire_d60_38;
	wire [WIDTH-1:0] wire_d60_39;
	wire [WIDTH-1:0] wire_d60_40;
	wire [WIDTH-1:0] wire_d60_41;
	wire [WIDTH-1:0] wire_d60_42;
	wire [WIDTH-1:0] wire_d60_43;
	wire [WIDTH-1:0] wire_d60_44;
	wire [WIDTH-1:0] wire_d60_45;
	wire [WIDTH-1:0] wire_d60_46;
	wire [WIDTH-1:0] wire_d60_47;
	wire [WIDTH-1:0] wire_d60_48;
	wire [WIDTH-1:0] wire_d60_49;
	wire [WIDTH-1:0] wire_d60_50;
	wire [WIDTH-1:0] wire_d60_51;
	wire [WIDTH-1:0] wire_d60_52;
	wire [WIDTH-1:0] wire_d60_53;
	wire [WIDTH-1:0] wire_d60_54;
	wire [WIDTH-1:0] wire_d60_55;
	wire [WIDTH-1:0] wire_d60_56;
	wire [WIDTH-1:0] wire_d60_57;
	wire [WIDTH-1:0] wire_d60_58;
	wire [WIDTH-1:0] wire_d60_59;
	wire [WIDTH-1:0] wire_d60_60;
	wire [WIDTH-1:0] wire_d60_61;
	wire [WIDTH-1:0] wire_d60_62;
	wire [WIDTH-1:0] wire_d60_63;
	wire [WIDTH-1:0] wire_d60_64;
	wire [WIDTH-1:0] wire_d60_65;
	wire [WIDTH-1:0] wire_d60_66;
	wire [WIDTH-1:0] wire_d60_67;
	wire [WIDTH-1:0] wire_d60_68;
	wire [WIDTH-1:0] wire_d60_69;
	wire [WIDTH-1:0] wire_d60_70;
	wire [WIDTH-1:0] wire_d60_71;
	wire [WIDTH-1:0] wire_d60_72;
	wire [WIDTH-1:0] wire_d60_73;
	wire [WIDTH-1:0] wire_d60_74;
	wire [WIDTH-1:0] wire_d60_75;
	wire [WIDTH-1:0] wire_d60_76;
	wire [WIDTH-1:0] wire_d60_77;
	wire [WIDTH-1:0] wire_d60_78;
	wire [WIDTH-1:0] wire_d61_0;
	wire [WIDTH-1:0] wire_d61_1;
	wire [WIDTH-1:0] wire_d61_2;
	wire [WIDTH-1:0] wire_d61_3;
	wire [WIDTH-1:0] wire_d61_4;
	wire [WIDTH-1:0] wire_d61_5;
	wire [WIDTH-1:0] wire_d61_6;
	wire [WIDTH-1:0] wire_d61_7;
	wire [WIDTH-1:0] wire_d61_8;
	wire [WIDTH-1:0] wire_d61_9;
	wire [WIDTH-1:0] wire_d61_10;
	wire [WIDTH-1:0] wire_d61_11;
	wire [WIDTH-1:0] wire_d61_12;
	wire [WIDTH-1:0] wire_d61_13;
	wire [WIDTH-1:0] wire_d61_14;
	wire [WIDTH-1:0] wire_d61_15;
	wire [WIDTH-1:0] wire_d61_16;
	wire [WIDTH-1:0] wire_d61_17;
	wire [WIDTH-1:0] wire_d61_18;
	wire [WIDTH-1:0] wire_d61_19;
	wire [WIDTH-1:0] wire_d61_20;
	wire [WIDTH-1:0] wire_d61_21;
	wire [WIDTH-1:0] wire_d61_22;
	wire [WIDTH-1:0] wire_d61_23;
	wire [WIDTH-1:0] wire_d61_24;
	wire [WIDTH-1:0] wire_d61_25;
	wire [WIDTH-1:0] wire_d61_26;
	wire [WIDTH-1:0] wire_d61_27;
	wire [WIDTH-1:0] wire_d61_28;
	wire [WIDTH-1:0] wire_d61_29;
	wire [WIDTH-1:0] wire_d61_30;
	wire [WIDTH-1:0] wire_d61_31;
	wire [WIDTH-1:0] wire_d61_32;
	wire [WIDTH-1:0] wire_d61_33;
	wire [WIDTH-1:0] wire_d61_34;
	wire [WIDTH-1:0] wire_d61_35;
	wire [WIDTH-1:0] wire_d61_36;
	wire [WIDTH-1:0] wire_d61_37;
	wire [WIDTH-1:0] wire_d61_38;
	wire [WIDTH-1:0] wire_d61_39;
	wire [WIDTH-1:0] wire_d61_40;
	wire [WIDTH-1:0] wire_d61_41;
	wire [WIDTH-1:0] wire_d61_42;
	wire [WIDTH-1:0] wire_d61_43;
	wire [WIDTH-1:0] wire_d61_44;
	wire [WIDTH-1:0] wire_d61_45;
	wire [WIDTH-1:0] wire_d61_46;
	wire [WIDTH-1:0] wire_d61_47;
	wire [WIDTH-1:0] wire_d61_48;
	wire [WIDTH-1:0] wire_d61_49;
	wire [WIDTH-1:0] wire_d61_50;
	wire [WIDTH-1:0] wire_d61_51;
	wire [WIDTH-1:0] wire_d61_52;
	wire [WIDTH-1:0] wire_d61_53;
	wire [WIDTH-1:0] wire_d61_54;
	wire [WIDTH-1:0] wire_d61_55;
	wire [WIDTH-1:0] wire_d61_56;
	wire [WIDTH-1:0] wire_d61_57;
	wire [WIDTH-1:0] wire_d61_58;
	wire [WIDTH-1:0] wire_d61_59;
	wire [WIDTH-1:0] wire_d61_60;
	wire [WIDTH-1:0] wire_d61_61;
	wire [WIDTH-1:0] wire_d61_62;
	wire [WIDTH-1:0] wire_d61_63;
	wire [WIDTH-1:0] wire_d61_64;
	wire [WIDTH-1:0] wire_d61_65;
	wire [WIDTH-1:0] wire_d61_66;
	wire [WIDTH-1:0] wire_d61_67;
	wire [WIDTH-1:0] wire_d61_68;
	wire [WIDTH-1:0] wire_d61_69;
	wire [WIDTH-1:0] wire_d61_70;
	wire [WIDTH-1:0] wire_d61_71;
	wire [WIDTH-1:0] wire_d61_72;
	wire [WIDTH-1:0] wire_d61_73;
	wire [WIDTH-1:0] wire_d61_74;
	wire [WIDTH-1:0] wire_d61_75;
	wire [WIDTH-1:0] wire_d61_76;
	wire [WIDTH-1:0] wire_d61_77;
	wire [WIDTH-1:0] wire_d61_78;
	wire [WIDTH-1:0] wire_d62_0;
	wire [WIDTH-1:0] wire_d62_1;
	wire [WIDTH-1:0] wire_d62_2;
	wire [WIDTH-1:0] wire_d62_3;
	wire [WIDTH-1:0] wire_d62_4;
	wire [WIDTH-1:0] wire_d62_5;
	wire [WIDTH-1:0] wire_d62_6;
	wire [WIDTH-1:0] wire_d62_7;
	wire [WIDTH-1:0] wire_d62_8;
	wire [WIDTH-1:0] wire_d62_9;
	wire [WIDTH-1:0] wire_d62_10;
	wire [WIDTH-1:0] wire_d62_11;
	wire [WIDTH-1:0] wire_d62_12;
	wire [WIDTH-1:0] wire_d62_13;
	wire [WIDTH-1:0] wire_d62_14;
	wire [WIDTH-1:0] wire_d62_15;
	wire [WIDTH-1:0] wire_d62_16;
	wire [WIDTH-1:0] wire_d62_17;
	wire [WIDTH-1:0] wire_d62_18;
	wire [WIDTH-1:0] wire_d62_19;
	wire [WIDTH-1:0] wire_d62_20;
	wire [WIDTH-1:0] wire_d62_21;
	wire [WIDTH-1:0] wire_d62_22;
	wire [WIDTH-1:0] wire_d62_23;
	wire [WIDTH-1:0] wire_d62_24;
	wire [WIDTH-1:0] wire_d62_25;
	wire [WIDTH-1:0] wire_d62_26;
	wire [WIDTH-1:0] wire_d62_27;
	wire [WIDTH-1:0] wire_d62_28;
	wire [WIDTH-1:0] wire_d62_29;
	wire [WIDTH-1:0] wire_d62_30;
	wire [WIDTH-1:0] wire_d62_31;
	wire [WIDTH-1:0] wire_d62_32;
	wire [WIDTH-1:0] wire_d62_33;
	wire [WIDTH-1:0] wire_d62_34;
	wire [WIDTH-1:0] wire_d62_35;
	wire [WIDTH-1:0] wire_d62_36;
	wire [WIDTH-1:0] wire_d62_37;
	wire [WIDTH-1:0] wire_d62_38;
	wire [WIDTH-1:0] wire_d62_39;
	wire [WIDTH-1:0] wire_d62_40;
	wire [WIDTH-1:0] wire_d62_41;
	wire [WIDTH-1:0] wire_d62_42;
	wire [WIDTH-1:0] wire_d62_43;
	wire [WIDTH-1:0] wire_d62_44;
	wire [WIDTH-1:0] wire_d62_45;
	wire [WIDTH-1:0] wire_d62_46;
	wire [WIDTH-1:0] wire_d62_47;
	wire [WIDTH-1:0] wire_d62_48;
	wire [WIDTH-1:0] wire_d62_49;
	wire [WIDTH-1:0] wire_d62_50;
	wire [WIDTH-1:0] wire_d62_51;
	wire [WIDTH-1:0] wire_d62_52;
	wire [WIDTH-1:0] wire_d62_53;
	wire [WIDTH-1:0] wire_d62_54;
	wire [WIDTH-1:0] wire_d62_55;
	wire [WIDTH-1:0] wire_d62_56;
	wire [WIDTH-1:0] wire_d62_57;
	wire [WIDTH-1:0] wire_d62_58;
	wire [WIDTH-1:0] wire_d62_59;
	wire [WIDTH-1:0] wire_d62_60;
	wire [WIDTH-1:0] wire_d62_61;
	wire [WIDTH-1:0] wire_d62_62;
	wire [WIDTH-1:0] wire_d62_63;
	wire [WIDTH-1:0] wire_d62_64;
	wire [WIDTH-1:0] wire_d62_65;
	wire [WIDTH-1:0] wire_d62_66;
	wire [WIDTH-1:0] wire_d62_67;
	wire [WIDTH-1:0] wire_d62_68;
	wire [WIDTH-1:0] wire_d62_69;
	wire [WIDTH-1:0] wire_d62_70;
	wire [WIDTH-1:0] wire_d62_71;
	wire [WIDTH-1:0] wire_d62_72;
	wire [WIDTH-1:0] wire_d62_73;
	wire [WIDTH-1:0] wire_d62_74;
	wire [WIDTH-1:0] wire_d62_75;
	wire [WIDTH-1:0] wire_d62_76;
	wire [WIDTH-1:0] wire_d62_77;
	wire [WIDTH-1:0] wire_d62_78;
	wire [WIDTH-1:0] wire_d63_0;
	wire [WIDTH-1:0] wire_d63_1;
	wire [WIDTH-1:0] wire_d63_2;
	wire [WIDTH-1:0] wire_d63_3;
	wire [WIDTH-1:0] wire_d63_4;
	wire [WIDTH-1:0] wire_d63_5;
	wire [WIDTH-1:0] wire_d63_6;
	wire [WIDTH-1:0] wire_d63_7;
	wire [WIDTH-1:0] wire_d63_8;
	wire [WIDTH-1:0] wire_d63_9;
	wire [WIDTH-1:0] wire_d63_10;
	wire [WIDTH-1:0] wire_d63_11;
	wire [WIDTH-1:0] wire_d63_12;
	wire [WIDTH-1:0] wire_d63_13;
	wire [WIDTH-1:0] wire_d63_14;
	wire [WIDTH-1:0] wire_d63_15;
	wire [WIDTH-1:0] wire_d63_16;
	wire [WIDTH-1:0] wire_d63_17;
	wire [WIDTH-1:0] wire_d63_18;
	wire [WIDTH-1:0] wire_d63_19;
	wire [WIDTH-1:0] wire_d63_20;
	wire [WIDTH-1:0] wire_d63_21;
	wire [WIDTH-1:0] wire_d63_22;
	wire [WIDTH-1:0] wire_d63_23;
	wire [WIDTH-1:0] wire_d63_24;
	wire [WIDTH-1:0] wire_d63_25;
	wire [WIDTH-1:0] wire_d63_26;
	wire [WIDTH-1:0] wire_d63_27;
	wire [WIDTH-1:0] wire_d63_28;
	wire [WIDTH-1:0] wire_d63_29;
	wire [WIDTH-1:0] wire_d63_30;
	wire [WIDTH-1:0] wire_d63_31;
	wire [WIDTH-1:0] wire_d63_32;
	wire [WIDTH-1:0] wire_d63_33;
	wire [WIDTH-1:0] wire_d63_34;
	wire [WIDTH-1:0] wire_d63_35;
	wire [WIDTH-1:0] wire_d63_36;
	wire [WIDTH-1:0] wire_d63_37;
	wire [WIDTH-1:0] wire_d63_38;
	wire [WIDTH-1:0] wire_d63_39;
	wire [WIDTH-1:0] wire_d63_40;
	wire [WIDTH-1:0] wire_d63_41;
	wire [WIDTH-1:0] wire_d63_42;
	wire [WIDTH-1:0] wire_d63_43;
	wire [WIDTH-1:0] wire_d63_44;
	wire [WIDTH-1:0] wire_d63_45;
	wire [WIDTH-1:0] wire_d63_46;
	wire [WIDTH-1:0] wire_d63_47;
	wire [WIDTH-1:0] wire_d63_48;
	wire [WIDTH-1:0] wire_d63_49;
	wire [WIDTH-1:0] wire_d63_50;
	wire [WIDTH-1:0] wire_d63_51;
	wire [WIDTH-1:0] wire_d63_52;
	wire [WIDTH-1:0] wire_d63_53;
	wire [WIDTH-1:0] wire_d63_54;
	wire [WIDTH-1:0] wire_d63_55;
	wire [WIDTH-1:0] wire_d63_56;
	wire [WIDTH-1:0] wire_d63_57;
	wire [WIDTH-1:0] wire_d63_58;
	wire [WIDTH-1:0] wire_d63_59;
	wire [WIDTH-1:0] wire_d63_60;
	wire [WIDTH-1:0] wire_d63_61;
	wire [WIDTH-1:0] wire_d63_62;
	wire [WIDTH-1:0] wire_d63_63;
	wire [WIDTH-1:0] wire_d63_64;
	wire [WIDTH-1:0] wire_d63_65;
	wire [WIDTH-1:0] wire_d63_66;
	wire [WIDTH-1:0] wire_d63_67;
	wire [WIDTH-1:0] wire_d63_68;
	wire [WIDTH-1:0] wire_d63_69;
	wire [WIDTH-1:0] wire_d63_70;
	wire [WIDTH-1:0] wire_d63_71;
	wire [WIDTH-1:0] wire_d63_72;
	wire [WIDTH-1:0] wire_d63_73;
	wire [WIDTH-1:0] wire_d63_74;
	wire [WIDTH-1:0] wire_d63_75;
	wire [WIDTH-1:0] wire_d63_76;
	wire [WIDTH-1:0] wire_d63_77;
	wire [WIDTH-1:0] wire_d63_78;
	wire [WIDTH-1:0] wire_d64_0;
	wire [WIDTH-1:0] wire_d64_1;
	wire [WIDTH-1:0] wire_d64_2;
	wire [WIDTH-1:0] wire_d64_3;
	wire [WIDTH-1:0] wire_d64_4;
	wire [WIDTH-1:0] wire_d64_5;
	wire [WIDTH-1:0] wire_d64_6;
	wire [WIDTH-1:0] wire_d64_7;
	wire [WIDTH-1:0] wire_d64_8;
	wire [WIDTH-1:0] wire_d64_9;
	wire [WIDTH-1:0] wire_d64_10;
	wire [WIDTH-1:0] wire_d64_11;
	wire [WIDTH-1:0] wire_d64_12;
	wire [WIDTH-1:0] wire_d64_13;
	wire [WIDTH-1:0] wire_d64_14;
	wire [WIDTH-1:0] wire_d64_15;
	wire [WIDTH-1:0] wire_d64_16;
	wire [WIDTH-1:0] wire_d64_17;
	wire [WIDTH-1:0] wire_d64_18;
	wire [WIDTH-1:0] wire_d64_19;
	wire [WIDTH-1:0] wire_d64_20;
	wire [WIDTH-1:0] wire_d64_21;
	wire [WIDTH-1:0] wire_d64_22;
	wire [WIDTH-1:0] wire_d64_23;
	wire [WIDTH-1:0] wire_d64_24;
	wire [WIDTH-1:0] wire_d64_25;
	wire [WIDTH-1:0] wire_d64_26;
	wire [WIDTH-1:0] wire_d64_27;
	wire [WIDTH-1:0] wire_d64_28;
	wire [WIDTH-1:0] wire_d64_29;
	wire [WIDTH-1:0] wire_d64_30;
	wire [WIDTH-1:0] wire_d64_31;
	wire [WIDTH-1:0] wire_d64_32;
	wire [WIDTH-1:0] wire_d64_33;
	wire [WIDTH-1:0] wire_d64_34;
	wire [WIDTH-1:0] wire_d64_35;
	wire [WIDTH-1:0] wire_d64_36;
	wire [WIDTH-1:0] wire_d64_37;
	wire [WIDTH-1:0] wire_d64_38;
	wire [WIDTH-1:0] wire_d64_39;
	wire [WIDTH-1:0] wire_d64_40;
	wire [WIDTH-1:0] wire_d64_41;
	wire [WIDTH-1:0] wire_d64_42;
	wire [WIDTH-1:0] wire_d64_43;
	wire [WIDTH-1:0] wire_d64_44;
	wire [WIDTH-1:0] wire_d64_45;
	wire [WIDTH-1:0] wire_d64_46;
	wire [WIDTH-1:0] wire_d64_47;
	wire [WIDTH-1:0] wire_d64_48;
	wire [WIDTH-1:0] wire_d64_49;
	wire [WIDTH-1:0] wire_d64_50;
	wire [WIDTH-1:0] wire_d64_51;
	wire [WIDTH-1:0] wire_d64_52;
	wire [WIDTH-1:0] wire_d64_53;
	wire [WIDTH-1:0] wire_d64_54;
	wire [WIDTH-1:0] wire_d64_55;
	wire [WIDTH-1:0] wire_d64_56;
	wire [WIDTH-1:0] wire_d64_57;
	wire [WIDTH-1:0] wire_d64_58;
	wire [WIDTH-1:0] wire_d64_59;
	wire [WIDTH-1:0] wire_d64_60;
	wire [WIDTH-1:0] wire_d64_61;
	wire [WIDTH-1:0] wire_d64_62;
	wire [WIDTH-1:0] wire_d64_63;
	wire [WIDTH-1:0] wire_d64_64;
	wire [WIDTH-1:0] wire_d64_65;
	wire [WIDTH-1:0] wire_d64_66;
	wire [WIDTH-1:0] wire_d64_67;
	wire [WIDTH-1:0] wire_d64_68;
	wire [WIDTH-1:0] wire_d64_69;
	wire [WIDTH-1:0] wire_d64_70;
	wire [WIDTH-1:0] wire_d64_71;
	wire [WIDTH-1:0] wire_d64_72;
	wire [WIDTH-1:0] wire_d64_73;
	wire [WIDTH-1:0] wire_d64_74;
	wire [WIDTH-1:0] wire_d64_75;
	wire [WIDTH-1:0] wire_d64_76;
	wire [WIDTH-1:0] wire_d64_77;
	wire [WIDTH-1:0] wire_d64_78;
	wire [WIDTH-1:0] wire_d65_0;
	wire [WIDTH-1:0] wire_d65_1;
	wire [WIDTH-1:0] wire_d65_2;
	wire [WIDTH-1:0] wire_d65_3;
	wire [WIDTH-1:0] wire_d65_4;
	wire [WIDTH-1:0] wire_d65_5;
	wire [WIDTH-1:0] wire_d65_6;
	wire [WIDTH-1:0] wire_d65_7;
	wire [WIDTH-1:0] wire_d65_8;
	wire [WIDTH-1:0] wire_d65_9;
	wire [WIDTH-1:0] wire_d65_10;
	wire [WIDTH-1:0] wire_d65_11;
	wire [WIDTH-1:0] wire_d65_12;
	wire [WIDTH-1:0] wire_d65_13;
	wire [WIDTH-1:0] wire_d65_14;
	wire [WIDTH-1:0] wire_d65_15;
	wire [WIDTH-1:0] wire_d65_16;
	wire [WIDTH-1:0] wire_d65_17;
	wire [WIDTH-1:0] wire_d65_18;
	wire [WIDTH-1:0] wire_d65_19;
	wire [WIDTH-1:0] wire_d65_20;
	wire [WIDTH-1:0] wire_d65_21;
	wire [WIDTH-1:0] wire_d65_22;
	wire [WIDTH-1:0] wire_d65_23;
	wire [WIDTH-1:0] wire_d65_24;
	wire [WIDTH-1:0] wire_d65_25;
	wire [WIDTH-1:0] wire_d65_26;
	wire [WIDTH-1:0] wire_d65_27;
	wire [WIDTH-1:0] wire_d65_28;
	wire [WIDTH-1:0] wire_d65_29;
	wire [WIDTH-1:0] wire_d65_30;
	wire [WIDTH-1:0] wire_d65_31;
	wire [WIDTH-1:0] wire_d65_32;
	wire [WIDTH-1:0] wire_d65_33;
	wire [WIDTH-1:0] wire_d65_34;
	wire [WIDTH-1:0] wire_d65_35;
	wire [WIDTH-1:0] wire_d65_36;
	wire [WIDTH-1:0] wire_d65_37;
	wire [WIDTH-1:0] wire_d65_38;
	wire [WIDTH-1:0] wire_d65_39;
	wire [WIDTH-1:0] wire_d65_40;
	wire [WIDTH-1:0] wire_d65_41;
	wire [WIDTH-1:0] wire_d65_42;
	wire [WIDTH-1:0] wire_d65_43;
	wire [WIDTH-1:0] wire_d65_44;
	wire [WIDTH-1:0] wire_d65_45;
	wire [WIDTH-1:0] wire_d65_46;
	wire [WIDTH-1:0] wire_d65_47;
	wire [WIDTH-1:0] wire_d65_48;
	wire [WIDTH-1:0] wire_d65_49;
	wire [WIDTH-1:0] wire_d65_50;
	wire [WIDTH-1:0] wire_d65_51;
	wire [WIDTH-1:0] wire_d65_52;
	wire [WIDTH-1:0] wire_d65_53;
	wire [WIDTH-1:0] wire_d65_54;
	wire [WIDTH-1:0] wire_d65_55;
	wire [WIDTH-1:0] wire_d65_56;
	wire [WIDTH-1:0] wire_d65_57;
	wire [WIDTH-1:0] wire_d65_58;
	wire [WIDTH-1:0] wire_d65_59;
	wire [WIDTH-1:0] wire_d65_60;
	wire [WIDTH-1:0] wire_d65_61;
	wire [WIDTH-1:0] wire_d65_62;
	wire [WIDTH-1:0] wire_d65_63;
	wire [WIDTH-1:0] wire_d65_64;
	wire [WIDTH-1:0] wire_d65_65;
	wire [WIDTH-1:0] wire_d65_66;
	wire [WIDTH-1:0] wire_d65_67;
	wire [WIDTH-1:0] wire_d65_68;
	wire [WIDTH-1:0] wire_d65_69;
	wire [WIDTH-1:0] wire_d65_70;
	wire [WIDTH-1:0] wire_d65_71;
	wire [WIDTH-1:0] wire_d65_72;
	wire [WIDTH-1:0] wire_d65_73;
	wire [WIDTH-1:0] wire_d65_74;
	wire [WIDTH-1:0] wire_d65_75;
	wire [WIDTH-1:0] wire_d65_76;
	wire [WIDTH-1:0] wire_d65_77;
	wire [WIDTH-1:0] wire_d65_78;
	wire [WIDTH-1:0] wire_d66_0;
	wire [WIDTH-1:0] wire_d66_1;
	wire [WIDTH-1:0] wire_d66_2;
	wire [WIDTH-1:0] wire_d66_3;
	wire [WIDTH-1:0] wire_d66_4;
	wire [WIDTH-1:0] wire_d66_5;
	wire [WIDTH-1:0] wire_d66_6;
	wire [WIDTH-1:0] wire_d66_7;
	wire [WIDTH-1:0] wire_d66_8;
	wire [WIDTH-1:0] wire_d66_9;
	wire [WIDTH-1:0] wire_d66_10;
	wire [WIDTH-1:0] wire_d66_11;
	wire [WIDTH-1:0] wire_d66_12;
	wire [WIDTH-1:0] wire_d66_13;
	wire [WIDTH-1:0] wire_d66_14;
	wire [WIDTH-1:0] wire_d66_15;
	wire [WIDTH-1:0] wire_d66_16;
	wire [WIDTH-1:0] wire_d66_17;
	wire [WIDTH-1:0] wire_d66_18;
	wire [WIDTH-1:0] wire_d66_19;
	wire [WIDTH-1:0] wire_d66_20;
	wire [WIDTH-1:0] wire_d66_21;
	wire [WIDTH-1:0] wire_d66_22;
	wire [WIDTH-1:0] wire_d66_23;
	wire [WIDTH-1:0] wire_d66_24;
	wire [WIDTH-1:0] wire_d66_25;
	wire [WIDTH-1:0] wire_d66_26;
	wire [WIDTH-1:0] wire_d66_27;
	wire [WIDTH-1:0] wire_d66_28;
	wire [WIDTH-1:0] wire_d66_29;
	wire [WIDTH-1:0] wire_d66_30;
	wire [WIDTH-1:0] wire_d66_31;
	wire [WIDTH-1:0] wire_d66_32;
	wire [WIDTH-1:0] wire_d66_33;
	wire [WIDTH-1:0] wire_d66_34;
	wire [WIDTH-1:0] wire_d66_35;
	wire [WIDTH-1:0] wire_d66_36;
	wire [WIDTH-1:0] wire_d66_37;
	wire [WIDTH-1:0] wire_d66_38;
	wire [WIDTH-1:0] wire_d66_39;
	wire [WIDTH-1:0] wire_d66_40;
	wire [WIDTH-1:0] wire_d66_41;
	wire [WIDTH-1:0] wire_d66_42;
	wire [WIDTH-1:0] wire_d66_43;
	wire [WIDTH-1:0] wire_d66_44;
	wire [WIDTH-1:0] wire_d66_45;
	wire [WIDTH-1:0] wire_d66_46;
	wire [WIDTH-1:0] wire_d66_47;
	wire [WIDTH-1:0] wire_d66_48;
	wire [WIDTH-1:0] wire_d66_49;
	wire [WIDTH-1:0] wire_d66_50;
	wire [WIDTH-1:0] wire_d66_51;
	wire [WIDTH-1:0] wire_d66_52;
	wire [WIDTH-1:0] wire_d66_53;
	wire [WIDTH-1:0] wire_d66_54;
	wire [WIDTH-1:0] wire_d66_55;
	wire [WIDTH-1:0] wire_d66_56;
	wire [WIDTH-1:0] wire_d66_57;
	wire [WIDTH-1:0] wire_d66_58;
	wire [WIDTH-1:0] wire_d66_59;
	wire [WIDTH-1:0] wire_d66_60;
	wire [WIDTH-1:0] wire_d66_61;
	wire [WIDTH-1:0] wire_d66_62;
	wire [WIDTH-1:0] wire_d66_63;
	wire [WIDTH-1:0] wire_d66_64;
	wire [WIDTH-1:0] wire_d66_65;
	wire [WIDTH-1:0] wire_d66_66;
	wire [WIDTH-1:0] wire_d66_67;
	wire [WIDTH-1:0] wire_d66_68;
	wire [WIDTH-1:0] wire_d66_69;
	wire [WIDTH-1:0] wire_d66_70;
	wire [WIDTH-1:0] wire_d66_71;
	wire [WIDTH-1:0] wire_d66_72;
	wire [WIDTH-1:0] wire_d66_73;
	wire [WIDTH-1:0] wire_d66_74;
	wire [WIDTH-1:0] wire_d66_75;
	wire [WIDTH-1:0] wire_d66_76;
	wire [WIDTH-1:0] wire_d66_77;
	wire [WIDTH-1:0] wire_d66_78;
	wire [WIDTH-1:0] wire_d67_0;
	wire [WIDTH-1:0] wire_d67_1;
	wire [WIDTH-1:0] wire_d67_2;
	wire [WIDTH-1:0] wire_d67_3;
	wire [WIDTH-1:0] wire_d67_4;
	wire [WIDTH-1:0] wire_d67_5;
	wire [WIDTH-1:0] wire_d67_6;
	wire [WIDTH-1:0] wire_d67_7;
	wire [WIDTH-1:0] wire_d67_8;
	wire [WIDTH-1:0] wire_d67_9;
	wire [WIDTH-1:0] wire_d67_10;
	wire [WIDTH-1:0] wire_d67_11;
	wire [WIDTH-1:0] wire_d67_12;
	wire [WIDTH-1:0] wire_d67_13;
	wire [WIDTH-1:0] wire_d67_14;
	wire [WIDTH-1:0] wire_d67_15;
	wire [WIDTH-1:0] wire_d67_16;
	wire [WIDTH-1:0] wire_d67_17;
	wire [WIDTH-1:0] wire_d67_18;
	wire [WIDTH-1:0] wire_d67_19;
	wire [WIDTH-1:0] wire_d67_20;
	wire [WIDTH-1:0] wire_d67_21;
	wire [WIDTH-1:0] wire_d67_22;
	wire [WIDTH-1:0] wire_d67_23;
	wire [WIDTH-1:0] wire_d67_24;
	wire [WIDTH-1:0] wire_d67_25;
	wire [WIDTH-1:0] wire_d67_26;
	wire [WIDTH-1:0] wire_d67_27;
	wire [WIDTH-1:0] wire_d67_28;
	wire [WIDTH-1:0] wire_d67_29;
	wire [WIDTH-1:0] wire_d67_30;
	wire [WIDTH-1:0] wire_d67_31;
	wire [WIDTH-1:0] wire_d67_32;
	wire [WIDTH-1:0] wire_d67_33;
	wire [WIDTH-1:0] wire_d67_34;
	wire [WIDTH-1:0] wire_d67_35;
	wire [WIDTH-1:0] wire_d67_36;
	wire [WIDTH-1:0] wire_d67_37;
	wire [WIDTH-1:0] wire_d67_38;
	wire [WIDTH-1:0] wire_d67_39;
	wire [WIDTH-1:0] wire_d67_40;
	wire [WIDTH-1:0] wire_d67_41;
	wire [WIDTH-1:0] wire_d67_42;
	wire [WIDTH-1:0] wire_d67_43;
	wire [WIDTH-1:0] wire_d67_44;
	wire [WIDTH-1:0] wire_d67_45;
	wire [WIDTH-1:0] wire_d67_46;
	wire [WIDTH-1:0] wire_d67_47;
	wire [WIDTH-1:0] wire_d67_48;
	wire [WIDTH-1:0] wire_d67_49;
	wire [WIDTH-1:0] wire_d67_50;
	wire [WIDTH-1:0] wire_d67_51;
	wire [WIDTH-1:0] wire_d67_52;
	wire [WIDTH-1:0] wire_d67_53;
	wire [WIDTH-1:0] wire_d67_54;
	wire [WIDTH-1:0] wire_d67_55;
	wire [WIDTH-1:0] wire_d67_56;
	wire [WIDTH-1:0] wire_d67_57;
	wire [WIDTH-1:0] wire_d67_58;
	wire [WIDTH-1:0] wire_d67_59;
	wire [WIDTH-1:0] wire_d67_60;
	wire [WIDTH-1:0] wire_d67_61;
	wire [WIDTH-1:0] wire_d67_62;
	wire [WIDTH-1:0] wire_d67_63;
	wire [WIDTH-1:0] wire_d67_64;
	wire [WIDTH-1:0] wire_d67_65;
	wire [WIDTH-1:0] wire_d67_66;
	wire [WIDTH-1:0] wire_d67_67;
	wire [WIDTH-1:0] wire_d67_68;
	wire [WIDTH-1:0] wire_d67_69;
	wire [WIDTH-1:0] wire_d67_70;
	wire [WIDTH-1:0] wire_d67_71;
	wire [WIDTH-1:0] wire_d67_72;
	wire [WIDTH-1:0] wire_d67_73;
	wire [WIDTH-1:0] wire_d67_74;
	wire [WIDTH-1:0] wire_d67_75;
	wire [WIDTH-1:0] wire_d67_76;
	wire [WIDTH-1:0] wire_d67_77;
	wire [WIDTH-1:0] wire_d67_78;
	wire [WIDTH-1:0] wire_d68_0;
	wire [WIDTH-1:0] wire_d68_1;
	wire [WIDTH-1:0] wire_d68_2;
	wire [WIDTH-1:0] wire_d68_3;
	wire [WIDTH-1:0] wire_d68_4;
	wire [WIDTH-1:0] wire_d68_5;
	wire [WIDTH-1:0] wire_d68_6;
	wire [WIDTH-1:0] wire_d68_7;
	wire [WIDTH-1:0] wire_d68_8;
	wire [WIDTH-1:0] wire_d68_9;
	wire [WIDTH-1:0] wire_d68_10;
	wire [WIDTH-1:0] wire_d68_11;
	wire [WIDTH-1:0] wire_d68_12;
	wire [WIDTH-1:0] wire_d68_13;
	wire [WIDTH-1:0] wire_d68_14;
	wire [WIDTH-1:0] wire_d68_15;
	wire [WIDTH-1:0] wire_d68_16;
	wire [WIDTH-1:0] wire_d68_17;
	wire [WIDTH-1:0] wire_d68_18;
	wire [WIDTH-1:0] wire_d68_19;
	wire [WIDTH-1:0] wire_d68_20;
	wire [WIDTH-1:0] wire_d68_21;
	wire [WIDTH-1:0] wire_d68_22;
	wire [WIDTH-1:0] wire_d68_23;
	wire [WIDTH-1:0] wire_d68_24;
	wire [WIDTH-1:0] wire_d68_25;
	wire [WIDTH-1:0] wire_d68_26;
	wire [WIDTH-1:0] wire_d68_27;
	wire [WIDTH-1:0] wire_d68_28;
	wire [WIDTH-1:0] wire_d68_29;
	wire [WIDTH-1:0] wire_d68_30;
	wire [WIDTH-1:0] wire_d68_31;
	wire [WIDTH-1:0] wire_d68_32;
	wire [WIDTH-1:0] wire_d68_33;
	wire [WIDTH-1:0] wire_d68_34;
	wire [WIDTH-1:0] wire_d68_35;
	wire [WIDTH-1:0] wire_d68_36;
	wire [WIDTH-1:0] wire_d68_37;
	wire [WIDTH-1:0] wire_d68_38;
	wire [WIDTH-1:0] wire_d68_39;
	wire [WIDTH-1:0] wire_d68_40;
	wire [WIDTH-1:0] wire_d68_41;
	wire [WIDTH-1:0] wire_d68_42;
	wire [WIDTH-1:0] wire_d68_43;
	wire [WIDTH-1:0] wire_d68_44;
	wire [WIDTH-1:0] wire_d68_45;
	wire [WIDTH-1:0] wire_d68_46;
	wire [WIDTH-1:0] wire_d68_47;
	wire [WIDTH-1:0] wire_d68_48;
	wire [WIDTH-1:0] wire_d68_49;
	wire [WIDTH-1:0] wire_d68_50;
	wire [WIDTH-1:0] wire_d68_51;
	wire [WIDTH-1:0] wire_d68_52;
	wire [WIDTH-1:0] wire_d68_53;
	wire [WIDTH-1:0] wire_d68_54;
	wire [WIDTH-1:0] wire_d68_55;
	wire [WIDTH-1:0] wire_d68_56;
	wire [WIDTH-1:0] wire_d68_57;
	wire [WIDTH-1:0] wire_d68_58;
	wire [WIDTH-1:0] wire_d68_59;
	wire [WIDTH-1:0] wire_d68_60;
	wire [WIDTH-1:0] wire_d68_61;
	wire [WIDTH-1:0] wire_d68_62;
	wire [WIDTH-1:0] wire_d68_63;
	wire [WIDTH-1:0] wire_d68_64;
	wire [WIDTH-1:0] wire_d68_65;
	wire [WIDTH-1:0] wire_d68_66;
	wire [WIDTH-1:0] wire_d68_67;
	wire [WIDTH-1:0] wire_d68_68;
	wire [WIDTH-1:0] wire_d68_69;
	wire [WIDTH-1:0] wire_d68_70;
	wire [WIDTH-1:0] wire_d68_71;
	wire [WIDTH-1:0] wire_d68_72;
	wire [WIDTH-1:0] wire_d68_73;
	wire [WIDTH-1:0] wire_d68_74;
	wire [WIDTH-1:0] wire_d68_75;
	wire [WIDTH-1:0] wire_d68_76;
	wire [WIDTH-1:0] wire_d68_77;
	wire [WIDTH-1:0] wire_d68_78;
	wire [WIDTH-1:0] wire_d69_0;
	wire [WIDTH-1:0] wire_d69_1;
	wire [WIDTH-1:0] wire_d69_2;
	wire [WIDTH-1:0] wire_d69_3;
	wire [WIDTH-1:0] wire_d69_4;
	wire [WIDTH-1:0] wire_d69_5;
	wire [WIDTH-1:0] wire_d69_6;
	wire [WIDTH-1:0] wire_d69_7;
	wire [WIDTH-1:0] wire_d69_8;
	wire [WIDTH-1:0] wire_d69_9;
	wire [WIDTH-1:0] wire_d69_10;
	wire [WIDTH-1:0] wire_d69_11;
	wire [WIDTH-1:0] wire_d69_12;
	wire [WIDTH-1:0] wire_d69_13;
	wire [WIDTH-1:0] wire_d69_14;
	wire [WIDTH-1:0] wire_d69_15;
	wire [WIDTH-1:0] wire_d69_16;
	wire [WIDTH-1:0] wire_d69_17;
	wire [WIDTH-1:0] wire_d69_18;
	wire [WIDTH-1:0] wire_d69_19;
	wire [WIDTH-1:0] wire_d69_20;
	wire [WIDTH-1:0] wire_d69_21;
	wire [WIDTH-1:0] wire_d69_22;
	wire [WIDTH-1:0] wire_d69_23;
	wire [WIDTH-1:0] wire_d69_24;
	wire [WIDTH-1:0] wire_d69_25;
	wire [WIDTH-1:0] wire_d69_26;
	wire [WIDTH-1:0] wire_d69_27;
	wire [WIDTH-1:0] wire_d69_28;
	wire [WIDTH-1:0] wire_d69_29;
	wire [WIDTH-1:0] wire_d69_30;
	wire [WIDTH-1:0] wire_d69_31;
	wire [WIDTH-1:0] wire_d69_32;
	wire [WIDTH-1:0] wire_d69_33;
	wire [WIDTH-1:0] wire_d69_34;
	wire [WIDTH-1:0] wire_d69_35;
	wire [WIDTH-1:0] wire_d69_36;
	wire [WIDTH-1:0] wire_d69_37;
	wire [WIDTH-1:0] wire_d69_38;
	wire [WIDTH-1:0] wire_d69_39;
	wire [WIDTH-1:0] wire_d69_40;
	wire [WIDTH-1:0] wire_d69_41;
	wire [WIDTH-1:0] wire_d69_42;
	wire [WIDTH-1:0] wire_d69_43;
	wire [WIDTH-1:0] wire_d69_44;
	wire [WIDTH-1:0] wire_d69_45;
	wire [WIDTH-1:0] wire_d69_46;
	wire [WIDTH-1:0] wire_d69_47;
	wire [WIDTH-1:0] wire_d69_48;
	wire [WIDTH-1:0] wire_d69_49;
	wire [WIDTH-1:0] wire_d69_50;
	wire [WIDTH-1:0] wire_d69_51;
	wire [WIDTH-1:0] wire_d69_52;
	wire [WIDTH-1:0] wire_d69_53;
	wire [WIDTH-1:0] wire_d69_54;
	wire [WIDTH-1:0] wire_d69_55;
	wire [WIDTH-1:0] wire_d69_56;
	wire [WIDTH-1:0] wire_d69_57;
	wire [WIDTH-1:0] wire_d69_58;
	wire [WIDTH-1:0] wire_d69_59;
	wire [WIDTH-1:0] wire_d69_60;
	wire [WIDTH-1:0] wire_d69_61;
	wire [WIDTH-1:0] wire_d69_62;
	wire [WIDTH-1:0] wire_d69_63;
	wire [WIDTH-1:0] wire_d69_64;
	wire [WIDTH-1:0] wire_d69_65;
	wire [WIDTH-1:0] wire_d69_66;
	wire [WIDTH-1:0] wire_d69_67;
	wire [WIDTH-1:0] wire_d69_68;
	wire [WIDTH-1:0] wire_d69_69;
	wire [WIDTH-1:0] wire_d69_70;
	wire [WIDTH-1:0] wire_d69_71;
	wire [WIDTH-1:0] wire_d69_72;
	wire [WIDTH-1:0] wire_d69_73;
	wire [WIDTH-1:0] wire_d69_74;
	wire [WIDTH-1:0] wire_d69_75;
	wire [WIDTH-1:0] wire_d69_76;
	wire [WIDTH-1:0] wire_d69_77;
	wire [WIDTH-1:0] wire_d69_78;
	wire [WIDTH-1:0] wire_d70_0;
	wire [WIDTH-1:0] wire_d70_1;
	wire [WIDTH-1:0] wire_d70_2;
	wire [WIDTH-1:0] wire_d70_3;
	wire [WIDTH-1:0] wire_d70_4;
	wire [WIDTH-1:0] wire_d70_5;
	wire [WIDTH-1:0] wire_d70_6;
	wire [WIDTH-1:0] wire_d70_7;
	wire [WIDTH-1:0] wire_d70_8;
	wire [WIDTH-1:0] wire_d70_9;
	wire [WIDTH-1:0] wire_d70_10;
	wire [WIDTH-1:0] wire_d70_11;
	wire [WIDTH-1:0] wire_d70_12;
	wire [WIDTH-1:0] wire_d70_13;
	wire [WIDTH-1:0] wire_d70_14;
	wire [WIDTH-1:0] wire_d70_15;
	wire [WIDTH-1:0] wire_d70_16;
	wire [WIDTH-1:0] wire_d70_17;
	wire [WIDTH-1:0] wire_d70_18;
	wire [WIDTH-1:0] wire_d70_19;
	wire [WIDTH-1:0] wire_d70_20;
	wire [WIDTH-1:0] wire_d70_21;
	wire [WIDTH-1:0] wire_d70_22;
	wire [WIDTH-1:0] wire_d70_23;
	wire [WIDTH-1:0] wire_d70_24;
	wire [WIDTH-1:0] wire_d70_25;
	wire [WIDTH-1:0] wire_d70_26;
	wire [WIDTH-1:0] wire_d70_27;
	wire [WIDTH-1:0] wire_d70_28;
	wire [WIDTH-1:0] wire_d70_29;
	wire [WIDTH-1:0] wire_d70_30;
	wire [WIDTH-1:0] wire_d70_31;
	wire [WIDTH-1:0] wire_d70_32;
	wire [WIDTH-1:0] wire_d70_33;
	wire [WIDTH-1:0] wire_d70_34;
	wire [WIDTH-1:0] wire_d70_35;
	wire [WIDTH-1:0] wire_d70_36;
	wire [WIDTH-1:0] wire_d70_37;
	wire [WIDTH-1:0] wire_d70_38;
	wire [WIDTH-1:0] wire_d70_39;
	wire [WIDTH-1:0] wire_d70_40;
	wire [WIDTH-1:0] wire_d70_41;
	wire [WIDTH-1:0] wire_d70_42;
	wire [WIDTH-1:0] wire_d70_43;
	wire [WIDTH-1:0] wire_d70_44;
	wire [WIDTH-1:0] wire_d70_45;
	wire [WIDTH-1:0] wire_d70_46;
	wire [WIDTH-1:0] wire_d70_47;
	wire [WIDTH-1:0] wire_d70_48;
	wire [WIDTH-1:0] wire_d70_49;
	wire [WIDTH-1:0] wire_d70_50;
	wire [WIDTH-1:0] wire_d70_51;
	wire [WIDTH-1:0] wire_d70_52;
	wire [WIDTH-1:0] wire_d70_53;
	wire [WIDTH-1:0] wire_d70_54;
	wire [WIDTH-1:0] wire_d70_55;
	wire [WIDTH-1:0] wire_d70_56;
	wire [WIDTH-1:0] wire_d70_57;
	wire [WIDTH-1:0] wire_d70_58;
	wire [WIDTH-1:0] wire_d70_59;
	wire [WIDTH-1:0] wire_d70_60;
	wire [WIDTH-1:0] wire_d70_61;
	wire [WIDTH-1:0] wire_d70_62;
	wire [WIDTH-1:0] wire_d70_63;
	wire [WIDTH-1:0] wire_d70_64;
	wire [WIDTH-1:0] wire_d70_65;
	wire [WIDTH-1:0] wire_d70_66;
	wire [WIDTH-1:0] wire_d70_67;
	wire [WIDTH-1:0] wire_d70_68;
	wire [WIDTH-1:0] wire_d70_69;
	wire [WIDTH-1:0] wire_d70_70;
	wire [WIDTH-1:0] wire_d70_71;
	wire [WIDTH-1:0] wire_d70_72;
	wire [WIDTH-1:0] wire_d70_73;
	wire [WIDTH-1:0] wire_d70_74;
	wire [WIDTH-1:0] wire_d70_75;
	wire [WIDTH-1:0] wire_d70_76;
	wire [WIDTH-1:0] wire_d70_77;
	wire [WIDTH-1:0] wire_d70_78;
	wire [WIDTH-1:0] wire_d71_0;
	wire [WIDTH-1:0] wire_d71_1;
	wire [WIDTH-1:0] wire_d71_2;
	wire [WIDTH-1:0] wire_d71_3;
	wire [WIDTH-1:0] wire_d71_4;
	wire [WIDTH-1:0] wire_d71_5;
	wire [WIDTH-1:0] wire_d71_6;
	wire [WIDTH-1:0] wire_d71_7;
	wire [WIDTH-1:0] wire_d71_8;
	wire [WIDTH-1:0] wire_d71_9;
	wire [WIDTH-1:0] wire_d71_10;
	wire [WIDTH-1:0] wire_d71_11;
	wire [WIDTH-1:0] wire_d71_12;
	wire [WIDTH-1:0] wire_d71_13;
	wire [WIDTH-1:0] wire_d71_14;
	wire [WIDTH-1:0] wire_d71_15;
	wire [WIDTH-1:0] wire_d71_16;
	wire [WIDTH-1:0] wire_d71_17;
	wire [WIDTH-1:0] wire_d71_18;
	wire [WIDTH-1:0] wire_d71_19;
	wire [WIDTH-1:0] wire_d71_20;
	wire [WIDTH-1:0] wire_d71_21;
	wire [WIDTH-1:0] wire_d71_22;
	wire [WIDTH-1:0] wire_d71_23;
	wire [WIDTH-1:0] wire_d71_24;
	wire [WIDTH-1:0] wire_d71_25;
	wire [WIDTH-1:0] wire_d71_26;
	wire [WIDTH-1:0] wire_d71_27;
	wire [WIDTH-1:0] wire_d71_28;
	wire [WIDTH-1:0] wire_d71_29;
	wire [WIDTH-1:0] wire_d71_30;
	wire [WIDTH-1:0] wire_d71_31;
	wire [WIDTH-1:0] wire_d71_32;
	wire [WIDTH-1:0] wire_d71_33;
	wire [WIDTH-1:0] wire_d71_34;
	wire [WIDTH-1:0] wire_d71_35;
	wire [WIDTH-1:0] wire_d71_36;
	wire [WIDTH-1:0] wire_d71_37;
	wire [WIDTH-1:0] wire_d71_38;
	wire [WIDTH-1:0] wire_d71_39;
	wire [WIDTH-1:0] wire_d71_40;
	wire [WIDTH-1:0] wire_d71_41;
	wire [WIDTH-1:0] wire_d71_42;
	wire [WIDTH-1:0] wire_d71_43;
	wire [WIDTH-1:0] wire_d71_44;
	wire [WIDTH-1:0] wire_d71_45;
	wire [WIDTH-1:0] wire_d71_46;
	wire [WIDTH-1:0] wire_d71_47;
	wire [WIDTH-1:0] wire_d71_48;
	wire [WIDTH-1:0] wire_d71_49;
	wire [WIDTH-1:0] wire_d71_50;
	wire [WIDTH-1:0] wire_d71_51;
	wire [WIDTH-1:0] wire_d71_52;
	wire [WIDTH-1:0] wire_d71_53;
	wire [WIDTH-1:0] wire_d71_54;
	wire [WIDTH-1:0] wire_d71_55;
	wire [WIDTH-1:0] wire_d71_56;
	wire [WIDTH-1:0] wire_d71_57;
	wire [WIDTH-1:0] wire_d71_58;
	wire [WIDTH-1:0] wire_d71_59;
	wire [WIDTH-1:0] wire_d71_60;
	wire [WIDTH-1:0] wire_d71_61;
	wire [WIDTH-1:0] wire_d71_62;
	wire [WIDTH-1:0] wire_d71_63;
	wire [WIDTH-1:0] wire_d71_64;
	wire [WIDTH-1:0] wire_d71_65;
	wire [WIDTH-1:0] wire_d71_66;
	wire [WIDTH-1:0] wire_d71_67;
	wire [WIDTH-1:0] wire_d71_68;
	wire [WIDTH-1:0] wire_d71_69;
	wire [WIDTH-1:0] wire_d71_70;
	wire [WIDTH-1:0] wire_d71_71;
	wire [WIDTH-1:0] wire_d71_72;
	wire [WIDTH-1:0] wire_d71_73;
	wire [WIDTH-1:0] wire_d71_74;
	wire [WIDTH-1:0] wire_d71_75;
	wire [WIDTH-1:0] wire_d71_76;
	wire [WIDTH-1:0] wire_d71_77;
	wire [WIDTH-1:0] wire_d71_78;
	wire [WIDTH-1:0] wire_d72_0;
	wire [WIDTH-1:0] wire_d72_1;
	wire [WIDTH-1:0] wire_d72_2;
	wire [WIDTH-1:0] wire_d72_3;
	wire [WIDTH-1:0] wire_d72_4;
	wire [WIDTH-1:0] wire_d72_5;
	wire [WIDTH-1:0] wire_d72_6;
	wire [WIDTH-1:0] wire_d72_7;
	wire [WIDTH-1:0] wire_d72_8;
	wire [WIDTH-1:0] wire_d72_9;
	wire [WIDTH-1:0] wire_d72_10;
	wire [WIDTH-1:0] wire_d72_11;
	wire [WIDTH-1:0] wire_d72_12;
	wire [WIDTH-1:0] wire_d72_13;
	wire [WIDTH-1:0] wire_d72_14;
	wire [WIDTH-1:0] wire_d72_15;
	wire [WIDTH-1:0] wire_d72_16;
	wire [WIDTH-1:0] wire_d72_17;
	wire [WIDTH-1:0] wire_d72_18;
	wire [WIDTH-1:0] wire_d72_19;
	wire [WIDTH-1:0] wire_d72_20;
	wire [WIDTH-1:0] wire_d72_21;
	wire [WIDTH-1:0] wire_d72_22;
	wire [WIDTH-1:0] wire_d72_23;
	wire [WIDTH-1:0] wire_d72_24;
	wire [WIDTH-1:0] wire_d72_25;
	wire [WIDTH-1:0] wire_d72_26;
	wire [WIDTH-1:0] wire_d72_27;
	wire [WIDTH-1:0] wire_d72_28;
	wire [WIDTH-1:0] wire_d72_29;
	wire [WIDTH-1:0] wire_d72_30;
	wire [WIDTH-1:0] wire_d72_31;
	wire [WIDTH-1:0] wire_d72_32;
	wire [WIDTH-1:0] wire_d72_33;
	wire [WIDTH-1:0] wire_d72_34;
	wire [WIDTH-1:0] wire_d72_35;
	wire [WIDTH-1:0] wire_d72_36;
	wire [WIDTH-1:0] wire_d72_37;
	wire [WIDTH-1:0] wire_d72_38;
	wire [WIDTH-1:0] wire_d72_39;
	wire [WIDTH-1:0] wire_d72_40;
	wire [WIDTH-1:0] wire_d72_41;
	wire [WIDTH-1:0] wire_d72_42;
	wire [WIDTH-1:0] wire_d72_43;
	wire [WIDTH-1:0] wire_d72_44;
	wire [WIDTH-1:0] wire_d72_45;
	wire [WIDTH-1:0] wire_d72_46;
	wire [WIDTH-1:0] wire_d72_47;
	wire [WIDTH-1:0] wire_d72_48;
	wire [WIDTH-1:0] wire_d72_49;
	wire [WIDTH-1:0] wire_d72_50;
	wire [WIDTH-1:0] wire_d72_51;
	wire [WIDTH-1:0] wire_d72_52;
	wire [WIDTH-1:0] wire_d72_53;
	wire [WIDTH-1:0] wire_d72_54;
	wire [WIDTH-1:0] wire_d72_55;
	wire [WIDTH-1:0] wire_d72_56;
	wire [WIDTH-1:0] wire_d72_57;
	wire [WIDTH-1:0] wire_d72_58;
	wire [WIDTH-1:0] wire_d72_59;
	wire [WIDTH-1:0] wire_d72_60;
	wire [WIDTH-1:0] wire_d72_61;
	wire [WIDTH-1:0] wire_d72_62;
	wire [WIDTH-1:0] wire_d72_63;
	wire [WIDTH-1:0] wire_d72_64;
	wire [WIDTH-1:0] wire_d72_65;
	wire [WIDTH-1:0] wire_d72_66;
	wire [WIDTH-1:0] wire_d72_67;
	wire [WIDTH-1:0] wire_d72_68;
	wire [WIDTH-1:0] wire_d72_69;
	wire [WIDTH-1:0] wire_d72_70;
	wire [WIDTH-1:0] wire_d72_71;
	wire [WIDTH-1:0] wire_d72_72;
	wire [WIDTH-1:0] wire_d72_73;
	wire [WIDTH-1:0] wire_d72_74;
	wire [WIDTH-1:0] wire_d72_75;
	wire [WIDTH-1:0] wire_d72_76;
	wire [WIDTH-1:0] wire_d72_77;
	wire [WIDTH-1:0] wire_d72_78;
	wire [WIDTH-1:0] wire_d73_0;
	wire [WIDTH-1:0] wire_d73_1;
	wire [WIDTH-1:0] wire_d73_2;
	wire [WIDTH-1:0] wire_d73_3;
	wire [WIDTH-1:0] wire_d73_4;
	wire [WIDTH-1:0] wire_d73_5;
	wire [WIDTH-1:0] wire_d73_6;
	wire [WIDTH-1:0] wire_d73_7;
	wire [WIDTH-1:0] wire_d73_8;
	wire [WIDTH-1:0] wire_d73_9;
	wire [WIDTH-1:0] wire_d73_10;
	wire [WIDTH-1:0] wire_d73_11;
	wire [WIDTH-1:0] wire_d73_12;
	wire [WIDTH-1:0] wire_d73_13;
	wire [WIDTH-1:0] wire_d73_14;
	wire [WIDTH-1:0] wire_d73_15;
	wire [WIDTH-1:0] wire_d73_16;
	wire [WIDTH-1:0] wire_d73_17;
	wire [WIDTH-1:0] wire_d73_18;
	wire [WIDTH-1:0] wire_d73_19;
	wire [WIDTH-1:0] wire_d73_20;
	wire [WIDTH-1:0] wire_d73_21;
	wire [WIDTH-1:0] wire_d73_22;
	wire [WIDTH-1:0] wire_d73_23;
	wire [WIDTH-1:0] wire_d73_24;
	wire [WIDTH-1:0] wire_d73_25;
	wire [WIDTH-1:0] wire_d73_26;
	wire [WIDTH-1:0] wire_d73_27;
	wire [WIDTH-1:0] wire_d73_28;
	wire [WIDTH-1:0] wire_d73_29;
	wire [WIDTH-1:0] wire_d73_30;
	wire [WIDTH-1:0] wire_d73_31;
	wire [WIDTH-1:0] wire_d73_32;
	wire [WIDTH-1:0] wire_d73_33;
	wire [WIDTH-1:0] wire_d73_34;
	wire [WIDTH-1:0] wire_d73_35;
	wire [WIDTH-1:0] wire_d73_36;
	wire [WIDTH-1:0] wire_d73_37;
	wire [WIDTH-1:0] wire_d73_38;
	wire [WIDTH-1:0] wire_d73_39;
	wire [WIDTH-1:0] wire_d73_40;
	wire [WIDTH-1:0] wire_d73_41;
	wire [WIDTH-1:0] wire_d73_42;
	wire [WIDTH-1:0] wire_d73_43;
	wire [WIDTH-1:0] wire_d73_44;
	wire [WIDTH-1:0] wire_d73_45;
	wire [WIDTH-1:0] wire_d73_46;
	wire [WIDTH-1:0] wire_d73_47;
	wire [WIDTH-1:0] wire_d73_48;
	wire [WIDTH-1:0] wire_d73_49;
	wire [WIDTH-1:0] wire_d73_50;
	wire [WIDTH-1:0] wire_d73_51;
	wire [WIDTH-1:0] wire_d73_52;
	wire [WIDTH-1:0] wire_d73_53;
	wire [WIDTH-1:0] wire_d73_54;
	wire [WIDTH-1:0] wire_d73_55;
	wire [WIDTH-1:0] wire_d73_56;
	wire [WIDTH-1:0] wire_d73_57;
	wire [WIDTH-1:0] wire_d73_58;
	wire [WIDTH-1:0] wire_d73_59;
	wire [WIDTH-1:0] wire_d73_60;
	wire [WIDTH-1:0] wire_d73_61;
	wire [WIDTH-1:0] wire_d73_62;
	wire [WIDTH-1:0] wire_d73_63;
	wire [WIDTH-1:0] wire_d73_64;
	wire [WIDTH-1:0] wire_d73_65;
	wire [WIDTH-1:0] wire_d73_66;
	wire [WIDTH-1:0] wire_d73_67;
	wire [WIDTH-1:0] wire_d73_68;
	wire [WIDTH-1:0] wire_d73_69;
	wire [WIDTH-1:0] wire_d73_70;
	wire [WIDTH-1:0] wire_d73_71;
	wire [WIDTH-1:0] wire_d73_72;
	wire [WIDTH-1:0] wire_d73_73;
	wire [WIDTH-1:0] wire_d73_74;
	wire [WIDTH-1:0] wire_d73_75;
	wire [WIDTH-1:0] wire_d73_76;
	wire [WIDTH-1:0] wire_d73_77;
	wire [WIDTH-1:0] wire_d73_78;
	wire [WIDTH-1:0] wire_d74_0;
	wire [WIDTH-1:0] wire_d74_1;
	wire [WIDTH-1:0] wire_d74_2;
	wire [WIDTH-1:0] wire_d74_3;
	wire [WIDTH-1:0] wire_d74_4;
	wire [WIDTH-1:0] wire_d74_5;
	wire [WIDTH-1:0] wire_d74_6;
	wire [WIDTH-1:0] wire_d74_7;
	wire [WIDTH-1:0] wire_d74_8;
	wire [WIDTH-1:0] wire_d74_9;
	wire [WIDTH-1:0] wire_d74_10;
	wire [WIDTH-1:0] wire_d74_11;
	wire [WIDTH-1:0] wire_d74_12;
	wire [WIDTH-1:0] wire_d74_13;
	wire [WIDTH-1:0] wire_d74_14;
	wire [WIDTH-1:0] wire_d74_15;
	wire [WIDTH-1:0] wire_d74_16;
	wire [WIDTH-1:0] wire_d74_17;
	wire [WIDTH-1:0] wire_d74_18;
	wire [WIDTH-1:0] wire_d74_19;
	wire [WIDTH-1:0] wire_d74_20;
	wire [WIDTH-1:0] wire_d74_21;
	wire [WIDTH-1:0] wire_d74_22;
	wire [WIDTH-1:0] wire_d74_23;
	wire [WIDTH-1:0] wire_d74_24;
	wire [WIDTH-1:0] wire_d74_25;
	wire [WIDTH-1:0] wire_d74_26;
	wire [WIDTH-1:0] wire_d74_27;
	wire [WIDTH-1:0] wire_d74_28;
	wire [WIDTH-1:0] wire_d74_29;
	wire [WIDTH-1:0] wire_d74_30;
	wire [WIDTH-1:0] wire_d74_31;
	wire [WIDTH-1:0] wire_d74_32;
	wire [WIDTH-1:0] wire_d74_33;
	wire [WIDTH-1:0] wire_d74_34;
	wire [WIDTH-1:0] wire_d74_35;
	wire [WIDTH-1:0] wire_d74_36;
	wire [WIDTH-1:0] wire_d74_37;
	wire [WIDTH-1:0] wire_d74_38;
	wire [WIDTH-1:0] wire_d74_39;
	wire [WIDTH-1:0] wire_d74_40;
	wire [WIDTH-1:0] wire_d74_41;
	wire [WIDTH-1:0] wire_d74_42;
	wire [WIDTH-1:0] wire_d74_43;
	wire [WIDTH-1:0] wire_d74_44;
	wire [WIDTH-1:0] wire_d74_45;
	wire [WIDTH-1:0] wire_d74_46;
	wire [WIDTH-1:0] wire_d74_47;
	wire [WIDTH-1:0] wire_d74_48;
	wire [WIDTH-1:0] wire_d74_49;
	wire [WIDTH-1:0] wire_d74_50;
	wire [WIDTH-1:0] wire_d74_51;
	wire [WIDTH-1:0] wire_d74_52;
	wire [WIDTH-1:0] wire_d74_53;
	wire [WIDTH-1:0] wire_d74_54;
	wire [WIDTH-1:0] wire_d74_55;
	wire [WIDTH-1:0] wire_d74_56;
	wire [WIDTH-1:0] wire_d74_57;
	wire [WIDTH-1:0] wire_d74_58;
	wire [WIDTH-1:0] wire_d74_59;
	wire [WIDTH-1:0] wire_d74_60;
	wire [WIDTH-1:0] wire_d74_61;
	wire [WIDTH-1:0] wire_d74_62;
	wire [WIDTH-1:0] wire_d74_63;
	wire [WIDTH-1:0] wire_d74_64;
	wire [WIDTH-1:0] wire_d74_65;
	wire [WIDTH-1:0] wire_d74_66;
	wire [WIDTH-1:0] wire_d74_67;
	wire [WIDTH-1:0] wire_d74_68;
	wire [WIDTH-1:0] wire_d74_69;
	wire [WIDTH-1:0] wire_d74_70;
	wire [WIDTH-1:0] wire_d74_71;
	wire [WIDTH-1:0] wire_d74_72;
	wire [WIDTH-1:0] wire_d74_73;
	wire [WIDTH-1:0] wire_d74_74;
	wire [WIDTH-1:0] wire_d74_75;
	wire [WIDTH-1:0] wire_d74_76;
	wire [WIDTH-1:0] wire_d74_77;
	wire [WIDTH-1:0] wire_d74_78;
	wire [WIDTH-1:0] wire_d75_0;
	wire [WIDTH-1:0] wire_d75_1;
	wire [WIDTH-1:0] wire_d75_2;
	wire [WIDTH-1:0] wire_d75_3;
	wire [WIDTH-1:0] wire_d75_4;
	wire [WIDTH-1:0] wire_d75_5;
	wire [WIDTH-1:0] wire_d75_6;
	wire [WIDTH-1:0] wire_d75_7;
	wire [WIDTH-1:0] wire_d75_8;
	wire [WIDTH-1:0] wire_d75_9;
	wire [WIDTH-1:0] wire_d75_10;
	wire [WIDTH-1:0] wire_d75_11;
	wire [WIDTH-1:0] wire_d75_12;
	wire [WIDTH-1:0] wire_d75_13;
	wire [WIDTH-1:0] wire_d75_14;
	wire [WIDTH-1:0] wire_d75_15;
	wire [WIDTH-1:0] wire_d75_16;
	wire [WIDTH-1:0] wire_d75_17;
	wire [WIDTH-1:0] wire_d75_18;
	wire [WIDTH-1:0] wire_d75_19;
	wire [WIDTH-1:0] wire_d75_20;
	wire [WIDTH-1:0] wire_d75_21;
	wire [WIDTH-1:0] wire_d75_22;
	wire [WIDTH-1:0] wire_d75_23;
	wire [WIDTH-1:0] wire_d75_24;
	wire [WIDTH-1:0] wire_d75_25;
	wire [WIDTH-1:0] wire_d75_26;
	wire [WIDTH-1:0] wire_d75_27;
	wire [WIDTH-1:0] wire_d75_28;
	wire [WIDTH-1:0] wire_d75_29;
	wire [WIDTH-1:0] wire_d75_30;
	wire [WIDTH-1:0] wire_d75_31;
	wire [WIDTH-1:0] wire_d75_32;
	wire [WIDTH-1:0] wire_d75_33;
	wire [WIDTH-1:0] wire_d75_34;
	wire [WIDTH-1:0] wire_d75_35;
	wire [WIDTH-1:0] wire_d75_36;
	wire [WIDTH-1:0] wire_d75_37;
	wire [WIDTH-1:0] wire_d75_38;
	wire [WIDTH-1:0] wire_d75_39;
	wire [WIDTH-1:0] wire_d75_40;
	wire [WIDTH-1:0] wire_d75_41;
	wire [WIDTH-1:0] wire_d75_42;
	wire [WIDTH-1:0] wire_d75_43;
	wire [WIDTH-1:0] wire_d75_44;
	wire [WIDTH-1:0] wire_d75_45;
	wire [WIDTH-1:0] wire_d75_46;
	wire [WIDTH-1:0] wire_d75_47;
	wire [WIDTH-1:0] wire_d75_48;
	wire [WIDTH-1:0] wire_d75_49;
	wire [WIDTH-1:0] wire_d75_50;
	wire [WIDTH-1:0] wire_d75_51;
	wire [WIDTH-1:0] wire_d75_52;
	wire [WIDTH-1:0] wire_d75_53;
	wire [WIDTH-1:0] wire_d75_54;
	wire [WIDTH-1:0] wire_d75_55;
	wire [WIDTH-1:0] wire_d75_56;
	wire [WIDTH-1:0] wire_d75_57;
	wire [WIDTH-1:0] wire_d75_58;
	wire [WIDTH-1:0] wire_d75_59;
	wire [WIDTH-1:0] wire_d75_60;
	wire [WIDTH-1:0] wire_d75_61;
	wire [WIDTH-1:0] wire_d75_62;
	wire [WIDTH-1:0] wire_d75_63;
	wire [WIDTH-1:0] wire_d75_64;
	wire [WIDTH-1:0] wire_d75_65;
	wire [WIDTH-1:0] wire_d75_66;
	wire [WIDTH-1:0] wire_d75_67;
	wire [WIDTH-1:0] wire_d75_68;
	wire [WIDTH-1:0] wire_d75_69;
	wire [WIDTH-1:0] wire_d75_70;
	wire [WIDTH-1:0] wire_d75_71;
	wire [WIDTH-1:0] wire_d75_72;
	wire [WIDTH-1:0] wire_d75_73;
	wire [WIDTH-1:0] wire_d75_74;
	wire [WIDTH-1:0] wire_d75_75;
	wire [WIDTH-1:0] wire_d75_76;
	wire [WIDTH-1:0] wire_d75_77;
	wire [WIDTH-1:0] wire_d75_78;
	wire [WIDTH-1:0] wire_d76_0;
	wire [WIDTH-1:0] wire_d76_1;
	wire [WIDTH-1:0] wire_d76_2;
	wire [WIDTH-1:0] wire_d76_3;
	wire [WIDTH-1:0] wire_d76_4;
	wire [WIDTH-1:0] wire_d76_5;
	wire [WIDTH-1:0] wire_d76_6;
	wire [WIDTH-1:0] wire_d76_7;
	wire [WIDTH-1:0] wire_d76_8;
	wire [WIDTH-1:0] wire_d76_9;
	wire [WIDTH-1:0] wire_d76_10;
	wire [WIDTH-1:0] wire_d76_11;
	wire [WIDTH-1:0] wire_d76_12;
	wire [WIDTH-1:0] wire_d76_13;
	wire [WIDTH-1:0] wire_d76_14;
	wire [WIDTH-1:0] wire_d76_15;
	wire [WIDTH-1:0] wire_d76_16;
	wire [WIDTH-1:0] wire_d76_17;
	wire [WIDTH-1:0] wire_d76_18;
	wire [WIDTH-1:0] wire_d76_19;
	wire [WIDTH-1:0] wire_d76_20;
	wire [WIDTH-1:0] wire_d76_21;
	wire [WIDTH-1:0] wire_d76_22;
	wire [WIDTH-1:0] wire_d76_23;
	wire [WIDTH-1:0] wire_d76_24;
	wire [WIDTH-1:0] wire_d76_25;
	wire [WIDTH-1:0] wire_d76_26;
	wire [WIDTH-1:0] wire_d76_27;
	wire [WIDTH-1:0] wire_d76_28;
	wire [WIDTH-1:0] wire_d76_29;
	wire [WIDTH-1:0] wire_d76_30;
	wire [WIDTH-1:0] wire_d76_31;
	wire [WIDTH-1:0] wire_d76_32;
	wire [WIDTH-1:0] wire_d76_33;
	wire [WIDTH-1:0] wire_d76_34;
	wire [WIDTH-1:0] wire_d76_35;
	wire [WIDTH-1:0] wire_d76_36;
	wire [WIDTH-1:0] wire_d76_37;
	wire [WIDTH-1:0] wire_d76_38;
	wire [WIDTH-1:0] wire_d76_39;
	wire [WIDTH-1:0] wire_d76_40;
	wire [WIDTH-1:0] wire_d76_41;
	wire [WIDTH-1:0] wire_d76_42;
	wire [WIDTH-1:0] wire_d76_43;
	wire [WIDTH-1:0] wire_d76_44;
	wire [WIDTH-1:0] wire_d76_45;
	wire [WIDTH-1:0] wire_d76_46;
	wire [WIDTH-1:0] wire_d76_47;
	wire [WIDTH-1:0] wire_d76_48;
	wire [WIDTH-1:0] wire_d76_49;
	wire [WIDTH-1:0] wire_d76_50;
	wire [WIDTH-1:0] wire_d76_51;
	wire [WIDTH-1:0] wire_d76_52;
	wire [WIDTH-1:0] wire_d76_53;
	wire [WIDTH-1:0] wire_d76_54;
	wire [WIDTH-1:0] wire_d76_55;
	wire [WIDTH-1:0] wire_d76_56;
	wire [WIDTH-1:0] wire_d76_57;
	wire [WIDTH-1:0] wire_d76_58;
	wire [WIDTH-1:0] wire_d76_59;
	wire [WIDTH-1:0] wire_d76_60;
	wire [WIDTH-1:0] wire_d76_61;
	wire [WIDTH-1:0] wire_d76_62;
	wire [WIDTH-1:0] wire_d76_63;
	wire [WIDTH-1:0] wire_d76_64;
	wire [WIDTH-1:0] wire_d76_65;
	wire [WIDTH-1:0] wire_d76_66;
	wire [WIDTH-1:0] wire_d76_67;
	wire [WIDTH-1:0] wire_d76_68;
	wire [WIDTH-1:0] wire_d76_69;
	wire [WIDTH-1:0] wire_d76_70;
	wire [WIDTH-1:0] wire_d76_71;
	wire [WIDTH-1:0] wire_d76_72;
	wire [WIDTH-1:0] wire_d76_73;
	wire [WIDTH-1:0] wire_d76_74;
	wire [WIDTH-1:0] wire_d76_75;
	wire [WIDTH-1:0] wire_d76_76;
	wire [WIDTH-1:0] wire_d76_77;
	wire [WIDTH-1:0] wire_d76_78;
	wire [WIDTH-1:0] wire_d77_0;
	wire [WIDTH-1:0] wire_d77_1;
	wire [WIDTH-1:0] wire_d77_2;
	wire [WIDTH-1:0] wire_d77_3;
	wire [WIDTH-1:0] wire_d77_4;
	wire [WIDTH-1:0] wire_d77_5;
	wire [WIDTH-1:0] wire_d77_6;
	wire [WIDTH-1:0] wire_d77_7;
	wire [WIDTH-1:0] wire_d77_8;
	wire [WIDTH-1:0] wire_d77_9;
	wire [WIDTH-1:0] wire_d77_10;
	wire [WIDTH-1:0] wire_d77_11;
	wire [WIDTH-1:0] wire_d77_12;
	wire [WIDTH-1:0] wire_d77_13;
	wire [WIDTH-1:0] wire_d77_14;
	wire [WIDTH-1:0] wire_d77_15;
	wire [WIDTH-1:0] wire_d77_16;
	wire [WIDTH-1:0] wire_d77_17;
	wire [WIDTH-1:0] wire_d77_18;
	wire [WIDTH-1:0] wire_d77_19;
	wire [WIDTH-1:0] wire_d77_20;
	wire [WIDTH-1:0] wire_d77_21;
	wire [WIDTH-1:0] wire_d77_22;
	wire [WIDTH-1:0] wire_d77_23;
	wire [WIDTH-1:0] wire_d77_24;
	wire [WIDTH-1:0] wire_d77_25;
	wire [WIDTH-1:0] wire_d77_26;
	wire [WIDTH-1:0] wire_d77_27;
	wire [WIDTH-1:0] wire_d77_28;
	wire [WIDTH-1:0] wire_d77_29;
	wire [WIDTH-1:0] wire_d77_30;
	wire [WIDTH-1:0] wire_d77_31;
	wire [WIDTH-1:0] wire_d77_32;
	wire [WIDTH-1:0] wire_d77_33;
	wire [WIDTH-1:0] wire_d77_34;
	wire [WIDTH-1:0] wire_d77_35;
	wire [WIDTH-1:0] wire_d77_36;
	wire [WIDTH-1:0] wire_d77_37;
	wire [WIDTH-1:0] wire_d77_38;
	wire [WIDTH-1:0] wire_d77_39;
	wire [WIDTH-1:0] wire_d77_40;
	wire [WIDTH-1:0] wire_d77_41;
	wire [WIDTH-1:0] wire_d77_42;
	wire [WIDTH-1:0] wire_d77_43;
	wire [WIDTH-1:0] wire_d77_44;
	wire [WIDTH-1:0] wire_d77_45;
	wire [WIDTH-1:0] wire_d77_46;
	wire [WIDTH-1:0] wire_d77_47;
	wire [WIDTH-1:0] wire_d77_48;
	wire [WIDTH-1:0] wire_d77_49;
	wire [WIDTH-1:0] wire_d77_50;
	wire [WIDTH-1:0] wire_d77_51;
	wire [WIDTH-1:0] wire_d77_52;
	wire [WIDTH-1:0] wire_d77_53;
	wire [WIDTH-1:0] wire_d77_54;
	wire [WIDTH-1:0] wire_d77_55;
	wire [WIDTH-1:0] wire_d77_56;
	wire [WIDTH-1:0] wire_d77_57;
	wire [WIDTH-1:0] wire_d77_58;
	wire [WIDTH-1:0] wire_d77_59;
	wire [WIDTH-1:0] wire_d77_60;
	wire [WIDTH-1:0] wire_d77_61;
	wire [WIDTH-1:0] wire_d77_62;
	wire [WIDTH-1:0] wire_d77_63;
	wire [WIDTH-1:0] wire_d77_64;
	wire [WIDTH-1:0] wire_d77_65;
	wire [WIDTH-1:0] wire_d77_66;
	wire [WIDTH-1:0] wire_d77_67;
	wire [WIDTH-1:0] wire_d77_68;
	wire [WIDTH-1:0] wire_d77_69;
	wire [WIDTH-1:0] wire_d77_70;
	wire [WIDTH-1:0] wire_d77_71;
	wire [WIDTH-1:0] wire_d77_72;
	wire [WIDTH-1:0] wire_d77_73;
	wire [WIDTH-1:0] wire_d77_74;
	wire [WIDTH-1:0] wire_d77_75;
	wire [WIDTH-1:0] wire_d77_76;
	wire [WIDTH-1:0] wire_d77_77;
	wire [WIDTH-1:0] wire_d77_78;
	wire [WIDTH-1:0] wire_d78_0;
	wire [WIDTH-1:0] wire_d78_1;
	wire [WIDTH-1:0] wire_d78_2;
	wire [WIDTH-1:0] wire_d78_3;
	wire [WIDTH-1:0] wire_d78_4;
	wire [WIDTH-1:0] wire_d78_5;
	wire [WIDTH-1:0] wire_d78_6;
	wire [WIDTH-1:0] wire_d78_7;
	wire [WIDTH-1:0] wire_d78_8;
	wire [WIDTH-1:0] wire_d78_9;
	wire [WIDTH-1:0] wire_d78_10;
	wire [WIDTH-1:0] wire_d78_11;
	wire [WIDTH-1:0] wire_d78_12;
	wire [WIDTH-1:0] wire_d78_13;
	wire [WIDTH-1:0] wire_d78_14;
	wire [WIDTH-1:0] wire_d78_15;
	wire [WIDTH-1:0] wire_d78_16;
	wire [WIDTH-1:0] wire_d78_17;
	wire [WIDTH-1:0] wire_d78_18;
	wire [WIDTH-1:0] wire_d78_19;
	wire [WIDTH-1:0] wire_d78_20;
	wire [WIDTH-1:0] wire_d78_21;
	wire [WIDTH-1:0] wire_d78_22;
	wire [WIDTH-1:0] wire_d78_23;
	wire [WIDTH-1:0] wire_d78_24;
	wire [WIDTH-1:0] wire_d78_25;
	wire [WIDTH-1:0] wire_d78_26;
	wire [WIDTH-1:0] wire_d78_27;
	wire [WIDTH-1:0] wire_d78_28;
	wire [WIDTH-1:0] wire_d78_29;
	wire [WIDTH-1:0] wire_d78_30;
	wire [WIDTH-1:0] wire_d78_31;
	wire [WIDTH-1:0] wire_d78_32;
	wire [WIDTH-1:0] wire_d78_33;
	wire [WIDTH-1:0] wire_d78_34;
	wire [WIDTH-1:0] wire_d78_35;
	wire [WIDTH-1:0] wire_d78_36;
	wire [WIDTH-1:0] wire_d78_37;
	wire [WIDTH-1:0] wire_d78_38;
	wire [WIDTH-1:0] wire_d78_39;
	wire [WIDTH-1:0] wire_d78_40;
	wire [WIDTH-1:0] wire_d78_41;
	wire [WIDTH-1:0] wire_d78_42;
	wire [WIDTH-1:0] wire_d78_43;
	wire [WIDTH-1:0] wire_d78_44;
	wire [WIDTH-1:0] wire_d78_45;
	wire [WIDTH-1:0] wire_d78_46;
	wire [WIDTH-1:0] wire_d78_47;
	wire [WIDTH-1:0] wire_d78_48;
	wire [WIDTH-1:0] wire_d78_49;
	wire [WIDTH-1:0] wire_d78_50;
	wire [WIDTH-1:0] wire_d78_51;
	wire [WIDTH-1:0] wire_d78_52;
	wire [WIDTH-1:0] wire_d78_53;
	wire [WIDTH-1:0] wire_d78_54;
	wire [WIDTH-1:0] wire_d78_55;
	wire [WIDTH-1:0] wire_d78_56;
	wire [WIDTH-1:0] wire_d78_57;
	wire [WIDTH-1:0] wire_d78_58;
	wire [WIDTH-1:0] wire_d78_59;
	wire [WIDTH-1:0] wire_d78_60;
	wire [WIDTH-1:0] wire_d78_61;
	wire [WIDTH-1:0] wire_d78_62;
	wire [WIDTH-1:0] wire_d78_63;
	wire [WIDTH-1:0] wire_d78_64;
	wire [WIDTH-1:0] wire_d78_65;
	wire [WIDTH-1:0] wire_d78_66;
	wire [WIDTH-1:0] wire_d78_67;
	wire [WIDTH-1:0] wire_d78_68;
	wire [WIDTH-1:0] wire_d78_69;
	wire [WIDTH-1:0] wire_d78_70;
	wire [WIDTH-1:0] wire_d78_71;
	wire [WIDTH-1:0] wire_d78_72;
	wire [WIDTH-1:0] wire_d78_73;
	wire [WIDTH-1:0] wire_d78_74;
	wire [WIDTH-1:0] wire_d78_75;
	wire [WIDTH-1:0] wire_d78_76;
	wire [WIDTH-1:0] wire_d78_77;
	wire [WIDTH-1:0] wire_d78_78;
	wire [WIDTH-1:0] wire_d79_0;
	wire [WIDTH-1:0] wire_d79_1;
	wire [WIDTH-1:0] wire_d79_2;
	wire [WIDTH-1:0] wire_d79_3;
	wire [WIDTH-1:0] wire_d79_4;
	wire [WIDTH-1:0] wire_d79_5;
	wire [WIDTH-1:0] wire_d79_6;
	wire [WIDTH-1:0] wire_d79_7;
	wire [WIDTH-1:0] wire_d79_8;
	wire [WIDTH-1:0] wire_d79_9;
	wire [WIDTH-1:0] wire_d79_10;
	wire [WIDTH-1:0] wire_d79_11;
	wire [WIDTH-1:0] wire_d79_12;
	wire [WIDTH-1:0] wire_d79_13;
	wire [WIDTH-1:0] wire_d79_14;
	wire [WIDTH-1:0] wire_d79_15;
	wire [WIDTH-1:0] wire_d79_16;
	wire [WIDTH-1:0] wire_d79_17;
	wire [WIDTH-1:0] wire_d79_18;
	wire [WIDTH-1:0] wire_d79_19;
	wire [WIDTH-1:0] wire_d79_20;
	wire [WIDTH-1:0] wire_d79_21;
	wire [WIDTH-1:0] wire_d79_22;
	wire [WIDTH-1:0] wire_d79_23;
	wire [WIDTH-1:0] wire_d79_24;
	wire [WIDTH-1:0] wire_d79_25;
	wire [WIDTH-1:0] wire_d79_26;
	wire [WIDTH-1:0] wire_d79_27;
	wire [WIDTH-1:0] wire_d79_28;
	wire [WIDTH-1:0] wire_d79_29;
	wire [WIDTH-1:0] wire_d79_30;
	wire [WIDTH-1:0] wire_d79_31;
	wire [WIDTH-1:0] wire_d79_32;
	wire [WIDTH-1:0] wire_d79_33;
	wire [WIDTH-1:0] wire_d79_34;
	wire [WIDTH-1:0] wire_d79_35;
	wire [WIDTH-1:0] wire_d79_36;
	wire [WIDTH-1:0] wire_d79_37;
	wire [WIDTH-1:0] wire_d79_38;
	wire [WIDTH-1:0] wire_d79_39;
	wire [WIDTH-1:0] wire_d79_40;
	wire [WIDTH-1:0] wire_d79_41;
	wire [WIDTH-1:0] wire_d79_42;
	wire [WIDTH-1:0] wire_d79_43;
	wire [WIDTH-1:0] wire_d79_44;
	wire [WIDTH-1:0] wire_d79_45;
	wire [WIDTH-1:0] wire_d79_46;
	wire [WIDTH-1:0] wire_d79_47;
	wire [WIDTH-1:0] wire_d79_48;
	wire [WIDTH-1:0] wire_d79_49;
	wire [WIDTH-1:0] wire_d79_50;
	wire [WIDTH-1:0] wire_d79_51;
	wire [WIDTH-1:0] wire_d79_52;
	wire [WIDTH-1:0] wire_d79_53;
	wire [WIDTH-1:0] wire_d79_54;
	wire [WIDTH-1:0] wire_d79_55;
	wire [WIDTH-1:0] wire_d79_56;
	wire [WIDTH-1:0] wire_d79_57;
	wire [WIDTH-1:0] wire_d79_58;
	wire [WIDTH-1:0] wire_d79_59;
	wire [WIDTH-1:0] wire_d79_60;
	wire [WIDTH-1:0] wire_d79_61;
	wire [WIDTH-1:0] wire_d79_62;
	wire [WIDTH-1:0] wire_d79_63;
	wire [WIDTH-1:0] wire_d79_64;
	wire [WIDTH-1:0] wire_d79_65;
	wire [WIDTH-1:0] wire_d79_66;
	wire [WIDTH-1:0] wire_d79_67;
	wire [WIDTH-1:0] wire_d79_68;
	wire [WIDTH-1:0] wire_d79_69;
	wire [WIDTH-1:0] wire_d79_70;
	wire [WIDTH-1:0] wire_d79_71;
	wire [WIDTH-1:0] wire_d79_72;
	wire [WIDTH-1:0] wire_d79_73;
	wire [WIDTH-1:0] wire_d79_74;
	wire [WIDTH-1:0] wire_d79_75;
	wire [WIDTH-1:0] wire_d79_76;
	wire [WIDTH-1:0] wire_d79_77;
	wire [WIDTH-1:0] wire_d79_78;
	wire [WIDTH-1:0] wire_d80_0;
	wire [WIDTH-1:0] wire_d80_1;
	wire [WIDTH-1:0] wire_d80_2;
	wire [WIDTH-1:0] wire_d80_3;
	wire [WIDTH-1:0] wire_d80_4;
	wire [WIDTH-1:0] wire_d80_5;
	wire [WIDTH-1:0] wire_d80_6;
	wire [WIDTH-1:0] wire_d80_7;
	wire [WIDTH-1:0] wire_d80_8;
	wire [WIDTH-1:0] wire_d80_9;
	wire [WIDTH-1:0] wire_d80_10;
	wire [WIDTH-1:0] wire_d80_11;
	wire [WIDTH-1:0] wire_d80_12;
	wire [WIDTH-1:0] wire_d80_13;
	wire [WIDTH-1:0] wire_d80_14;
	wire [WIDTH-1:0] wire_d80_15;
	wire [WIDTH-1:0] wire_d80_16;
	wire [WIDTH-1:0] wire_d80_17;
	wire [WIDTH-1:0] wire_d80_18;
	wire [WIDTH-1:0] wire_d80_19;
	wire [WIDTH-1:0] wire_d80_20;
	wire [WIDTH-1:0] wire_d80_21;
	wire [WIDTH-1:0] wire_d80_22;
	wire [WIDTH-1:0] wire_d80_23;
	wire [WIDTH-1:0] wire_d80_24;
	wire [WIDTH-1:0] wire_d80_25;
	wire [WIDTH-1:0] wire_d80_26;
	wire [WIDTH-1:0] wire_d80_27;
	wire [WIDTH-1:0] wire_d80_28;
	wire [WIDTH-1:0] wire_d80_29;
	wire [WIDTH-1:0] wire_d80_30;
	wire [WIDTH-1:0] wire_d80_31;
	wire [WIDTH-1:0] wire_d80_32;
	wire [WIDTH-1:0] wire_d80_33;
	wire [WIDTH-1:0] wire_d80_34;
	wire [WIDTH-1:0] wire_d80_35;
	wire [WIDTH-1:0] wire_d80_36;
	wire [WIDTH-1:0] wire_d80_37;
	wire [WIDTH-1:0] wire_d80_38;
	wire [WIDTH-1:0] wire_d80_39;
	wire [WIDTH-1:0] wire_d80_40;
	wire [WIDTH-1:0] wire_d80_41;
	wire [WIDTH-1:0] wire_d80_42;
	wire [WIDTH-1:0] wire_d80_43;
	wire [WIDTH-1:0] wire_d80_44;
	wire [WIDTH-1:0] wire_d80_45;
	wire [WIDTH-1:0] wire_d80_46;
	wire [WIDTH-1:0] wire_d80_47;
	wire [WIDTH-1:0] wire_d80_48;
	wire [WIDTH-1:0] wire_d80_49;
	wire [WIDTH-1:0] wire_d80_50;
	wire [WIDTH-1:0] wire_d80_51;
	wire [WIDTH-1:0] wire_d80_52;
	wire [WIDTH-1:0] wire_d80_53;
	wire [WIDTH-1:0] wire_d80_54;
	wire [WIDTH-1:0] wire_d80_55;
	wire [WIDTH-1:0] wire_d80_56;
	wire [WIDTH-1:0] wire_d80_57;
	wire [WIDTH-1:0] wire_d80_58;
	wire [WIDTH-1:0] wire_d80_59;
	wire [WIDTH-1:0] wire_d80_60;
	wire [WIDTH-1:0] wire_d80_61;
	wire [WIDTH-1:0] wire_d80_62;
	wire [WIDTH-1:0] wire_d80_63;
	wire [WIDTH-1:0] wire_d80_64;
	wire [WIDTH-1:0] wire_d80_65;
	wire [WIDTH-1:0] wire_d80_66;
	wire [WIDTH-1:0] wire_d80_67;
	wire [WIDTH-1:0] wire_d80_68;
	wire [WIDTH-1:0] wire_d80_69;
	wire [WIDTH-1:0] wire_d80_70;
	wire [WIDTH-1:0] wire_d80_71;
	wire [WIDTH-1:0] wire_d80_72;
	wire [WIDTH-1:0] wire_d80_73;
	wire [WIDTH-1:0] wire_d80_74;
	wire [WIDTH-1:0] wire_d80_75;
	wire [WIDTH-1:0] wire_d80_76;
	wire [WIDTH-1:0] wire_d80_77;
	wire [WIDTH-1:0] wire_d80_78;
	wire [WIDTH-1:0] wire_d81_0;
	wire [WIDTH-1:0] wire_d81_1;
	wire [WIDTH-1:0] wire_d81_2;
	wire [WIDTH-1:0] wire_d81_3;
	wire [WIDTH-1:0] wire_d81_4;
	wire [WIDTH-1:0] wire_d81_5;
	wire [WIDTH-1:0] wire_d81_6;
	wire [WIDTH-1:0] wire_d81_7;
	wire [WIDTH-1:0] wire_d81_8;
	wire [WIDTH-1:0] wire_d81_9;
	wire [WIDTH-1:0] wire_d81_10;
	wire [WIDTH-1:0] wire_d81_11;
	wire [WIDTH-1:0] wire_d81_12;
	wire [WIDTH-1:0] wire_d81_13;
	wire [WIDTH-1:0] wire_d81_14;
	wire [WIDTH-1:0] wire_d81_15;
	wire [WIDTH-1:0] wire_d81_16;
	wire [WIDTH-1:0] wire_d81_17;
	wire [WIDTH-1:0] wire_d81_18;
	wire [WIDTH-1:0] wire_d81_19;
	wire [WIDTH-1:0] wire_d81_20;
	wire [WIDTH-1:0] wire_d81_21;
	wire [WIDTH-1:0] wire_d81_22;
	wire [WIDTH-1:0] wire_d81_23;
	wire [WIDTH-1:0] wire_d81_24;
	wire [WIDTH-1:0] wire_d81_25;
	wire [WIDTH-1:0] wire_d81_26;
	wire [WIDTH-1:0] wire_d81_27;
	wire [WIDTH-1:0] wire_d81_28;
	wire [WIDTH-1:0] wire_d81_29;
	wire [WIDTH-1:0] wire_d81_30;
	wire [WIDTH-1:0] wire_d81_31;
	wire [WIDTH-1:0] wire_d81_32;
	wire [WIDTH-1:0] wire_d81_33;
	wire [WIDTH-1:0] wire_d81_34;
	wire [WIDTH-1:0] wire_d81_35;
	wire [WIDTH-1:0] wire_d81_36;
	wire [WIDTH-1:0] wire_d81_37;
	wire [WIDTH-1:0] wire_d81_38;
	wire [WIDTH-1:0] wire_d81_39;
	wire [WIDTH-1:0] wire_d81_40;
	wire [WIDTH-1:0] wire_d81_41;
	wire [WIDTH-1:0] wire_d81_42;
	wire [WIDTH-1:0] wire_d81_43;
	wire [WIDTH-1:0] wire_d81_44;
	wire [WIDTH-1:0] wire_d81_45;
	wire [WIDTH-1:0] wire_d81_46;
	wire [WIDTH-1:0] wire_d81_47;
	wire [WIDTH-1:0] wire_d81_48;
	wire [WIDTH-1:0] wire_d81_49;
	wire [WIDTH-1:0] wire_d81_50;
	wire [WIDTH-1:0] wire_d81_51;
	wire [WIDTH-1:0] wire_d81_52;
	wire [WIDTH-1:0] wire_d81_53;
	wire [WIDTH-1:0] wire_d81_54;
	wire [WIDTH-1:0] wire_d81_55;
	wire [WIDTH-1:0] wire_d81_56;
	wire [WIDTH-1:0] wire_d81_57;
	wire [WIDTH-1:0] wire_d81_58;
	wire [WIDTH-1:0] wire_d81_59;
	wire [WIDTH-1:0] wire_d81_60;
	wire [WIDTH-1:0] wire_d81_61;
	wire [WIDTH-1:0] wire_d81_62;
	wire [WIDTH-1:0] wire_d81_63;
	wire [WIDTH-1:0] wire_d81_64;
	wire [WIDTH-1:0] wire_d81_65;
	wire [WIDTH-1:0] wire_d81_66;
	wire [WIDTH-1:0] wire_d81_67;
	wire [WIDTH-1:0] wire_d81_68;
	wire [WIDTH-1:0] wire_d81_69;
	wire [WIDTH-1:0] wire_d81_70;
	wire [WIDTH-1:0] wire_d81_71;
	wire [WIDTH-1:0] wire_d81_72;
	wire [WIDTH-1:0] wire_d81_73;
	wire [WIDTH-1:0] wire_d81_74;
	wire [WIDTH-1:0] wire_d81_75;
	wire [WIDTH-1:0] wire_d81_76;
	wire [WIDTH-1:0] wire_d81_77;
	wire [WIDTH-1:0] wire_d81_78;
	wire [WIDTH-1:0] wire_d82_0;
	wire [WIDTH-1:0] wire_d82_1;
	wire [WIDTH-1:0] wire_d82_2;
	wire [WIDTH-1:0] wire_d82_3;
	wire [WIDTH-1:0] wire_d82_4;
	wire [WIDTH-1:0] wire_d82_5;
	wire [WIDTH-1:0] wire_d82_6;
	wire [WIDTH-1:0] wire_d82_7;
	wire [WIDTH-1:0] wire_d82_8;
	wire [WIDTH-1:0] wire_d82_9;
	wire [WIDTH-1:0] wire_d82_10;
	wire [WIDTH-1:0] wire_d82_11;
	wire [WIDTH-1:0] wire_d82_12;
	wire [WIDTH-1:0] wire_d82_13;
	wire [WIDTH-1:0] wire_d82_14;
	wire [WIDTH-1:0] wire_d82_15;
	wire [WIDTH-1:0] wire_d82_16;
	wire [WIDTH-1:0] wire_d82_17;
	wire [WIDTH-1:0] wire_d82_18;
	wire [WIDTH-1:0] wire_d82_19;
	wire [WIDTH-1:0] wire_d82_20;
	wire [WIDTH-1:0] wire_d82_21;
	wire [WIDTH-1:0] wire_d82_22;
	wire [WIDTH-1:0] wire_d82_23;
	wire [WIDTH-1:0] wire_d82_24;
	wire [WIDTH-1:0] wire_d82_25;
	wire [WIDTH-1:0] wire_d82_26;
	wire [WIDTH-1:0] wire_d82_27;
	wire [WIDTH-1:0] wire_d82_28;
	wire [WIDTH-1:0] wire_d82_29;
	wire [WIDTH-1:0] wire_d82_30;
	wire [WIDTH-1:0] wire_d82_31;
	wire [WIDTH-1:0] wire_d82_32;
	wire [WIDTH-1:0] wire_d82_33;
	wire [WIDTH-1:0] wire_d82_34;
	wire [WIDTH-1:0] wire_d82_35;
	wire [WIDTH-1:0] wire_d82_36;
	wire [WIDTH-1:0] wire_d82_37;
	wire [WIDTH-1:0] wire_d82_38;
	wire [WIDTH-1:0] wire_d82_39;
	wire [WIDTH-1:0] wire_d82_40;
	wire [WIDTH-1:0] wire_d82_41;
	wire [WIDTH-1:0] wire_d82_42;
	wire [WIDTH-1:0] wire_d82_43;
	wire [WIDTH-1:0] wire_d82_44;
	wire [WIDTH-1:0] wire_d82_45;
	wire [WIDTH-1:0] wire_d82_46;
	wire [WIDTH-1:0] wire_d82_47;
	wire [WIDTH-1:0] wire_d82_48;
	wire [WIDTH-1:0] wire_d82_49;
	wire [WIDTH-1:0] wire_d82_50;
	wire [WIDTH-1:0] wire_d82_51;
	wire [WIDTH-1:0] wire_d82_52;
	wire [WIDTH-1:0] wire_d82_53;
	wire [WIDTH-1:0] wire_d82_54;
	wire [WIDTH-1:0] wire_d82_55;
	wire [WIDTH-1:0] wire_d82_56;
	wire [WIDTH-1:0] wire_d82_57;
	wire [WIDTH-1:0] wire_d82_58;
	wire [WIDTH-1:0] wire_d82_59;
	wire [WIDTH-1:0] wire_d82_60;
	wire [WIDTH-1:0] wire_d82_61;
	wire [WIDTH-1:0] wire_d82_62;
	wire [WIDTH-1:0] wire_d82_63;
	wire [WIDTH-1:0] wire_d82_64;
	wire [WIDTH-1:0] wire_d82_65;
	wire [WIDTH-1:0] wire_d82_66;
	wire [WIDTH-1:0] wire_d82_67;
	wire [WIDTH-1:0] wire_d82_68;
	wire [WIDTH-1:0] wire_d82_69;
	wire [WIDTH-1:0] wire_d82_70;
	wire [WIDTH-1:0] wire_d82_71;
	wire [WIDTH-1:0] wire_d82_72;
	wire [WIDTH-1:0] wire_d82_73;
	wire [WIDTH-1:0] wire_d82_74;
	wire [WIDTH-1:0] wire_d82_75;
	wire [WIDTH-1:0] wire_d82_76;
	wire [WIDTH-1:0] wire_d82_77;
	wire [WIDTH-1:0] wire_d82_78;
	wire [WIDTH-1:0] wire_d83_0;
	wire [WIDTH-1:0] wire_d83_1;
	wire [WIDTH-1:0] wire_d83_2;
	wire [WIDTH-1:0] wire_d83_3;
	wire [WIDTH-1:0] wire_d83_4;
	wire [WIDTH-1:0] wire_d83_5;
	wire [WIDTH-1:0] wire_d83_6;
	wire [WIDTH-1:0] wire_d83_7;
	wire [WIDTH-1:0] wire_d83_8;
	wire [WIDTH-1:0] wire_d83_9;
	wire [WIDTH-1:0] wire_d83_10;
	wire [WIDTH-1:0] wire_d83_11;
	wire [WIDTH-1:0] wire_d83_12;
	wire [WIDTH-1:0] wire_d83_13;
	wire [WIDTH-1:0] wire_d83_14;
	wire [WIDTH-1:0] wire_d83_15;
	wire [WIDTH-1:0] wire_d83_16;
	wire [WIDTH-1:0] wire_d83_17;
	wire [WIDTH-1:0] wire_d83_18;
	wire [WIDTH-1:0] wire_d83_19;
	wire [WIDTH-1:0] wire_d83_20;
	wire [WIDTH-1:0] wire_d83_21;
	wire [WIDTH-1:0] wire_d83_22;
	wire [WIDTH-1:0] wire_d83_23;
	wire [WIDTH-1:0] wire_d83_24;
	wire [WIDTH-1:0] wire_d83_25;
	wire [WIDTH-1:0] wire_d83_26;
	wire [WIDTH-1:0] wire_d83_27;
	wire [WIDTH-1:0] wire_d83_28;
	wire [WIDTH-1:0] wire_d83_29;
	wire [WIDTH-1:0] wire_d83_30;
	wire [WIDTH-1:0] wire_d83_31;
	wire [WIDTH-1:0] wire_d83_32;
	wire [WIDTH-1:0] wire_d83_33;
	wire [WIDTH-1:0] wire_d83_34;
	wire [WIDTH-1:0] wire_d83_35;
	wire [WIDTH-1:0] wire_d83_36;
	wire [WIDTH-1:0] wire_d83_37;
	wire [WIDTH-1:0] wire_d83_38;
	wire [WIDTH-1:0] wire_d83_39;
	wire [WIDTH-1:0] wire_d83_40;
	wire [WIDTH-1:0] wire_d83_41;
	wire [WIDTH-1:0] wire_d83_42;
	wire [WIDTH-1:0] wire_d83_43;
	wire [WIDTH-1:0] wire_d83_44;
	wire [WIDTH-1:0] wire_d83_45;
	wire [WIDTH-1:0] wire_d83_46;
	wire [WIDTH-1:0] wire_d83_47;
	wire [WIDTH-1:0] wire_d83_48;
	wire [WIDTH-1:0] wire_d83_49;
	wire [WIDTH-1:0] wire_d83_50;
	wire [WIDTH-1:0] wire_d83_51;
	wire [WIDTH-1:0] wire_d83_52;
	wire [WIDTH-1:0] wire_d83_53;
	wire [WIDTH-1:0] wire_d83_54;
	wire [WIDTH-1:0] wire_d83_55;
	wire [WIDTH-1:0] wire_d83_56;
	wire [WIDTH-1:0] wire_d83_57;
	wire [WIDTH-1:0] wire_d83_58;
	wire [WIDTH-1:0] wire_d83_59;
	wire [WIDTH-1:0] wire_d83_60;
	wire [WIDTH-1:0] wire_d83_61;
	wire [WIDTH-1:0] wire_d83_62;
	wire [WIDTH-1:0] wire_d83_63;
	wire [WIDTH-1:0] wire_d83_64;
	wire [WIDTH-1:0] wire_d83_65;
	wire [WIDTH-1:0] wire_d83_66;
	wire [WIDTH-1:0] wire_d83_67;
	wire [WIDTH-1:0] wire_d83_68;
	wire [WIDTH-1:0] wire_d83_69;
	wire [WIDTH-1:0] wire_d83_70;
	wire [WIDTH-1:0] wire_d83_71;
	wire [WIDTH-1:0] wire_d83_72;
	wire [WIDTH-1:0] wire_d83_73;
	wire [WIDTH-1:0] wire_d83_74;
	wire [WIDTH-1:0] wire_d83_75;
	wire [WIDTH-1:0] wire_d83_76;
	wire [WIDTH-1:0] wire_d83_77;
	wire [WIDTH-1:0] wire_d83_78;
	wire [WIDTH-1:0] wire_d84_0;
	wire [WIDTH-1:0] wire_d84_1;
	wire [WIDTH-1:0] wire_d84_2;
	wire [WIDTH-1:0] wire_d84_3;
	wire [WIDTH-1:0] wire_d84_4;
	wire [WIDTH-1:0] wire_d84_5;
	wire [WIDTH-1:0] wire_d84_6;
	wire [WIDTH-1:0] wire_d84_7;
	wire [WIDTH-1:0] wire_d84_8;
	wire [WIDTH-1:0] wire_d84_9;
	wire [WIDTH-1:0] wire_d84_10;
	wire [WIDTH-1:0] wire_d84_11;
	wire [WIDTH-1:0] wire_d84_12;
	wire [WIDTH-1:0] wire_d84_13;
	wire [WIDTH-1:0] wire_d84_14;
	wire [WIDTH-1:0] wire_d84_15;
	wire [WIDTH-1:0] wire_d84_16;
	wire [WIDTH-1:0] wire_d84_17;
	wire [WIDTH-1:0] wire_d84_18;
	wire [WIDTH-1:0] wire_d84_19;
	wire [WIDTH-1:0] wire_d84_20;
	wire [WIDTH-1:0] wire_d84_21;
	wire [WIDTH-1:0] wire_d84_22;
	wire [WIDTH-1:0] wire_d84_23;
	wire [WIDTH-1:0] wire_d84_24;
	wire [WIDTH-1:0] wire_d84_25;
	wire [WIDTH-1:0] wire_d84_26;
	wire [WIDTH-1:0] wire_d84_27;
	wire [WIDTH-1:0] wire_d84_28;
	wire [WIDTH-1:0] wire_d84_29;
	wire [WIDTH-1:0] wire_d84_30;
	wire [WIDTH-1:0] wire_d84_31;
	wire [WIDTH-1:0] wire_d84_32;
	wire [WIDTH-1:0] wire_d84_33;
	wire [WIDTH-1:0] wire_d84_34;
	wire [WIDTH-1:0] wire_d84_35;
	wire [WIDTH-1:0] wire_d84_36;
	wire [WIDTH-1:0] wire_d84_37;
	wire [WIDTH-1:0] wire_d84_38;
	wire [WIDTH-1:0] wire_d84_39;
	wire [WIDTH-1:0] wire_d84_40;
	wire [WIDTH-1:0] wire_d84_41;
	wire [WIDTH-1:0] wire_d84_42;
	wire [WIDTH-1:0] wire_d84_43;
	wire [WIDTH-1:0] wire_d84_44;
	wire [WIDTH-1:0] wire_d84_45;
	wire [WIDTH-1:0] wire_d84_46;
	wire [WIDTH-1:0] wire_d84_47;
	wire [WIDTH-1:0] wire_d84_48;
	wire [WIDTH-1:0] wire_d84_49;
	wire [WIDTH-1:0] wire_d84_50;
	wire [WIDTH-1:0] wire_d84_51;
	wire [WIDTH-1:0] wire_d84_52;
	wire [WIDTH-1:0] wire_d84_53;
	wire [WIDTH-1:0] wire_d84_54;
	wire [WIDTH-1:0] wire_d84_55;
	wire [WIDTH-1:0] wire_d84_56;
	wire [WIDTH-1:0] wire_d84_57;
	wire [WIDTH-1:0] wire_d84_58;
	wire [WIDTH-1:0] wire_d84_59;
	wire [WIDTH-1:0] wire_d84_60;
	wire [WIDTH-1:0] wire_d84_61;
	wire [WIDTH-1:0] wire_d84_62;
	wire [WIDTH-1:0] wire_d84_63;
	wire [WIDTH-1:0] wire_d84_64;
	wire [WIDTH-1:0] wire_d84_65;
	wire [WIDTH-1:0] wire_d84_66;
	wire [WIDTH-1:0] wire_d84_67;
	wire [WIDTH-1:0] wire_d84_68;
	wire [WIDTH-1:0] wire_d84_69;
	wire [WIDTH-1:0] wire_d84_70;
	wire [WIDTH-1:0] wire_d84_71;
	wire [WIDTH-1:0] wire_d84_72;
	wire [WIDTH-1:0] wire_d84_73;
	wire [WIDTH-1:0] wire_d84_74;
	wire [WIDTH-1:0] wire_d84_75;
	wire [WIDTH-1:0] wire_d84_76;
	wire [WIDTH-1:0] wire_d84_77;
	wire [WIDTH-1:0] wire_d84_78;
	wire [WIDTH-1:0] wire_d85_0;
	wire [WIDTH-1:0] wire_d85_1;
	wire [WIDTH-1:0] wire_d85_2;
	wire [WIDTH-1:0] wire_d85_3;
	wire [WIDTH-1:0] wire_d85_4;
	wire [WIDTH-1:0] wire_d85_5;
	wire [WIDTH-1:0] wire_d85_6;
	wire [WIDTH-1:0] wire_d85_7;
	wire [WIDTH-1:0] wire_d85_8;
	wire [WIDTH-1:0] wire_d85_9;
	wire [WIDTH-1:0] wire_d85_10;
	wire [WIDTH-1:0] wire_d85_11;
	wire [WIDTH-1:0] wire_d85_12;
	wire [WIDTH-1:0] wire_d85_13;
	wire [WIDTH-1:0] wire_d85_14;
	wire [WIDTH-1:0] wire_d85_15;
	wire [WIDTH-1:0] wire_d85_16;
	wire [WIDTH-1:0] wire_d85_17;
	wire [WIDTH-1:0] wire_d85_18;
	wire [WIDTH-1:0] wire_d85_19;
	wire [WIDTH-1:0] wire_d85_20;
	wire [WIDTH-1:0] wire_d85_21;
	wire [WIDTH-1:0] wire_d85_22;
	wire [WIDTH-1:0] wire_d85_23;
	wire [WIDTH-1:0] wire_d85_24;
	wire [WIDTH-1:0] wire_d85_25;
	wire [WIDTH-1:0] wire_d85_26;
	wire [WIDTH-1:0] wire_d85_27;
	wire [WIDTH-1:0] wire_d85_28;
	wire [WIDTH-1:0] wire_d85_29;
	wire [WIDTH-1:0] wire_d85_30;
	wire [WIDTH-1:0] wire_d85_31;
	wire [WIDTH-1:0] wire_d85_32;
	wire [WIDTH-1:0] wire_d85_33;
	wire [WIDTH-1:0] wire_d85_34;
	wire [WIDTH-1:0] wire_d85_35;
	wire [WIDTH-1:0] wire_d85_36;
	wire [WIDTH-1:0] wire_d85_37;
	wire [WIDTH-1:0] wire_d85_38;
	wire [WIDTH-1:0] wire_d85_39;
	wire [WIDTH-1:0] wire_d85_40;
	wire [WIDTH-1:0] wire_d85_41;
	wire [WIDTH-1:0] wire_d85_42;
	wire [WIDTH-1:0] wire_d85_43;
	wire [WIDTH-1:0] wire_d85_44;
	wire [WIDTH-1:0] wire_d85_45;
	wire [WIDTH-1:0] wire_d85_46;
	wire [WIDTH-1:0] wire_d85_47;
	wire [WIDTH-1:0] wire_d85_48;
	wire [WIDTH-1:0] wire_d85_49;
	wire [WIDTH-1:0] wire_d85_50;
	wire [WIDTH-1:0] wire_d85_51;
	wire [WIDTH-1:0] wire_d85_52;
	wire [WIDTH-1:0] wire_d85_53;
	wire [WIDTH-1:0] wire_d85_54;
	wire [WIDTH-1:0] wire_d85_55;
	wire [WIDTH-1:0] wire_d85_56;
	wire [WIDTH-1:0] wire_d85_57;
	wire [WIDTH-1:0] wire_d85_58;
	wire [WIDTH-1:0] wire_d85_59;
	wire [WIDTH-1:0] wire_d85_60;
	wire [WIDTH-1:0] wire_d85_61;
	wire [WIDTH-1:0] wire_d85_62;
	wire [WIDTH-1:0] wire_d85_63;
	wire [WIDTH-1:0] wire_d85_64;
	wire [WIDTH-1:0] wire_d85_65;
	wire [WIDTH-1:0] wire_d85_66;
	wire [WIDTH-1:0] wire_d85_67;
	wire [WIDTH-1:0] wire_d85_68;
	wire [WIDTH-1:0] wire_d85_69;
	wire [WIDTH-1:0] wire_d85_70;
	wire [WIDTH-1:0] wire_d85_71;
	wire [WIDTH-1:0] wire_d85_72;
	wire [WIDTH-1:0] wire_d85_73;
	wire [WIDTH-1:0] wire_d85_74;
	wire [WIDTH-1:0] wire_d85_75;
	wire [WIDTH-1:0] wire_d85_76;
	wire [WIDTH-1:0] wire_d85_77;
	wire [WIDTH-1:0] wire_d85_78;
	wire [WIDTH-1:0] wire_d86_0;
	wire [WIDTH-1:0] wire_d86_1;
	wire [WIDTH-1:0] wire_d86_2;
	wire [WIDTH-1:0] wire_d86_3;
	wire [WIDTH-1:0] wire_d86_4;
	wire [WIDTH-1:0] wire_d86_5;
	wire [WIDTH-1:0] wire_d86_6;
	wire [WIDTH-1:0] wire_d86_7;
	wire [WIDTH-1:0] wire_d86_8;
	wire [WIDTH-1:0] wire_d86_9;
	wire [WIDTH-1:0] wire_d86_10;
	wire [WIDTH-1:0] wire_d86_11;
	wire [WIDTH-1:0] wire_d86_12;
	wire [WIDTH-1:0] wire_d86_13;
	wire [WIDTH-1:0] wire_d86_14;
	wire [WIDTH-1:0] wire_d86_15;
	wire [WIDTH-1:0] wire_d86_16;
	wire [WIDTH-1:0] wire_d86_17;
	wire [WIDTH-1:0] wire_d86_18;
	wire [WIDTH-1:0] wire_d86_19;
	wire [WIDTH-1:0] wire_d86_20;
	wire [WIDTH-1:0] wire_d86_21;
	wire [WIDTH-1:0] wire_d86_22;
	wire [WIDTH-1:0] wire_d86_23;
	wire [WIDTH-1:0] wire_d86_24;
	wire [WIDTH-1:0] wire_d86_25;
	wire [WIDTH-1:0] wire_d86_26;
	wire [WIDTH-1:0] wire_d86_27;
	wire [WIDTH-1:0] wire_d86_28;
	wire [WIDTH-1:0] wire_d86_29;
	wire [WIDTH-1:0] wire_d86_30;
	wire [WIDTH-1:0] wire_d86_31;
	wire [WIDTH-1:0] wire_d86_32;
	wire [WIDTH-1:0] wire_d86_33;
	wire [WIDTH-1:0] wire_d86_34;
	wire [WIDTH-1:0] wire_d86_35;
	wire [WIDTH-1:0] wire_d86_36;
	wire [WIDTH-1:0] wire_d86_37;
	wire [WIDTH-1:0] wire_d86_38;
	wire [WIDTH-1:0] wire_d86_39;
	wire [WIDTH-1:0] wire_d86_40;
	wire [WIDTH-1:0] wire_d86_41;
	wire [WIDTH-1:0] wire_d86_42;
	wire [WIDTH-1:0] wire_d86_43;
	wire [WIDTH-1:0] wire_d86_44;
	wire [WIDTH-1:0] wire_d86_45;
	wire [WIDTH-1:0] wire_d86_46;
	wire [WIDTH-1:0] wire_d86_47;
	wire [WIDTH-1:0] wire_d86_48;
	wire [WIDTH-1:0] wire_d86_49;
	wire [WIDTH-1:0] wire_d86_50;
	wire [WIDTH-1:0] wire_d86_51;
	wire [WIDTH-1:0] wire_d86_52;
	wire [WIDTH-1:0] wire_d86_53;
	wire [WIDTH-1:0] wire_d86_54;
	wire [WIDTH-1:0] wire_d86_55;
	wire [WIDTH-1:0] wire_d86_56;
	wire [WIDTH-1:0] wire_d86_57;
	wire [WIDTH-1:0] wire_d86_58;
	wire [WIDTH-1:0] wire_d86_59;
	wire [WIDTH-1:0] wire_d86_60;
	wire [WIDTH-1:0] wire_d86_61;
	wire [WIDTH-1:0] wire_d86_62;
	wire [WIDTH-1:0] wire_d86_63;
	wire [WIDTH-1:0] wire_d86_64;
	wire [WIDTH-1:0] wire_d86_65;
	wire [WIDTH-1:0] wire_d86_66;
	wire [WIDTH-1:0] wire_d86_67;
	wire [WIDTH-1:0] wire_d86_68;
	wire [WIDTH-1:0] wire_d86_69;
	wire [WIDTH-1:0] wire_d86_70;
	wire [WIDTH-1:0] wire_d86_71;
	wire [WIDTH-1:0] wire_d86_72;
	wire [WIDTH-1:0] wire_d86_73;
	wire [WIDTH-1:0] wire_d86_74;
	wire [WIDTH-1:0] wire_d86_75;
	wire [WIDTH-1:0] wire_d86_76;
	wire [WIDTH-1:0] wire_d86_77;
	wire [WIDTH-1:0] wire_d86_78;
	wire [WIDTH-1:0] wire_d87_0;
	wire [WIDTH-1:0] wire_d87_1;
	wire [WIDTH-1:0] wire_d87_2;
	wire [WIDTH-1:0] wire_d87_3;
	wire [WIDTH-1:0] wire_d87_4;
	wire [WIDTH-1:0] wire_d87_5;
	wire [WIDTH-1:0] wire_d87_6;
	wire [WIDTH-1:0] wire_d87_7;
	wire [WIDTH-1:0] wire_d87_8;
	wire [WIDTH-1:0] wire_d87_9;
	wire [WIDTH-1:0] wire_d87_10;
	wire [WIDTH-1:0] wire_d87_11;
	wire [WIDTH-1:0] wire_d87_12;
	wire [WIDTH-1:0] wire_d87_13;
	wire [WIDTH-1:0] wire_d87_14;
	wire [WIDTH-1:0] wire_d87_15;
	wire [WIDTH-1:0] wire_d87_16;
	wire [WIDTH-1:0] wire_d87_17;
	wire [WIDTH-1:0] wire_d87_18;
	wire [WIDTH-1:0] wire_d87_19;
	wire [WIDTH-1:0] wire_d87_20;
	wire [WIDTH-1:0] wire_d87_21;
	wire [WIDTH-1:0] wire_d87_22;
	wire [WIDTH-1:0] wire_d87_23;
	wire [WIDTH-1:0] wire_d87_24;
	wire [WIDTH-1:0] wire_d87_25;
	wire [WIDTH-1:0] wire_d87_26;
	wire [WIDTH-1:0] wire_d87_27;
	wire [WIDTH-1:0] wire_d87_28;
	wire [WIDTH-1:0] wire_d87_29;
	wire [WIDTH-1:0] wire_d87_30;
	wire [WIDTH-1:0] wire_d87_31;
	wire [WIDTH-1:0] wire_d87_32;
	wire [WIDTH-1:0] wire_d87_33;
	wire [WIDTH-1:0] wire_d87_34;
	wire [WIDTH-1:0] wire_d87_35;
	wire [WIDTH-1:0] wire_d87_36;
	wire [WIDTH-1:0] wire_d87_37;
	wire [WIDTH-1:0] wire_d87_38;
	wire [WIDTH-1:0] wire_d87_39;
	wire [WIDTH-1:0] wire_d87_40;
	wire [WIDTH-1:0] wire_d87_41;
	wire [WIDTH-1:0] wire_d87_42;
	wire [WIDTH-1:0] wire_d87_43;
	wire [WIDTH-1:0] wire_d87_44;
	wire [WIDTH-1:0] wire_d87_45;
	wire [WIDTH-1:0] wire_d87_46;
	wire [WIDTH-1:0] wire_d87_47;
	wire [WIDTH-1:0] wire_d87_48;
	wire [WIDTH-1:0] wire_d87_49;
	wire [WIDTH-1:0] wire_d87_50;
	wire [WIDTH-1:0] wire_d87_51;
	wire [WIDTH-1:0] wire_d87_52;
	wire [WIDTH-1:0] wire_d87_53;
	wire [WIDTH-1:0] wire_d87_54;
	wire [WIDTH-1:0] wire_d87_55;
	wire [WIDTH-1:0] wire_d87_56;
	wire [WIDTH-1:0] wire_d87_57;
	wire [WIDTH-1:0] wire_d87_58;
	wire [WIDTH-1:0] wire_d87_59;
	wire [WIDTH-1:0] wire_d87_60;
	wire [WIDTH-1:0] wire_d87_61;
	wire [WIDTH-1:0] wire_d87_62;
	wire [WIDTH-1:0] wire_d87_63;
	wire [WIDTH-1:0] wire_d87_64;
	wire [WIDTH-1:0] wire_d87_65;
	wire [WIDTH-1:0] wire_d87_66;
	wire [WIDTH-1:0] wire_d87_67;
	wire [WIDTH-1:0] wire_d87_68;
	wire [WIDTH-1:0] wire_d87_69;
	wire [WIDTH-1:0] wire_d87_70;
	wire [WIDTH-1:0] wire_d87_71;
	wire [WIDTH-1:0] wire_d87_72;
	wire [WIDTH-1:0] wire_d87_73;
	wire [WIDTH-1:0] wire_d87_74;
	wire [WIDTH-1:0] wire_d87_75;
	wire [WIDTH-1:0] wire_d87_76;
	wire [WIDTH-1:0] wire_d87_77;
	wire [WIDTH-1:0] wire_d87_78;
	wire [WIDTH-1:0] wire_d88_0;
	wire [WIDTH-1:0] wire_d88_1;
	wire [WIDTH-1:0] wire_d88_2;
	wire [WIDTH-1:0] wire_d88_3;
	wire [WIDTH-1:0] wire_d88_4;
	wire [WIDTH-1:0] wire_d88_5;
	wire [WIDTH-1:0] wire_d88_6;
	wire [WIDTH-1:0] wire_d88_7;
	wire [WIDTH-1:0] wire_d88_8;
	wire [WIDTH-1:0] wire_d88_9;
	wire [WIDTH-1:0] wire_d88_10;
	wire [WIDTH-1:0] wire_d88_11;
	wire [WIDTH-1:0] wire_d88_12;
	wire [WIDTH-1:0] wire_d88_13;
	wire [WIDTH-1:0] wire_d88_14;
	wire [WIDTH-1:0] wire_d88_15;
	wire [WIDTH-1:0] wire_d88_16;
	wire [WIDTH-1:0] wire_d88_17;
	wire [WIDTH-1:0] wire_d88_18;
	wire [WIDTH-1:0] wire_d88_19;
	wire [WIDTH-1:0] wire_d88_20;
	wire [WIDTH-1:0] wire_d88_21;
	wire [WIDTH-1:0] wire_d88_22;
	wire [WIDTH-1:0] wire_d88_23;
	wire [WIDTH-1:0] wire_d88_24;
	wire [WIDTH-1:0] wire_d88_25;
	wire [WIDTH-1:0] wire_d88_26;
	wire [WIDTH-1:0] wire_d88_27;
	wire [WIDTH-1:0] wire_d88_28;
	wire [WIDTH-1:0] wire_d88_29;
	wire [WIDTH-1:0] wire_d88_30;
	wire [WIDTH-1:0] wire_d88_31;
	wire [WIDTH-1:0] wire_d88_32;
	wire [WIDTH-1:0] wire_d88_33;
	wire [WIDTH-1:0] wire_d88_34;
	wire [WIDTH-1:0] wire_d88_35;
	wire [WIDTH-1:0] wire_d88_36;
	wire [WIDTH-1:0] wire_d88_37;
	wire [WIDTH-1:0] wire_d88_38;
	wire [WIDTH-1:0] wire_d88_39;
	wire [WIDTH-1:0] wire_d88_40;
	wire [WIDTH-1:0] wire_d88_41;
	wire [WIDTH-1:0] wire_d88_42;
	wire [WIDTH-1:0] wire_d88_43;
	wire [WIDTH-1:0] wire_d88_44;
	wire [WIDTH-1:0] wire_d88_45;
	wire [WIDTH-1:0] wire_d88_46;
	wire [WIDTH-1:0] wire_d88_47;
	wire [WIDTH-1:0] wire_d88_48;
	wire [WIDTH-1:0] wire_d88_49;
	wire [WIDTH-1:0] wire_d88_50;
	wire [WIDTH-1:0] wire_d88_51;
	wire [WIDTH-1:0] wire_d88_52;
	wire [WIDTH-1:0] wire_d88_53;
	wire [WIDTH-1:0] wire_d88_54;
	wire [WIDTH-1:0] wire_d88_55;
	wire [WIDTH-1:0] wire_d88_56;
	wire [WIDTH-1:0] wire_d88_57;
	wire [WIDTH-1:0] wire_d88_58;
	wire [WIDTH-1:0] wire_d88_59;
	wire [WIDTH-1:0] wire_d88_60;
	wire [WIDTH-1:0] wire_d88_61;
	wire [WIDTH-1:0] wire_d88_62;
	wire [WIDTH-1:0] wire_d88_63;
	wire [WIDTH-1:0] wire_d88_64;
	wire [WIDTH-1:0] wire_d88_65;
	wire [WIDTH-1:0] wire_d88_66;
	wire [WIDTH-1:0] wire_d88_67;
	wire [WIDTH-1:0] wire_d88_68;
	wire [WIDTH-1:0] wire_d88_69;
	wire [WIDTH-1:0] wire_d88_70;
	wire [WIDTH-1:0] wire_d88_71;
	wire [WIDTH-1:0] wire_d88_72;
	wire [WIDTH-1:0] wire_d88_73;
	wire [WIDTH-1:0] wire_d88_74;
	wire [WIDTH-1:0] wire_d88_75;
	wire [WIDTH-1:0] wire_d88_76;
	wire [WIDTH-1:0] wire_d88_77;
	wire [WIDTH-1:0] wire_d88_78;
	wire [WIDTH-1:0] wire_d89_0;
	wire [WIDTH-1:0] wire_d89_1;
	wire [WIDTH-1:0] wire_d89_2;
	wire [WIDTH-1:0] wire_d89_3;
	wire [WIDTH-1:0] wire_d89_4;
	wire [WIDTH-1:0] wire_d89_5;
	wire [WIDTH-1:0] wire_d89_6;
	wire [WIDTH-1:0] wire_d89_7;
	wire [WIDTH-1:0] wire_d89_8;
	wire [WIDTH-1:0] wire_d89_9;
	wire [WIDTH-1:0] wire_d89_10;
	wire [WIDTH-1:0] wire_d89_11;
	wire [WIDTH-1:0] wire_d89_12;
	wire [WIDTH-1:0] wire_d89_13;
	wire [WIDTH-1:0] wire_d89_14;
	wire [WIDTH-1:0] wire_d89_15;
	wire [WIDTH-1:0] wire_d89_16;
	wire [WIDTH-1:0] wire_d89_17;
	wire [WIDTH-1:0] wire_d89_18;
	wire [WIDTH-1:0] wire_d89_19;
	wire [WIDTH-1:0] wire_d89_20;
	wire [WIDTH-1:0] wire_d89_21;
	wire [WIDTH-1:0] wire_d89_22;
	wire [WIDTH-1:0] wire_d89_23;
	wire [WIDTH-1:0] wire_d89_24;
	wire [WIDTH-1:0] wire_d89_25;
	wire [WIDTH-1:0] wire_d89_26;
	wire [WIDTH-1:0] wire_d89_27;
	wire [WIDTH-1:0] wire_d89_28;
	wire [WIDTH-1:0] wire_d89_29;
	wire [WIDTH-1:0] wire_d89_30;
	wire [WIDTH-1:0] wire_d89_31;
	wire [WIDTH-1:0] wire_d89_32;
	wire [WIDTH-1:0] wire_d89_33;
	wire [WIDTH-1:0] wire_d89_34;
	wire [WIDTH-1:0] wire_d89_35;
	wire [WIDTH-1:0] wire_d89_36;
	wire [WIDTH-1:0] wire_d89_37;
	wire [WIDTH-1:0] wire_d89_38;
	wire [WIDTH-1:0] wire_d89_39;
	wire [WIDTH-1:0] wire_d89_40;
	wire [WIDTH-1:0] wire_d89_41;
	wire [WIDTH-1:0] wire_d89_42;
	wire [WIDTH-1:0] wire_d89_43;
	wire [WIDTH-1:0] wire_d89_44;
	wire [WIDTH-1:0] wire_d89_45;
	wire [WIDTH-1:0] wire_d89_46;
	wire [WIDTH-1:0] wire_d89_47;
	wire [WIDTH-1:0] wire_d89_48;
	wire [WIDTH-1:0] wire_d89_49;
	wire [WIDTH-1:0] wire_d89_50;
	wire [WIDTH-1:0] wire_d89_51;
	wire [WIDTH-1:0] wire_d89_52;
	wire [WIDTH-1:0] wire_d89_53;
	wire [WIDTH-1:0] wire_d89_54;
	wire [WIDTH-1:0] wire_d89_55;
	wire [WIDTH-1:0] wire_d89_56;
	wire [WIDTH-1:0] wire_d89_57;
	wire [WIDTH-1:0] wire_d89_58;
	wire [WIDTH-1:0] wire_d89_59;
	wire [WIDTH-1:0] wire_d89_60;
	wire [WIDTH-1:0] wire_d89_61;
	wire [WIDTH-1:0] wire_d89_62;
	wire [WIDTH-1:0] wire_d89_63;
	wire [WIDTH-1:0] wire_d89_64;
	wire [WIDTH-1:0] wire_d89_65;
	wire [WIDTH-1:0] wire_d89_66;
	wire [WIDTH-1:0] wire_d89_67;
	wire [WIDTH-1:0] wire_d89_68;
	wire [WIDTH-1:0] wire_d89_69;
	wire [WIDTH-1:0] wire_d89_70;
	wire [WIDTH-1:0] wire_d89_71;
	wire [WIDTH-1:0] wire_d89_72;
	wire [WIDTH-1:0] wire_d89_73;
	wire [WIDTH-1:0] wire_d89_74;
	wire [WIDTH-1:0] wire_d89_75;
	wire [WIDTH-1:0] wire_d89_76;
	wire [WIDTH-1:0] wire_d89_77;
	wire [WIDTH-1:0] wire_d89_78;
	wire [WIDTH-1:0] wire_d90_0;
	wire [WIDTH-1:0] wire_d90_1;
	wire [WIDTH-1:0] wire_d90_2;
	wire [WIDTH-1:0] wire_d90_3;
	wire [WIDTH-1:0] wire_d90_4;
	wire [WIDTH-1:0] wire_d90_5;
	wire [WIDTH-1:0] wire_d90_6;
	wire [WIDTH-1:0] wire_d90_7;
	wire [WIDTH-1:0] wire_d90_8;
	wire [WIDTH-1:0] wire_d90_9;
	wire [WIDTH-1:0] wire_d90_10;
	wire [WIDTH-1:0] wire_d90_11;
	wire [WIDTH-1:0] wire_d90_12;
	wire [WIDTH-1:0] wire_d90_13;
	wire [WIDTH-1:0] wire_d90_14;
	wire [WIDTH-1:0] wire_d90_15;
	wire [WIDTH-1:0] wire_d90_16;
	wire [WIDTH-1:0] wire_d90_17;
	wire [WIDTH-1:0] wire_d90_18;
	wire [WIDTH-1:0] wire_d90_19;
	wire [WIDTH-1:0] wire_d90_20;
	wire [WIDTH-1:0] wire_d90_21;
	wire [WIDTH-1:0] wire_d90_22;
	wire [WIDTH-1:0] wire_d90_23;
	wire [WIDTH-1:0] wire_d90_24;
	wire [WIDTH-1:0] wire_d90_25;
	wire [WIDTH-1:0] wire_d90_26;
	wire [WIDTH-1:0] wire_d90_27;
	wire [WIDTH-1:0] wire_d90_28;
	wire [WIDTH-1:0] wire_d90_29;
	wire [WIDTH-1:0] wire_d90_30;
	wire [WIDTH-1:0] wire_d90_31;
	wire [WIDTH-1:0] wire_d90_32;
	wire [WIDTH-1:0] wire_d90_33;
	wire [WIDTH-1:0] wire_d90_34;
	wire [WIDTH-1:0] wire_d90_35;
	wire [WIDTH-1:0] wire_d90_36;
	wire [WIDTH-1:0] wire_d90_37;
	wire [WIDTH-1:0] wire_d90_38;
	wire [WIDTH-1:0] wire_d90_39;
	wire [WIDTH-1:0] wire_d90_40;
	wire [WIDTH-1:0] wire_d90_41;
	wire [WIDTH-1:0] wire_d90_42;
	wire [WIDTH-1:0] wire_d90_43;
	wire [WIDTH-1:0] wire_d90_44;
	wire [WIDTH-1:0] wire_d90_45;
	wire [WIDTH-1:0] wire_d90_46;
	wire [WIDTH-1:0] wire_d90_47;
	wire [WIDTH-1:0] wire_d90_48;
	wire [WIDTH-1:0] wire_d90_49;
	wire [WIDTH-1:0] wire_d90_50;
	wire [WIDTH-1:0] wire_d90_51;
	wire [WIDTH-1:0] wire_d90_52;
	wire [WIDTH-1:0] wire_d90_53;
	wire [WIDTH-1:0] wire_d90_54;
	wire [WIDTH-1:0] wire_d90_55;
	wire [WIDTH-1:0] wire_d90_56;
	wire [WIDTH-1:0] wire_d90_57;
	wire [WIDTH-1:0] wire_d90_58;
	wire [WIDTH-1:0] wire_d90_59;
	wire [WIDTH-1:0] wire_d90_60;
	wire [WIDTH-1:0] wire_d90_61;
	wire [WIDTH-1:0] wire_d90_62;
	wire [WIDTH-1:0] wire_d90_63;
	wire [WIDTH-1:0] wire_d90_64;
	wire [WIDTH-1:0] wire_d90_65;
	wire [WIDTH-1:0] wire_d90_66;
	wire [WIDTH-1:0] wire_d90_67;
	wire [WIDTH-1:0] wire_d90_68;
	wire [WIDTH-1:0] wire_d90_69;
	wire [WIDTH-1:0] wire_d90_70;
	wire [WIDTH-1:0] wire_d90_71;
	wire [WIDTH-1:0] wire_d90_72;
	wire [WIDTH-1:0] wire_d90_73;
	wire [WIDTH-1:0] wire_d90_74;
	wire [WIDTH-1:0] wire_d90_75;
	wire [WIDTH-1:0] wire_d90_76;
	wire [WIDTH-1:0] wire_d90_77;
	wire [WIDTH-1:0] wire_d90_78;
	wire [WIDTH-1:0] wire_d91_0;
	wire [WIDTH-1:0] wire_d91_1;
	wire [WIDTH-1:0] wire_d91_2;
	wire [WIDTH-1:0] wire_d91_3;
	wire [WIDTH-1:0] wire_d91_4;
	wire [WIDTH-1:0] wire_d91_5;
	wire [WIDTH-1:0] wire_d91_6;
	wire [WIDTH-1:0] wire_d91_7;
	wire [WIDTH-1:0] wire_d91_8;
	wire [WIDTH-1:0] wire_d91_9;
	wire [WIDTH-1:0] wire_d91_10;
	wire [WIDTH-1:0] wire_d91_11;
	wire [WIDTH-1:0] wire_d91_12;
	wire [WIDTH-1:0] wire_d91_13;
	wire [WIDTH-1:0] wire_d91_14;
	wire [WIDTH-1:0] wire_d91_15;
	wire [WIDTH-1:0] wire_d91_16;
	wire [WIDTH-1:0] wire_d91_17;
	wire [WIDTH-1:0] wire_d91_18;
	wire [WIDTH-1:0] wire_d91_19;
	wire [WIDTH-1:0] wire_d91_20;
	wire [WIDTH-1:0] wire_d91_21;
	wire [WIDTH-1:0] wire_d91_22;
	wire [WIDTH-1:0] wire_d91_23;
	wire [WIDTH-1:0] wire_d91_24;
	wire [WIDTH-1:0] wire_d91_25;
	wire [WIDTH-1:0] wire_d91_26;
	wire [WIDTH-1:0] wire_d91_27;
	wire [WIDTH-1:0] wire_d91_28;
	wire [WIDTH-1:0] wire_d91_29;
	wire [WIDTH-1:0] wire_d91_30;
	wire [WIDTH-1:0] wire_d91_31;
	wire [WIDTH-1:0] wire_d91_32;
	wire [WIDTH-1:0] wire_d91_33;
	wire [WIDTH-1:0] wire_d91_34;
	wire [WIDTH-1:0] wire_d91_35;
	wire [WIDTH-1:0] wire_d91_36;
	wire [WIDTH-1:0] wire_d91_37;
	wire [WIDTH-1:0] wire_d91_38;
	wire [WIDTH-1:0] wire_d91_39;
	wire [WIDTH-1:0] wire_d91_40;
	wire [WIDTH-1:0] wire_d91_41;
	wire [WIDTH-1:0] wire_d91_42;
	wire [WIDTH-1:0] wire_d91_43;
	wire [WIDTH-1:0] wire_d91_44;
	wire [WIDTH-1:0] wire_d91_45;
	wire [WIDTH-1:0] wire_d91_46;
	wire [WIDTH-1:0] wire_d91_47;
	wire [WIDTH-1:0] wire_d91_48;
	wire [WIDTH-1:0] wire_d91_49;
	wire [WIDTH-1:0] wire_d91_50;
	wire [WIDTH-1:0] wire_d91_51;
	wire [WIDTH-1:0] wire_d91_52;
	wire [WIDTH-1:0] wire_d91_53;
	wire [WIDTH-1:0] wire_d91_54;
	wire [WIDTH-1:0] wire_d91_55;
	wire [WIDTH-1:0] wire_d91_56;
	wire [WIDTH-1:0] wire_d91_57;
	wire [WIDTH-1:0] wire_d91_58;
	wire [WIDTH-1:0] wire_d91_59;
	wire [WIDTH-1:0] wire_d91_60;
	wire [WIDTH-1:0] wire_d91_61;
	wire [WIDTH-1:0] wire_d91_62;
	wire [WIDTH-1:0] wire_d91_63;
	wire [WIDTH-1:0] wire_d91_64;
	wire [WIDTH-1:0] wire_d91_65;
	wire [WIDTH-1:0] wire_d91_66;
	wire [WIDTH-1:0] wire_d91_67;
	wire [WIDTH-1:0] wire_d91_68;
	wire [WIDTH-1:0] wire_d91_69;
	wire [WIDTH-1:0] wire_d91_70;
	wire [WIDTH-1:0] wire_d91_71;
	wire [WIDTH-1:0] wire_d91_72;
	wire [WIDTH-1:0] wire_d91_73;
	wire [WIDTH-1:0] wire_d91_74;
	wire [WIDTH-1:0] wire_d91_75;
	wire [WIDTH-1:0] wire_d91_76;
	wire [WIDTH-1:0] wire_d91_77;
	wire [WIDTH-1:0] wire_d91_78;
	wire [WIDTH-1:0] wire_d92_0;
	wire [WIDTH-1:0] wire_d92_1;
	wire [WIDTH-1:0] wire_d92_2;
	wire [WIDTH-1:0] wire_d92_3;
	wire [WIDTH-1:0] wire_d92_4;
	wire [WIDTH-1:0] wire_d92_5;
	wire [WIDTH-1:0] wire_d92_6;
	wire [WIDTH-1:0] wire_d92_7;
	wire [WIDTH-1:0] wire_d92_8;
	wire [WIDTH-1:0] wire_d92_9;
	wire [WIDTH-1:0] wire_d92_10;
	wire [WIDTH-1:0] wire_d92_11;
	wire [WIDTH-1:0] wire_d92_12;
	wire [WIDTH-1:0] wire_d92_13;
	wire [WIDTH-1:0] wire_d92_14;
	wire [WIDTH-1:0] wire_d92_15;
	wire [WIDTH-1:0] wire_d92_16;
	wire [WIDTH-1:0] wire_d92_17;
	wire [WIDTH-1:0] wire_d92_18;
	wire [WIDTH-1:0] wire_d92_19;
	wire [WIDTH-1:0] wire_d92_20;
	wire [WIDTH-1:0] wire_d92_21;
	wire [WIDTH-1:0] wire_d92_22;
	wire [WIDTH-1:0] wire_d92_23;
	wire [WIDTH-1:0] wire_d92_24;
	wire [WIDTH-1:0] wire_d92_25;
	wire [WIDTH-1:0] wire_d92_26;
	wire [WIDTH-1:0] wire_d92_27;
	wire [WIDTH-1:0] wire_d92_28;
	wire [WIDTH-1:0] wire_d92_29;
	wire [WIDTH-1:0] wire_d92_30;
	wire [WIDTH-1:0] wire_d92_31;
	wire [WIDTH-1:0] wire_d92_32;
	wire [WIDTH-1:0] wire_d92_33;
	wire [WIDTH-1:0] wire_d92_34;
	wire [WIDTH-1:0] wire_d92_35;
	wire [WIDTH-1:0] wire_d92_36;
	wire [WIDTH-1:0] wire_d92_37;
	wire [WIDTH-1:0] wire_d92_38;
	wire [WIDTH-1:0] wire_d92_39;
	wire [WIDTH-1:0] wire_d92_40;
	wire [WIDTH-1:0] wire_d92_41;
	wire [WIDTH-1:0] wire_d92_42;
	wire [WIDTH-1:0] wire_d92_43;
	wire [WIDTH-1:0] wire_d92_44;
	wire [WIDTH-1:0] wire_d92_45;
	wire [WIDTH-1:0] wire_d92_46;
	wire [WIDTH-1:0] wire_d92_47;
	wire [WIDTH-1:0] wire_d92_48;
	wire [WIDTH-1:0] wire_d92_49;
	wire [WIDTH-1:0] wire_d92_50;
	wire [WIDTH-1:0] wire_d92_51;
	wire [WIDTH-1:0] wire_d92_52;
	wire [WIDTH-1:0] wire_d92_53;
	wire [WIDTH-1:0] wire_d92_54;
	wire [WIDTH-1:0] wire_d92_55;
	wire [WIDTH-1:0] wire_d92_56;
	wire [WIDTH-1:0] wire_d92_57;
	wire [WIDTH-1:0] wire_d92_58;
	wire [WIDTH-1:0] wire_d92_59;
	wire [WIDTH-1:0] wire_d92_60;
	wire [WIDTH-1:0] wire_d92_61;
	wire [WIDTH-1:0] wire_d92_62;
	wire [WIDTH-1:0] wire_d92_63;
	wire [WIDTH-1:0] wire_d92_64;
	wire [WIDTH-1:0] wire_d92_65;
	wire [WIDTH-1:0] wire_d92_66;
	wire [WIDTH-1:0] wire_d92_67;
	wire [WIDTH-1:0] wire_d92_68;
	wire [WIDTH-1:0] wire_d92_69;
	wire [WIDTH-1:0] wire_d92_70;
	wire [WIDTH-1:0] wire_d92_71;
	wire [WIDTH-1:0] wire_d92_72;
	wire [WIDTH-1:0] wire_d92_73;
	wire [WIDTH-1:0] wire_d92_74;
	wire [WIDTH-1:0] wire_d92_75;
	wire [WIDTH-1:0] wire_d92_76;
	wire [WIDTH-1:0] wire_d92_77;
	wire [WIDTH-1:0] wire_d92_78;
	wire [WIDTH-1:0] wire_d93_0;
	wire [WIDTH-1:0] wire_d93_1;
	wire [WIDTH-1:0] wire_d93_2;
	wire [WIDTH-1:0] wire_d93_3;
	wire [WIDTH-1:0] wire_d93_4;
	wire [WIDTH-1:0] wire_d93_5;
	wire [WIDTH-1:0] wire_d93_6;
	wire [WIDTH-1:0] wire_d93_7;
	wire [WIDTH-1:0] wire_d93_8;
	wire [WIDTH-1:0] wire_d93_9;
	wire [WIDTH-1:0] wire_d93_10;
	wire [WIDTH-1:0] wire_d93_11;
	wire [WIDTH-1:0] wire_d93_12;
	wire [WIDTH-1:0] wire_d93_13;
	wire [WIDTH-1:0] wire_d93_14;
	wire [WIDTH-1:0] wire_d93_15;
	wire [WIDTH-1:0] wire_d93_16;
	wire [WIDTH-1:0] wire_d93_17;
	wire [WIDTH-1:0] wire_d93_18;
	wire [WIDTH-1:0] wire_d93_19;
	wire [WIDTH-1:0] wire_d93_20;
	wire [WIDTH-1:0] wire_d93_21;
	wire [WIDTH-1:0] wire_d93_22;
	wire [WIDTH-1:0] wire_d93_23;
	wire [WIDTH-1:0] wire_d93_24;
	wire [WIDTH-1:0] wire_d93_25;
	wire [WIDTH-1:0] wire_d93_26;
	wire [WIDTH-1:0] wire_d93_27;
	wire [WIDTH-1:0] wire_d93_28;
	wire [WIDTH-1:0] wire_d93_29;
	wire [WIDTH-1:0] wire_d93_30;
	wire [WIDTH-1:0] wire_d93_31;
	wire [WIDTH-1:0] wire_d93_32;
	wire [WIDTH-1:0] wire_d93_33;
	wire [WIDTH-1:0] wire_d93_34;
	wire [WIDTH-1:0] wire_d93_35;
	wire [WIDTH-1:0] wire_d93_36;
	wire [WIDTH-1:0] wire_d93_37;
	wire [WIDTH-1:0] wire_d93_38;
	wire [WIDTH-1:0] wire_d93_39;
	wire [WIDTH-1:0] wire_d93_40;
	wire [WIDTH-1:0] wire_d93_41;
	wire [WIDTH-1:0] wire_d93_42;
	wire [WIDTH-1:0] wire_d93_43;
	wire [WIDTH-1:0] wire_d93_44;
	wire [WIDTH-1:0] wire_d93_45;
	wire [WIDTH-1:0] wire_d93_46;
	wire [WIDTH-1:0] wire_d93_47;
	wire [WIDTH-1:0] wire_d93_48;
	wire [WIDTH-1:0] wire_d93_49;
	wire [WIDTH-1:0] wire_d93_50;
	wire [WIDTH-1:0] wire_d93_51;
	wire [WIDTH-1:0] wire_d93_52;
	wire [WIDTH-1:0] wire_d93_53;
	wire [WIDTH-1:0] wire_d93_54;
	wire [WIDTH-1:0] wire_d93_55;
	wire [WIDTH-1:0] wire_d93_56;
	wire [WIDTH-1:0] wire_d93_57;
	wire [WIDTH-1:0] wire_d93_58;
	wire [WIDTH-1:0] wire_d93_59;
	wire [WIDTH-1:0] wire_d93_60;
	wire [WIDTH-1:0] wire_d93_61;
	wire [WIDTH-1:0] wire_d93_62;
	wire [WIDTH-1:0] wire_d93_63;
	wire [WIDTH-1:0] wire_d93_64;
	wire [WIDTH-1:0] wire_d93_65;
	wire [WIDTH-1:0] wire_d93_66;
	wire [WIDTH-1:0] wire_d93_67;
	wire [WIDTH-1:0] wire_d93_68;
	wire [WIDTH-1:0] wire_d93_69;
	wire [WIDTH-1:0] wire_d93_70;
	wire [WIDTH-1:0] wire_d93_71;
	wire [WIDTH-1:0] wire_d93_72;
	wire [WIDTH-1:0] wire_d93_73;
	wire [WIDTH-1:0] wire_d93_74;
	wire [WIDTH-1:0] wire_d93_75;
	wire [WIDTH-1:0] wire_d93_76;
	wire [WIDTH-1:0] wire_d93_77;
	wire [WIDTH-1:0] wire_d93_78;
	wire [WIDTH-1:0] wire_d94_0;
	wire [WIDTH-1:0] wire_d94_1;
	wire [WIDTH-1:0] wire_d94_2;
	wire [WIDTH-1:0] wire_d94_3;
	wire [WIDTH-1:0] wire_d94_4;
	wire [WIDTH-1:0] wire_d94_5;
	wire [WIDTH-1:0] wire_d94_6;
	wire [WIDTH-1:0] wire_d94_7;
	wire [WIDTH-1:0] wire_d94_8;
	wire [WIDTH-1:0] wire_d94_9;
	wire [WIDTH-1:0] wire_d94_10;
	wire [WIDTH-1:0] wire_d94_11;
	wire [WIDTH-1:0] wire_d94_12;
	wire [WIDTH-1:0] wire_d94_13;
	wire [WIDTH-1:0] wire_d94_14;
	wire [WIDTH-1:0] wire_d94_15;
	wire [WIDTH-1:0] wire_d94_16;
	wire [WIDTH-1:0] wire_d94_17;
	wire [WIDTH-1:0] wire_d94_18;
	wire [WIDTH-1:0] wire_d94_19;
	wire [WIDTH-1:0] wire_d94_20;
	wire [WIDTH-1:0] wire_d94_21;
	wire [WIDTH-1:0] wire_d94_22;
	wire [WIDTH-1:0] wire_d94_23;
	wire [WIDTH-1:0] wire_d94_24;
	wire [WIDTH-1:0] wire_d94_25;
	wire [WIDTH-1:0] wire_d94_26;
	wire [WIDTH-1:0] wire_d94_27;
	wire [WIDTH-1:0] wire_d94_28;
	wire [WIDTH-1:0] wire_d94_29;
	wire [WIDTH-1:0] wire_d94_30;
	wire [WIDTH-1:0] wire_d94_31;
	wire [WIDTH-1:0] wire_d94_32;
	wire [WIDTH-1:0] wire_d94_33;
	wire [WIDTH-1:0] wire_d94_34;
	wire [WIDTH-1:0] wire_d94_35;
	wire [WIDTH-1:0] wire_d94_36;
	wire [WIDTH-1:0] wire_d94_37;
	wire [WIDTH-1:0] wire_d94_38;
	wire [WIDTH-1:0] wire_d94_39;
	wire [WIDTH-1:0] wire_d94_40;
	wire [WIDTH-1:0] wire_d94_41;
	wire [WIDTH-1:0] wire_d94_42;
	wire [WIDTH-1:0] wire_d94_43;
	wire [WIDTH-1:0] wire_d94_44;
	wire [WIDTH-1:0] wire_d94_45;
	wire [WIDTH-1:0] wire_d94_46;
	wire [WIDTH-1:0] wire_d94_47;
	wire [WIDTH-1:0] wire_d94_48;
	wire [WIDTH-1:0] wire_d94_49;
	wire [WIDTH-1:0] wire_d94_50;
	wire [WIDTH-1:0] wire_d94_51;
	wire [WIDTH-1:0] wire_d94_52;
	wire [WIDTH-1:0] wire_d94_53;
	wire [WIDTH-1:0] wire_d94_54;
	wire [WIDTH-1:0] wire_d94_55;
	wire [WIDTH-1:0] wire_d94_56;
	wire [WIDTH-1:0] wire_d94_57;
	wire [WIDTH-1:0] wire_d94_58;
	wire [WIDTH-1:0] wire_d94_59;
	wire [WIDTH-1:0] wire_d94_60;
	wire [WIDTH-1:0] wire_d94_61;
	wire [WIDTH-1:0] wire_d94_62;
	wire [WIDTH-1:0] wire_d94_63;
	wire [WIDTH-1:0] wire_d94_64;
	wire [WIDTH-1:0] wire_d94_65;
	wire [WIDTH-1:0] wire_d94_66;
	wire [WIDTH-1:0] wire_d94_67;
	wire [WIDTH-1:0] wire_d94_68;
	wire [WIDTH-1:0] wire_d94_69;
	wire [WIDTH-1:0] wire_d94_70;
	wire [WIDTH-1:0] wire_d94_71;
	wire [WIDTH-1:0] wire_d94_72;
	wire [WIDTH-1:0] wire_d94_73;
	wire [WIDTH-1:0] wire_d94_74;
	wire [WIDTH-1:0] wire_d94_75;
	wire [WIDTH-1:0] wire_d94_76;
	wire [WIDTH-1:0] wire_d94_77;
	wire [WIDTH-1:0] wire_d94_78;
	wire [WIDTH-1:0] wire_d95_0;
	wire [WIDTH-1:0] wire_d95_1;
	wire [WIDTH-1:0] wire_d95_2;
	wire [WIDTH-1:0] wire_d95_3;
	wire [WIDTH-1:0] wire_d95_4;
	wire [WIDTH-1:0] wire_d95_5;
	wire [WIDTH-1:0] wire_d95_6;
	wire [WIDTH-1:0] wire_d95_7;
	wire [WIDTH-1:0] wire_d95_8;
	wire [WIDTH-1:0] wire_d95_9;
	wire [WIDTH-1:0] wire_d95_10;
	wire [WIDTH-1:0] wire_d95_11;
	wire [WIDTH-1:0] wire_d95_12;
	wire [WIDTH-1:0] wire_d95_13;
	wire [WIDTH-1:0] wire_d95_14;
	wire [WIDTH-1:0] wire_d95_15;
	wire [WIDTH-1:0] wire_d95_16;
	wire [WIDTH-1:0] wire_d95_17;
	wire [WIDTH-1:0] wire_d95_18;
	wire [WIDTH-1:0] wire_d95_19;
	wire [WIDTH-1:0] wire_d95_20;
	wire [WIDTH-1:0] wire_d95_21;
	wire [WIDTH-1:0] wire_d95_22;
	wire [WIDTH-1:0] wire_d95_23;
	wire [WIDTH-1:0] wire_d95_24;
	wire [WIDTH-1:0] wire_d95_25;
	wire [WIDTH-1:0] wire_d95_26;
	wire [WIDTH-1:0] wire_d95_27;
	wire [WIDTH-1:0] wire_d95_28;
	wire [WIDTH-1:0] wire_d95_29;
	wire [WIDTH-1:0] wire_d95_30;
	wire [WIDTH-1:0] wire_d95_31;
	wire [WIDTH-1:0] wire_d95_32;
	wire [WIDTH-1:0] wire_d95_33;
	wire [WIDTH-1:0] wire_d95_34;
	wire [WIDTH-1:0] wire_d95_35;
	wire [WIDTH-1:0] wire_d95_36;
	wire [WIDTH-1:0] wire_d95_37;
	wire [WIDTH-1:0] wire_d95_38;
	wire [WIDTH-1:0] wire_d95_39;
	wire [WIDTH-1:0] wire_d95_40;
	wire [WIDTH-1:0] wire_d95_41;
	wire [WIDTH-1:0] wire_d95_42;
	wire [WIDTH-1:0] wire_d95_43;
	wire [WIDTH-1:0] wire_d95_44;
	wire [WIDTH-1:0] wire_d95_45;
	wire [WIDTH-1:0] wire_d95_46;
	wire [WIDTH-1:0] wire_d95_47;
	wire [WIDTH-1:0] wire_d95_48;
	wire [WIDTH-1:0] wire_d95_49;
	wire [WIDTH-1:0] wire_d95_50;
	wire [WIDTH-1:0] wire_d95_51;
	wire [WIDTH-1:0] wire_d95_52;
	wire [WIDTH-1:0] wire_d95_53;
	wire [WIDTH-1:0] wire_d95_54;
	wire [WIDTH-1:0] wire_d95_55;
	wire [WIDTH-1:0] wire_d95_56;
	wire [WIDTH-1:0] wire_d95_57;
	wire [WIDTH-1:0] wire_d95_58;
	wire [WIDTH-1:0] wire_d95_59;
	wire [WIDTH-1:0] wire_d95_60;
	wire [WIDTH-1:0] wire_d95_61;
	wire [WIDTH-1:0] wire_d95_62;
	wire [WIDTH-1:0] wire_d95_63;
	wire [WIDTH-1:0] wire_d95_64;
	wire [WIDTH-1:0] wire_d95_65;
	wire [WIDTH-1:0] wire_d95_66;
	wire [WIDTH-1:0] wire_d95_67;
	wire [WIDTH-1:0] wire_d95_68;
	wire [WIDTH-1:0] wire_d95_69;
	wire [WIDTH-1:0] wire_d95_70;
	wire [WIDTH-1:0] wire_d95_71;
	wire [WIDTH-1:0] wire_d95_72;
	wire [WIDTH-1:0] wire_d95_73;
	wire [WIDTH-1:0] wire_d95_74;
	wire [WIDTH-1:0] wire_d95_75;
	wire [WIDTH-1:0] wire_d95_76;
	wire [WIDTH-1:0] wire_d95_77;
	wire [WIDTH-1:0] wire_d95_78;
	wire [WIDTH-1:0] wire_d96_0;
	wire [WIDTH-1:0] wire_d96_1;
	wire [WIDTH-1:0] wire_d96_2;
	wire [WIDTH-1:0] wire_d96_3;
	wire [WIDTH-1:0] wire_d96_4;
	wire [WIDTH-1:0] wire_d96_5;
	wire [WIDTH-1:0] wire_d96_6;
	wire [WIDTH-1:0] wire_d96_7;
	wire [WIDTH-1:0] wire_d96_8;
	wire [WIDTH-1:0] wire_d96_9;
	wire [WIDTH-1:0] wire_d96_10;
	wire [WIDTH-1:0] wire_d96_11;
	wire [WIDTH-1:0] wire_d96_12;
	wire [WIDTH-1:0] wire_d96_13;
	wire [WIDTH-1:0] wire_d96_14;
	wire [WIDTH-1:0] wire_d96_15;
	wire [WIDTH-1:0] wire_d96_16;
	wire [WIDTH-1:0] wire_d96_17;
	wire [WIDTH-1:0] wire_d96_18;
	wire [WIDTH-1:0] wire_d96_19;
	wire [WIDTH-1:0] wire_d96_20;
	wire [WIDTH-1:0] wire_d96_21;
	wire [WIDTH-1:0] wire_d96_22;
	wire [WIDTH-1:0] wire_d96_23;
	wire [WIDTH-1:0] wire_d96_24;
	wire [WIDTH-1:0] wire_d96_25;
	wire [WIDTH-1:0] wire_d96_26;
	wire [WIDTH-1:0] wire_d96_27;
	wire [WIDTH-1:0] wire_d96_28;
	wire [WIDTH-1:0] wire_d96_29;
	wire [WIDTH-1:0] wire_d96_30;
	wire [WIDTH-1:0] wire_d96_31;
	wire [WIDTH-1:0] wire_d96_32;
	wire [WIDTH-1:0] wire_d96_33;
	wire [WIDTH-1:0] wire_d96_34;
	wire [WIDTH-1:0] wire_d96_35;
	wire [WIDTH-1:0] wire_d96_36;
	wire [WIDTH-1:0] wire_d96_37;
	wire [WIDTH-1:0] wire_d96_38;
	wire [WIDTH-1:0] wire_d96_39;
	wire [WIDTH-1:0] wire_d96_40;
	wire [WIDTH-1:0] wire_d96_41;
	wire [WIDTH-1:0] wire_d96_42;
	wire [WIDTH-1:0] wire_d96_43;
	wire [WIDTH-1:0] wire_d96_44;
	wire [WIDTH-1:0] wire_d96_45;
	wire [WIDTH-1:0] wire_d96_46;
	wire [WIDTH-1:0] wire_d96_47;
	wire [WIDTH-1:0] wire_d96_48;
	wire [WIDTH-1:0] wire_d96_49;
	wire [WIDTH-1:0] wire_d96_50;
	wire [WIDTH-1:0] wire_d96_51;
	wire [WIDTH-1:0] wire_d96_52;
	wire [WIDTH-1:0] wire_d96_53;
	wire [WIDTH-1:0] wire_d96_54;
	wire [WIDTH-1:0] wire_d96_55;
	wire [WIDTH-1:0] wire_d96_56;
	wire [WIDTH-1:0] wire_d96_57;
	wire [WIDTH-1:0] wire_d96_58;
	wire [WIDTH-1:0] wire_d96_59;
	wire [WIDTH-1:0] wire_d96_60;
	wire [WIDTH-1:0] wire_d96_61;
	wire [WIDTH-1:0] wire_d96_62;
	wire [WIDTH-1:0] wire_d96_63;
	wire [WIDTH-1:0] wire_d96_64;
	wire [WIDTH-1:0] wire_d96_65;
	wire [WIDTH-1:0] wire_d96_66;
	wire [WIDTH-1:0] wire_d96_67;
	wire [WIDTH-1:0] wire_d96_68;
	wire [WIDTH-1:0] wire_d96_69;
	wire [WIDTH-1:0] wire_d96_70;
	wire [WIDTH-1:0] wire_d96_71;
	wire [WIDTH-1:0] wire_d96_72;
	wire [WIDTH-1:0] wire_d96_73;
	wire [WIDTH-1:0] wire_d96_74;
	wire [WIDTH-1:0] wire_d96_75;
	wire [WIDTH-1:0] wire_d96_76;
	wire [WIDTH-1:0] wire_d96_77;
	wire [WIDTH-1:0] wire_d96_78;
	wire [WIDTH-1:0] wire_d97_0;
	wire [WIDTH-1:0] wire_d97_1;
	wire [WIDTH-1:0] wire_d97_2;
	wire [WIDTH-1:0] wire_d97_3;
	wire [WIDTH-1:0] wire_d97_4;
	wire [WIDTH-1:0] wire_d97_5;
	wire [WIDTH-1:0] wire_d97_6;
	wire [WIDTH-1:0] wire_d97_7;
	wire [WIDTH-1:0] wire_d97_8;
	wire [WIDTH-1:0] wire_d97_9;
	wire [WIDTH-1:0] wire_d97_10;
	wire [WIDTH-1:0] wire_d97_11;
	wire [WIDTH-1:0] wire_d97_12;
	wire [WIDTH-1:0] wire_d97_13;
	wire [WIDTH-1:0] wire_d97_14;
	wire [WIDTH-1:0] wire_d97_15;
	wire [WIDTH-1:0] wire_d97_16;
	wire [WIDTH-1:0] wire_d97_17;
	wire [WIDTH-1:0] wire_d97_18;
	wire [WIDTH-1:0] wire_d97_19;
	wire [WIDTH-1:0] wire_d97_20;
	wire [WIDTH-1:0] wire_d97_21;
	wire [WIDTH-1:0] wire_d97_22;
	wire [WIDTH-1:0] wire_d97_23;
	wire [WIDTH-1:0] wire_d97_24;
	wire [WIDTH-1:0] wire_d97_25;
	wire [WIDTH-1:0] wire_d97_26;
	wire [WIDTH-1:0] wire_d97_27;
	wire [WIDTH-1:0] wire_d97_28;
	wire [WIDTH-1:0] wire_d97_29;
	wire [WIDTH-1:0] wire_d97_30;
	wire [WIDTH-1:0] wire_d97_31;
	wire [WIDTH-1:0] wire_d97_32;
	wire [WIDTH-1:0] wire_d97_33;
	wire [WIDTH-1:0] wire_d97_34;
	wire [WIDTH-1:0] wire_d97_35;
	wire [WIDTH-1:0] wire_d97_36;
	wire [WIDTH-1:0] wire_d97_37;
	wire [WIDTH-1:0] wire_d97_38;
	wire [WIDTH-1:0] wire_d97_39;
	wire [WIDTH-1:0] wire_d97_40;
	wire [WIDTH-1:0] wire_d97_41;
	wire [WIDTH-1:0] wire_d97_42;
	wire [WIDTH-1:0] wire_d97_43;
	wire [WIDTH-1:0] wire_d97_44;
	wire [WIDTH-1:0] wire_d97_45;
	wire [WIDTH-1:0] wire_d97_46;
	wire [WIDTH-1:0] wire_d97_47;
	wire [WIDTH-1:0] wire_d97_48;
	wire [WIDTH-1:0] wire_d97_49;
	wire [WIDTH-1:0] wire_d97_50;
	wire [WIDTH-1:0] wire_d97_51;
	wire [WIDTH-1:0] wire_d97_52;
	wire [WIDTH-1:0] wire_d97_53;
	wire [WIDTH-1:0] wire_d97_54;
	wire [WIDTH-1:0] wire_d97_55;
	wire [WIDTH-1:0] wire_d97_56;
	wire [WIDTH-1:0] wire_d97_57;
	wire [WIDTH-1:0] wire_d97_58;
	wire [WIDTH-1:0] wire_d97_59;
	wire [WIDTH-1:0] wire_d97_60;
	wire [WIDTH-1:0] wire_d97_61;
	wire [WIDTH-1:0] wire_d97_62;
	wire [WIDTH-1:0] wire_d97_63;
	wire [WIDTH-1:0] wire_d97_64;
	wire [WIDTH-1:0] wire_d97_65;
	wire [WIDTH-1:0] wire_d97_66;
	wire [WIDTH-1:0] wire_d97_67;
	wire [WIDTH-1:0] wire_d97_68;
	wire [WIDTH-1:0] wire_d97_69;
	wire [WIDTH-1:0] wire_d97_70;
	wire [WIDTH-1:0] wire_d97_71;
	wire [WIDTH-1:0] wire_d97_72;
	wire [WIDTH-1:0] wire_d97_73;
	wire [WIDTH-1:0] wire_d97_74;
	wire [WIDTH-1:0] wire_d97_75;
	wire [WIDTH-1:0] wire_d97_76;
	wire [WIDTH-1:0] wire_d97_77;
	wire [WIDTH-1:0] wire_d97_78;
	wire [WIDTH-1:0] wire_d98_0;
	wire [WIDTH-1:0] wire_d98_1;
	wire [WIDTH-1:0] wire_d98_2;
	wire [WIDTH-1:0] wire_d98_3;
	wire [WIDTH-1:0] wire_d98_4;
	wire [WIDTH-1:0] wire_d98_5;
	wire [WIDTH-1:0] wire_d98_6;
	wire [WIDTH-1:0] wire_d98_7;
	wire [WIDTH-1:0] wire_d98_8;
	wire [WIDTH-1:0] wire_d98_9;
	wire [WIDTH-1:0] wire_d98_10;
	wire [WIDTH-1:0] wire_d98_11;
	wire [WIDTH-1:0] wire_d98_12;
	wire [WIDTH-1:0] wire_d98_13;
	wire [WIDTH-1:0] wire_d98_14;
	wire [WIDTH-1:0] wire_d98_15;
	wire [WIDTH-1:0] wire_d98_16;
	wire [WIDTH-1:0] wire_d98_17;
	wire [WIDTH-1:0] wire_d98_18;
	wire [WIDTH-1:0] wire_d98_19;
	wire [WIDTH-1:0] wire_d98_20;
	wire [WIDTH-1:0] wire_d98_21;
	wire [WIDTH-1:0] wire_d98_22;
	wire [WIDTH-1:0] wire_d98_23;
	wire [WIDTH-1:0] wire_d98_24;
	wire [WIDTH-1:0] wire_d98_25;
	wire [WIDTH-1:0] wire_d98_26;
	wire [WIDTH-1:0] wire_d98_27;
	wire [WIDTH-1:0] wire_d98_28;
	wire [WIDTH-1:0] wire_d98_29;
	wire [WIDTH-1:0] wire_d98_30;
	wire [WIDTH-1:0] wire_d98_31;
	wire [WIDTH-1:0] wire_d98_32;
	wire [WIDTH-1:0] wire_d98_33;
	wire [WIDTH-1:0] wire_d98_34;
	wire [WIDTH-1:0] wire_d98_35;
	wire [WIDTH-1:0] wire_d98_36;
	wire [WIDTH-1:0] wire_d98_37;
	wire [WIDTH-1:0] wire_d98_38;
	wire [WIDTH-1:0] wire_d98_39;
	wire [WIDTH-1:0] wire_d98_40;
	wire [WIDTH-1:0] wire_d98_41;
	wire [WIDTH-1:0] wire_d98_42;
	wire [WIDTH-1:0] wire_d98_43;
	wire [WIDTH-1:0] wire_d98_44;
	wire [WIDTH-1:0] wire_d98_45;
	wire [WIDTH-1:0] wire_d98_46;
	wire [WIDTH-1:0] wire_d98_47;
	wire [WIDTH-1:0] wire_d98_48;
	wire [WIDTH-1:0] wire_d98_49;
	wire [WIDTH-1:0] wire_d98_50;
	wire [WIDTH-1:0] wire_d98_51;
	wire [WIDTH-1:0] wire_d98_52;
	wire [WIDTH-1:0] wire_d98_53;
	wire [WIDTH-1:0] wire_d98_54;
	wire [WIDTH-1:0] wire_d98_55;
	wire [WIDTH-1:0] wire_d98_56;
	wire [WIDTH-1:0] wire_d98_57;
	wire [WIDTH-1:0] wire_d98_58;
	wire [WIDTH-1:0] wire_d98_59;
	wire [WIDTH-1:0] wire_d98_60;
	wire [WIDTH-1:0] wire_d98_61;
	wire [WIDTH-1:0] wire_d98_62;
	wire [WIDTH-1:0] wire_d98_63;
	wire [WIDTH-1:0] wire_d98_64;
	wire [WIDTH-1:0] wire_d98_65;
	wire [WIDTH-1:0] wire_d98_66;
	wire [WIDTH-1:0] wire_d98_67;
	wire [WIDTH-1:0] wire_d98_68;
	wire [WIDTH-1:0] wire_d98_69;
	wire [WIDTH-1:0] wire_d98_70;
	wire [WIDTH-1:0] wire_d98_71;
	wire [WIDTH-1:0] wire_d98_72;
	wire [WIDTH-1:0] wire_d98_73;
	wire [WIDTH-1:0] wire_d98_74;
	wire [WIDTH-1:0] wire_d98_75;
	wire [WIDTH-1:0] wire_d98_76;
	wire [WIDTH-1:0] wire_d98_77;
	wire [WIDTH-1:0] wire_d98_78;
	wire [WIDTH-1:0] wire_d99_0;
	wire [WIDTH-1:0] wire_d99_1;
	wire [WIDTH-1:0] wire_d99_2;
	wire [WIDTH-1:0] wire_d99_3;
	wire [WIDTH-1:0] wire_d99_4;
	wire [WIDTH-1:0] wire_d99_5;
	wire [WIDTH-1:0] wire_d99_6;
	wire [WIDTH-1:0] wire_d99_7;
	wire [WIDTH-1:0] wire_d99_8;
	wire [WIDTH-1:0] wire_d99_9;
	wire [WIDTH-1:0] wire_d99_10;
	wire [WIDTH-1:0] wire_d99_11;
	wire [WIDTH-1:0] wire_d99_12;
	wire [WIDTH-1:0] wire_d99_13;
	wire [WIDTH-1:0] wire_d99_14;
	wire [WIDTH-1:0] wire_d99_15;
	wire [WIDTH-1:0] wire_d99_16;
	wire [WIDTH-1:0] wire_d99_17;
	wire [WIDTH-1:0] wire_d99_18;
	wire [WIDTH-1:0] wire_d99_19;
	wire [WIDTH-1:0] wire_d99_20;
	wire [WIDTH-1:0] wire_d99_21;
	wire [WIDTH-1:0] wire_d99_22;
	wire [WIDTH-1:0] wire_d99_23;
	wire [WIDTH-1:0] wire_d99_24;
	wire [WIDTH-1:0] wire_d99_25;
	wire [WIDTH-1:0] wire_d99_26;
	wire [WIDTH-1:0] wire_d99_27;
	wire [WIDTH-1:0] wire_d99_28;
	wire [WIDTH-1:0] wire_d99_29;
	wire [WIDTH-1:0] wire_d99_30;
	wire [WIDTH-1:0] wire_d99_31;
	wire [WIDTH-1:0] wire_d99_32;
	wire [WIDTH-1:0] wire_d99_33;
	wire [WIDTH-1:0] wire_d99_34;
	wire [WIDTH-1:0] wire_d99_35;
	wire [WIDTH-1:0] wire_d99_36;
	wire [WIDTH-1:0] wire_d99_37;
	wire [WIDTH-1:0] wire_d99_38;
	wire [WIDTH-1:0] wire_d99_39;
	wire [WIDTH-1:0] wire_d99_40;
	wire [WIDTH-1:0] wire_d99_41;
	wire [WIDTH-1:0] wire_d99_42;
	wire [WIDTH-1:0] wire_d99_43;
	wire [WIDTH-1:0] wire_d99_44;
	wire [WIDTH-1:0] wire_d99_45;
	wire [WIDTH-1:0] wire_d99_46;
	wire [WIDTH-1:0] wire_d99_47;
	wire [WIDTH-1:0] wire_d99_48;
	wire [WIDTH-1:0] wire_d99_49;
	wire [WIDTH-1:0] wire_d99_50;
	wire [WIDTH-1:0] wire_d99_51;
	wire [WIDTH-1:0] wire_d99_52;
	wire [WIDTH-1:0] wire_d99_53;
	wire [WIDTH-1:0] wire_d99_54;
	wire [WIDTH-1:0] wire_d99_55;
	wire [WIDTH-1:0] wire_d99_56;
	wire [WIDTH-1:0] wire_d99_57;
	wire [WIDTH-1:0] wire_d99_58;
	wire [WIDTH-1:0] wire_d99_59;
	wire [WIDTH-1:0] wire_d99_60;
	wire [WIDTH-1:0] wire_d99_61;
	wire [WIDTH-1:0] wire_d99_62;
	wire [WIDTH-1:0] wire_d99_63;
	wire [WIDTH-1:0] wire_d99_64;
	wire [WIDTH-1:0] wire_d99_65;
	wire [WIDTH-1:0] wire_d99_66;
	wire [WIDTH-1:0] wire_d99_67;
	wire [WIDTH-1:0] wire_d99_68;
	wire [WIDTH-1:0] wire_d99_69;
	wire [WIDTH-1:0] wire_d99_70;
	wire [WIDTH-1:0] wire_d99_71;
	wire [WIDTH-1:0] wire_d99_72;
	wire [WIDTH-1:0] wire_d99_73;
	wire [WIDTH-1:0] wire_d99_74;
	wire [WIDTH-1:0] wire_d99_75;
	wire [WIDTH-1:0] wire_d99_76;
	wire [WIDTH-1:0] wire_d99_77;
	wire [WIDTH-1:0] wire_d99_78;

	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100(.data_in(d_in0),.data_out(wire_d0_0),.clk(clk),.rst(rst));            //channel 1
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance101(.data_in(wire_d0_0),.data_out(wire_d0_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance102(.data_in(wire_d0_1),.data_out(wire_d0_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance103(.data_in(wire_d0_2),.data_out(wire_d0_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance104(.data_in(wire_d0_3),.data_out(wire_d0_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance105(.data_in(wire_d0_4),.data_out(wire_d0_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance106(.data_in(wire_d0_5),.data_out(wire_d0_6),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance107(.data_in(wire_d0_6),.data_out(wire_d0_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance108(.data_in(wire_d0_7),.data_out(wire_d0_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance109(.data_in(wire_d0_8),.data_out(wire_d0_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1010(.data_in(wire_d0_9),.data_out(wire_d0_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1011(.data_in(wire_d0_10),.data_out(wire_d0_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1012(.data_in(wire_d0_11),.data_out(wire_d0_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1013(.data_in(wire_d0_12),.data_out(wire_d0_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1014(.data_in(wire_d0_13),.data_out(wire_d0_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1015(.data_in(wire_d0_14),.data_out(wire_d0_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1016(.data_in(wire_d0_15),.data_out(wire_d0_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1017(.data_in(wire_d0_16),.data_out(wire_d0_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1018(.data_in(wire_d0_17),.data_out(wire_d0_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1019(.data_in(wire_d0_18),.data_out(wire_d0_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1020(.data_in(wire_d0_19),.data_out(wire_d0_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1021(.data_in(wire_d0_20),.data_out(wire_d0_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1022(.data_in(wire_d0_21),.data_out(wire_d0_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1023(.data_in(wire_d0_22),.data_out(wire_d0_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1024(.data_in(wire_d0_23),.data_out(wire_d0_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1025(.data_in(wire_d0_24),.data_out(wire_d0_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1026(.data_in(wire_d0_25),.data_out(wire_d0_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1027(.data_in(wire_d0_26),.data_out(wire_d0_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1028(.data_in(wire_d0_27),.data_out(wire_d0_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1029(.data_in(wire_d0_28),.data_out(wire_d0_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1030(.data_in(wire_d0_29),.data_out(wire_d0_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1031(.data_in(wire_d0_30),.data_out(wire_d0_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1032(.data_in(wire_d0_31),.data_out(wire_d0_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1033(.data_in(wire_d0_32),.data_out(wire_d0_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1034(.data_in(wire_d0_33),.data_out(wire_d0_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1035(.data_in(wire_d0_34),.data_out(wire_d0_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1036(.data_in(wire_d0_35),.data_out(wire_d0_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1037(.data_in(wire_d0_36),.data_out(wire_d0_37),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1038(.data_in(wire_d0_37),.data_out(wire_d0_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1039(.data_in(wire_d0_38),.data_out(wire_d0_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1040(.data_in(wire_d0_39),.data_out(wire_d0_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1041(.data_in(wire_d0_40),.data_out(wire_d0_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1042(.data_in(wire_d0_41),.data_out(wire_d0_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1043(.data_in(wire_d0_42),.data_out(wire_d0_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1044(.data_in(wire_d0_43),.data_out(wire_d0_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1045(.data_in(wire_d0_44),.data_out(wire_d0_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1046(.data_in(wire_d0_45),.data_out(wire_d0_46),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1047(.data_in(wire_d0_46),.data_out(wire_d0_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1048(.data_in(wire_d0_47),.data_out(wire_d0_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1049(.data_in(wire_d0_48),.data_out(wire_d0_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1050(.data_in(wire_d0_49),.data_out(wire_d0_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1051(.data_in(wire_d0_50),.data_out(wire_d0_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1052(.data_in(wire_d0_51),.data_out(wire_d0_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1053(.data_in(wire_d0_52),.data_out(wire_d0_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1054(.data_in(wire_d0_53),.data_out(wire_d0_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1055(.data_in(wire_d0_54),.data_out(wire_d0_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1056(.data_in(wire_d0_55),.data_out(wire_d0_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1057(.data_in(wire_d0_56),.data_out(wire_d0_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1058(.data_in(wire_d0_57),.data_out(wire_d0_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1059(.data_in(wire_d0_58),.data_out(wire_d0_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1060(.data_in(wire_d0_59),.data_out(wire_d0_60),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1061(.data_in(wire_d0_60),.data_out(wire_d0_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1062(.data_in(wire_d0_61),.data_out(wire_d0_62),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1063(.data_in(wire_d0_62),.data_out(wire_d0_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1064(.data_in(wire_d0_63),.data_out(wire_d0_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1065(.data_in(wire_d0_64),.data_out(wire_d0_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1066(.data_in(wire_d0_65),.data_out(wire_d0_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1067(.data_in(wire_d0_66),.data_out(wire_d0_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1068(.data_in(wire_d0_67),.data_out(wire_d0_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1069(.data_in(wire_d0_68),.data_out(wire_d0_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1070(.data_in(wire_d0_69),.data_out(wire_d0_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1071(.data_in(wire_d0_70),.data_out(wire_d0_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1072(.data_in(wire_d0_71),.data_out(wire_d0_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1073(.data_in(wire_d0_72),.data_out(wire_d0_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1074(.data_in(wire_d0_73),.data_out(wire_d0_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1075(.data_in(wire_d0_74),.data_out(wire_d0_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1076(.data_in(wire_d0_75),.data_out(wire_d0_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1077(.data_in(wire_d0_76),.data_out(wire_d0_77),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1078(.data_in(wire_d0_77),.data_out(wire_d0_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1079(.data_in(wire_d0_78),.data_out(d_out0),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance210(.data_in(d_in1),.data_out(wire_d1_0),.clk(clk),.rst(rst));            //channel 2
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance211(.data_in(wire_d1_0),.data_out(wire_d1_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance212(.data_in(wire_d1_1),.data_out(wire_d1_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance213(.data_in(wire_d1_2),.data_out(wire_d1_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance214(.data_in(wire_d1_3),.data_out(wire_d1_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance215(.data_in(wire_d1_4),.data_out(wire_d1_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance216(.data_in(wire_d1_5),.data_out(wire_d1_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance217(.data_in(wire_d1_6),.data_out(wire_d1_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance218(.data_in(wire_d1_7),.data_out(wire_d1_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance219(.data_in(wire_d1_8),.data_out(wire_d1_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2110(.data_in(wire_d1_9),.data_out(wire_d1_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2111(.data_in(wire_d1_10),.data_out(wire_d1_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2112(.data_in(wire_d1_11),.data_out(wire_d1_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2113(.data_in(wire_d1_12),.data_out(wire_d1_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2114(.data_in(wire_d1_13),.data_out(wire_d1_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2115(.data_in(wire_d1_14),.data_out(wire_d1_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2116(.data_in(wire_d1_15),.data_out(wire_d1_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2117(.data_in(wire_d1_16),.data_out(wire_d1_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2118(.data_in(wire_d1_17),.data_out(wire_d1_18),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2119(.data_in(wire_d1_18),.data_out(wire_d1_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2120(.data_in(wire_d1_19),.data_out(wire_d1_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2121(.data_in(wire_d1_20),.data_out(wire_d1_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2122(.data_in(wire_d1_21),.data_out(wire_d1_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2123(.data_in(wire_d1_22),.data_out(wire_d1_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2124(.data_in(wire_d1_23),.data_out(wire_d1_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2125(.data_in(wire_d1_24),.data_out(wire_d1_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2126(.data_in(wire_d1_25),.data_out(wire_d1_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2127(.data_in(wire_d1_26),.data_out(wire_d1_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2128(.data_in(wire_d1_27),.data_out(wire_d1_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2129(.data_in(wire_d1_28),.data_out(wire_d1_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2130(.data_in(wire_d1_29),.data_out(wire_d1_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2131(.data_in(wire_d1_30),.data_out(wire_d1_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2132(.data_in(wire_d1_31),.data_out(wire_d1_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2133(.data_in(wire_d1_32),.data_out(wire_d1_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2134(.data_in(wire_d1_33),.data_out(wire_d1_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2135(.data_in(wire_d1_34),.data_out(wire_d1_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2136(.data_in(wire_d1_35),.data_out(wire_d1_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2137(.data_in(wire_d1_36),.data_out(wire_d1_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2138(.data_in(wire_d1_37),.data_out(wire_d1_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2139(.data_in(wire_d1_38),.data_out(wire_d1_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2140(.data_in(wire_d1_39),.data_out(wire_d1_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2141(.data_in(wire_d1_40),.data_out(wire_d1_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2142(.data_in(wire_d1_41),.data_out(wire_d1_42),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2143(.data_in(wire_d1_42),.data_out(wire_d1_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2144(.data_in(wire_d1_43),.data_out(wire_d1_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2145(.data_in(wire_d1_44),.data_out(wire_d1_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2146(.data_in(wire_d1_45),.data_out(wire_d1_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2147(.data_in(wire_d1_46),.data_out(wire_d1_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2148(.data_in(wire_d1_47),.data_out(wire_d1_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2149(.data_in(wire_d1_48),.data_out(wire_d1_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2150(.data_in(wire_d1_49),.data_out(wire_d1_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2151(.data_in(wire_d1_50),.data_out(wire_d1_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2152(.data_in(wire_d1_51),.data_out(wire_d1_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2153(.data_in(wire_d1_52),.data_out(wire_d1_53),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2154(.data_in(wire_d1_53),.data_out(wire_d1_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2155(.data_in(wire_d1_54),.data_out(wire_d1_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2156(.data_in(wire_d1_55),.data_out(wire_d1_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2157(.data_in(wire_d1_56),.data_out(wire_d1_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2158(.data_in(wire_d1_57),.data_out(wire_d1_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2159(.data_in(wire_d1_58),.data_out(wire_d1_59),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2160(.data_in(wire_d1_59),.data_out(wire_d1_60),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2161(.data_in(wire_d1_60),.data_out(wire_d1_61),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2162(.data_in(wire_d1_61),.data_out(wire_d1_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2163(.data_in(wire_d1_62),.data_out(wire_d1_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2164(.data_in(wire_d1_63),.data_out(wire_d1_64),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2165(.data_in(wire_d1_64),.data_out(wire_d1_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2166(.data_in(wire_d1_65),.data_out(wire_d1_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2167(.data_in(wire_d1_66),.data_out(wire_d1_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2168(.data_in(wire_d1_67),.data_out(wire_d1_68),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2169(.data_in(wire_d1_68),.data_out(wire_d1_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2170(.data_in(wire_d1_69),.data_out(wire_d1_70),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2171(.data_in(wire_d1_70),.data_out(wire_d1_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2172(.data_in(wire_d1_71),.data_out(wire_d1_72),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2173(.data_in(wire_d1_72),.data_out(wire_d1_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2174(.data_in(wire_d1_73),.data_out(wire_d1_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2175(.data_in(wire_d1_74),.data_out(wire_d1_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2176(.data_in(wire_d1_75),.data_out(wire_d1_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2177(.data_in(wire_d1_76),.data_out(wire_d1_77),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2178(.data_in(wire_d1_77),.data_out(wire_d1_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2179(.data_in(wire_d1_78),.data_out(d_out1),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance320(.data_in(d_in2),.data_out(wire_d2_0),.clk(clk),.rst(rst));            //channel 3
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance321(.data_in(wire_d2_0),.data_out(wire_d2_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance322(.data_in(wire_d2_1),.data_out(wire_d2_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance323(.data_in(wire_d2_2),.data_out(wire_d2_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance324(.data_in(wire_d2_3),.data_out(wire_d2_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance325(.data_in(wire_d2_4),.data_out(wire_d2_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance326(.data_in(wire_d2_5),.data_out(wire_d2_6),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance327(.data_in(wire_d2_6),.data_out(wire_d2_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance328(.data_in(wire_d2_7),.data_out(wire_d2_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance329(.data_in(wire_d2_8),.data_out(wire_d2_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3210(.data_in(wire_d2_9),.data_out(wire_d2_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3211(.data_in(wire_d2_10),.data_out(wire_d2_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3212(.data_in(wire_d2_11),.data_out(wire_d2_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3213(.data_in(wire_d2_12),.data_out(wire_d2_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3214(.data_in(wire_d2_13),.data_out(wire_d2_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3215(.data_in(wire_d2_14),.data_out(wire_d2_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3216(.data_in(wire_d2_15),.data_out(wire_d2_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3217(.data_in(wire_d2_16),.data_out(wire_d2_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3218(.data_in(wire_d2_17),.data_out(wire_d2_18),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3219(.data_in(wire_d2_18),.data_out(wire_d2_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3220(.data_in(wire_d2_19),.data_out(wire_d2_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3221(.data_in(wire_d2_20),.data_out(wire_d2_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3222(.data_in(wire_d2_21),.data_out(wire_d2_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3223(.data_in(wire_d2_22),.data_out(wire_d2_23),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3224(.data_in(wire_d2_23),.data_out(wire_d2_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3225(.data_in(wire_d2_24),.data_out(wire_d2_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3226(.data_in(wire_d2_25),.data_out(wire_d2_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3227(.data_in(wire_d2_26),.data_out(wire_d2_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3228(.data_in(wire_d2_27),.data_out(wire_d2_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3229(.data_in(wire_d2_28),.data_out(wire_d2_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3230(.data_in(wire_d2_29),.data_out(wire_d2_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3231(.data_in(wire_d2_30),.data_out(wire_d2_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3232(.data_in(wire_d2_31),.data_out(wire_d2_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3233(.data_in(wire_d2_32),.data_out(wire_d2_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3234(.data_in(wire_d2_33),.data_out(wire_d2_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3235(.data_in(wire_d2_34),.data_out(wire_d2_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3236(.data_in(wire_d2_35),.data_out(wire_d2_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3237(.data_in(wire_d2_36),.data_out(wire_d2_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3238(.data_in(wire_d2_37),.data_out(wire_d2_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3239(.data_in(wire_d2_38),.data_out(wire_d2_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3240(.data_in(wire_d2_39),.data_out(wire_d2_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3241(.data_in(wire_d2_40),.data_out(wire_d2_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3242(.data_in(wire_d2_41),.data_out(wire_d2_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3243(.data_in(wire_d2_42),.data_out(wire_d2_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3244(.data_in(wire_d2_43),.data_out(wire_d2_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3245(.data_in(wire_d2_44),.data_out(wire_d2_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3246(.data_in(wire_d2_45),.data_out(wire_d2_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3247(.data_in(wire_d2_46),.data_out(wire_d2_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3248(.data_in(wire_d2_47),.data_out(wire_d2_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3249(.data_in(wire_d2_48),.data_out(wire_d2_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3250(.data_in(wire_d2_49),.data_out(wire_d2_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3251(.data_in(wire_d2_50),.data_out(wire_d2_51),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3252(.data_in(wire_d2_51),.data_out(wire_d2_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3253(.data_in(wire_d2_52),.data_out(wire_d2_53),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3254(.data_in(wire_d2_53),.data_out(wire_d2_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3255(.data_in(wire_d2_54),.data_out(wire_d2_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3256(.data_in(wire_d2_55),.data_out(wire_d2_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3257(.data_in(wire_d2_56),.data_out(wire_d2_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3258(.data_in(wire_d2_57),.data_out(wire_d2_58),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3259(.data_in(wire_d2_58),.data_out(wire_d2_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3260(.data_in(wire_d2_59),.data_out(wire_d2_60),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3261(.data_in(wire_d2_60),.data_out(wire_d2_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3262(.data_in(wire_d2_61),.data_out(wire_d2_62),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3263(.data_in(wire_d2_62),.data_out(wire_d2_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3264(.data_in(wire_d2_63),.data_out(wire_d2_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3265(.data_in(wire_d2_64),.data_out(wire_d2_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3266(.data_in(wire_d2_65),.data_out(wire_d2_66),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3267(.data_in(wire_d2_66),.data_out(wire_d2_67),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3268(.data_in(wire_d2_67),.data_out(wire_d2_68),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3269(.data_in(wire_d2_68),.data_out(wire_d2_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3270(.data_in(wire_d2_69),.data_out(wire_d2_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3271(.data_in(wire_d2_70),.data_out(wire_d2_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3272(.data_in(wire_d2_71),.data_out(wire_d2_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3273(.data_in(wire_d2_72),.data_out(wire_d2_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3274(.data_in(wire_d2_73),.data_out(wire_d2_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3275(.data_in(wire_d2_74),.data_out(wire_d2_75),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3276(.data_in(wire_d2_75),.data_out(wire_d2_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3277(.data_in(wire_d2_76),.data_out(wire_d2_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3278(.data_in(wire_d2_77),.data_out(wire_d2_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3279(.data_in(wire_d2_78),.data_out(d_out2),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance430(.data_in(d_in3),.data_out(wire_d3_0),.clk(clk),.rst(rst));            //channel 4
	large_mux #(.WIDTH(WIDTH)) large_mux_instance431(.data_in(wire_d3_0),.data_out(wire_d3_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance432(.data_in(wire_d3_1),.data_out(wire_d3_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance433(.data_in(wire_d3_2),.data_out(wire_d3_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance434(.data_in(wire_d3_3),.data_out(wire_d3_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance435(.data_in(wire_d3_4),.data_out(wire_d3_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance436(.data_in(wire_d3_5),.data_out(wire_d3_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance437(.data_in(wire_d3_6),.data_out(wire_d3_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance438(.data_in(wire_d3_7),.data_out(wire_d3_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance439(.data_in(wire_d3_8),.data_out(wire_d3_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4310(.data_in(wire_d3_9),.data_out(wire_d3_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4311(.data_in(wire_d3_10),.data_out(wire_d3_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4312(.data_in(wire_d3_11),.data_out(wire_d3_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4313(.data_in(wire_d3_12),.data_out(wire_d3_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4314(.data_in(wire_d3_13),.data_out(wire_d3_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4315(.data_in(wire_d3_14),.data_out(wire_d3_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4316(.data_in(wire_d3_15),.data_out(wire_d3_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4317(.data_in(wire_d3_16),.data_out(wire_d3_17),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4318(.data_in(wire_d3_17),.data_out(wire_d3_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4319(.data_in(wire_d3_18),.data_out(wire_d3_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4320(.data_in(wire_d3_19),.data_out(wire_d3_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4321(.data_in(wire_d3_20),.data_out(wire_d3_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4322(.data_in(wire_d3_21),.data_out(wire_d3_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4323(.data_in(wire_d3_22),.data_out(wire_d3_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4324(.data_in(wire_d3_23),.data_out(wire_d3_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4325(.data_in(wire_d3_24),.data_out(wire_d3_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4326(.data_in(wire_d3_25),.data_out(wire_d3_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4327(.data_in(wire_d3_26),.data_out(wire_d3_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4328(.data_in(wire_d3_27),.data_out(wire_d3_28),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4329(.data_in(wire_d3_28),.data_out(wire_d3_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4330(.data_in(wire_d3_29),.data_out(wire_d3_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4331(.data_in(wire_d3_30),.data_out(wire_d3_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4332(.data_in(wire_d3_31),.data_out(wire_d3_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4333(.data_in(wire_d3_32),.data_out(wire_d3_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4334(.data_in(wire_d3_33),.data_out(wire_d3_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4335(.data_in(wire_d3_34),.data_out(wire_d3_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4336(.data_in(wire_d3_35),.data_out(wire_d3_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4337(.data_in(wire_d3_36),.data_out(wire_d3_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4338(.data_in(wire_d3_37),.data_out(wire_d3_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4339(.data_in(wire_d3_38),.data_out(wire_d3_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4340(.data_in(wire_d3_39),.data_out(wire_d3_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4341(.data_in(wire_d3_40),.data_out(wire_d3_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4342(.data_in(wire_d3_41),.data_out(wire_d3_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4343(.data_in(wire_d3_42),.data_out(wire_d3_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4344(.data_in(wire_d3_43),.data_out(wire_d3_44),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4345(.data_in(wire_d3_44),.data_out(wire_d3_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4346(.data_in(wire_d3_45),.data_out(wire_d3_46),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4347(.data_in(wire_d3_46),.data_out(wire_d3_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4348(.data_in(wire_d3_47),.data_out(wire_d3_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4349(.data_in(wire_d3_48),.data_out(wire_d3_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4350(.data_in(wire_d3_49),.data_out(wire_d3_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4351(.data_in(wire_d3_50),.data_out(wire_d3_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4352(.data_in(wire_d3_51),.data_out(wire_d3_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4353(.data_in(wire_d3_52),.data_out(wire_d3_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4354(.data_in(wire_d3_53),.data_out(wire_d3_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4355(.data_in(wire_d3_54),.data_out(wire_d3_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4356(.data_in(wire_d3_55),.data_out(wire_d3_56),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4357(.data_in(wire_d3_56),.data_out(wire_d3_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4358(.data_in(wire_d3_57),.data_out(wire_d3_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4359(.data_in(wire_d3_58),.data_out(wire_d3_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4360(.data_in(wire_d3_59),.data_out(wire_d3_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4361(.data_in(wire_d3_60),.data_out(wire_d3_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4362(.data_in(wire_d3_61),.data_out(wire_d3_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4363(.data_in(wire_d3_62),.data_out(wire_d3_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4364(.data_in(wire_d3_63),.data_out(wire_d3_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4365(.data_in(wire_d3_64),.data_out(wire_d3_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4366(.data_in(wire_d3_65),.data_out(wire_d3_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4367(.data_in(wire_d3_66),.data_out(wire_d3_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4368(.data_in(wire_d3_67),.data_out(wire_d3_68),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4369(.data_in(wire_d3_68),.data_out(wire_d3_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4370(.data_in(wire_d3_69),.data_out(wire_d3_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4371(.data_in(wire_d3_70),.data_out(wire_d3_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4372(.data_in(wire_d3_71),.data_out(wire_d3_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4373(.data_in(wire_d3_72),.data_out(wire_d3_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4374(.data_in(wire_d3_73),.data_out(wire_d3_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4375(.data_in(wire_d3_74),.data_out(wire_d3_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4376(.data_in(wire_d3_75),.data_out(wire_d3_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4377(.data_in(wire_d3_76),.data_out(wire_d3_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4378(.data_in(wire_d3_77),.data_out(wire_d3_78),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4379(.data_in(wire_d3_78),.data_out(d_out3),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance540(.data_in(d_in4),.data_out(wire_d4_0),.clk(clk),.rst(rst));            //channel 5
	register #(.WIDTH(WIDTH)) register_instance541(.data_in(wire_d4_0),.data_out(wire_d4_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance542(.data_in(wire_d4_1),.data_out(wire_d4_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance543(.data_in(wire_d4_2),.data_out(wire_d4_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance544(.data_in(wire_d4_3),.data_out(wire_d4_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance545(.data_in(wire_d4_4),.data_out(wire_d4_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance546(.data_in(wire_d4_5),.data_out(wire_d4_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance547(.data_in(wire_d4_6),.data_out(wire_d4_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance548(.data_in(wire_d4_7),.data_out(wire_d4_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance549(.data_in(wire_d4_8),.data_out(wire_d4_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5410(.data_in(wire_d4_9),.data_out(wire_d4_10),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5411(.data_in(wire_d4_10),.data_out(wire_d4_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5412(.data_in(wire_d4_11),.data_out(wire_d4_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5413(.data_in(wire_d4_12),.data_out(wire_d4_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5414(.data_in(wire_d4_13),.data_out(wire_d4_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5415(.data_in(wire_d4_14),.data_out(wire_d4_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5416(.data_in(wire_d4_15),.data_out(wire_d4_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5417(.data_in(wire_d4_16),.data_out(wire_d4_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5418(.data_in(wire_d4_17),.data_out(wire_d4_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5419(.data_in(wire_d4_18),.data_out(wire_d4_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5420(.data_in(wire_d4_19),.data_out(wire_d4_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5421(.data_in(wire_d4_20),.data_out(wire_d4_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5422(.data_in(wire_d4_21),.data_out(wire_d4_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5423(.data_in(wire_d4_22),.data_out(wire_d4_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5424(.data_in(wire_d4_23),.data_out(wire_d4_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5425(.data_in(wire_d4_24),.data_out(wire_d4_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5426(.data_in(wire_d4_25),.data_out(wire_d4_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5427(.data_in(wire_d4_26),.data_out(wire_d4_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5428(.data_in(wire_d4_27),.data_out(wire_d4_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5429(.data_in(wire_d4_28),.data_out(wire_d4_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5430(.data_in(wire_d4_29),.data_out(wire_d4_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5431(.data_in(wire_d4_30),.data_out(wire_d4_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5432(.data_in(wire_d4_31),.data_out(wire_d4_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5433(.data_in(wire_d4_32),.data_out(wire_d4_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5434(.data_in(wire_d4_33),.data_out(wire_d4_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5435(.data_in(wire_d4_34),.data_out(wire_d4_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5436(.data_in(wire_d4_35),.data_out(wire_d4_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5437(.data_in(wire_d4_36),.data_out(wire_d4_37),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5438(.data_in(wire_d4_37),.data_out(wire_d4_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5439(.data_in(wire_d4_38),.data_out(wire_d4_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5440(.data_in(wire_d4_39),.data_out(wire_d4_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5441(.data_in(wire_d4_40),.data_out(wire_d4_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5442(.data_in(wire_d4_41),.data_out(wire_d4_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5443(.data_in(wire_d4_42),.data_out(wire_d4_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5444(.data_in(wire_d4_43),.data_out(wire_d4_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5445(.data_in(wire_d4_44),.data_out(wire_d4_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5446(.data_in(wire_d4_45),.data_out(wire_d4_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5447(.data_in(wire_d4_46),.data_out(wire_d4_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5448(.data_in(wire_d4_47),.data_out(wire_d4_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5449(.data_in(wire_d4_48),.data_out(wire_d4_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5450(.data_in(wire_d4_49),.data_out(wire_d4_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5451(.data_in(wire_d4_50),.data_out(wire_d4_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5452(.data_in(wire_d4_51),.data_out(wire_d4_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5453(.data_in(wire_d4_52),.data_out(wire_d4_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5454(.data_in(wire_d4_53),.data_out(wire_d4_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5455(.data_in(wire_d4_54),.data_out(wire_d4_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5456(.data_in(wire_d4_55),.data_out(wire_d4_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5457(.data_in(wire_d4_56),.data_out(wire_d4_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5458(.data_in(wire_d4_57),.data_out(wire_d4_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5459(.data_in(wire_d4_58),.data_out(wire_d4_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5460(.data_in(wire_d4_59),.data_out(wire_d4_60),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5461(.data_in(wire_d4_60),.data_out(wire_d4_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5462(.data_in(wire_d4_61),.data_out(wire_d4_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5463(.data_in(wire_d4_62),.data_out(wire_d4_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5464(.data_in(wire_d4_63),.data_out(wire_d4_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5465(.data_in(wire_d4_64),.data_out(wire_d4_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5466(.data_in(wire_d4_65),.data_out(wire_d4_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5467(.data_in(wire_d4_66),.data_out(wire_d4_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5468(.data_in(wire_d4_67),.data_out(wire_d4_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5469(.data_in(wire_d4_68),.data_out(wire_d4_69),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5470(.data_in(wire_d4_69),.data_out(wire_d4_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5471(.data_in(wire_d4_70),.data_out(wire_d4_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5472(.data_in(wire_d4_71),.data_out(wire_d4_72),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5473(.data_in(wire_d4_72),.data_out(wire_d4_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5474(.data_in(wire_d4_73),.data_out(wire_d4_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5475(.data_in(wire_d4_74),.data_out(wire_d4_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5476(.data_in(wire_d4_75),.data_out(wire_d4_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5477(.data_in(wire_d4_76),.data_out(wire_d4_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5478(.data_in(wire_d4_77),.data_out(wire_d4_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5479(.data_in(wire_d4_78),.data_out(d_out4),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance650(.data_in(d_in5),.data_out(wire_d5_0),.clk(clk),.rst(rst));            //channel 6
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance651(.data_in(wire_d5_0),.data_out(wire_d5_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance652(.data_in(wire_d5_1),.data_out(wire_d5_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance653(.data_in(wire_d5_2),.data_out(wire_d5_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance654(.data_in(wire_d5_3),.data_out(wire_d5_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance655(.data_in(wire_d5_4),.data_out(wire_d5_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance656(.data_in(wire_d5_5),.data_out(wire_d5_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance657(.data_in(wire_d5_6),.data_out(wire_d5_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance658(.data_in(wire_d5_7),.data_out(wire_d5_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance659(.data_in(wire_d5_8),.data_out(wire_d5_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6510(.data_in(wire_d5_9),.data_out(wire_d5_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6511(.data_in(wire_d5_10),.data_out(wire_d5_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6512(.data_in(wire_d5_11),.data_out(wire_d5_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6513(.data_in(wire_d5_12),.data_out(wire_d5_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6514(.data_in(wire_d5_13),.data_out(wire_d5_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6515(.data_in(wire_d5_14),.data_out(wire_d5_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6516(.data_in(wire_d5_15),.data_out(wire_d5_16),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6517(.data_in(wire_d5_16),.data_out(wire_d5_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6518(.data_in(wire_d5_17),.data_out(wire_d5_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6519(.data_in(wire_d5_18),.data_out(wire_d5_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6520(.data_in(wire_d5_19),.data_out(wire_d5_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6521(.data_in(wire_d5_20),.data_out(wire_d5_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6522(.data_in(wire_d5_21),.data_out(wire_d5_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6523(.data_in(wire_d5_22),.data_out(wire_d5_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6524(.data_in(wire_d5_23),.data_out(wire_d5_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6525(.data_in(wire_d5_24),.data_out(wire_d5_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6526(.data_in(wire_d5_25),.data_out(wire_d5_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6527(.data_in(wire_d5_26),.data_out(wire_d5_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6528(.data_in(wire_d5_27),.data_out(wire_d5_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6529(.data_in(wire_d5_28),.data_out(wire_d5_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6530(.data_in(wire_d5_29),.data_out(wire_d5_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6531(.data_in(wire_d5_30),.data_out(wire_d5_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6532(.data_in(wire_d5_31),.data_out(wire_d5_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6533(.data_in(wire_d5_32),.data_out(wire_d5_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6534(.data_in(wire_d5_33),.data_out(wire_d5_34),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6535(.data_in(wire_d5_34),.data_out(wire_d5_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6536(.data_in(wire_d5_35),.data_out(wire_d5_36),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6537(.data_in(wire_d5_36),.data_out(wire_d5_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6538(.data_in(wire_d5_37),.data_out(wire_d5_38),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6539(.data_in(wire_d5_38),.data_out(wire_d5_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6540(.data_in(wire_d5_39),.data_out(wire_d5_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6541(.data_in(wire_d5_40),.data_out(wire_d5_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6542(.data_in(wire_d5_41),.data_out(wire_d5_42),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6543(.data_in(wire_d5_42),.data_out(wire_d5_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6544(.data_in(wire_d5_43),.data_out(wire_d5_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6545(.data_in(wire_d5_44),.data_out(wire_d5_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6546(.data_in(wire_d5_45),.data_out(wire_d5_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6547(.data_in(wire_d5_46),.data_out(wire_d5_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6548(.data_in(wire_d5_47),.data_out(wire_d5_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6549(.data_in(wire_d5_48),.data_out(wire_d5_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6550(.data_in(wire_d5_49),.data_out(wire_d5_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6551(.data_in(wire_d5_50),.data_out(wire_d5_51),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6552(.data_in(wire_d5_51),.data_out(wire_d5_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6553(.data_in(wire_d5_52),.data_out(wire_d5_53),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6554(.data_in(wire_d5_53),.data_out(wire_d5_54),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6555(.data_in(wire_d5_54),.data_out(wire_d5_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6556(.data_in(wire_d5_55),.data_out(wire_d5_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6557(.data_in(wire_d5_56),.data_out(wire_d5_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6558(.data_in(wire_d5_57),.data_out(wire_d5_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6559(.data_in(wire_d5_58),.data_out(wire_d5_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6560(.data_in(wire_d5_59),.data_out(wire_d5_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6561(.data_in(wire_d5_60),.data_out(wire_d5_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6562(.data_in(wire_d5_61),.data_out(wire_d5_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6563(.data_in(wire_d5_62),.data_out(wire_d5_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6564(.data_in(wire_d5_63),.data_out(wire_d5_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6565(.data_in(wire_d5_64),.data_out(wire_d5_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6566(.data_in(wire_d5_65),.data_out(wire_d5_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6567(.data_in(wire_d5_66),.data_out(wire_d5_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6568(.data_in(wire_d5_67),.data_out(wire_d5_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6569(.data_in(wire_d5_68),.data_out(wire_d5_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6570(.data_in(wire_d5_69),.data_out(wire_d5_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6571(.data_in(wire_d5_70),.data_out(wire_d5_71),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6572(.data_in(wire_d5_71),.data_out(wire_d5_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6573(.data_in(wire_d5_72),.data_out(wire_d5_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6574(.data_in(wire_d5_73),.data_out(wire_d5_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6575(.data_in(wire_d5_74),.data_out(wire_d5_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6576(.data_in(wire_d5_75),.data_out(wire_d5_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6577(.data_in(wire_d5_76),.data_out(wire_d5_77),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6578(.data_in(wire_d5_77),.data_out(wire_d5_78),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6579(.data_in(wire_d5_78),.data_out(d_out5),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance760(.data_in(d_in6),.data_out(wire_d6_0),.clk(clk),.rst(rst));            //channel 7
	decoder_top #(.WIDTH(WIDTH)) decoder_instance761(.data_in(wire_d6_0),.data_out(wire_d6_1),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance762(.data_in(wire_d6_1),.data_out(wire_d6_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance763(.data_in(wire_d6_2),.data_out(wire_d6_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance764(.data_in(wire_d6_3),.data_out(wire_d6_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance765(.data_in(wire_d6_4),.data_out(wire_d6_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance766(.data_in(wire_d6_5),.data_out(wire_d6_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767(.data_in(wire_d6_6),.data_out(wire_d6_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance768(.data_in(wire_d6_7),.data_out(wire_d6_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance769(.data_in(wire_d6_8),.data_out(wire_d6_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7610(.data_in(wire_d6_9),.data_out(wire_d6_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7611(.data_in(wire_d6_10),.data_out(wire_d6_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7612(.data_in(wire_d6_11),.data_out(wire_d6_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7613(.data_in(wire_d6_12),.data_out(wire_d6_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7614(.data_in(wire_d6_13),.data_out(wire_d6_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7615(.data_in(wire_d6_14),.data_out(wire_d6_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7616(.data_in(wire_d6_15),.data_out(wire_d6_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7617(.data_in(wire_d6_16),.data_out(wire_d6_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7618(.data_in(wire_d6_17),.data_out(wire_d6_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7619(.data_in(wire_d6_18),.data_out(wire_d6_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7620(.data_in(wire_d6_19),.data_out(wire_d6_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7621(.data_in(wire_d6_20),.data_out(wire_d6_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7622(.data_in(wire_d6_21),.data_out(wire_d6_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7623(.data_in(wire_d6_22),.data_out(wire_d6_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7624(.data_in(wire_d6_23),.data_out(wire_d6_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7625(.data_in(wire_d6_24),.data_out(wire_d6_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7626(.data_in(wire_d6_25),.data_out(wire_d6_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7627(.data_in(wire_d6_26),.data_out(wire_d6_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7628(.data_in(wire_d6_27),.data_out(wire_d6_28),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7629(.data_in(wire_d6_28),.data_out(wire_d6_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7630(.data_in(wire_d6_29),.data_out(wire_d6_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7631(.data_in(wire_d6_30),.data_out(wire_d6_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7632(.data_in(wire_d6_31),.data_out(wire_d6_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7633(.data_in(wire_d6_32),.data_out(wire_d6_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7634(.data_in(wire_d6_33),.data_out(wire_d6_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7635(.data_in(wire_d6_34),.data_out(wire_d6_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7636(.data_in(wire_d6_35),.data_out(wire_d6_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7637(.data_in(wire_d6_36),.data_out(wire_d6_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7638(.data_in(wire_d6_37),.data_out(wire_d6_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7639(.data_in(wire_d6_38),.data_out(wire_d6_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7640(.data_in(wire_d6_39),.data_out(wire_d6_40),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7641(.data_in(wire_d6_40),.data_out(wire_d6_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7642(.data_in(wire_d6_41),.data_out(wire_d6_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7643(.data_in(wire_d6_42),.data_out(wire_d6_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7644(.data_in(wire_d6_43),.data_out(wire_d6_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7645(.data_in(wire_d6_44),.data_out(wire_d6_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7646(.data_in(wire_d6_45),.data_out(wire_d6_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7647(.data_in(wire_d6_46),.data_out(wire_d6_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7648(.data_in(wire_d6_47),.data_out(wire_d6_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7649(.data_in(wire_d6_48),.data_out(wire_d6_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7650(.data_in(wire_d6_49),.data_out(wire_d6_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7651(.data_in(wire_d6_50),.data_out(wire_d6_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7652(.data_in(wire_d6_51),.data_out(wire_d6_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7653(.data_in(wire_d6_52),.data_out(wire_d6_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7654(.data_in(wire_d6_53),.data_out(wire_d6_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7655(.data_in(wire_d6_54),.data_out(wire_d6_55),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7656(.data_in(wire_d6_55),.data_out(wire_d6_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7657(.data_in(wire_d6_56),.data_out(wire_d6_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7658(.data_in(wire_d6_57),.data_out(wire_d6_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7659(.data_in(wire_d6_58),.data_out(wire_d6_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7660(.data_in(wire_d6_59),.data_out(wire_d6_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7661(.data_in(wire_d6_60),.data_out(wire_d6_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7662(.data_in(wire_d6_61),.data_out(wire_d6_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7663(.data_in(wire_d6_62),.data_out(wire_d6_63),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7664(.data_in(wire_d6_63),.data_out(wire_d6_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7665(.data_in(wire_d6_64),.data_out(wire_d6_65),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7666(.data_in(wire_d6_65),.data_out(wire_d6_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7667(.data_in(wire_d6_66),.data_out(wire_d6_67),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7668(.data_in(wire_d6_67),.data_out(wire_d6_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7669(.data_in(wire_d6_68),.data_out(wire_d6_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7670(.data_in(wire_d6_69),.data_out(wire_d6_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7671(.data_in(wire_d6_70),.data_out(wire_d6_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7672(.data_in(wire_d6_71),.data_out(wire_d6_72),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7673(.data_in(wire_d6_72),.data_out(wire_d6_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7674(.data_in(wire_d6_73),.data_out(wire_d6_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7675(.data_in(wire_d6_74),.data_out(wire_d6_75),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7676(.data_in(wire_d6_75),.data_out(wire_d6_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7677(.data_in(wire_d6_76),.data_out(wire_d6_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7678(.data_in(wire_d6_77),.data_out(wire_d6_78),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7679(.data_in(wire_d6_78),.data_out(d_out6),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance870(.data_in(d_in7),.data_out(wire_d7_0),.clk(clk),.rst(rst));            //channel 8
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance871(.data_in(wire_d7_0),.data_out(wire_d7_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance872(.data_in(wire_d7_1),.data_out(wire_d7_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance873(.data_in(wire_d7_2),.data_out(wire_d7_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance874(.data_in(wire_d7_3),.data_out(wire_d7_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance875(.data_in(wire_d7_4),.data_out(wire_d7_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance876(.data_in(wire_d7_5),.data_out(wire_d7_6),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance877(.data_in(wire_d7_6),.data_out(wire_d7_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance878(.data_in(wire_d7_7),.data_out(wire_d7_8),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance879(.data_in(wire_d7_8),.data_out(wire_d7_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8710(.data_in(wire_d7_9),.data_out(wire_d7_10),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8711(.data_in(wire_d7_10),.data_out(wire_d7_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8712(.data_in(wire_d7_11),.data_out(wire_d7_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8713(.data_in(wire_d7_12),.data_out(wire_d7_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8714(.data_in(wire_d7_13),.data_out(wire_d7_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8715(.data_in(wire_d7_14),.data_out(wire_d7_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8716(.data_in(wire_d7_15),.data_out(wire_d7_16),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8717(.data_in(wire_d7_16),.data_out(wire_d7_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8718(.data_in(wire_d7_17),.data_out(wire_d7_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8719(.data_in(wire_d7_18),.data_out(wire_d7_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8720(.data_in(wire_d7_19),.data_out(wire_d7_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8721(.data_in(wire_d7_20),.data_out(wire_d7_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8722(.data_in(wire_d7_21),.data_out(wire_d7_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8723(.data_in(wire_d7_22),.data_out(wire_d7_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8724(.data_in(wire_d7_23),.data_out(wire_d7_24),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8725(.data_in(wire_d7_24),.data_out(wire_d7_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8726(.data_in(wire_d7_25),.data_out(wire_d7_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8727(.data_in(wire_d7_26),.data_out(wire_d7_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8728(.data_in(wire_d7_27),.data_out(wire_d7_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8729(.data_in(wire_d7_28),.data_out(wire_d7_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8730(.data_in(wire_d7_29),.data_out(wire_d7_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8731(.data_in(wire_d7_30),.data_out(wire_d7_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8732(.data_in(wire_d7_31),.data_out(wire_d7_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8733(.data_in(wire_d7_32),.data_out(wire_d7_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8734(.data_in(wire_d7_33),.data_out(wire_d7_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8735(.data_in(wire_d7_34),.data_out(wire_d7_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8736(.data_in(wire_d7_35),.data_out(wire_d7_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8737(.data_in(wire_d7_36),.data_out(wire_d7_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8738(.data_in(wire_d7_37),.data_out(wire_d7_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8739(.data_in(wire_d7_38),.data_out(wire_d7_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8740(.data_in(wire_d7_39),.data_out(wire_d7_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8741(.data_in(wire_d7_40),.data_out(wire_d7_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8742(.data_in(wire_d7_41),.data_out(wire_d7_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8743(.data_in(wire_d7_42),.data_out(wire_d7_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8744(.data_in(wire_d7_43),.data_out(wire_d7_44),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8745(.data_in(wire_d7_44),.data_out(wire_d7_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8746(.data_in(wire_d7_45),.data_out(wire_d7_46),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8747(.data_in(wire_d7_46),.data_out(wire_d7_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8748(.data_in(wire_d7_47),.data_out(wire_d7_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8749(.data_in(wire_d7_48),.data_out(wire_d7_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8750(.data_in(wire_d7_49),.data_out(wire_d7_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8751(.data_in(wire_d7_50),.data_out(wire_d7_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8752(.data_in(wire_d7_51),.data_out(wire_d7_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8753(.data_in(wire_d7_52),.data_out(wire_d7_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8754(.data_in(wire_d7_53),.data_out(wire_d7_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8755(.data_in(wire_d7_54),.data_out(wire_d7_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8756(.data_in(wire_d7_55),.data_out(wire_d7_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8757(.data_in(wire_d7_56),.data_out(wire_d7_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8758(.data_in(wire_d7_57),.data_out(wire_d7_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8759(.data_in(wire_d7_58),.data_out(wire_d7_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8760(.data_in(wire_d7_59),.data_out(wire_d7_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8761(.data_in(wire_d7_60),.data_out(wire_d7_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8762(.data_in(wire_d7_61),.data_out(wire_d7_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8763(.data_in(wire_d7_62),.data_out(wire_d7_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8764(.data_in(wire_d7_63),.data_out(wire_d7_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8765(.data_in(wire_d7_64),.data_out(wire_d7_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8766(.data_in(wire_d7_65),.data_out(wire_d7_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8767(.data_in(wire_d7_66),.data_out(wire_d7_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8768(.data_in(wire_d7_67),.data_out(wire_d7_68),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8769(.data_in(wire_d7_68),.data_out(wire_d7_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8770(.data_in(wire_d7_69),.data_out(wire_d7_70),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8771(.data_in(wire_d7_70),.data_out(wire_d7_71),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8772(.data_in(wire_d7_71),.data_out(wire_d7_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8773(.data_in(wire_d7_72),.data_out(wire_d7_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8774(.data_in(wire_d7_73),.data_out(wire_d7_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8775(.data_in(wire_d7_74),.data_out(wire_d7_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8776(.data_in(wire_d7_75),.data_out(wire_d7_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8777(.data_in(wire_d7_76),.data_out(wire_d7_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8778(.data_in(wire_d7_77),.data_out(wire_d7_78),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8779(.data_in(wire_d7_78),.data_out(d_out7),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance980(.data_in(d_in8),.data_out(wire_d8_0),.clk(clk),.rst(rst));            //channel 9
	large_mux #(.WIDTH(WIDTH)) large_mux_instance981(.data_in(wire_d8_0),.data_out(wire_d8_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance982(.data_in(wire_d8_1),.data_out(wire_d8_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance983(.data_in(wire_d8_2),.data_out(wire_d8_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance984(.data_in(wire_d8_3),.data_out(wire_d8_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance985(.data_in(wire_d8_4),.data_out(wire_d8_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance986(.data_in(wire_d8_5),.data_out(wire_d8_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance987(.data_in(wire_d8_6),.data_out(wire_d8_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance988(.data_in(wire_d8_7),.data_out(wire_d8_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance989(.data_in(wire_d8_8),.data_out(wire_d8_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9810(.data_in(wire_d8_9),.data_out(wire_d8_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9811(.data_in(wire_d8_10),.data_out(wire_d8_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9812(.data_in(wire_d8_11),.data_out(wire_d8_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9813(.data_in(wire_d8_12),.data_out(wire_d8_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9814(.data_in(wire_d8_13),.data_out(wire_d8_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9815(.data_in(wire_d8_14),.data_out(wire_d8_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9816(.data_in(wire_d8_15),.data_out(wire_d8_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9817(.data_in(wire_d8_16),.data_out(wire_d8_17),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9818(.data_in(wire_d8_17),.data_out(wire_d8_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9819(.data_in(wire_d8_18),.data_out(wire_d8_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9820(.data_in(wire_d8_19),.data_out(wire_d8_20),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9821(.data_in(wire_d8_20),.data_out(wire_d8_21),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9822(.data_in(wire_d8_21),.data_out(wire_d8_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9823(.data_in(wire_d8_22),.data_out(wire_d8_23),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9824(.data_in(wire_d8_23),.data_out(wire_d8_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9825(.data_in(wire_d8_24),.data_out(wire_d8_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9826(.data_in(wire_d8_25),.data_out(wire_d8_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9827(.data_in(wire_d8_26),.data_out(wire_d8_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9828(.data_in(wire_d8_27),.data_out(wire_d8_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9829(.data_in(wire_d8_28),.data_out(wire_d8_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9830(.data_in(wire_d8_29),.data_out(wire_d8_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9831(.data_in(wire_d8_30),.data_out(wire_d8_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9832(.data_in(wire_d8_31),.data_out(wire_d8_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9833(.data_in(wire_d8_32),.data_out(wire_d8_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9834(.data_in(wire_d8_33),.data_out(wire_d8_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9835(.data_in(wire_d8_34),.data_out(wire_d8_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9836(.data_in(wire_d8_35),.data_out(wire_d8_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9837(.data_in(wire_d8_36),.data_out(wire_d8_37),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9838(.data_in(wire_d8_37),.data_out(wire_d8_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9839(.data_in(wire_d8_38),.data_out(wire_d8_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9840(.data_in(wire_d8_39),.data_out(wire_d8_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9841(.data_in(wire_d8_40),.data_out(wire_d8_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9842(.data_in(wire_d8_41),.data_out(wire_d8_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9843(.data_in(wire_d8_42),.data_out(wire_d8_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9844(.data_in(wire_d8_43),.data_out(wire_d8_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9845(.data_in(wire_d8_44),.data_out(wire_d8_45),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9846(.data_in(wire_d8_45),.data_out(wire_d8_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9847(.data_in(wire_d8_46),.data_out(wire_d8_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9848(.data_in(wire_d8_47),.data_out(wire_d8_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9849(.data_in(wire_d8_48),.data_out(wire_d8_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9850(.data_in(wire_d8_49),.data_out(wire_d8_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9851(.data_in(wire_d8_50),.data_out(wire_d8_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9852(.data_in(wire_d8_51),.data_out(wire_d8_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9853(.data_in(wire_d8_52),.data_out(wire_d8_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9854(.data_in(wire_d8_53),.data_out(wire_d8_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9855(.data_in(wire_d8_54),.data_out(wire_d8_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9856(.data_in(wire_d8_55),.data_out(wire_d8_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9857(.data_in(wire_d8_56),.data_out(wire_d8_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9858(.data_in(wire_d8_57),.data_out(wire_d8_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9859(.data_in(wire_d8_58),.data_out(wire_d8_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9860(.data_in(wire_d8_59),.data_out(wire_d8_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9861(.data_in(wire_d8_60),.data_out(wire_d8_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9862(.data_in(wire_d8_61),.data_out(wire_d8_62),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9863(.data_in(wire_d8_62),.data_out(wire_d8_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9864(.data_in(wire_d8_63),.data_out(wire_d8_64),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9865(.data_in(wire_d8_64),.data_out(wire_d8_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9866(.data_in(wire_d8_65),.data_out(wire_d8_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9867(.data_in(wire_d8_66),.data_out(wire_d8_67),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9868(.data_in(wire_d8_67),.data_out(wire_d8_68),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9869(.data_in(wire_d8_68),.data_out(wire_d8_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9870(.data_in(wire_d8_69),.data_out(wire_d8_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9871(.data_in(wire_d8_70),.data_out(wire_d8_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9872(.data_in(wire_d8_71),.data_out(wire_d8_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9873(.data_in(wire_d8_72),.data_out(wire_d8_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9874(.data_in(wire_d8_73),.data_out(wire_d8_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9875(.data_in(wire_d8_74),.data_out(wire_d8_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9876(.data_in(wire_d8_75),.data_out(wire_d8_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9877(.data_in(wire_d8_76),.data_out(wire_d8_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9878(.data_in(wire_d8_77),.data_out(wire_d8_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9879(.data_in(wire_d8_78),.data_out(d_out8),.clk(clk),.rst(rst));

	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance10090(.data_in(d_in9),.data_out(wire_d9_0),.clk(clk),.rst(rst));            //channel 10
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10091(.data_in(wire_d9_0),.data_out(wire_d9_1),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10092(.data_in(wire_d9_1),.data_out(wire_d9_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance10093(.data_in(wire_d9_2),.data_out(wire_d9_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance10094(.data_in(wire_d9_3),.data_out(wire_d9_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10095(.data_in(wire_d9_4),.data_out(wire_d9_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10096(.data_in(wire_d9_5),.data_out(wire_d9_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10097(.data_in(wire_d9_6),.data_out(wire_d9_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance10098(.data_in(wire_d9_7),.data_out(wire_d9_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10099(.data_in(wire_d9_8),.data_out(wire_d9_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100910(.data_in(wire_d9_9),.data_out(wire_d9_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100911(.data_in(wire_d9_10),.data_out(wire_d9_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100912(.data_in(wire_d9_11),.data_out(wire_d9_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100913(.data_in(wire_d9_12),.data_out(wire_d9_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100914(.data_in(wire_d9_13),.data_out(wire_d9_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100915(.data_in(wire_d9_14),.data_out(wire_d9_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100916(.data_in(wire_d9_15),.data_out(wire_d9_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100917(.data_in(wire_d9_16),.data_out(wire_d9_17),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100918(.data_in(wire_d9_17),.data_out(wire_d9_18),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100919(.data_in(wire_d9_18),.data_out(wire_d9_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100920(.data_in(wire_d9_19),.data_out(wire_d9_20),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100921(.data_in(wire_d9_20),.data_out(wire_d9_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100922(.data_in(wire_d9_21),.data_out(wire_d9_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100923(.data_in(wire_d9_22),.data_out(wire_d9_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100924(.data_in(wire_d9_23),.data_out(wire_d9_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100925(.data_in(wire_d9_24),.data_out(wire_d9_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100926(.data_in(wire_d9_25),.data_out(wire_d9_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100927(.data_in(wire_d9_26),.data_out(wire_d9_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance100928(.data_in(wire_d9_27),.data_out(wire_d9_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100929(.data_in(wire_d9_28),.data_out(wire_d9_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100930(.data_in(wire_d9_29),.data_out(wire_d9_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100931(.data_in(wire_d9_30),.data_out(wire_d9_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100932(.data_in(wire_d9_31),.data_out(wire_d9_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100933(.data_in(wire_d9_32),.data_out(wire_d9_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100934(.data_in(wire_d9_33),.data_out(wire_d9_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100935(.data_in(wire_d9_34),.data_out(wire_d9_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100936(.data_in(wire_d9_35),.data_out(wire_d9_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100937(.data_in(wire_d9_36),.data_out(wire_d9_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100938(.data_in(wire_d9_37),.data_out(wire_d9_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100939(.data_in(wire_d9_38),.data_out(wire_d9_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100940(.data_in(wire_d9_39),.data_out(wire_d9_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100941(.data_in(wire_d9_40),.data_out(wire_d9_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100942(.data_in(wire_d9_41),.data_out(wire_d9_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100943(.data_in(wire_d9_42),.data_out(wire_d9_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100944(.data_in(wire_d9_43),.data_out(wire_d9_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100945(.data_in(wire_d9_44),.data_out(wire_d9_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100946(.data_in(wire_d9_45),.data_out(wire_d9_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100947(.data_in(wire_d9_46),.data_out(wire_d9_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100948(.data_in(wire_d9_47),.data_out(wire_d9_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100949(.data_in(wire_d9_48),.data_out(wire_d9_49),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100950(.data_in(wire_d9_49),.data_out(wire_d9_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100951(.data_in(wire_d9_50),.data_out(wire_d9_51),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100952(.data_in(wire_d9_51),.data_out(wire_d9_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance100953(.data_in(wire_d9_52),.data_out(wire_d9_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100954(.data_in(wire_d9_53),.data_out(wire_d9_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100955(.data_in(wire_d9_54),.data_out(wire_d9_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100956(.data_in(wire_d9_55),.data_out(wire_d9_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100957(.data_in(wire_d9_56),.data_out(wire_d9_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance100958(.data_in(wire_d9_57),.data_out(wire_d9_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100959(.data_in(wire_d9_58),.data_out(wire_d9_59),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100960(.data_in(wire_d9_59),.data_out(wire_d9_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100961(.data_in(wire_d9_60),.data_out(wire_d9_61),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100962(.data_in(wire_d9_61),.data_out(wire_d9_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100963(.data_in(wire_d9_62),.data_out(wire_d9_63),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100964(.data_in(wire_d9_63),.data_out(wire_d9_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100965(.data_in(wire_d9_64),.data_out(wire_d9_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100966(.data_in(wire_d9_65),.data_out(wire_d9_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100967(.data_in(wire_d9_66),.data_out(wire_d9_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100968(.data_in(wire_d9_67),.data_out(wire_d9_68),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance100969(.data_in(wire_d9_68),.data_out(wire_d9_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100970(.data_in(wire_d9_69),.data_out(wire_d9_70),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance100971(.data_in(wire_d9_70),.data_out(wire_d9_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100972(.data_in(wire_d9_71),.data_out(wire_d9_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100973(.data_in(wire_d9_72),.data_out(wire_d9_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100974(.data_in(wire_d9_73),.data_out(wire_d9_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100975(.data_in(wire_d9_74),.data_out(wire_d9_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100976(.data_in(wire_d9_75),.data_out(wire_d9_76),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100977(.data_in(wire_d9_76),.data_out(wire_d9_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100978(.data_in(wire_d9_77),.data_out(wire_d9_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100979(.data_in(wire_d9_78),.data_out(d_out9),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance110100(.data_in(d_in10),.data_out(wire_d10_0),.clk(clk),.rst(rst));            //channel 11
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance110101(.data_in(wire_d10_0),.data_out(wire_d10_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance110102(.data_in(wire_d10_1),.data_out(wire_d10_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance110103(.data_in(wire_d10_2),.data_out(wire_d10_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance110104(.data_in(wire_d10_3),.data_out(wire_d10_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance110105(.data_in(wire_d10_4),.data_out(wire_d10_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance110106(.data_in(wire_d10_5),.data_out(wire_d10_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance110107(.data_in(wire_d10_6),.data_out(wire_d10_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance110108(.data_in(wire_d10_7),.data_out(wire_d10_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance110109(.data_in(wire_d10_8),.data_out(wire_d10_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101010(.data_in(wire_d10_9),.data_out(wire_d10_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101011(.data_in(wire_d10_10),.data_out(wire_d10_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101012(.data_in(wire_d10_11),.data_out(wire_d10_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101013(.data_in(wire_d10_12),.data_out(wire_d10_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1101014(.data_in(wire_d10_13),.data_out(wire_d10_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101015(.data_in(wire_d10_14),.data_out(wire_d10_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101016(.data_in(wire_d10_15),.data_out(wire_d10_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101017(.data_in(wire_d10_16),.data_out(wire_d10_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1101018(.data_in(wire_d10_17),.data_out(wire_d10_18),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101019(.data_in(wire_d10_18),.data_out(wire_d10_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101020(.data_in(wire_d10_19),.data_out(wire_d10_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101021(.data_in(wire_d10_20),.data_out(wire_d10_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1101022(.data_in(wire_d10_21),.data_out(wire_d10_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101023(.data_in(wire_d10_22),.data_out(wire_d10_23),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101024(.data_in(wire_d10_23),.data_out(wire_d10_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101025(.data_in(wire_d10_24),.data_out(wire_d10_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101026(.data_in(wire_d10_25),.data_out(wire_d10_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101027(.data_in(wire_d10_26),.data_out(wire_d10_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101028(.data_in(wire_d10_27),.data_out(wire_d10_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101029(.data_in(wire_d10_28),.data_out(wire_d10_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101030(.data_in(wire_d10_29),.data_out(wire_d10_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101031(.data_in(wire_d10_30),.data_out(wire_d10_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1101032(.data_in(wire_d10_31),.data_out(wire_d10_32),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101033(.data_in(wire_d10_32),.data_out(wire_d10_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101034(.data_in(wire_d10_33),.data_out(wire_d10_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101035(.data_in(wire_d10_34),.data_out(wire_d10_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101036(.data_in(wire_d10_35),.data_out(wire_d10_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1101037(.data_in(wire_d10_36),.data_out(wire_d10_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101038(.data_in(wire_d10_37),.data_out(wire_d10_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101039(.data_in(wire_d10_38),.data_out(wire_d10_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101040(.data_in(wire_d10_39),.data_out(wire_d10_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101041(.data_in(wire_d10_40),.data_out(wire_d10_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101042(.data_in(wire_d10_41),.data_out(wire_d10_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101043(.data_in(wire_d10_42),.data_out(wire_d10_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101044(.data_in(wire_d10_43),.data_out(wire_d10_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101045(.data_in(wire_d10_44),.data_out(wire_d10_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1101046(.data_in(wire_d10_45),.data_out(wire_d10_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101047(.data_in(wire_d10_46),.data_out(wire_d10_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101048(.data_in(wire_d10_47),.data_out(wire_d10_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1101049(.data_in(wire_d10_48),.data_out(wire_d10_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101050(.data_in(wire_d10_49),.data_out(wire_d10_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101051(.data_in(wire_d10_50),.data_out(wire_d10_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1101052(.data_in(wire_d10_51),.data_out(wire_d10_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101053(.data_in(wire_d10_52),.data_out(wire_d10_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101054(.data_in(wire_d10_53),.data_out(wire_d10_54),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101055(.data_in(wire_d10_54),.data_out(wire_d10_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101056(.data_in(wire_d10_55),.data_out(wire_d10_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101057(.data_in(wire_d10_56),.data_out(wire_d10_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1101058(.data_in(wire_d10_57),.data_out(wire_d10_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101059(.data_in(wire_d10_58),.data_out(wire_d10_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101060(.data_in(wire_d10_59),.data_out(wire_d10_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101061(.data_in(wire_d10_60),.data_out(wire_d10_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1101062(.data_in(wire_d10_61),.data_out(wire_d10_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101063(.data_in(wire_d10_62),.data_out(wire_d10_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101064(.data_in(wire_d10_63),.data_out(wire_d10_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101065(.data_in(wire_d10_64),.data_out(wire_d10_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101066(.data_in(wire_d10_65),.data_out(wire_d10_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1101067(.data_in(wire_d10_66),.data_out(wire_d10_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1101068(.data_in(wire_d10_67),.data_out(wire_d10_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1101069(.data_in(wire_d10_68),.data_out(wire_d10_69),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101070(.data_in(wire_d10_69),.data_out(wire_d10_70),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101071(.data_in(wire_d10_70),.data_out(wire_d10_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101072(.data_in(wire_d10_71),.data_out(wire_d10_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101073(.data_in(wire_d10_72),.data_out(wire_d10_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101074(.data_in(wire_d10_73),.data_out(wire_d10_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101075(.data_in(wire_d10_74),.data_out(wire_d10_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101076(.data_in(wire_d10_75),.data_out(wire_d10_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101077(.data_in(wire_d10_76),.data_out(wire_d10_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101078(.data_in(wire_d10_77),.data_out(wire_d10_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1101079(.data_in(wire_d10_78),.data_out(d_out10),.clk(clk),.rst(rst));

	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance120110(.data_in(d_in11),.data_out(wire_d11_0),.clk(clk),.rst(rst));            //channel 12
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance120111(.data_in(wire_d11_0),.data_out(wire_d11_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance120112(.data_in(wire_d11_1),.data_out(wire_d11_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance120113(.data_in(wire_d11_2),.data_out(wire_d11_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance120114(.data_in(wire_d11_3),.data_out(wire_d11_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance120115(.data_in(wire_d11_4),.data_out(wire_d11_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance120116(.data_in(wire_d11_5),.data_out(wire_d11_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance120117(.data_in(wire_d11_6),.data_out(wire_d11_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance120118(.data_in(wire_d11_7),.data_out(wire_d11_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance120119(.data_in(wire_d11_8),.data_out(wire_d11_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201110(.data_in(wire_d11_9),.data_out(wire_d11_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201111(.data_in(wire_d11_10),.data_out(wire_d11_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201112(.data_in(wire_d11_11),.data_out(wire_d11_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201113(.data_in(wire_d11_12),.data_out(wire_d11_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201114(.data_in(wire_d11_13),.data_out(wire_d11_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201115(.data_in(wire_d11_14),.data_out(wire_d11_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201116(.data_in(wire_d11_15),.data_out(wire_d11_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201117(.data_in(wire_d11_16),.data_out(wire_d11_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201118(.data_in(wire_d11_17),.data_out(wire_d11_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201119(.data_in(wire_d11_18),.data_out(wire_d11_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1201120(.data_in(wire_d11_19),.data_out(wire_d11_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201121(.data_in(wire_d11_20),.data_out(wire_d11_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201122(.data_in(wire_d11_21),.data_out(wire_d11_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201123(.data_in(wire_d11_22),.data_out(wire_d11_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201124(.data_in(wire_d11_23),.data_out(wire_d11_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201125(.data_in(wire_d11_24),.data_out(wire_d11_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201126(.data_in(wire_d11_25),.data_out(wire_d11_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201127(.data_in(wire_d11_26),.data_out(wire_d11_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201128(.data_in(wire_d11_27),.data_out(wire_d11_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201129(.data_in(wire_d11_28),.data_out(wire_d11_29),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201130(.data_in(wire_d11_29),.data_out(wire_d11_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1201131(.data_in(wire_d11_30),.data_out(wire_d11_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201132(.data_in(wire_d11_31),.data_out(wire_d11_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201133(.data_in(wire_d11_32),.data_out(wire_d11_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201134(.data_in(wire_d11_33),.data_out(wire_d11_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1201135(.data_in(wire_d11_34),.data_out(wire_d11_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201136(.data_in(wire_d11_35),.data_out(wire_d11_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201137(.data_in(wire_d11_36),.data_out(wire_d11_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201138(.data_in(wire_d11_37),.data_out(wire_d11_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201139(.data_in(wire_d11_38),.data_out(wire_d11_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201140(.data_in(wire_d11_39),.data_out(wire_d11_40),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201141(.data_in(wire_d11_40),.data_out(wire_d11_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201142(.data_in(wire_d11_41),.data_out(wire_d11_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201143(.data_in(wire_d11_42),.data_out(wire_d11_43),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201144(.data_in(wire_d11_43),.data_out(wire_d11_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201145(.data_in(wire_d11_44),.data_out(wire_d11_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201146(.data_in(wire_d11_45),.data_out(wire_d11_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201147(.data_in(wire_d11_46),.data_out(wire_d11_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201148(.data_in(wire_d11_47),.data_out(wire_d11_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201149(.data_in(wire_d11_48),.data_out(wire_d11_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201150(.data_in(wire_d11_49),.data_out(wire_d11_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201151(.data_in(wire_d11_50),.data_out(wire_d11_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201152(.data_in(wire_d11_51),.data_out(wire_d11_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201153(.data_in(wire_d11_52),.data_out(wire_d11_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201154(.data_in(wire_d11_53),.data_out(wire_d11_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1201155(.data_in(wire_d11_54),.data_out(wire_d11_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201156(.data_in(wire_d11_55),.data_out(wire_d11_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201157(.data_in(wire_d11_56),.data_out(wire_d11_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201158(.data_in(wire_d11_57),.data_out(wire_d11_58),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1201159(.data_in(wire_d11_58),.data_out(wire_d11_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201160(.data_in(wire_d11_59),.data_out(wire_d11_60),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201161(.data_in(wire_d11_60),.data_out(wire_d11_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201162(.data_in(wire_d11_61),.data_out(wire_d11_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201163(.data_in(wire_d11_62),.data_out(wire_d11_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201164(.data_in(wire_d11_63),.data_out(wire_d11_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201165(.data_in(wire_d11_64),.data_out(wire_d11_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1201166(.data_in(wire_d11_65),.data_out(wire_d11_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201167(.data_in(wire_d11_66),.data_out(wire_d11_67),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201168(.data_in(wire_d11_67),.data_out(wire_d11_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201169(.data_in(wire_d11_68),.data_out(wire_d11_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1201170(.data_in(wire_d11_69),.data_out(wire_d11_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201171(.data_in(wire_d11_70),.data_out(wire_d11_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201172(.data_in(wire_d11_71),.data_out(wire_d11_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201173(.data_in(wire_d11_72),.data_out(wire_d11_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201174(.data_in(wire_d11_73),.data_out(wire_d11_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201175(.data_in(wire_d11_74),.data_out(wire_d11_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201176(.data_in(wire_d11_75),.data_out(wire_d11_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201177(.data_in(wire_d11_76),.data_out(wire_d11_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201178(.data_in(wire_d11_77),.data_out(wire_d11_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201179(.data_in(wire_d11_78),.data_out(d_out11),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance130120(.data_in(d_in12),.data_out(wire_d12_0),.clk(clk),.rst(rst));            //channel 13
	decoder_top #(.WIDTH(WIDTH)) decoder_instance130121(.data_in(wire_d12_0),.data_out(wire_d12_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance130122(.data_in(wire_d12_1),.data_out(wire_d12_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance130123(.data_in(wire_d12_2),.data_out(wire_d12_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance130124(.data_in(wire_d12_3),.data_out(wire_d12_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance130125(.data_in(wire_d12_4),.data_out(wire_d12_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance130126(.data_in(wire_d12_5),.data_out(wire_d12_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance130127(.data_in(wire_d12_6),.data_out(wire_d12_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance130128(.data_in(wire_d12_7),.data_out(wire_d12_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance130129(.data_in(wire_d12_8),.data_out(wire_d12_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301210(.data_in(wire_d12_9),.data_out(wire_d12_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301211(.data_in(wire_d12_10),.data_out(wire_d12_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301212(.data_in(wire_d12_11),.data_out(wire_d12_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301213(.data_in(wire_d12_12),.data_out(wire_d12_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301214(.data_in(wire_d12_13),.data_out(wire_d12_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301215(.data_in(wire_d12_14),.data_out(wire_d12_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301216(.data_in(wire_d12_15),.data_out(wire_d12_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301217(.data_in(wire_d12_16),.data_out(wire_d12_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301218(.data_in(wire_d12_17),.data_out(wire_d12_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301219(.data_in(wire_d12_18),.data_out(wire_d12_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1301220(.data_in(wire_d12_19),.data_out(wire_d12_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301221(.data_in(wire_d12_20),.data_out(wire_d12_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1301222(.data_in(wire_d12_21),.data_out(wire_d12_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301223(.data_in(wire_d12_22),.data_out(wire_d12_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1301224(.data_in(wire_d12_23),.data_out(wire_d12_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301225(.data_in(wire_d12_24),.data_out(wire_d12_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301226(.data_in(wire_d12_25),.data_out(wire_d12_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301227(.data_in(wire_d12_26),.data_out(wire_d12_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1301228(.data_in(wire_d12_27),.data_out(wire_d12_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301229(.data_in(wire_d12_28),.data_out(wire_d12_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301230(.data_in(wire_d12_29),.data_out(wire_d12_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1301231(.data_in(wire_d12_30),.data_out(wire_d12_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1301232(.data_in(wire_d12_31),.data_out(wire_d12_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301233(.data_in(wire_d12_32),.data_out(wire_d12_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301234(.data_in(wire_d12_33),.data_out(wire_d12_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301235(.data_in(wire_d12_34),.data_out(wire_d12_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301236(.data_in(wire_d12_35),.data_out(wire_d12_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301237(.data_in(wire_d12_36),.data_out(wire_d12_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1301238(.data_in(wire_d12_37),.data_out(wire_d12_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301239(.data_in(wire_d12_38),.data_out(wire_d12_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301240(.data_in(wire_d12_39),.data_out(wire_d12_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301241(.data_in(wire_d12_40),.data_out(wire_d12_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301242(.data_in(wire_d12_41),.data_out(wire_d12_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1301243(.data_in(wire_d12_42),.data_out(wire_d12_43),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1301244(.data_in(wire_d12_43),.data_out(wire_d12_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301245(.data_in(wire_d12_44),.data_out(wire_d12_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301246(.data_in(wire_d12_45),.data_out(wire_d12_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301247(.data_in(wire_d12_46),.data_out(wire_d12_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301248(.data_in(wire_d12_47),.data_out(wire_d12_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301249(.data_in(wire_d12_48),.data_out(wire_d12_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301250(.data_in(wire_d12_49),.data_out(wire_d12_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301251(.data_in(wire_d12_50),.data_out(wire_d12_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1301252(.data_in(wire_d12_51),.data_out(wire_d12_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301253(.data_in(wire_d12_52),.data_out(wire_d12_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301254(.data_in(wire_d12_53),.data_out(wire_d12_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1301255(.data_in(wire_d12_54),.data_out(wire_d12_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301256(.data_in(wire_d12_55),.data_out(wire_d12_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1301257(.data_in(wire_d12_56),.data_out(wire_d12_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301258(.data_in(wire_d12_57),.data_out(wire_d12_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301259(.data_in(wire_d12_58),.data_out(wire_d12_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301260(.data_in(wire_d12_59),.data_out(wire_d12_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301261(.data_in(wire_d12_60),.data_out(wire_d12_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301262(.data_in(wire_d12_61),.data_out(wire_d12_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301263(.data_in(wire_d12_62),.data_out(wire_d12_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301264(.data_in(wire_d12_63),.data_out(wire_d12_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301265(.data_in(wire_d12_64),.data_out(wire_d12_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301266(.data_in(wire_d12_65),.data_out(wire_d12_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1301267(.data_in(wire_d12_66),.data_out(wire_d12_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301268(.data_in(wire_d12_67),.data_out(wire_d12_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301269(.data_in(wire_d12_68),.data_out(wire_d12_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301270(.data_in(wire_d12_69),.data_out(wire_d12_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301271(.data_in(wire_d12_70),.data_out(wire_d12_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1301272(.data_in(wire_d12_71),.data_out(wire_d12_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301273(.data_in(wire_d12_72),.data_out(wire_d12_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301274(.data_in(wire_d12_73),.data_out(wire_d12_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301275(.data_in(wire_d12_74),.data_out(wire_d12_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1301276(.data_in(wire_d12_75),.data_out(wire_d12_76),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301277(.data_in(wire_d12_76),.data_out(wire_d12_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301278(.data_in(wire_d12_77),.data_out(wire_d12_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301279(.data_in(wire_d12_78),.data_out(d_out12),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance140130(.data_in(d_in13),.data_out(wire_d13_0),.clk(clk),.rst(rst));            //channel 14
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance140131(.data_in(wire_d13_0),.data_out(wire_d13_1),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance140132(.data_in(wire_d13_1),.data_out(wire_d13_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance140133(.data_in(wire_d13_2),.data_out(wire_d13_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance140134(.data_in(wire_d13_3),.data_out(wire_d13_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance140135(.data_in(wire_d13_4),.data_out(wire_d13_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance140136(.data_in(wire_d13_5),.data_out(wire_d13_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance140137(.data_in(wire_d13_6),.data_out(wire_d13_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance140138(.data_in(wire_d13_7),.data_out(wire_d13_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance140139(.data_in(wire_d13_8),.data_out(wire_d13_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401310(.data_in(wire_d13_9),.data_out(wire_d13_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1401311(.data_in(wire_d13_10),.data_out(wire_d13_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401312(.data_in(wire_d13_11),.data_out(wire_d13_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401313(.data_in(wire_d13_12),.data_out(wire_d13_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401314(.data_in(wire_d13_13),.data_out(wire_d13_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401315(.data_in(wire_d13_14),.data_out(wire_d13_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401316(.data_in(wire_d13_15),.data_out(wire_d13_16),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1401317(.data_in(wire_d13_16),.data_out(wire_d13_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1401318(.data_in(wire_d13_17),.data_out(wire_d13_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401319(.data_in(wire_d13_18),.data_out(wire_d13_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1401320(.data_in(wire_d13_19),.data_out(wire_d13_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401321(.data_in(wire_d13_20),.data_out(wire_d13_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401322(.data_in(wire_d13_21),.data_out(wire_d13_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401323(.data_in(wire_d13_22),.data_out(wire_d13_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1401324(.data_in(wire_d13_23),.data_out(wire_d13_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401325(.data_in(wire_d13_24),.data_out(wire_d13_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1401326(.data_in(wire_d13_25),.data_out(wire_d13_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401327(.data_in(wire_d13_26),.data_out(wire_d13_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1401328(.data_in(wire_d13_27),.data_out(wire_d13_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401329(.data_in(wire_d13_28),.data_out(wire_d13_29),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401330(.data_in(wire_d13_29),.data_out(wire_d13_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1401331(.data_in(wire_d13_30),.data_out(wire_d13_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401332(.data_in(wire_d13_31),.data_out(wire_d13_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401333(.data_in(wire_d13_32),.data_out(wire_d13_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401334(.data_in(wire_d13_33),.data_out(wire_d13_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401335(.data_in(wire_d13_34),.data_out(wire_d13_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401336(.data_in(wire_d13_35),.data_out(wire_d13_36),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401337(.data_in(wire_d13_36),.data_out(wire_d13_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401338(.data_in(wire_d13_37),.data_out(wire_d13_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401339(.data_in(wire_d13_38),.data_out(wire_d13_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401340(.data_in(wire_d13_39),.data_out(wire_d13_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401341(.data_in(wire_d13_40),.data_out(wire_d13_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1401342(.data_in(wire_d13_41),.data_out(wire_d13_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401343(.data_in(wire_d13_42),.data_out(wire_d13_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401344(.data_in(wire_d13_43),.data_out(wire_d13_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1401345(.data_in(wire_d13_44),.data_out(wire_d13_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401346(.data_in(wire_d13_45),.data_out(wire_d13_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401347(.data_in(wire_d13_46),.data_out(wire_d13_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1401348(.data_in(wire_d13_47),.data_out(wire_d13_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401349(.data_in(wire_d13_48),.data_out(wire_d13_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401350(.data_in(wire_d13_49),.data_out(wire_d13_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401351(.data_in(wire_d13_50),.data_out(wire_d13_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1401352(.data_in(wire_d13_51),.data_out(wire_d13_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401353(.data_in(wire_d13_52),.data_out(wire_d13_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401354(.data_in(wire_d13_53),.data_out(wire_d13_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401355(.data_in(wire_d13_54),.data_out(wire_d13_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1401356(.data_in(wire_d13_55),.data_out(wire_d13_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401357(.data_in(wire_d13_56),.data_out(wire_d13_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401358(.data_in(wire_d13_57),.data_out(wire_d13_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401359(.data_in(wire_d13_58),.data_out(wire_d13_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401360(.data_in(wire_d13_59),.data_out(wire_d13_60),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401361(.data_in(wire_d13_60),.data_out(wire_d13_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1401362(.data_in(wire_d13_61),.data_out(wire_d13_62),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401363(.data_in(wire_d13_62),.data_out(wire_d13_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401364(.data_in(wire_d13_63),.data_out(wire_d13_64),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401365(.data_in(wire_d13_64),.data_out(wire_d13_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401366(.data_in(wire_d13_65),.data_out(wire_d13_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401367(.data_in(wire_d13_66),.data_out(wire_d13_67),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401368(.data_in(wire_d13_67),.data_out(wire_d13_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401369(.data_in(wire_d13_68),.data_out(wire_d13_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401370(.data_in(wire_d13_69),.data_out(wire_d13_70),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401371(.data_in(wire_d13_70),.data_out(wire_d13_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401372(.data_in(wire_d13_71),.data_out(wire_d13_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1401373(.data_in(wire_d13_72),.data_out(wire_d13_73),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401374(.data_in(wire_d13_73),.data_out(wire_d13_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401375(.data_in(wire_d13_74),.data_out(wire_d13_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1401376(.data_in(wire_d13_75),.data_out(wire_d13_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401377(.data_in(wire_d13_76),.data_out(wire_d13_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401378(.data_in(wire_d13_77),.data_out(wire_d13_78),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401379(.data_in(wire_d13_78),.data_out(d_out13),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance150140(.data_in(d_in14),.data_out(wire_d14_0),.clk(clk),.rst(rst));            //channel 15
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance150141(.data_in(wire_d14_0),.data_out(wire_d14_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance150142(.data_in(wire_d14_1),.data_out(wire_d14_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance150143(.data_in(wire_d14_2),.data_out(wire_d14_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance150144(.data_in(wire_d14_3),.data_out(wire_d14_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance150145(.data_in(wire_d14_4),.data_out(wire_d14_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance150146(.data_in(wire_d14_5),.data_out(wire_d14_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance150147(.data_in(wire_d14_6),.data_out(wire_d14_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance150148(.data_in(wire_d14_7),.data_out(wire_d14_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance150149(.data_in(wire_d14_8),.data_out(wire_d14_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501410(.data_in(wire_d14_9),.data_out(wire_d14_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501411(.data_in(wire_d14_10),.data_out(wire_d14_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501412(.data_in(wire_d14_11),.data_out(wire_d14_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501413(.data_in(wire_d14_12),.data_out(wire_d14_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501414(.data_in(wire_d14_13),.data_out(wire_d14_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1501415(.data_in(wire_d14_14),.data_out(wire_d14_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501416(.data_in(wire_d14_15),.data_out(wire_d14_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501417(.data_in(wire_d14_16),.data_out(wire_d14_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501418(.data_in(wire_d14_17),.data_out(wire_d14_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501419(.data_in(wire_d14_18),.data_out(wire_d14_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501420(.data_in(wire_d14_19),.data_out(wire_d14_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501421(.data_in(wire_d14_20),.data_out(wire_d14_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1501422(.data_in(wire_d14_21),.data_out(wire_d14_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501423(.data_in(wire_d14_22),.data_out(wire_d14_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501424(.data_in(wire_d14_23),.data_out(wire_d14_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501425(.data_in(wire_d14_24),.data_out(wire_d14_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501426(.data_in(wire_d14_25),.data_out(wire_d14_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501427(.data_in(wire_d14_26),.data_out(wire_d14_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1501428(.data_in(wire_d14_27),.data_out(wire_d14_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501429(.data_in(wire_d14_28),.data_out(wire_d14_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501430(.data_in(wire_d14_29),.data_out(wire_d14_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501431(.data_in(wire_d14_30),.data_out(wire_d14_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1501432(.data_in(wire_d14_31),.data_out(wire_d14_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501433(.data_in(wire_d14_32),.data_out(wire_d14_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1501434(.data_in(wire_d14_33),.data_out(wire_d14_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501435(.data_in(wire_d14_34),.data_out(wire_d14_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1501436(.data_in(wire_d14_35),.data_out(wire_d14_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501437(.data_in(wire_d14_36),.data_out(wire_d14_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501438(.data_in(wire_d14_37),.data_out(wire_d14_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1501439(.data_in(wire_d14_38),.data_out(wire_d14_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1501440(.data_in(wire_d14_39),.data_out(wire_d14_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501441(.data_in(wire_d14_40),.data_out(wire_d14_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501442(.data_in(wire_d14_41),.data_out(wire_d14_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501443(.data_in(wire_d14_42),.data_out(wire_d14_43),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501444(.data_in(wire_d14_43),.data_out(wire_d14_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1501445(.data_in(wire_d14_44),.data_out(wire_d14_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501446(.data_in(wire_d14_45),.data_out(wire_d14_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1501447(.data_in(wire_d14_46),.data_out(wire_d14_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501448(.data_in(wire_d14_47),.data_out(wire_d14_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501449(.data_in(wire_d14_48),.data_out(wire_d14_49),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501450(.data_in(wire_d14_49),.data_out(wire_d14_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1501451(.data_in(wire_d14_50),.data_out(wire_d14_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501452(.data_in(wire_d14_51),.data_out(wire_d14_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1501453(.data_in(wire_d14_52),.data_out(wire_d14_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1501454(.data_in(wire_d14_53),.data_out(wire_d14_54),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501455(.data_in(wire_d14_54),.data_out(wire_d14_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501456(.data_in(wire_d14_55),.data_out(wire_d14_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501457(.data_in(wire_d14_56),.data_out(wire_d14_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501458(.data_in(wire_d14_57),.data_out(wire_d14_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1501459(.data_in(wire_d14_58),.data_out(wire_d14_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501460(.data_in(wire_d14_59),.data_out(wire_d14_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501461(.data_in(wire_d14_60),.data_out(wire_d14_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501462(.data_in(wire_d14_61),.data_out(wire_d14_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1501463(.data_in(wire_d14_62),.data_out(wire_d14_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501464(.data_in(wire_d14_63),.data_out(wire_d14_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501465(.data_in(wire_d14_64),.data_out(wire_d14_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501466(.data_in(wire_d14_65),.data_out(wire_d14_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501467(.data_in(wire_d14_66),.data_out(wire_d14_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1501468(.data_in(wire_d14_67),.data_out(wire_d14_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501469(.data_in(wire_d14_68),.data_out(wire_d14_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501470(.data_in(wire_d14_69),.data_out(wire_d14_70),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501471(.data_in(wire_d14_70),.data_out(wire_d14_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1501472(.data_in(wire_d14_71),.data_out(wire_d14_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501473(.data_in(wire_d14_72),.data_out(wire_d14_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501474(.data_in(wire_d14_73),.data_out(wire_d14_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501475(.data_in(wire_d14_74),.data_out(wire_d14_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501476(.data_in(wire_d14_75),.data_out(wire_d14_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501477(.data_in(wire_d14_76),.data_out(wire_d14_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501478(.data_in(wire_d14_77),.data_out(wire_d14_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501479(.data_in(wire_d14_78),.data_out(d_out14),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance160150(.data_in(d_in15),.data_out(wire_d15_0),.clk(clk),.rst(rst));            //channel 16
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance160151(.data_in(wire_d15_0),.data_out(wire_d15_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance160152(.data_in(wire_d15_1),.data_out(wire_d15_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance160153(.data_in(wire_d15_2),.data_out(wire_d15_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance160154(.data_in(wire_d15_3),.data_out(wire_d15_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance160155(.data_in(wire_d15_4),.data_out(wire_d15_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance160156(.data_in(wire_d15_5),.data_out(wire_d15_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance160157(.data_in(wire_d15_6),.data_out(wire_d15_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance160158(.data_in(wire_d15_7),.data_out(wire_d15_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance160159(.data_in(wire_d15_8),.data_out(wire_d15_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601510(.data_in(wire_d15_9),.data_out(wire_d15_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601511(.data_in(wire_d15_10),.data_out(wire_d15_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601512(.data_in(wire_d15_11),.data_out(wire_d15_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601513(.data_in(wire_d15_12),.data_out(wire_d15_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601514(.data_in(wire_d15_13),.data_out(wire_d15_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601515(.data_in(wire_d15_14),.data_out(wire_d15_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601516(.data_in(wire_d15_15),.data_out(wire_d15_16),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601517(.data_in(wire_d15_16),.data_out(wire_d15_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601518(.data_in(wire_d15_17),.data_out(wire_d15_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601519(.data_in(wire_d15_18),.data_out(wire_d15_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601520(.data_in(wire_d15_19),.data_out(wire_d15_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1601521(.data_in(wire_d15_20),.data_out(wire_d15_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601522(.data_in(wire_d15_21),.data_out(wire_d15_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1601523(.data_in(wire_d15_22),.data_out(wire_d15_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601524(.data_in(wire_d15_23),.data_out(wire_d15_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601525(.data_in(wire_d15_24),.data_out(wire_d15_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601526(.data_in(wire_d15_25),.data_out(wire_d15_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601527(.data_in(wire_d15_26),.data_out(wire_d15_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601528(.data_in(wire_d15_27),.data_out(wire_d15_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601529(.data_in(wire_d15_28),.data_out(wire_d15_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601530(.data_in(wire_d15_29),.data_out(wire_d15_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601531(.data_in(wire_d15_30),.data_out(wire_d15_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601532(.data_in(wire_d15_31),.data_out(wire_d15_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601533(.data_in(wire_d15_32),.data_out(wire_d15_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1601534(.data_in(wire_d15_33),.data_out(wire_d15_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601535(.data_in(wire_d15_34),.data_out(wire_d15_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601536(.data_in(wire_d15_35),.data_out(wire_d15_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1601537(.data_in(wire_d15_36),.data_out(wire_d15_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601538(.data_in(wire_d15_37),.data_out(wire_d15_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1601539(.data_in(wire_d15_38),.data_out(wire_d15_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601540(.data_in(wire_d15_39),.data_out(wire_d15_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601541(.data_in(wire_d15_40),.data_out(wire_d15_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601542(.data_in(wire_d15_41),.data_out(wire_d15_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601543(.data_in(wire_d15_42),.data_out(wire_d15_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601544(.data_in(wire_d15_43),.data_out(wire_d15_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601545(.data_in(wire_d15_44),.data_out(wire_d15_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601546(.data_in(wire_d15_45),.data_out(wire_d15_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601547(.data_in(wire_d15_46),.data_out(wire_d15_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1601548(.data_in(wire_d15_47),.data_out(wire_d15_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601549(.data_in(wire_d15_48),.data_out(wire_d15_49),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601550(.data_in(wire_d15_49),.data_out(wire_d15_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601551(.data_in(wire_d15_50),.data_out(wire_d15_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1601552(.data_in(wire_d15_51),.data_out(wire_d15_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1601553(.data_in(wire_d15_52),.data_out(wire_d15_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601554(.data_in(wire_d15_53),.data_out(wire_d15_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1601555(.data_in(wire_d15_54),.data_out(wire_d15_55),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601556(.data_in(wire_d15_55),.data_out(wire_d15_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601557(.data_in(wire_d15_56),.data_out(wire_d15_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601558(.data_in(wire_d15_57),.data_out(wire_d15_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601559(.data_in(wire_d15_58),.data_out(wire_d15_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601560(.data_in(wire_d15_59),.data_out(wire_d15_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601561(.data_in(wire_d15_60),.data_out(wire_d15_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601562(.data_in(wire_d15_61),.data_out(wire_d15_62),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601563(.data_in(wire_d15_62),.data_out(wire_d15_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1601564(.data_in(wire_d15_63),.data_out(wire_d15_64),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601565(.data_in(wire_d15_64),.data_out(wire_d15_65),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601566(.data_in(wire_d15_65),.data_out(wire_d15_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1601567(.data_in(wire_d15_66),.data_out(wire_d15_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601568(.data_in(wire_d15_67),.data_out(wire_d15_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601569(.data_in(wire_d15_68),.data_out(wire_d15_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601570(.data_in(wire_d15_69),.data_out(wire_d15_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601571(.data_in(wire_d15_70),.data_out(wire_d15_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601572(.data_in(wire_d15_71),.data_out(wire_d15_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601573(.data_in(wire_d15_72),.data_out(wire_d15_73),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601574(.data_in(wire_d15_73),.data_out(wire_d15_74),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1601575(.data_in(wire_d15_74),.data_out(wire_d15_75),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601576(.data_in(wire_d15_75),.data_out(wire_d15_76),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601577(.data_in(wire_d15_76),.data_out(wire_d15_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601578(.data_in(wire_d15_77),.data_out(wire_d15_78),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601579(.data_in(wire_d15_78),.data_out(d_out15),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance170160(.data_in(d_in16),.data_out(wire_d16_0),.clk(clk),.rst(rst));            //channel 17
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance170161(.data_in(wire_d16_0),.data_out(wire_d16_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance170162(.data_in(wire_d16_1),.data_out(wire_d16_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance170163(.data_in(wire_d16_2),.data_out(wire_d16_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance170164(.data_in(wire_d16_3),.data_out(wire_d16_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance170165(.data_in(wire_d16_4),.data_out(wire_d16_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance170166(.data_in(wire_d16_5),.data_out(wire_d16_6),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance170167(.data_in(wire_d16_6),.data_out(wire_d16_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance170168(.data_in(wire_d16_7),.data_out(wire_d16_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance170169(.data_in(wire_d16_8),.data_out(wire_d16_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701610(.data_in(wire_d16_9),.data_out(wire_d16_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1701611(.data_in(wire_d16_10),.data_out(wire_d16_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701612(.data_in(wire_d16_11),.data_out(wire_d16_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701613(.data_in(wire_d16_12),.data_out(wire_d16_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701614(.data_in(wire_d16_13),.data_out(wire_d16_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1701615(.data_in(wire_d16_14),.data_out(wire_d16_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701616(.data_in(wire_d16_15),.data_out(wire_d16_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701617(.data_in(wire_d16_16),.data_out(wire_d16_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1701618(.data_in(wire_d16_17),.data_out(wire_d16_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1701619(.data_in(wire_d16_18),.data_out(wire_d16_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1701620(.data_in(wire_d16_19),.data_out(wire_d16_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701621(.data_in(wire_d16_20),.data_out(wire_d16_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701622(.data_in(wire_d16_21),.data_out(wire_d16_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701623(.data_in(wire_d16_22),.data_out(wire_d16_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701624(.data_in(wire_d16_23),.data_out(wire_d16_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1701625(.data_in(wire_d16_24),.data_out(wire_d16_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701626(.data_in(wire_d16_25),.data_out(wire_d16_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701627(.data_in(wire_d16_26),.data_out(wire_d16_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701628(.data_in(wire_d16_27),.data_out(wire_d16_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701629(.data_in(wire_d16_28),.data_out(wire_d16_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1701630(.data_in(wire_d16_29),.data_out(wire_d16_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701631(.data_in(wire_d16_30),.data_out(wire_d16_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701632(.data_in(wire_d16_31),.data_out(wire_d16_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701633(.data_in(wire_d16_32),.data_out(wire_d16_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701634(.data_in(wire_d16_33),.data_out(wire_d16_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701635(.data_in(wire_d16_34),.data_out(wire_d16_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701636(.data_in(wire_d16_35),.data_out(wire_d16_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701637(.data_in(wire_d16_36),.data_out(wire_d16_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1701638(.data_in(wire_d16_37),.data_out(wire_d16_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701639(.data_in(wire_d16_38),.data_out(wire_d16_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701640(.data_in(wire_d16_39),.data_out(wire_d16_40),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701641(.data_in(wire_d16_40),.data_out(wire_d16_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701642(.data_in(wire_d16_41),.data_out(wire_d16_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701643(.data_in(wire_d16_42),.data_out(wire_d16_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701644(.data_in(wire_d16_43),.data_out(wire_d16_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701645(.data_in(wire_d16_44),.data_out(wire_d16_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1701646(.data_in(wire_d16_45),.data_out(wire_d16_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701647(.data_in(wire_d16_46),.data_out(wire_d16_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701648(.data_in(wire_d16_47),.data_out(wire_d16_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701649(.data_in(wire_d16_48),.data_out(wire_d16_49),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1701650(.data_in(wire_d16_49),.data_out(wire_d16_50),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1701651(.data_in(wire_d16_50),.data_out(wire_d16_51),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701652(.data_in(wire_d16_51),.data_out(wire_d16_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701653(.data_in(wire_d16_52),.data_out(wire_d16_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701654(.data_in(wire_d16_53),.data_out(wire_d16_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701655(.data_in(wire_d16_54),.data_out(wire_d16_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701656(.data_in(wire_d16_55),.data_out(wire_d16_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701657(.data_in(wire_d16_56),.data_out(wire_d16_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701658(.data_in(wire_d16_57),.data_out(wire_d16_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701659(.data_in(wire_d16_58),.data_out(wire_d16_59),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1701660(.data_in(wire_d16_59),.data_out(wire_d16_60),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701661(.data_in(wire_d16_60),.data_out(wire_d16_61),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1701662(.data_in(wire_d16_61),.data_out(wire_d16_62),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701663(.data_in(wire_d16_62),.data_out(wire_d16_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1701664(.data_in(wire_d16_63),.data_out(wire_d16_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701665(.data_in(wire_d16_64),.data_out(wire_d16_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701666(.data_in(wire_d16_65),.data_out(wire_d16_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701667(.data_in(wire_d16_66),.data_out(wire_d16_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701668(.data_in(wire_d16_67),.data_out(wire_d16_68),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701669(.data_in(wire_d16_68),.data_out(wire_d16_69),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701670(.data_in(wire_d16_69),.data_out(wire_d16_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701671(.data_in(wire_d16_70),.data_out(wire_d16_71),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701672(.data_in(wire_d16_71),.data_out(wire_d16_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701673(.data_in(wire_d16_72),.data_out(wire_d16_73),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701674(.data_in(wire_d16_73),.data_out(wire_d16_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701675(.data_in(wire_d16_74),.data_out(wire_d16_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701676(.data_in(wire_d16_75),.data_out(wire_d16_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701677(.data_in(wire_d16_76),.data_out(wire_d16_77),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701678(.data_in(wire_d16_77),.data_out(wire_d16_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701679(.data_in(wire_d16_78),.data_out(d_out16),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance180170(.data_in(d_in17),.data_out(wire_d17_0),.clk(clk),.rst(rst));            //channel 18
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance180171(.data_in(wire_d17_0),.data_out(wire_d17_1),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance180172(.data_in(wire_d17_1),.data_out(wire_d17_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance180173(.data_in(wire_d17_2),.data_out(wire_d17_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance180174(.data_in(wire_d17_3),.data_out(wire_d17_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance180175(.data_in(wire_d17_4),.data_out(wire_d17_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance180176(.data_in(wire_d17_5),.data_out(wire_d17_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance180177(.data_in(wire_d17_6),.data_out(wire_d17_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance180178(.data_in(wire_d17_7),.data_out(wire_d17_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance180179(.data_in(wire_d17_8),.data_out(wire_d17_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801710(.data_in(wire_d17_9),.data_out(wire_d17_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801711(.data_in(wire_d17_10),.data_out(wire_d17_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801712(.data_in(wire_d17_11),.data_out(wire_d17_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801713(.data_in(wire_d17_12),.data_out(wire_d17_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801714(.data_in(wire_d17_13),.data_out(wire_d17_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801715(.data_in(wire_d17_14),.data_out(wire_d17_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1801716(.data_in(wire_d17_15),.data_out(wire_d17_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1801717(.data_in(wire_d17_16),.data_out(wire_d17_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801718(.data_in(wire_d17_17),.data_out(wire_d17_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801719(.data_in(wire_d17_18),.data_out(wire_d17_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1801720(.data_in(wire_d17_19),.data_out(wire_d17_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801721(.data_in(wire_d17_20),.data_out(wire_d17_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801722(.data_in(wire_d17_21),.data_out(wire_d17_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1801723(.data_in(wire_d17_22),.data_out(wire_d17_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801724(.data_in(wire_d17_23),.data_out(wire_d17_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801725(.data_in(wire_d17_24),.data_out(wire_d17_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801726(.data_in(wire_d17_25),.data_out(wire_d17_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801727(.data_in(wire_d17_26),.data_out(wire_d17_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801728(.data_in(wire_d17_27),.data_out(wire_d17_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801729(.data_in(wire_d17_28),.data_out(wire_d17_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801730(.data_in(wire_d17_29),.data_out(wire_d17_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801731(.data_in(wire_d17_30),.data_out(wire_d17_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801732(.data_in(wire_d17_31),.data_out(wire_d17_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801733(.data_in(wire_d17_32),.data_out(wire_d17_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801734(.data_in(wire_d17_33),.data_out(wire_d17_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801735(.data_in(wire_d17_34),.data_out(wire_d17_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801736(.data_in(wire_d17_35),.data_out(wire_d17_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801737(.data_in(wire_d17_36),.data_out(wire_d17_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801738(.data_in(wire_d17_37),.data_out(wire_d17_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801739(.data_in(wire_d17_38),.data_out(wire_d17_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801740(.data_in(wire_d17_39),.data_out(wire_d17_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801741(.data_in(wire_d17_40),.data_out(wire_d17_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801742(.data_in(wire_d17_41),.data_out(wire_d17_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801743(.data_in(wire_d17_42),.data_out(wire_d17_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801744(.data_in(wire_d17_43),.data_out(wire_d17_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801745(.data_in(wire_d17_44),.data_out(wire_d17_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1801746(.data_in(wire_d17_45),.data_out(wire_d17_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801747(.data_in(wire_d17_46),.data_out(wire_d17_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801748(.data_in(wire_d17_47),.data_out(wire_d17_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801749(.data_in(wire_d17_48),.data_out(wire_d17_49),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801750(.data_in(wire_d17_49),.data_out(wire_d17_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801751(.data_in(wire_d17_50),.data_out(wire_d17_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801752(.data_in(wire_d17_51),.data_out(wire_d17_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801753(.data_in(wire_d17_52),.data_out(wire_d17_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801754(.data_in(wire_d17_53),.data_out(wire_d17_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801755(.data_in(wire_d17_54),.data_out(wire_d17_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801756(.data_in(wire_d17_55),.data_out(wire_d17_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801757(.data_in(wire_d17_56),.data_out(wire_d17_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801758(.data_in(wire_d17_57),.data_out(wire_d17_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801759(.data_in(wire_d17_58),.data_out(wire_d17_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801760(.data_in(wire_d17_59),.data_out(wire_d17_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801761(.data_in(wire_d17_60),.data_out(wire_d17_61),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801762(.data_in(wire_d17_61),.data_out(wire_d17_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801763(.data_in(wire_d17_62),.data_out(wire_d17_63),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801764(.data_in(wire_d17_63),.data_out(wire_d17_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801765(.data_in(wire_d17_64),.data_out(wire_d17_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801766(.data_in(wire_d17_65),.data_out(wire_d17_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1801767(.data_in(wire_d17_66),.data_out(wire_d17_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801768(.data_in(wire_d17_67),.data_out(wire_d17_68),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801769(.data_in(wire_d17_68),.data_out(wire_d17_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801770(.data_in(wire_d17_69),.data_out(wire_d17_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801771(.data_in(wire_d17_70),.data_out(wire_d17_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1801772(.data_in(wire_d17_71),.data_out(wire_d17_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801773(.data_in(wire_d17_72),.data_out(wire_d17_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801774(.data_in(wire_d17_73),.data_out(wire_d17_74),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801775(.data_in(wire_d17_74),.data_out(wire_d17_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1801776(.data_in(wire_d17_75),.data_out(wire_d17_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801777(.data_in(wire_d17_76),.data_out(wire_d17_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801778(.data_in(wire_d17_77),.data_out(wire_d17_78),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801779(.data_in(wire_d17_78),.data_out(d_out17),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance190180(.data_in(d_in18),.data_out(wire_d18_0),.clk(clk),.rst(rst));            //channel 19
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance190181(.data_in(wire_d18_0),.data_out(wire_d18_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance190182(.data_in(wire_d18_1),.data_out(wire_d18_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance190183(.data_in(wire_d18_2),.data_out(wire_d18_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance190184(.data_in(wire_d18_3),.data_out(wire_d18_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance190185(.data_in(wire_d18_4),.data_out(wire_d18_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance190186(.data_in(wire_d18_5),.data_out(wire_d18_6),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance190187(.data_in(wire_d18_6),.data_out(wire_d18_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance190188(.data_in(wire_d18_7),.data_out(wire_d18_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance190189(.data_in(wire_d18_8),.data_out(wire_d18_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901810(.data_in(wire_d18_9),.data_out(wire_d18_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1901811(.data_in(wire_d18_10),.data_out(wire_d18_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901812(.data_in(wire_d18_11),.data_out(wire_d18_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901813(.data_in(wire_d18_12),.data_out(wire_d18_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901814(.data_in(wire_d18_13),.data_out(wire_d18_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901815(.data_in(wire_d18_14),.data_out(wire_d18_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901816(.data_in(wire_d18_15),.data_out(wire_d18_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901817(.data_in(wire_d18_16),.data_out(wire_d18_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901818(.data_in(wire_d18_17),.data_out(wire_d18_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901819(.data_in(wire_d18_18),.data_out(wire_d18_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901820(.data_in(wire_d18_19),.data_out(wire_d18_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901821(.data_in(wire_d18_20),.data_out(wire_d18_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901822(.data_in(wire_d18_21),.data_out(wire_d18_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901823(.data_in(wire_d18_22),.data_out(wire_d18_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901824(.data_in(wire_d18_23),.data_out(wire_d18_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901825(.data_in(wire_d18_24),.data_out(wire_d18_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901826(.data_in(wire_d18_25),.data_out(wire_d18_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901827(.data_in(wire_d18_26),.data_out(wire_d18_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901828(.data_in(wire_d18_27),.data_out(wire_d18_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901829(.data_in(wire_d18_28),.data_out(wire_d18_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901830(.data_in(wire_d18_29),.data_out(wire_d18_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901831(.data_in(wire_d18_30),.data_out(wire_d18_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901832(.data_in(wire_d18_31),.data_out(wire_d18_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901833(.data_in(wire_d18_32),.data_out(wire_d18_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1901834(.data_in(wire_d18_33),.data_out(wire_d18_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901835(.data_in(wire_d18_34),.data_out(wire_d18_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901836(.data_in(wire_d18_35),.data_out(wire_d18_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901837(.data_in(wire_d18_36),.data_out(wire_d18_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901838(.data_in(wire_d18_37),.data_out(wire_d18_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901839(.data_in(wire_d18_38),.data_out(wire_d18_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901840(.data_in(wire_d18_39),.data_out(wire_d18_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1901841(.data_in(wire_d18_40),.data_out(wire_d18_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901842(.data_in(wire_d18_41),.data_out(wire_d18_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901843(.data_in(wire_d18_42),.data_out(wire_d18_43),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901844(.data_in(wire_d18_43),.data_out(wire_d18_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901845(.data_in(wire_d18_44),.data_out(wire_d18_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901846(.data_in(wire_d18_45),.data_out(wire_d18_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901847(.data_in(wire_d18_46),.data_out(wire_d18_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901848(.data_in(wire_d18_47),.data_out(wire_d18_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1901849(.data_in(wire_d18_48),.data_out(wire_d18_49),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901850(.data_in(wire_d18_49),.data_out(wire_d18_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901851(.data_in(wire_d18_50),.data_out(wire_d18_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901852(.data_in(wire_d18_51),.data_out(wire_d18_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901853(.data_in(wire_d18_52),.data_out(wire_d18_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901854(.data_in(wire_d18_53),.data_out(wire_d18_54),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1901855(.data_in(wire_d18_54),.data_out(wire_d18_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901856(.data_in(wire_d18_55),.data_out(wire_d18_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901857(.data_in(wire_d18_56),.data_out(wire_d18_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901858(.data_in(wire_d18_57),.data_out(wire_d18_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901859(.data_in(wire_d18_58),.data_out(wire_d18_59),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901860(.data_in(wire_d18_59),.data_out(wire_d18_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1901861(.data_in(wire_d18_60),.data_out(wire_d18_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901862(.data_in(wire_d18_61),.data_out(wire_d18_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901863(.data_in(wire_d18_62),.data_out(wire_d18_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901864(.data_in(wire_d18_63),.data_out(wire_d18_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901865(.data_in(wire_d18_64),.data_out(wire_d18_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901866(.data_in(wire_d18_65),.data_out(wire_d18_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901867(.data_in(wire_d18_66),.data_out(wire_d18_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901868(.data_in(wire_d18_67),.data_out(wire_d18_68),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901869(.data_in(wire_d18_68),.data_out(wire_d18_69),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901870(.data_in(wire_d18_69),.data_out(wire_d18_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901871(.data_in(wire_d18_70),.data_out(wire_d18_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901872(.data_in(wire_d18_71),.data_out(wire_d18_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901873(.data_in(wire_d18_72),.data_out(wire_d18_73),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901874(.data_in(wire_d18_73),.data_out(wire_d18_74),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901875(.data_in(wire_d18_74),.data_out(wire_d18_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901876(.data_in(wire_d18_75),.data_out(wire_d18_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901877(.data_in(wire_d18_76),.data_out(wire_d18_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901878(.data_in(wire_d18_77),.data_out(wire_d18_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901879(.data_in(wire_d18_78),.data_out(d_out18),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance200190(.data_in(d_in19),.data_out(wire_d19_0),.clk(clk),.rst(rst));            //channel 20
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance200191(.data_in(wire_d19_0),.data_out(wire_d19_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance200192(.data_in(wire_d19_1),.data_out(wire_d19_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance200193(.data_in(wire_d19_2),.data_out(wire_d19_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance200194(.data_in(wire_d19_3),.data_out(wire_d19_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance200195(.data_in(wire_d19_4),.data_out(wire_d19_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance200196(.data_in(wire_d19_5),.data_out(wire_d19_6),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance200197(.data_in(wire_d19_6),.data_out(wire_d19_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance200198(.data_in(wire_d19_7),.data_out(wire_d19_8),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance200199(.data_in(wire_d19_8),.data_out(wire_d19_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2001910(.data_in(wire_d19_9),.data_out(wire_d19_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2001911(.data_in(wire_d19_10),.data_out(wire_d19_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001912(.data_in(wire_d19_11),.data_out(wire_d19_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001913(.data_in(wire_d19_12),.data_out(wire_d19_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001914(.data_in(wire_d19_13),.data_out(wire_d19_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001915(.data_in(wire_d19_14),.data_out(wire_d19_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2001916(.data_in(wire_d19_15),.data_out(wire_d19_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2001917(.data_in(wire_d19_16),.data_out(wire_d19_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2001918(.data_in(wire_d19_17),.data_out(wire_d19_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001919(.data_in(wire_d19_18),.data_out(wire_d19_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001920(.data_in(wire_d19_19),.data_out(wire_d19_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001921(.data_in(wire_d19_20),.data_out(wire_d19_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001922(.data_in(wire_d19_21),.data_out(wire_d19_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001923(.data_in(wire_d19_22),.data_out(wire_d19_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2001924(.data_in(wire_d19_23),.data_out(wire_d19_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2001925(.data_in(wire_d19_24),.data_out(wire_d19_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001926(.data_in(wire_d19_25),.data_out(wire_d19_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2001927(.data_in(wire_d19_26),.data_out(wire_d19_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001928(.data_in(wire_d19_27),.data_out(wire_d19_28),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001929(.data_in(wire_d19_28),.data_out(wire_d19_29),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001930(.data_in(wire_d19_29),.data_out(wire_d19_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001931(.data_in(wire_d19_30),.data_out(wire_d19_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001932(.data_in(wire_d19_31),.data_out(wire_d19_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2001933(.data_in(wire_d19_32),.data_out(wire_d19_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001934(.data_in(wire_d19_33),.data_out(wire_d19_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001935(.data_in(wire_d19_34),.data_out(wire_d19_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2001936(.data_in(wire_d19_35),.data_out(wire_d19_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001937(.data_in(wire_d19_36),.data_out(wire_d19_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2001938(.data_in(wire_d19_37),.data_out(wire_d19_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001939(.data_in(wire_d19_38),.data_out(wire_d19_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2001940(.data_in(wire_d19_39),.data_out(wire_d19_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001941(.data_in(wire_d19_40),.data_out(wire_d19_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2001942(.data_in(wire_d19_41),.data_out(wire_d19_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2001943(.data_in(wire_d19_42),.data_out(wire_d19_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001944(.data_in(wire_d19_43),.data_out(wire_d19_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001945(.data_in(wire_d19_44),.data_out(wire_d19_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001946(.data_in(wire_d19_45),.data_out(wire_d19_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001947(.data_in(wire_d19_46),.data_out(wire_d19_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001948(.data_in(wire_d19_47),.data_out(wire_d19_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001949(.data_in(wire_d19_48),.data_out(wire_d19_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001950(.data_in(wire_d19_49),.data_out(wire_d19_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001951(.data_in(wire_d19_50),.data_out(wire_d19_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001952(.data_in(wire_d19_51),.data_out(wire_d19_52),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2001953(.data_in(wire_d19_52),.data_out(wire_d19_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001954(.data_in(wire_d19_53),.data_out(wire_d19_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001955(.data_in(wire_d19_54),.data_out(wire_d19_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001956(.data_in(wire_d19_55),.data_out(wire_d19_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001957(.data_in(wire_d19_56),.data_out(wire_d19_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001958(.data_in(wire_d19_57),.data_out(wire_d19_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2001959(.data_in(wire_d19_58),.data_out(wire_d19_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001960(.data_in(wire_d19_59),.data_out(wire_d19_60),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001961(.data_in(wire_d19_60),.data_out(wire_d19_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2001962(.data_in(wire_d19_61),.data_out(wire_d19_62),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001963(.data_in(wire_d19_62),.data_out(wire_d19_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001964(.data_in(wire_d19_63),.data_out(wire_d19_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2001965(.data_in(wire_d19_64),.data_out(wire_d19_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001966(.data_in(wire_d19_65),.data_out(wire_d19_66),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001967(.data_in(wire_d19_66),.data_out(wire_d19_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001968(.data_in(wire_d19_67),.data_out(wire_d19_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2001969(.data_in(wire_d19_68),.data_out(wire_d19_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001970(.data_in(wire_d19_69),.data_out(wire_d19_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2001971(.data_in(wire_d19_70),.data_out(wire_d19_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001972(.data_in(wire_d19_71),.data_out(wire_d19_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001973(.data_in(wire_d19_72),.data_out(wire_d19_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001974(.data_in(wire_d19_73),.data_out(wire_d19_74),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001975(.data_in(wire_d19_74),.data_out(wire_d19_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001976(.data_in(wire_d19_75),.data_out(wire_d19_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2001977(.data_in(wire_d19_76),.data_out(wire_d19_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001978(.data_in(wire_d19_77),.data_out(wire_d19_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2001979(.data_in(wire_d19_78),.data_out(d_out19),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance210200(.data_in(d_in20),.data_out(wire_d20_0),.clk(clk),.rst(rst));            //channel 21
	decoder_top #(.WIDTH(WIDTH)) decoder_instance210201(.data_in(wire_d20_0),.data_out(wire_d20_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance210202(.data_in(wire_d20_1),.data_out(wire_d20_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance210203(.data_in(wire_d20_2),.data_out(wire_d20_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance210204(.data_in(wire_d20_3),.data_out(wire_d20_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance210205(.data_in(wire_d20_4),.data_out(wire_d20_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance210206(.data_in(wire_d20_5),.data_out(wire_d20_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance210207(.data_in(wire_d20_6),.data_out(wire_d20_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance210208(.data_in(wire_d20_7),.data_out(wire_d20_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance210209(.data_in(wire_d20_8),.data_out(wire_d20_9),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2102010(.data_in(wire_d20_9),.data_out(wire_d20_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102011(.data_in(wire_d20_10),.data_out(wire_d20_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102012(.data_in(wire_d20_11),.data_out(wire_d20_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102013(.data_in(wire_d20_12),.data_out(wire_d20_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102014(.data_in(wire_d20_13),.data_out(wire_d20_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102015(.data_in(wire_d20_14),.data_out(wire_d20_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102016(.data_in(wire_d20_15),.data_out(wire_d20_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102017(.data_in(wire_d20_16),.data_out(wire_d20_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102018(.data_in(wire_d20_17),.data_out(wire_d20_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102019(.data_in(wire_d20_18),.data_out(wire_d20_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2102020(.data_in(wire_d20_19),.data_out(wire_d20_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102021(.data_in(wire_d20_20),.data_out(wire_d20_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2102022(.data_in(wire_d20_21),.data_out(wire_d20_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102023(.data_in(wire_d20_22),.data_out(wire_d20_23),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102024(.data_in(wire_d20_23),.data_out(wire_d20_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2102025(.data_in(wire_d20_24),.data_out(wire_d20_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102026(.data_in(wire_d20_25),.data_out(wire_d20_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102027(.data_in(wire_d20_26),.data_out(wire_d20_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102028(.data_in(wire_d20_27),.data_out(wire_d20_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102029(.data_in(wire_d20_28),.data_out(wire_d20_29),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2102030(.data_in(wire_d20_29),.data_out(wire_d20_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102031(.data_in(wire_d20_30),.data_out(wire_d20_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102032(.data_in(wire_d20_31),.data_out(wire_d20_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102033(.data_in(wire_d20_32),.data_out(wire_d20_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102034(.data_in(wire_d20_33),.data_out(wire_d20_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2102035(.data_in(wire_d20_34),.data_out(wire_d20_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102036(.data_in(wire_d20_35),.data_out(wire_d20_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2102037(.data_in(wire_d20_36),.data_out(wire_d20_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102038(.data_in(wire_d20_37),.data_out(wire_d20_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102039(.data_in(wire_d20_38),.data_out(wire_d20_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102040(.data_in(wire_d20_39),.data_out(wire_d20_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102041(.data_in(wire_d20_40),.data_out(wire_d20_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102042(.data_in(wire_d20_41),.data_out(wire_d20_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102043(.data_in(wire_d20_42),.data_out(wire_d20_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102044(.data_in(wire_d20_43),.data_out(wire_d20_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102045(.data_in(wire_d20_44),.data_out(wire_d20_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2102046(.data_in(wire_d20_45),.data_out(wire_d20_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2102047(.data_in(wire_d20_46),.data_out(wire_d20_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102048(.data_in(wire_d20_47),.data_out(wire_d20_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102049(.data_in(wire_d20_48),.data_out(wire_d20_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102050(.data_in(wire_d20_49),.data_out(wire_d20_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102051(.data_in(wire_d20_50),.data_out(wire_d20_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2102052(.data_in(wire_d20_51),.data_out(wire_d20_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102053(.data_in(wire_d20_52),.data_out(wire_d20_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102054(.data_in(wire_d20_53),.data_out(wire_d20_54),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2102055(.data_in(wire_d20_54),.data_out(wire_d20_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102056(.data_in(wire_d20_55),.data_out(wire_d20_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102057(.data_in(wire_d20_56),.data_out(wire_d20_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102058(.data_in(wire_d20_57),.data_out(wire_d20_58),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102059(.data_in(wire_d20_58),.data_out(wire_d20_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102060(.data_in(wire_d20_59),.data_out(wire_d20_60),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102061(.data_in(wire_d20_60),.data_out(wire_d20_61),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102062(.data_in(wire_d20_61),.data_out(wire_d20_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2102063(.data_in(wire_d20_62),.data_out(wire_d20_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102064(.data_in(wire_d20_63),.data_out(wire_d20_64),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102065(.data_in(wire_d20_64),.data_out(wire_d20_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102066(.data_in(wire_d20_65),.data_out(wire_d20_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2102067(.data_in(wire_d20_66),.data_out(wire_d20_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102068(.data_in(wire_d20_67),.data_out(wire_d20_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102069(.data_in(wire_d20_68),.data_out(wire_d20_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102070(.data_in(wire_d20_69),.data_out(wire_d20_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2102071(.data_in(wire_d20_70),.data_out(wire_d20_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102072(.data_in(wire_d20_71),.data_out(wire_d20_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102073(.data_in(wire_d20_72),.data_out(wire_d20_73),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102074(.data_in(wire_d20_73),.data_out(wire_d20_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102075(.data_in(wire_d20_74),.data_out(wire_d20_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102076(.data_in(wire_d20_75),.data_out(wire_d20_76),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102077(.data_in(wire_d20_76),.data_out(wire_d20_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102078(.data_in(wire_d20_77),.data_out(wire_d20_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102079(.data_in(wire_d20_78),.data_out(d_out20),.clk(clk),.rst(rst));

	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance220210(.data_in(d_in21),.data_out(wire_d21_0),.clk(clk),.rst(rst));            //channel 22
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance220211(.data_in(wire_d21_0),.data_out(wire_d21_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance220212(.data_in(wire_d21_1),.data_out(wire_d21_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance220213(.data_in(wire_d21_2),.data_out(wire_d21_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance220214(.data_in(wire_d21_3),.data_out(wire_d21_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance220215(.data_in(wire_d21_4),.data_out(wire_d21_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance220216(.data_in(wire_d21_5),.data_out(wire_d21_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance220217(.data_in(wire_d21_6),.data_out(wire_d21_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance220218(.data_in(wire_d21_7),.data_out(wire_d21_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance220219(.data_in(wire_d21_8),.data_out(wire_d21_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202110(.data_in(wire_d21_9),.data_out(wire_d21_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202111(.data_in(wire_d21_10),.data_out(wire_d21_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202112(.data_in(wire_d21_11),.data_out(wire_d21_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2202113(.data_in(wire_d21_12),.data_out(wire_d21_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202114(.data_in(wire_d21_13),.data_out(wire_d21_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2202115(.data_in(wire_d21_14),.data_out(wire_d21_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2202116(.data_in(wire_d21_15),.data_out(wire_d21_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2202117(.data_in(wire_d21_16),.data_out(wire_d21_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202118(.data_in(wire_d21_17),.data_out(wire_d21_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202119(.data_in(wire_d21_18),.data_out(wire_d21_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202120(.data_in(wire_d21_19),.data_out(wire_d21_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2202121(.data_in(wire_d21_20),.data_out(wire_d21_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202122(.data_in(wire_d21_21),.data_out(wire_d21_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202123(.data_in(wire_d21_22),.data_out(wire_d21_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202124(.data_in(wire_d21_23),.data_out(wire_d21_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2202125(.data_in(wire_d21_24),.data_out(wire_d21_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202126(.data_in(wire_d21_25),.data_out(wire_d21_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2202127(.data_in(wire_d21_26),.data_out(wire_d21_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2202128(.data_in(wire_d21_27),.data_out(wire_d21_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202129(.data_in(wire_d21_28),.data_out(wire_d21_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202130(.data_in(wire_d21_29),.data_out(wire_d21_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2202131(.data_in(wire_d21_30),.data_out(wire_d21_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2202132(.data_in(wire_d21_31),.data_out(wire_d21_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2202133(.data_in(wire_d21_32),.data_out(wire_d21_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202134(.data_in(wire_d21_33),.data_out(wire_d21_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202135(.data_in(wire_d21_34),.data_out(wire_d21_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2202136(.data_in(wire_d21_35),.data_out(wire_d21_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2202137(.data_in(wire_d21_36),.data_out(wire_d21_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202138(.data_in(wire_d21_37),.data_out(wire_d21_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2202139(.data_in(wire_d21_38),.data_out(wire_d21_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202140(.data_in(wire_d21_39),.data_out(wire_d21_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202141(.data_in(wire_d21_40),.data_out(wire_d21_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202142(.data_in(wire_d21_41),.data_out(wire_d21_42),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2202143(.data_in(wire_d21_42),.data_out(wire_d21_43),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202144(.data_in(wire_d21_43),.data_out(wire_d21_44),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202145(.data_in(wire_d21_44),.data_out(wire_d21_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2202146(.data_in(wire_d21_45),.data_out(wire_d21_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2202147(.data_in(wire_d21_46),.data_out(wire_d21_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202148(.data_in(wire_d21_47),.data_out(wire_d21_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202149(.data_in(wire_d21_48),.data_out(wire_d21_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2202150(.data_in(wire_d21_49),.data_out(wire_d21_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202151(.data_in(wire_d21_50),.data_out(wire_d21_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202152(.data_in(wire_d21_51),.data_out(wire_d21_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202153(.data_in(wire_d21_52),.data_out(wire_d21_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202154(.data_in(wire_d21_53),.data_out(wire_d21_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2202155(.data_in(wire_d21_54),.data_out(wire_d21_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202156(.data_in(wire_d21_55),.data_out(wire_d21_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202157(.data_in(wire_d21_56),.data_out(wire_d21_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202158(.data_in(wire_d21_57),.data_out(wire_d21_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202159(.data_in(wire_d21_58),.data_out(wire_d21_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2202160(.data_in(wire_d21_59),.data_out(wire_d21_60),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202161(.data_in(wire_d21_60),.data_out(wire_d21_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202162(.data_in(wire_d21_61),.data_out(wire_d21_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202163(.data_in(wire_d21_62),.data_out(wire_d21_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202164(.data_in(wire_d21_63),.data_out(wire_d21_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202165(.data_in(wire_d21_64),.data_out(wire_d21_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202166(.data_in(wire_d21_65),.data_out(wire_d21_66),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202167(.data_in(wire_d21_66),.data_out(wire_d21_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202168(.data_in(wire_d21_67),.data_out(wire_d21_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202169(.data_in(wire_d21_68),.data_out(wire_d21_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202170(.data_in(wire_d21_69),.data_out(wire_d21_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202171(.data_in(wire_d21_70),.data_out(wire_d21_71),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202172(.data_in(wire_d21_71),.data_out(wire_d21_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202173(.data_in(wire_d21_72),.data_out(wire_d21_73),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202174(.data_in(wire_d21_73),.data_out(wire_d21_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202175(.data_in(wire_d21_74),.data_out(wire_d21_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202176(.data_in(wire_d21_75),.data_out(wire_d21_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2202177(.data_in(wire_d21_76),.data_out(wire_d21_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202178(.data_in(wire_d21_77),.data_out(wire_d21_78),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202179(.data_in(wire_d21_78),.data_out(d_out21),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance230220(.data_in(d_in22),.data_out(wire_d22_0),.clk(clk),.rst(rst));            //channel 23
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance230221(.data_in(wire_d22_0),.data_out(wire_d22_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance230222(.data_in(wire_d22_1),.data_out(wire_d22_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance230223(.data_in(wire_d22_2),.data_out(wire_d22_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance230224(.data_in(wire_d22_3),.data_out(wire_d22_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance230225(.data_in(wire_d22_4),.data_out(wire_d22_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance230226(.data_in(wire_d22_5),.data_out(wire_d22_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance230227(.data_in(wire_d22_6),.data_out(wire_d22_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance230228(.data_in(wire_d22_7),.data_out(wire_d22_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance230229(.data_in(wire_d22_8),.data_out(wire_d22_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2302210(.data_in(wire_d22_9),.data_out(wire_d22_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302211(.data_in(wire_d22_10),.data_out(wire_d22_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302212(.data_in(wire_d22_11),.data_out(wire_d22_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2302213(.data_in(wire_d22_12),.data_out(wire_d22_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302214(.data_in(wire_d22_13),.data_out(wire_d22_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302215(.data_in(wire_d22_14),.data_out(wire_d22_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302216(.data_in(wire_d22_15),.data_out(wire_d22_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302217(.data_in(wire_d22_16),.data_out(wire_d22_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302218(.data_in(wire_d22_17),.data_out(wire_d22_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302219(.data_in(wire_d22_18),.data_out(wire_d22_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302220(.data_in(wire_d22_19),.data_out(wire_d22_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302221(.data_in(wire_d22_20),.data_out(wire_d22_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302222(.data_in(wire_d22_21),.data_out(wire_d22_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2302223(.data_in(wire_d22_22),.data_out(wire_d22_23),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302224(.data_in(wire_d22_23),.data_out(wire_d22_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302225(.data_in(wire_d22_24),.data_out(wire_d22_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302226(.data_in(wire_d22_25),.data_out(wire_d22_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2302227(.data_in(wire_d22_26),.data_out(wire_d22_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302228(.data_in(wire_d22_27),.data_out(wire_d22_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2302229(.data_in(wire_d22_28),.data_out(wire_d22_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302230(.data_in(wire_d22_29),.data_out(wire_d22_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302231(.data_in(wire_d22_30),.data_out(wire_d22_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302232(.data_in(wire_d22_31),.data_out(wire_d22_32),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302233(.data_in(wire_d22_32),.data_out(wire_d22_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302234(.data_in(wire_d22_33),.data_out(wire_d22_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302235(.data_in(wire_d22_34),.data_out(wire_d22_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302236(.data_in(wire_d22_35),.data_out(wire_d22_36),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302237(.data_in(wire_d22_36),.data_out(wire_d22_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302238(.data_in(wire_d22_37),.data_out(wire_d22_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302239(.data_in(wire_d22_38),.data_out(wire_d22_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302240(.data_in(wire_d22_39),.data_out(wire_d22_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302241(.data_in(wire_d22_40),.data_out(wire_d22_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302242(.data_in(wire_d22_41),.data_out(wire_d22_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302243(.data_in(wire_d22_42),.data_out(wire_d22_43),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302244(.data_in(wire_d22_43),.data_out(wire_d22_44),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302245(.data_in(wire_d22_44),.data_out(wire_d22_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302246(.data_in(wire_d22_45),.data_out(wire_d22_46),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302247(.data_in(wire_d22_46),.data_out(wire_d22_47),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302248(.data_in(wire_d22_47),.data_out(wire_d22_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302249(.data_in(wire_d22_48),.data_out(wire_d22_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302250(.data_in(wire_d22_49),.data_out(wire_d22_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302251(.data_in(wire_d22_50),.data_out(wire_d22_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302252(.data_in(wire_d22_51),.data_out(wire_d22_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302253(.data_in(wire_d22_52),.data_out(wire_d22_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302254(.data_in(wire_d22_53),.data_out(wire_d22_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302255(.data_in(wire_d22_54),.data_out(wire_d22_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302256(.data_in(wire_d22_55),.data_out(wire_d22_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302257(.data_in(wire_d22_56),.data_out(wire_d22_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302258(.data_in(wire_d22_57),.data_out(wire_d22_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302259(.data_in(wire_d22_58),.data_out(wire_d22_59),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302260(.data_in(wire_d22_59),.data_out(wire_d22_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302261(.data_in(wire_d22_60),.data_out(wire_d22_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302262(.data_in(wire_d22_61),.data_out(wire_d22_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302263(.data_in(wire_d22_62),.data_out(wire_d22_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302264(.data_in(wire_d22_63),.data_out(wire_d22_64),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302265(.data_in(wire_d22_64),.data_out(wire_d22_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2302266(.data_in(wire_d22_65),.data_out(wire_d22_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302267(.data_in(wire_d22_66),.data_out(wire_d22_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302268(.data_in(wire_d22_67),.data_out(wire_d22_68),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302269(.data_in(wire_d22_68),.data_out(wire_d22_69),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302270(.data_in(wire_d22_69),.data_out(wire_d22_70),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302271(.data_in(wire_d22_70),.data_out(wire_d22_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2302272(.data_in(wire_d22_71),.data_out(wire_d22_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2302273(.data_in(wire_d22_72),.data_out(wire_d22_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302274(.data_in(wire_d22_73),.data_out(wire_d22_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302275(.data_in(wire_d22_74),.data_out(wire_d22_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302276(.data_in(wire_d22_75),.data_out(wire_d22_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2302277(.data_in(wire_d22_76),.data_out(wire_d22_77),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302278(.data_in(wire_d22_77),.data_out(wire_d22_78),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302279(.data_in(wire_d22_78),.data_out(d_out22),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance240230(.data_in(d_in23),.data_out(wire_d23_0),.clk(clk),.rst(rst));            //channel 24
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance240231(.data_in(wire_d23_0),.data_out(wire_d23_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance240232(.data_in(wire_d23_1),.data_out(wire_d23_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance240233(.data_in(wire_d23_2),.data_out(wire_d23_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance240234(.data_in(wire_d23_3),.data_out(wire_d23_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance240235(.data_in(wire_d23_4),.data_out(wire_d23_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance240236(.data_in(wire_d23_5),.data_out(wire_d23_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance240237(.data_in(wire_d23_6),.data_out(wire_d23_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance240238(.data_in(wire_d23_7),.data_out(wire_d23_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance240239(.data_in(wire_d23_8),.data_out(wire_d23_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402310(.data_in(wire_d23_9),.data_out(wire_d23_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402311(.data_in(wire_d23_10),.data_out(wire_d23_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2402312(.data_in(wire_d23_11),.data_out(wire_d23_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402313(.data_in(wire_d23_12),.data_out(wire_d23_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2402314(.data_in(wire_d23_13),.data_out(wire_d23_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402315(.data_in(wire_d23_14),.data_out(wire_d23_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2402316(.data_in(wire_d23_15),.data_out(wire_d23_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402317(.data_in(wire_d23_16),.data_out(wire_d23_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402318(.data_in(wire_d23_17),.data_out(wire_d23_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402319(.data_in(wire_d23_18),.data_out(wire_d23_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2402320(.data_in(wire_d23_19),.data_out(wire_d23_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402321(.data_in(wire_d23_20),.data_out(wire_d23_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402322(.data_in(wire_d23_21),.data_out(wire_d23_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402323(.data_in(wire_d23_22),.data_out(wire_d23_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402324(.data_in(wire_d23_23),.data_out(wire_d23_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402325(.data_in(wire_d23_24),.data_out(wire_d23_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402326(.data_in(wire_d23_25),.data_out(wire_d23_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402327(.data_in(wire_d23_26),.data_out(wire_d23_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402328(.data_in(wire_d23_27),.data_out(wire_d23_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402329(.data_in(wire_d23_28),.data_out(wire_d23_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402330(.data_in(wire_d23_29),.data_out(wire_d23_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402331(.data_in(wire_d23_30),.data_out(wire_d23_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402332(.data_in(wire_d23_31),.data_out(wire_d23_32),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402333(.data_in(wire_d23_32),.data_out(wire_d23_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402334(.data_in(wire_d23_33),.data_out(wire_d23_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402335(.data_in(wire_d23_34),.data_out(wire_d23_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2402336(.data_in(wire_d23_35),.data_out(wire_d23_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2402337(.data_in(wire_d23_36),.data_out(wire_d23_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402338(.data_in(wire_d23_37),.data_out(wire_d23_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402339(.data_in(wire_d23_38),.data_out(wire_d23_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402340(.data_in(wire_d23_39),.data_out(wire_d23_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402341(.data_in(wire_d23_40),.data_out(wire_d23_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2402342(.data_in(wire_d23_41),.data_out(wire_d23_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402343(.data_in(wire_d23_42),.data_out(wire_d23_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402344(.data_in(wire_d23_43),.data_out(wire_d23_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402345(.data_in(wire_d23_44),.data_out(wire_d23_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402346(.data_in(wire_d23_45),.data_out(wire_d23_46),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402347(.data_in(wire_d23_46),.data_out(wire_d23_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402348(.data_in(wire_d23_47),.data_out(wire_d23_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402349(.data_in(wire_d23_48),.data_out(wire_d23_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402350(.data_in(wire_d23_49),.data_out(wire_d23_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402351(.data_in(wire_d23_50),.data_out(wire_d23_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2402352(.data_in(wire_d23_51),.data_out(wire_d23_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2402353(.data_in(wire_d23_52),.data_out(wire_d23_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402354(.data_in(wire_d23_53),.data_out(wire_d23_54),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402355(.data_in(wire_d23_54),.data_out(wire_d23_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2402356(.data_in(wire_d23_55),.data_out(wire_d23_56),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402357(.data_in(wire_d23_56),.data_out(wire_d23_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2402358(.data_in(wire_d23_57),.data_out(wire_d23_58),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2402359(.data_in(wire_d23_58),.data_out(wire_d23_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402360(.data_in(wire_d23_59),.data_out(wire_d23_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402361(.data_in(wire_d23_60),.data_out(wire_d23_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402362(.data_in(wire_d23_61),.data_out(wire_d23_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402363(.data_in(wire_d23_62),.data_out(wire_d23_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2402364(.data_in(wire_d23_63),.data_out(wire_d23_64),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402365(.data_in(wire_d23_64),.data_out(wire_d23_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402366(.data_in(wire_d23_65),.data_out(wire_d23_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402367(.data_in(wire_d23_66),.data_out(wire_d23_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2402368(.data_in(wire_d23_67),.data_out(wire_d23_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402369(.data_in(wire_d23_68),.data_out(wire_d23_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402370(.data_in(wire_d23_69),.data_out(wire_d23_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402371(.data_in(wire_d23_70),.data_out(wire_d23_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2402372(.data_in(wire_d23_71),.data_out(wire_d23_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402373(.data_in(wire_d23_72),.data_out(wire_d23_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2402374(.data_in(wire_d23_73),.data_out(wire_d23_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402375(.data_in(wire_d23_74),.data_out(wire_d23_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402376(.data_in(wire_d23_75),.data_out(wire_d23_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402377(.data_in(wire_d23_76),.data_out(wire_d23_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402378(.data_in(wire_d23_77),.data_out(wire_d23_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402379(.data_in(wire_d23_78),.data_out(d_out23),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance250240(.data_in(d_in24),.data_out(wire_d24_0),.clk(clk),.rst(rst));            //channel 25
	register #(.WIDTH(WIDTH)) register_instance250241(.data_in(wire_d24_0),.data_out(wire_d24_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance250242(.data_in(wire_d24_1),.data_out(wire_d24_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance250243(.data_in(wire_d24_2),.data_out(wire_d24_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance250244(.data_in(wire_d24_3),.data_out(wire_d24_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance250245(.data_in(wire_d24_4),.data_out(wire_d24_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance250246(.data_in(wire_d24_5),.data_out(wire_d24_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance250247(.data_in(wire_d24_6),.data_out(wire_d24_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance250248(.data_in(wire_d24_7),.data_out(wire_d24_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance250249(.data_in(wire_d24_8),.data_out(wire_d24_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2502410(.data_in(wire_d24_9),.data_out(wire_d24_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502411(.data_in(wire_d24_10),.data_out(wire_d24_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2502412(.data_in(wire_d24_11),.data_out(wire_d24_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2502413(.data_in(wire_d24_12),.data_out(wire_d24_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502414(.data_in(wire_d24_13),.data_out(wire_d24_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502415(.data_in(wire_d24_14),.data_out(wire_d24_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502416(.data_in(wire_d24_15),.data_out(wire_d24_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502417(.data_in(wire_d24_16),.data_out(wire_d24_17),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2502418(.data_in(wire_d24_17),.data_out(wire_d24_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502419(.data_in(wire_d24_18),.data_out(wire_d24_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502420(.data_in(wire_d24_19),.data_out(wire_d24_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502421(.data_in(wire_d24_20),.data_out(wire_d24_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502422(.data_in(wire_d24_21),.data_out(wire_d24_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502423(.data_in(wire_d24_22),.data_out(wire_d24_23),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502424(.data_in(wire_d24_23),.data_out(wire_d24_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502425(.data_in(wire_d24_24),.data_out(wire_d24_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2502426(.data_in(wire_d24_25),.data_out(wire_d24_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2502427(.data_in(wire_d24_26),.data_out(wire_d24_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502428(.data_in(wire_d24_27),.data_out(wire_d24_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502429(.data_in(wire_d24_28),.data_out(wire_d24_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502430(.data_in(wire_d24_29),.data_out(wire_d24_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2502431(.data_in(wire_d24_30),.data_out(wire_d24_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502432(.data_in(wire_d24_31),.data_out(wire_d24_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502433(.data_in(wire_d24_32),.data_out(wire_d24_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502434(.data_in(wire_d24_33),.data_out(wire_d24_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502435(.data_in(wire_d24_34),.data_out(wire_d24_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502436(.data_in(wire_d24_35),.data_out(wire_d24_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2502437(.data_in(wire_d24_36),.data_out(wire_d24_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2502438(.data_in(wire_d24_37),.data_out(wire_d24_38),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502439(.data_in(wire_d24_38),.data_out(wire_d24_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502440(.data_in(wire_d24_39),.data_out(wire_d24_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2502441(.data_in(wire_d24_40),.data_out(wire_d24_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502442(.data_in(wire_d24_41),.data_out(wire_d24_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2502443(.data_in(wire_d24_42),.data_out(wire_d24_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502444(.data_in(wire_d24_43),.data_out(wire_d24_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2502445(.data_in(wire_d24_44),.data_out(wire_d24_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2502446(.data_in(wire_d24_45),.data_out(wire_d24_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502447(.data_in(wire_d24_46),.data_out(wire_d24_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2502448(.data_in(wire_d24_47),.data_out(wire_d24_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502449(.data_in(wire_d24_48),.data_out(wire_d24_49),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2502450(.data_in(wire_d24_49),.data_out(wire_d24_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502451(.data_in(wire_d24_50),.data_out(wire_d24_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502452(.data_in(wire_d24_51),.data_out(wire_d24_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502453(.data_in(wire_d24_52),.data_out(wire_d24_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502454(.data_in(wire_d24_53),.data_out(wire_d24_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502455(.data_in(wire_d24_54),.data_out(wire_d24_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502456(.data_in(wire_d24_55),.data_out(wire_d24_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502457(.data_in(wire_d24_56),.data_out(wire_d24_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502458(.data_in(wire_d24_57),.data_out(wire_d24_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2502459(.data_in(wire_d24_58),.data_out(wire_d24_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502460(.data_in(wire_d24_59),.data_out(wire_d24_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2502461(.data_in(wire_d24_60),.data_out(wire_d24_61),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502462(.data_in(wire_d24_61),.data_out(wire_d24_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502463(.data_in(wire_d24_62),.data_out(wire_d24_63),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502464(.data_in(wire_d24_63),.data_out(wire_d24_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502465(.data_in(wire_d24_64),.data_out(wire_d24_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2502466(.data_in(wire_d24_65),.data_out(wire_d24_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502467(.data_in(wire_d24_66),.data_out(wire_d24_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502468(.data_in(wire_d24_67),.data_out(wire_d24_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502469(.data_in(wire_d24_68),.data_out(wire_d24_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2502470(.data_in(wire_d24_69),.data_out(wire_d24_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502471(.data_in(wire_d24_70),.data_out(wire_d24_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2502472(.data_in(wire_d24_71),.data_out(wire_d24_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502473(.data_in(wire_d24_72),.data_out(wire_d24_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2502474(.data_in(wire_d24_73),.data_out(wire_d24_74),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502475(.data_in(wire_d24_74),.data_out(wire_d24_75),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502476(.data_in(wire_d24_75),.data_out(wire_d24_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502477(.data_in(wire_d24_76),.data_out(wire_d24_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2502478(.data_in(wire_d24_77),.data_out(wire_d24_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502479(.data_in(wire_d24_78),.data_out(d_out24),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance260250(.data_in(d_in25),.data_out(wire_d25_0),.clk(clk),.rst(rst));            //channel 26
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance260251(.data_in(wire_d25_0),.data_out(wire_d25_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance260252(.data_in(wire_d25_1),.data_out(wire_d25_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance260253(.data_in(wire_d25_2),.data_out(wire_d25_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance260254(.data_in(wire_d25_3),.data_out(wire_d25_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance260255(.data_in(wire_d25_4),.data_out(wire_d25_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance260256(.data_in(wire_d25_5),.data_out(wire_d25_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance260257(.data_in(wire_d25_6),.data_out(wire_d25_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance260258(.data_in(wire_d25_7),.data_out(wire_d25_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance260259(.data_in(wire_d25_8),.data_out(wire_d25_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602510(.data_in(wire_d25_9),.data_out(wire_d25_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2602511(.data_in(wire_d25_10),.data_out(wire_d25_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2602512(.data_in(wire_d25_11),.data_out(wire_d25_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2602513(.data_in(wire_d25_12),.data_out(wire_d25_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2602514(.data_in(wire_d25_13),.data_out(wire_d25_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602515(.data_in(wire_d25_14),.data_out(wire_d25_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602516(.data_in(wire_d25_15),.data_out(wire_d25_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602517(.data_in(wire_d25_16),.data_out(wire_d25_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2602518(.data_in(wire_d25_17),.data_out(wire_d25_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602519(.data_in(wire_d25_18),.data_out(wire_d25_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602520(.data_in(wire_d25_19),.data_out(wire_d25_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602521(.data_in(wire_d25_20),.data_out(wire_d25_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602522(.data_in(wire_d25_21),.data_out(wire_d25_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602523(.data_in(wire_d25_22),.data_out(wire_d25_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602524(.data_in(wire_d25_23),.data_out(wire_d25_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602525(.data_in(wire_d25_24),.data_out(wire_d25_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602526(.data_in(wire_d25_25),.data_out(wire_d25_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602527(.data_in(wire_d25_26),.data_out(wire_d25_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602528(.data_in(wire_d25_27),.data_out(wire_d25_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602529(.data_in(wire_d25_28),.data_out(wire_d25_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602530(.data_in(wire_d25_29),.data_out(wire_d25_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602531(.data_in(wire_d25_30),.data_out(wire_d25_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2602532(.data_in(wire_d25_31),.data_out(wire_d25_32),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602533(.data_in(wire_d25_32),.data_out(wire_d25_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602534(.data_in(wire_d25_33),.data_out(wire_d25_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602535(.data_in(wire_d25_34),.data_out(wire_d25_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602536(.data_in(wire_d25_35),.data_out(wire_d25_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602537(.data_in(wire_d25_36),.data_out(wire_d25_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602538(.data_in(wire_d25_37),.data_out(wire_d25_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602539(.data_in(wire_d25_38),.data_out(wire_d25_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2602540(.data_in(wire_d25_39),.data_out(wire_d25_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2602541(.data_in(wire_d25_40),.data_out(wire_d25_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602542(.data_in(wire_d25_41),.data_out(wire_d25_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2602543(.data_in(wire_d25_42),.data_out(wire_d25_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602544(.data_in(wire_d25_43),.data_out(wire_d25_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602545(.data_in(wire_d25_44),.data_out(wire_d25_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602546(.data_in(wire_d25_45),.data_out(wire_d25_46),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602547(.data_in(wire_d25_46),.data_out(wire_d25_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602548(.data_in(wire_d25_47),.data_out(wire_d25_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2602549(.data_in(wire_d25_48),.data_out(wire_d25_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602550(.data_in(wire_d25_49),.data_out(wire_d25_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602551(.data_in(wire_d25_50),.data_out(wire_d25_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602552(.data_in(wire_d25_51),.data_out(wire_d25_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602553(.data_in(wire_d25_52),.data_out(wire_d25_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602554(.data_in(wire_d25_53),.data_out(wire_d25_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2602555(.data_in(wire_d25_54),.data_out(wire_d25_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602556(.data_in(wire_d25_55),.data_out(wire_d25_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602557(.data_in(wire_d25_56),.data_out(wire_d25_57),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2602558(.data_in(wire_d25_57),.data_out(wire_d25_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602559(.data_in(wire_d25_58),.data_out(wire_d25_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602560(.data_in(wire_d25_59),.data_out(wire_d25_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602561(.data_in(wire_d25_60),.data_out(wire_d25_61),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602562(.data_in(wire_d25_61),.data_out(wire_d25_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602563(.data_in(wire_d25_62),.data_out(wire_d25_63),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602564(.data_in(wire_d25_63),.data_out(wire_d25_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602565(.data_in(wire_d25_64),.data_out(wire_d25_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602566(.data_in(wire_d25_65),.data_out(wire_d25_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2602567(.data_in(wire_d25_66),.data_out(wire_d25_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602568(.data_in(wire_d25_67),.data_out(wire_d25_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602569(.data_in(wire_d25_68),.data_out(wire_d25_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602570(.data_in(wire_d25_69),.data_out(wire_d25_70),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602571(.data_in(wire_d25_70),.data_out(wire_d25_71),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602572(.data_in(wire_d25_71),.data_out(wire_d25_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602573(.data_in(wire_d25_72),.data_out(wire_d25_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602574(.data_in(wire_d25_73),.data_out(wire_d25_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602575(.data_in(wire_d25_74),.data_out(wire_d25_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602576(.data_in(wire_d25_75),.data_out(wire_d25_76),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602577(.data_in(wire_d25_76),.data_out(wire_d25_77),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602578(.data_in(wire_d25_77),.data_out(wire_d25_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2602579(.data_in(wire_d25_78),.data_out(d_out25),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance270260(.data_in(d_in26),.data_out(wire_d26_0),.clk(clk),.rst(rst));            //channel 27
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance270261(.data_in(wire_d26_0),.data_out(wire_d26_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance270262(.data_in(wire_d26_1),.data_out(wire_d26_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance270263(.data_in(wire_d26_2),.data_out(wire_d26_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance270264(.data_in(wire_d26_3),.data_out(wire_d26_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance270265(.data_in(wire_d26_4),.data_out(wire_d26_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance270266(.data_in(wire_d26_5),.data_out(wire_d26_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance270267(.data_in(wire_d26_6),.data_out(wire_d26_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance270268(.data_in(wire_d26_7),.data_out(wire_d26_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance270269(.data_in(wire_d26_8),.data_out(wire_d26_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2702610(.data_in(wire_d26_9),.data_out(wire_d26_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702611(.data_in(wire_d26_10),.data_out(wire_d26_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702612(.data_in(wire_d26_11),.data_out(wire_d26_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702613(.data_in(wire_d26_12),.data_out(wire_d26_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702614(.data_in(wire_d26_13),.data_out(wire_d26_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2702615(.data_in(wire_d26_14),.data_out(wire_d26_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702616(.data_in(wire_d26_15),.data_out(wire_d26_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702617(.data_in(wire_d26_16),.data_out(wire_d26_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702618(.data_in(wire_d26_17),.data_out(wire_d26_18),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2702619(.data_in(wire_d26_18),.data_out(wire_d26_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702620(.data_in(wire_d26_19),.data_out(wire_d26_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702621(.data_in(wire_d26_20),.data_out(wire_d26_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702622(.data_in(wire_d26_21),.data_out(wire_d26_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702623(.data_in(wire_d26_22),.data_out(wire_d26_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702624(.data_in(wire_d26_23),.data_out(wire_d26_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702625(.data_in(wire_d26_24),.data_out(wire_d26_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702626(.data_in(wire_d26_25),.data_out(wire_d26_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702627(.data_in(wire_d26_26),.data_out(wire_d26_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702628(.data_in(wire_d26_27),.data_out(wire_d26_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702629(.data_in(wire_d26_28),.data_out(wire_d26_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702630(.data_in(wire_d26_29),.data_out(wire_d26_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702631(.data_in(wire_d26_30),.data_out(wire_d26_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702632(.data_in(wire_d26_31),.data_out(wire_d26_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702633(.data_in(wire_d26_32),.data_out(wire_d26_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702634(.data_in(wire_d26_33),.data_out(wire_d26_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702635(.data_in(wire_d26_34),.data_out(wire_d26_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702636(.data_in(wire_d26_35),.data_out(wire_d26_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702637(.data_in(wire_d26_36),.data_out(wire_d26_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2702638(.data_in(wire_d26_37),.data_out(wire_d26_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702639(.data_in(wire_d26_38),.data_out(wire_d26_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702640(.data_in(wire_d26_39),.data_out(wire_d26_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702641(.data_in(wire_d26_40),.data_out(wire_d26_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2702642(.data_in(wire_d26_41),.data_out(wire_d26_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702643(.data_in(wire_d26_42),.data_out(wire_d26_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702644(.data_in(wire_d26_43),.data_out(wire_d26_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702645(.data_in(wire_d26_44),.data_out(wire_d26_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702646(.data_in(wire_d26_45),.data_out(wire_d26_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702647(.data_in(wire_d26_46),.data_out(wire_d26_47),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2702648(.data_in(wire_d26_47),.data_out(wire_d26_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702649(.data_in(wire_d26_48),.data_out(wire_d26_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2702650(.data_in(wire_d26_49),.data_out(wire_d26_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702651(.data_in(wire_d26_50),.data_out(wire_d26_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702652(.data_in(wire_d26_51),.data_out(wire_d26_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702653(.data_in(wire_d26_52),.data_out(wire_d26_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702654(.data_in(wire_d26_53),.data_out(wire_d26_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702655(.data_in(wire_d26_54),.data_out(wire_d26_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2702656(.data_in(wire_d26_55),.data_out(wire_d26_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702657(.data_in(wire_d26_56),.data_out(wire_d26_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2702658(.data_in(wire_d26_57),.data_out(wire_d26_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702659(.data_in(wire_d26_58),.data_out(wire_d26_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702660(.data_in(wire_d26_59),.data_out(wire_d26_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702661(.data_in(wire_d26_60),.data_out(wire_d26_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702662(.data_in(wire_d26_61),.data_out(wire_d26_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702663(.data_in(wire_d26_62),.data_out(wire_d26_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2702664(.data_in(wire_d26_63),.data_out(wire_d26_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702665(.data_in(wire_d26_64),.data_out(wire_d26_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702666(.data_in(wire_d26_65),.data_out(wire_d26_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702667(.data_in(wire_d26_66),.data_out(wire_d26_67),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702668(.data_in(wire_d26_67),.data_out(wire_d26_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2702669(.data_in(wire_d26_68),.data_out(wire_d26_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702670(.data_in(wire_d26_69),.data_out(wire_d26_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2702671(.data_in(wire_d26_70),.data_out(wire_d26_71),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702672(.data_in(wire_d26_71),.data_out(wire_d26_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702673(.data_in(wire_d26_72),.data_out(wire_d26_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702674(.data_in(wire_d26_73),.data_out(wire_d26_74),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702675(.data_in(wire_d26_74),.data_out(wire_d26_75),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702676(.data_in(wire_d26_75),.data_out(wire_d26_76),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702677(.data_in(wire_d26_76),.data_out(wire_d26_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702678(.data_in(wire_d26_77),.data_out(wire_d26_78),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702679(.data_in(wire_d26_78),.data_out(d_out26),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance280270(.data_in(d_in27),.data_out(wire_d27_0),.clk(clk),.rst(rst));            //channel 28
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance280271(.data_in(wire_d27_0),.data_out(wire_d27_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance280272(.data_in(wire_d27_1),.data_out(wire_d27_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance280273(.data_in(wire_d27_2),.data_out(wire_d27_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance280274(.data_in(wire_d27_3),.data_out(wire_d27_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance280275(.data_in(wire_d27_4),.data_out(wire_d27_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance280276(.data_in(wire_d27_5),.data_out(wire_d27_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance280277(.data_in(wire_d27_6),.data_out(wire_d27_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance280278(.data_in(wire_d27_7),.data_out(wire_d27_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance280279(.data_in(wire_d27_8),.data_out(wire_d27_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802710(.data_in(wire_d27_9),.data_out(wire_d27_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802711(.data_in(wire_d27_10),.data_out(wire_d27_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802712(.data_in(wire_d27_11),.data_out(wire_d27_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802713(.data_in(wire_d27_12),.data_out(wire_d27_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802714(.data_in(wire_d27_13),.data_out(wire_d27_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802715(.data_in(wire_d27_14),.data_out(wire_d27_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802716(.data_in(wire_d27_15),.data_out(wire_d27_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802717(.data_in(wire_d27_16),.data_out(wire_d27_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802718(.data_in(wire_d27_17),.data_out(wire_d27_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802719(.data_in(wire_d27_18),.data_out(wire_d27_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802720(.data_in(wire_d27_19),.data_out(wire_d27_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802721(.data_in(wire_d27_20),.data_out(wire_d27_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802722(.data_in(wire_d27_21),.data_out(wire_d27_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802723(.data_in(wire_d27_22),.data_out(wire_d27_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802724(.data_in(wire_d27_23),.data_out(wire_d27_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802725(.data_in(wire_d27_24),.data_out(wire_d27_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802726(.data_in(wire_d27_25),.data_out(wire_d27_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802727(.data_in(wire_d27_26),.data_out(wire_d27_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802728(.data_in(wire_d27_27),.data_out(wire_d27_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802729(.data_in(wire_d27_28),.data_out(wire_d27_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802730(.data_in(wire_d27_29),.data_out(wire_d27_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802731(.data_in(wire_d27_30),.data_out(wire_d27_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802732(.data_in(wire_d27_31),.data_out(wire_d27_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802733(.data_in(wire_d27_32),.data_out(wire_d27_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802734(.data_in(wire_d27_33),.data_out(wire_d27_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802735(.data_in(wire_d27_34),.data_out(wire_d27_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802736(.data_in(wire_d27_35),.data_out(wire_d27_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802737(.data_in(wire_d27_36),.data_out(wire_d27_37),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802738(.data_in(wire_d27_37),.data_out(wire_d27_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802739(.data_in(wire_d27_38),.data_out(wire_d27_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802740(.data_in(wire_d27_39),.data_out(wire_d27_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802741(.data_in(wire_d27_40),.data_out(wire_d27_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802742(.data_in(wire_d27_41),.data_out(wire_d27_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802743(.data_in(wire_d27_42),.data_out(wire_d27_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802744(.data_in(wire_d27_43),.data_out(wire_d27_44),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802745(.data_in(wire_d27_44),.data_out(wire_d27_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802746(.data_in(wire_d27_45),.data_out(wire_d27_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802747(.data_in(wire_d27_46),.data_out(wire_d27_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802748(.data_in(wire_d27_47),.data_out(wire_d27_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802749(.data_in(wire_d27_48),.data_out(wire_d27_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802750(.data_in(wire_d27_49),.data_out(wire_d27_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802751(.data_in(wire_d27_50),.data_out(wire_d27_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802752(.data_in(wire_d27_51),.data_out(wire_d27_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802753(.data_in(wire_d27_52),.data_out(wire_d27_53),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802754(.data_in(wire_d27_53),.data_out(wire_d27_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802755(.data_in(wire_d27_54),.data_out(wire_d27_55),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802756(.data_in(wire_d27_55),.data_out(wire_d27_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802757(.data_in(wire_d27_56),.data_out(wire_d27_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802758(.data_in(wire_d27_57),.data_out(wire_d27_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802759(.data_in(wire_d27_58),.data_out(wire_d27_59),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802760(.data_in(wire_d27_59),.data_out(wire_d27_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802761(.data_in(wire_d27_60),.data_out(wire_d27_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802762(.data_in(wire_d27_61),.data_out(wire_d27_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802763(.data_in(wire_d27_62),.data_out(wire_d27_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802764(.data_in(wire_d27_63),.data_out(wire_d27_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802765(.data_in(wire_d27_64),.data_out(wire_d27_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802766(.data_in(wire_d27_65),.data_out(wire_d27_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802767(.data_in(wire_d27_66),.data_out(wire_d27_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802768(.data_in(wire_d27_67),.data_out(wire_d27_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802769(.data_in(wire_d27_68),.data_out(wire_d27_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802770(.data_in(wire_d27_69),.data_out(wire_d27_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802771(.data_in(wire_d27_70),.data_out(wire_d27_71),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802772(.data_in(wire_d27_71),.data_out(wire_d27_72),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802773(.data_in(wire_d27_72),.data_out(wire_d27_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802774(.data_in(wire_d27_73),.data_out(wire_d27_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802775(.data_in(wire_d27_74),.data_out(wire_d27_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802776(.data_in(wire_d27_75),.data_out(wire_d27_76),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802777(.data_in(wire_d27_76),.data_out(wire_d27_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802778(.data_in(wire_d27_77),.data_out(wire_d27_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802779(.data_in(wire_d27_78),.data_out(d_out27),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance290280(.data_in(d_in28),.data_out(wire_d28_0),.clk(clk),.rst(rst));            //channel 29
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance290281(.data_in(wire_d28_0),.data_out(wire_d28_1),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance290282(.data_in(wire_d28_1),.data_out(wire_d28_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance290283(.data_in(wire_d28_2),.data_out(wire_d28_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance290284(.data_in(wire_d28_3),.data_out(wire_d28_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance290285(.data_in(wire_d28_4),.data_out(wire_d28_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance290286(.data_in(wire_d28_5),.data_out(wire_d28_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance290287(.data_in(wire_d28_6),.data_out(wire_d28_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance290288(.data_in(wire_d28_7),.data_out(wire_d28_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance290289(.data_in(wire_d28_8),.data_out(wire_d28_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902810(.data_in(wire_d28_9),.data_out(wire_d28_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902811(.data_in(wire_d28_10),.data_out(wire_d28_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902812(.data_in(wire_d28_11),.data_out(wire_d28_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902813(.data_in(wire_d28_12),.data_out(wire_d28_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902814(.data_in(wire_d28_13),.data_out(wire_d28_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902815(.data_in(wire_d28_14),.data_out(wire_d28_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902816(.data_in(wire_d28_15),.data_out(wire_d28_16),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902817(.data_in(wire_d28_16),.data_out(wire_d28_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902818(.data_in(wire_d28_17),.data_out(wire_d28_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2902819(.data_in(wire_d28_18),.data_out(wire_d28_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902820(.data_in(wire_d28_19),.data_out(wire_d28_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902821(.data_in(wire_d28_20),.data_out(wire_d28_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902822(.data_in(wire_d28_21),.data_out(wire_d28_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902823(.data_in(wire_d28_22),.data_out(wire_d28_23),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902824(.data_in(wire_d28_23),.data_out(wire_d28_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902825(.data_in(wire_d28_24),.data_out(wire_d28_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902826(.data_in(wire_d28_25),.data_out(wire_d28_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902827(.data_in(wire_d28_26),.data_out(wire_d28_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902828(.data_in(wire_d28_27),.data_out(wire_d28_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902829(.data_in(wire_d28_28),.data_out(wire_d28_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902830(.data_in(wire_d28_29),.data_out(wire_d28_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902831(.data_in(wire_d28_30),.data_out(wire_d28_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2902832(.data_in(wire_d28_31),.data_out(wire_d28_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902833(.data_in(wire_d28_32),.data_out(wire_d28_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902834(.data_in(wire_d28_33),.data_out(wire_d28_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902835(.data_in(wire_d28_34),.data_out(wire_d28_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902836(.data_in(wire_d28_35),.data_out(wire_d28_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902837(.data_in(wire_d28_36),.data_out(wire_d28_37),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902838(.data_in(wire_d28_37),.data_out(wire_d28_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902839(.data_in(wire_d28_38),.data_out(wire_d28_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902840(.data_in(wire_d28_39),.data_out(wire_d28_40),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902841(.data_in(wire_d28_40),.data_out(wire_d28_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902842(.data_in(wire_d28_41),.data_out(wire_d28_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2902843(.data_in(wire_d28_42),.data_out(wire_d28_43),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902844(.data_in(wire_d28_43),.data_out(wire_d28_44),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902845(.data_in(wire_d28_44),.data_out(wire_d28_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902846(.data_in(wire_d28_45),.data_out(wire_d28_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902847(.data_in(wire_d28_46),.data_out(wire_d28_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902848(.data_in(wire_d28_47),.data_out(wire_d28_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902849(.data_in(wire_d28_48),.data_out(wire_d28_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2902850(.data_in(wire_d28_49),.data_out(wire_d28_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902851(.data_in(wire_d28_50),.data_out(wire_d28_51),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902852(.data_in(wire_d28_51),.data_out(wire_d28_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902853(.data_in(wire_d28_52),.data_out(wire_d28_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902854(.data_in(wire_d28_53),.data_out(wire_d28_54),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902855(.data_in(wire_d28_54),.data_out(wire_d28_55),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902856(.data_in(wire_d28_55),.data_out(wire_d28_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902857(.data_in(wire_d28_56),.data_out(wire_d28_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902858(.data_in(wire_d28_57),.data_out(wire_d28_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902859(.data_in(wire_d28_58),.data_out(wire_d28_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902860(.data_in(wire_d28_59),.data_out(wire_d28_60),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902861(.data_in(wire_d28_60),.data_out(wire_d28_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902862(.data_in(wire_d28_61),.data_out(wire_d28_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902863(.data_in(wire_d28_62),.data_out(wire_d28_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902864(.data_in(wire_d28_63),.data_out(wire_d28_64),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902865(.data_in(wire_d28_64),.data_out(wire_d28_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902866(.data_in(wire_d28_65),.data_out(wire_d28_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902867(.data_in(wire_d28_66),.data_out(wire_d28_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2902868(.data_in(wire_d28_67),.data_out(wire_d28_68),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902869(.data_in(wire_d28_68),.data_out(wire_d28_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2902870(.data_in(wire_d28_69),.data_out(wire_d28_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902871(.data_in(wire_d28_70),.data_out(wire_d28_71),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902872(.data_in(wire_d28_71),.data_out(wire_d28_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902873(.data_in(wire_d28_72),.data_out(wire_d28_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902874(.data_in(wire_d28_73),.data_out(wire_d28_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902875(.data_in(wire_d28_74),.data_out(wire_d28_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2902876(.data_in(wire_d28_75),.data_out(wire_d28_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902877(.data_in(wire_d28_76),.data_out(wire_d28_77),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902878(.data_in(wire_d28_77),.data_out(wire_d28_78),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902879(.data_in(wire_d28_78),.data_out(d_out28),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance300290(.data_in(d_in29),.data_out(wire_d29_0),.clk(clk),.rst(rst));            //channel 30
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance300291(.data_in(wire_d29_0),.data_out(wire_d29_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance300292(.data_in(wire_d29_1),.data_out(wire_d29_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance300293(.data_in(wire_d29_2),.data_out(wire_d29_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance300294(.data_in(wire_d29_3),.data_out(wire_d29_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance300295(.data_in(wire_d29_4),.data_out(wire_d29_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance300296(.data_in(wire_d29_5),.data_out(wire_d29_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance300297(.data_in(wire_d29_6),.data_out(wire_d29_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance300298(.data_in(wire_d29_7),.data_out(wire_d29_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance300299(.data_in(wire_d29_8),.data_out(wire_d29_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002910(.data_in(wire_d29_9),.data_out(wire_d29_10),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002911(.data_in(wire_d29_10),.data_out(wire_d29_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002912(.data_in(wire_d29_11),.data_out(wire_d29_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002913(.data_in(wire_d29_12),.data_out(wire_d29_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002914(.data_in(wire_d29_13),.data_out(wire_d29_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002915(.data_in(wire_d29_14),.data_out(wire_d29_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002916(.data_in(wire_d29_15),.data_out(wire_d29_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002917(.data_in(wire_d29_16),.data_out(wire_d29_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3002918(.data_in(wire_d29_17),.data_out(wire_d29_18),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002919(.data_in(wire_d29_18),.data_out(wire_d29_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3002920(.data_in(wire_d29_19),.data_out(wire_d29_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002921(.data_in(wire_d29_20),.data_out(wire_d29_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002922(.data_in(wire_d29_21),.data_out(wire_d29_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3002923(.data_in(wire_d29_22),.data_out(wire_d29_23),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002924(.data_in(wire_d29_23),.data_out(wire_d29_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002925(.data_in(wire_d29_24),.data_out(wire_d29_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002926(.data_in(wire_d29_25),.data_out(wire_d29_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002927(.data_in(wire_d29_26),.data_out(wire_d29_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002928(.data_in(wire_d29_27),.data_out(wire_d29_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002929(.data_in(wire_d29_28),.data_out(wire_d29_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002930(.data_in(wire_d29_29),.data_out(wire_d29_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3002931(.data_in(wire_d29_30),.data_out(wire_d29_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002932(.data_in(wire_d29_31),.data_out(wire_d29_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002933(.data_in(wire_d29_32),.data_out(wire_d29_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002934(.data_in(wire_d29_33),.data_out(wire_d29_34),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002935(.data_in(wire_d29_34),.data_out(wire_d29_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002936(.data_in(wire_d29_35),.data_out(wire_d29_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002937(.data_in(wire_d29_36),.data_out(wire_d29_37),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002938(.data_in(wire_d29_37),.data_out(wire_d29_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002939(.data_in(wire_d29_38),.data_out(wire_d29_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002940(.data_in(wire_d29_39),.data_out(wire_d29_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002941(.data_in(wire_d29_40),.data_out(wire_d29_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3002942(.data_in(wire_d29_41),.data_out(wire_d29_42),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002943(.data_in(wire_d29_42),.data_out(wire_d29_43),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002944(.data_in(wire_d29_43),.data_out(wire_d29_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002945(.data_in(wire_d29_44),.data_out(wire_d29_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002946(.data_in(wire_d29_45),.data_out(wire_d29_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002947(.data_in(wire_d29_46),.data_out(wire_d29_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002948(.data_in(wire_d29_47),.data_out(wire_d29_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002949(.data_in(wire_d29_48),.data_out(wire_d29_49),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3002950(.data_in(wire_d29_49),.data_out(wire_d29_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002951(.data_in(wire_d29_50),.data_out(wire_d29_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002952(.data_in(wire_d29_51),.data_out(wire_d29_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002953(.data_in(wire_d29_52),.data_out(wire_d29_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002954(.data_in(wire_d29_53),.data_out(wire_d29_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002955(.data_in(wire_d29_54),.data_out(wire_d29_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002956(.data_in(wire_d29_55),.data_out(wire_d29_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002957(.data_in(wire_d29_56),.data_out(wire_d29_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002958(.data_in(wire_d29_57),.data_out(wire_d29_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002959(.data_in(wire_d29_58),.data_out(wire_d29_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3002960(.data_in(wire_d29_59),.data_out(wire_d29_60),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002961(.data_in(wire_d29_60),.data_out(wire_d29_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002962(.data_in(wire_d29_61),.data_out(wire_d29_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002963(.data_in(wire_d29_62),.data_out(wire_d29_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002964(.data_in(wire_d29_63),.data_out(wire_d29_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002965(.data_in(wire_d29_64),.data_out(wire_d29_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002966(.data_in(wire_d29_65),.data_out(wire_d29_66),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002967(.data_in(wire_d29_66),.data_out(wire_d29_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002968(.data_in(wire_d29_67),.data_out(wire_d29_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002969(.data_in(wire_d29_68),.data_out(wire_d29_69),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3002970(.data_in(wire_d29_69),.data_out(wire_d29_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002971(.data_in(wire_d29_70),.data_out(wire_d29_71),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002972(.data_in(wire_d29_71),.data_out(wire_d29_72),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002973(.data_in(wire_d29_72),.data_out(wire_d29_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002974(.data_in(wire_d29_73),.data_out(wire_d29_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002975(.data_in(wire_d29_74),.data_out(wire_d29_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002976(.data_in(wire_d29_75),.data_out(wire_d29_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002977(.data_in(wire_d29_76),.data_out(wire_d29_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002978(.data_in(wire_d29_77),.data_out(wire_d29_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002979(.data_in(wire_d29_78),.data_out(d_out29),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance310300(.data_in(d_in30),.data_out(wire_d30_0),.clk(clk),.rst(rst));            //channel 31
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance310301(.data_in(wire_d30_0),.data_out(wire_d30_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance310302(.data_in(wire_d30_1),.data_out(wire_d30_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance310303(.data_in(wire_d30_2),.data_out(wire_d30_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance310304(.data_in(wire_d30_3),.data_out(wire_d30_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance310305(.data_in(wire_d30_4),.data_out(wire_d30_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance310306(.data_in(wire_d30_5),.data_out(wire_d30_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance310307(.data_in(wire_d30_6),.data_out(wire_d30_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance310308(.data_in(wire_d30_7),.data_out(wire_d30_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance310309(.data_in(wire_d30_8),.data_out(wire_d30_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103010(.data_in(wire_d30_9),.data_out(wire_d30_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3103011(.data_in(wire_d30_10),.data_out(wire_d30_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103012(.data_in(wire_d30_11),.data_out(wire_d30_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3103013(.data_in(wire_d30_12),.data_out(wire_d30_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103014(.data_in(wire_d30_13),.data_out(wire_d30_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3103015(.data_in(wire_d30_14),.data_out(wire_d30_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103016(.data_in(wire_d30_15),.data_out(wire_d30_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103017(.data_in(wire_d30_16),.data_out(wire_d30_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3103018(.data_in(wire_d30_17),.data_out(wire_d30_18),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103019(.data_in(wire_d30_18),.data_out(wire_d30_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3103020(.data_in(wire_d30_19),.data_out(wire_d30_20),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103021(.data_in(wire_d30_20),.data_out(wire_d30_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103022(.data_in(wire_d30_21),.data_out(wire_d30_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103023(.data_in(wire_d30_22),.data_out(wire_d30_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103024(.data_in(wire_d30_23),.data_out(wire_d30_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103025(.data_in(wire_d30_24),.data_out(wire_d30_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103026(.data_in(wire_d30_25),.data_out(wire_d30_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3103027(.data_in(wire_d30_26),.data_out(wire_d30_27),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3103028(.data_in(wire_d30_27),.data_out(wire_d30_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103029(.data_in(wire_d30_28),.data_out(wire_d30_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103030(.data_in(wire_d30_29),.data_out(wire_d30_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3103031(.data_in(wire_d30_30),.data_out(wire_d30_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103032(.data_in(wire_d30_31),.data_out(wire_d30_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103033(.data_in(wire_d30_32),.data_out(wire_d30_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3103034(.data_in(wire_d30_33),.data_out(wire_d30_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3103035(.data_in(wire_d30_34),.data_out(wire_d30_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103036(.data_in(wire_d30_35),.data_out(wire_d30_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103037(.data_in(wire_d30_36),.data_out(wire_d30_37),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103038(.data_in(wire_d30_37),.data_out(wire_d30_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103039(.data_in(wire_d30_38),.data_out(wire_d30_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103040(.data_in(wire_d30_39),.data_out(wire_d30_40),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103041(.data_in(wire_d30_40),.data_out(wire_d30_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103042(.data_in(wire_d30_41),.data_out(wire_d30_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3103043(.data_in(wire_d30_42),.data_out(wire_d30_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103044(.data_in(wire_d30_43),.data_out(wire_d30_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103045(.data_in(wire_d30_44),.data_out(wire_d30_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103046(.data_in(wire_d30_45),.data_out(wire_d30_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103047(.data_in(wire_d30_46),.data_out(wire_d30_47),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103048(.data_in(wire_d30_47),.data_out(wire_d30_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103049(.data_in(wire_d30_48),.data_out(wire_d30_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103050(.data_in(wire_d30_49),.data_out(wire_d30_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103051(.data_in(wire_d30_50),.data_out(wire_d30_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103052(.data_in(wire_d30_51),.data_out(wire_d30_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103053(.data_in(wire_d30_52),.data_out(wire_d30_53),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103054(.data_in(wire_d30_53),.data_out(wire_d30_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103055(.data_in(wire_d30_54),.data_out(wire_d30_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103056(.data_in(wire_d30_55),.data_out(wire_d30_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103057(.data_in(wire_d30_56),.data_out(wire_d30_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3103058(.data_in(wire_d30_57),.data_out(wire_d30_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103059(.data_in(wire_d30_58),.data_out(wire_d30_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103060(.data_in(wire_d30_59),.data_out(wire_d30_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3103061(.data_in(wire_d30_60),.data_out(wire_d30_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103062(.data_in(wire_d30_61),.data_out(wire_d30_62),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103063(.data_in(wire_d30_62),.data_out(wire_d30_63),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103064(.data_in(wire_d30_63),.data_out(wire_d30_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103065(.data_in(wire_d30_64),.data_out(wire_d30_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103066(.data_in(wire_d30_65),.data_out(wire_d30_66),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103067(.data_in(wire_d30_66),.data_out(wire_d30_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103068(.data_in(wire_d30_67),.data_out(wire_d30_68),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103069(.data_in(wire_d30_68),.data_out(wire_d30_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103070(.data_in(wire_d30_69),.data_out(wire_d30_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103071(.data_in(wire_d30_70),.data_out(wire_d30_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103072(.data_in(wire_d30_71),.data_out(wire_d30_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103073(.data_in(wire_d30_72),.data_out(wire_d30_73),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103074(.data_in(wire_d30_73),.data_out(wire_d30_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103075(.data_in(wire_d30_74),.data_out(wire_d30_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3103076(.data_in(wire_d30_75),.data_out(wire_d30_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103077(.data_in(wire_d30_76),.data_out(wire_d30_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103078(.data_in(wire_d30_77),.data_out(wire_d30_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103079(.data_in(wire_d30_78),.data_out(d_out30),.clk(clk),.rst(rst));

	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance320310(.data_in(d_in31),.data_out(wire_d31_0),.clk(clk),.rst(rst));            //channel 32
	decoder_top #(.WIDTH(WIDTH)) decoder_instance320311(.data_in(wire_d31_0),.data_out(wire_d31_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance320312(.data_in(wire_d31_1),.data_out(wire_d31_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance320313(.data_in(wire_d31_2),.data_out(wire_d31_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance320314(.data_in(wire_d31_3),.data_out(wire_d31_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance320315(.data_in(wire_d31_4),.data_out(wire_d31_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance320316(.data_in(wire_d31_5),.data_out(wire_d31_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance320317(.data_in(wire_d31_6),.data_out(wire_d31_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance320318(.data_in(wire_d31_7),.data_out(wire_d31_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance320319(.data_in(wire_d31_8),.data_out(wire_d31_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203110(.data_in(wire_d31_9),.data_out(wire_d31_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203111(.data_in(wire_d31_10),.data_out(wire_d31_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203112(.data_in(wire_d31_11),.data_out(wire_d31_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203113(.data_in(wire_d31_12),.data_out(wire_d31_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203114(.data_in(wire_d31_13),.data_out(wire_d31_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203115(.data_in(wire_d31_14),.data_out(wire_d31_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203116(.data_in(wire_d31_15),.data_out(wire_d31_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203117(.data_in(wire_d31_16),.data_out(wire_d31_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203118(.data_in(wire_d31_17),.data_out(wire_d31_18),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203119(.data_in(wire_d31_18),.data_out(wire_d31_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203120(.data_in(wire_d31_19),.data_out(wire_d31_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203121(.data_in(wire_d31_20),.data_out(wire_d31_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203122(.data_in(wire_d31_21),.data_out(wire_d31_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203123(.data_in(wire_d31_22),.data_out(wire_d31_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203124(.data_in(wire_d31_23),.data_out(wire_d31_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203125(.data_in(wire_d31_24),.data_out(wire_d31_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203126(.data_in(wire_d31_25),.data_out(wire_d31_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203127(.data_in(wire_d31_26),.data_out(wire_d31_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203128(.data_in(wire_d31_27),.data_out(wire_d31_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203129(.data_in(wire_d31_28),.data_out(wire_d31_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203130(.data_in(wire_d31_29),.data_out(wire_d31_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203131(.data_in(wire_d31_30),.data_out(wire_d31_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203132(.data_in(wire_d31_31),.data_out(wire_d31_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203133(.data_in(wire_d31_32),.data_out(wire_d31_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203134(.data_in(wire_d31_33),.data_out(wire_d31_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203135(.data_in(wire_d31_34),.data_out(wire_d31_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203136(.data_in(wire_d31_35),.data_out(wire_d31_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203137(.data_in(wire_d31_36),.data_out(wire_d31_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203138(.data_in(wire_d31_37),.data_out(wire_d31_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203139(.data_in(wire_d31_38),.data_out(wire_d31_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203140(.data_in(wire_d31_39),.data_out(wire_d31_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203141(.data_in(wire_d31_40),.data_out(wire_d31_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203142(.data_in(wire_d31_41),.data_out(wire_d31_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203143(.data_in(wire_d31_42),.data_out(wire_d31_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203144(.data_in(wire_d31_43),.data_out(wire_d31_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203145(.data_in(wire_d31_44),.data_out(wire_d31_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203146(.data_in(wire_d31_45),.data_out(wire_d31_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203147(.data_in(wire_d31_46),.data_out(wire_d31_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203148(.data_in(wire_d31_47),.data_out(wire_d31_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203149(.data_in(wire_d31_48),.data_out(wire_d31_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203150(.data_in(wire_d31_49),.data_out(wire_d31_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203151(.data_in(wire_d31_50),.data_out(wire_d31_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203152(.data_in(wire_d31_51),.data_out(wire_d31_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203153(.data_in(wire_d31_52),.data_out(wire_d31_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203154(.data_in(wire_d31_53),.data_out(wire_d31_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203155(.data_in(wire_d31_54),.data_out(wire_d31_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203156(.data_in(wire_d31_55),.data_out(wire_d31_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203157(.data_in(wire_d31_56),.data_out(wire_d31_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203158(.data_in(wire_d31_57),.data_out(wire_d31_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203159(.data_in(wire_d31_58),.data_out(wire_d31_59),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203160(.data_in(wire_d31_59),.data_out(wire_d31_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203161(.data_in(wire_d31_60),.data_out(wire_d31_61),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203162(.data_in(wire_d31_61),.data_out(wire_d31_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203163(.data_in(wire_d31_62),.data_out(wire_d31_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203164(.data_in(wire_d31_63),.data_out(wire_d31_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203165(.data_in(wire_d31_64),.data_out(wire_d31_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203166(.data_in(wire_d31_65),.data_out(wire_d31_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203167(.data_in(wire_d31_66),.data_out(wire_d31_67),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203168(.data_in(wire_d31_67),.data_out(wire_d31_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203169(.data_in(wire_d31_68),.data_out(wire_d31_69),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203170(.data_in(wire_d31_69),.data_out(wire_d31_70),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203171(.data_in(wire_d31_70),.data_out(wire_d31_71),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203172(.data_in(wire_d31_71),.data_out(wire_d31_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203173(.data_in(wire_d31_72),.data_out(wire_d31_73),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203174(.data_in(wire_d31_73),.data_out(wire_d31_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203175(.data_in(wire_d31_74),.data_out(wire_d31_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203176(.data_in(wire_d31_75),.data_out(wire_d31_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203177(.data_in(wire_d31_76),.data_out(wire_d31_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203178(.data_in(wire_d31_77),.data_out(wire_d31_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203179(.data_in(wire_d31_78),.data_out(d_out31),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance330320(.data_in(d_in32),.data_out(wire_d32_0),.clk(clk),.rst(rst));            //channel 33
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance330321(.data_in(wire_d32_0),.data_out(wire_d32_1),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance330322(.data_in(wire_d32_1),.data_out(wire_d32_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance330323(.data_in(wire_d32_2),.data_out(wire_d32_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance330324(.data_in(wire_d32_3),.data_out(wire_d32_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance330325(.data_in(wire_d32_4),.data_out(wire_d32_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance330326(.data_in(wire_d32_5),.data_out(wire_d32_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance330327(.data_in(wire_d32_6),.data_out(wire_d32_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance330328(.data_in(wire_d32_7),.data_out(wire_d32_8),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance330329(.data_in(wire_d32_8),.data_out(wire_d32_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303210(.data_in(wire_d32_9),.data_out(wire_d32_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303211(.data_in(wire_d32_10),.data_out(wire_d32_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303212(.data_in(wire_d32_11),.data_out(wire_d32_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303213(.data_in(wire_d32_12),.data_out(wire_d32_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303214(.data_in(wire_d32_13),.data_out(wire_d32_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303215(.data_in(wire_d32_14),.data_out(wire_d32_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303216(.data_in(wire_d32_15),.data_out(wire_d32_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303217(.data_in(wire_d32_16),.data_out(wire_d32_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303218(.data_in(wire_d32_17),.data_out(wire_d32_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303219(.data_in(wire_d32_18),.data_out(wire_d32_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303220(.data_in(wire_d32_19),.data_out(wire_d32_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303221(.data_in(wire_d32_20),.data_out(wire_d32_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303222(.data_in(wire_d32_21),.data_out(wire_d32_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303223(.data_in(wire_d32_22),.data_out(wire_d32_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303224(.data_in(wire_d32_23),.data_out(wire_d32_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3303225(.data_in(wire_d32_24),.data_out(wire_d32_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303226(.data_in(wire_d32_25),.data_out(wire_d32_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303227(.data_in(wire_d32_26),.data_out(wire_d32_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303228(.data_in(wire_d32_27),.data_out(wire_d32_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303229(.data_in(wire_d32_28),.data_out(wire_d32_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303230(.data_in(wire_d32_29),.data_out(wire_d32_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303231(.data_in(wire_d32_30),.data_out(wire_d32_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303232(.data_in(wire_d32_31),.data_out(wire_d32_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3303233(.data_in(wire_d32_32),.data_out(wire_d32_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3303234(.data_in(wire_d32_33),.data_out(wire_d32_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303235(.data_in(wire_d32_34),.data_out(wire_d32_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303236(.data_in(wire_d32_35),.data_out(wire_d32_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303237(.data_in(wire_d32_36),.data_out(wire_d32_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303238(.data_in(wire_d32_37),.data_out(wire_d32_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303239(.data_in(wire_d32_38),.data_out(wire_d32_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303240(.data_in(wire_d32_39),.data_out(wire_d32_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303241(.data_in(wire_d32_40),.data_out(wire_d32_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303242(.data_in(wire_d32_41),.data_out(wire_d32_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3303243(.data_in(wire_d32_42),.data_out(wire_d32_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303244(.data_in(wire_d32_43),.data_out(wire_d32_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303245(.data_in(wire_d32_44),.data_out(wire_d32_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303246(.data_in(wire_d32_45),.data_out(wire_d32_46),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303247(.data_in(wire_d32_46),.data_out(wire_d32_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303248(.data_in(wire_d32_47),.data_out(wire_d32_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3303249(.data_in(wire_d32_48),.data_out(wire_d32_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303250(.data_in(wire_d32_49),.data_out(wire_d32_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303251(.data_in(wire_d32_50),.data_out(wire_d32_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303252(.data_in(wire_d32_51),.data_out(wire_d32_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303253(.data_in(wire_d32_52),.data_out(wire_d32_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303254(.data_in(wire_d32_53),.data_out(wire_d32_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303255(.data_in(wire_d32_54),.data_out(wire_d32_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303256(.data_in(wire_d32_55),.data_out(wire_d32_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303257(.data_in(wire_d32_56),.data_out(wire_d32_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303258(.data_in(wire_d32_57),.data_out(wire_d32_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3303259(.data_in(wire_d32_58),.data_out(wire_d32_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303260(.data_in(wire_d32_59),.data_out(wire_d32_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303261(.data_in(wire_d32_60),.data_out(wire_d32_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303262(.data_in(wire_d32_61),.data_out(wire_d32_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303263(.data_in(wire_d32_62),.data_out(wire_d32_63),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303264(.data_in(wire_d32_63),.data_out(wire_d32_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303265(.data_in(wire_d32_64),.data_out(wire_d32_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303266(.data_in(wire_d32_65),.data_out(wire_d32_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303267(.data_in(wire_d32_66),.data_out(wire_d32_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303268(.data_in(wire_d32_67),.data_out(wire_d32_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303269(.data_in(wire_d32_68),.data_out(wire_d32_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303270(.data_in(wire_d32_69),.data_out(wire_d32_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303271(.data_in(wire_d32_70),.data_out(wire_d32_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303272(.data_in(wire_d32_71),.data_out(wire_d32_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303273(.data_in(wire_d32_72),.data_out(wire_d32_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3303274(.data_in(wire_d32_73),.data_out(wire_d32_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303275(.data_in(wire_d32_74),.data_out(wire_d32_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303276(.data_in(wire_d32_75),.data_out(wire_d32_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303277(.data_in(wire_d32_76),.data_out(wire_d32_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303278(.data_in(wire_d32_77),.data_out(wire_d32_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303279(.data_in(wire_d32_78),.data_out(d_out32),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance340330(.data_in(d_in33),.data_out(wire_d33_0),.clk(clk),.rst(rst));            //channel 34
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance340331(.data_in(wire_d33_0),.data_out(wire_d33_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance340332(.data_in(wire_d33_1),.data_out(wire_d33_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance340333(.data_in(wire_d33_2),.data_out(wire_d33_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance340334(.data_in(wire_d33_3),.data_out(wire_d33_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance340335(.data_in(wire_d33_4),.data_out(wire_d33_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance340336(.data_in(wire_d33_5),.data_out(wire_d33_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance340337(.data_in(wire_d33_6),.data_out(wire_d33_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance340338(.data_in(wire_d33_7),.data_out(wire_d33_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance340339(.data_in(wire_d33_8),.data_out(wire_d33_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3403310(.data_in(wire_d33_9),.data_out(wire_d33_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3403311(.data_in(wire_d33_10),.data_out(wire_d33_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403312(.data_in(wire_d33_11),.data_out(wire_d33_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403313(.data_in(wire_d33_12),.data_out(wire_d33_13),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403314(.data_in(wire_d33_13),.data_out(wire_d33_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403315(.data_in(wire_d33_14),.data_out(wire_d33_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3403316(.data_in(wire_d33_15),.data_out(wire_d33_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3403317(.data_in(wire_d33_16),.data_out(wire_d33_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3403318(.data_in(wire_d33_17),.data_out(wire_d33_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3403319(.data_in(wire_d33_18),.data_out(wire_d33_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3403320(.data_in(wire_d33_19),.data_out(wire_d33_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3403321(.data_in(wire_d33_20),.data_out(wire_d33_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3403322(.data_in(wire_d33_21),.data_out(wire_d33_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3403323(.data_in(wire_d33_22),.data_out(wire_d33_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3403324(.data_in(wire_d33_23),.data_out(wire_d33_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3403325(.data_in(wire_d33_24),.data_out(wire_d33_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403326(.data_in(wire_d33_25),.data_out(wire_d33_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3403327(.data_in(wire_d33_26),.data_out(wire_d33_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3403328(.data_in(wire_d33_27),.data_out(wire_d33_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403329(.data_in(wire_d33_28),.data_out(wire_d33_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403330(.data_in(wire_d33_29),.data_out(wire_d33_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403331(.data_in(wire_d33_30),.data_out(wire_d33_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403332(.data_in(wire_d33_31),.data_out(wire_d33_32),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403333(.data_in(wire_d33_32),.data_out(wire_d33_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403334(.data_in(wire_d33_33),.data_out(wire_d33_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3403335(.data_in(wire_d33_34),.data_out(wire_d33_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3403336(.data_in(wire_d33_35),.data_out(wire_d33_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403337(.data_in(wire_d33_36),.data_out(wire_d33_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403338(.data_in(wire_d33_37),.data_out(wire_d33_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403339(.data_in(wire_d33_38),.data_out(wire_d33_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403340(.data_in(wire_d33_39),.data_out(wire_d33_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3403341(.data_in(wire_d33_40),.data_out(wire_d33_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3403342(.data_in(wire_d33_41),.data_out(wire_d33_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403343(.data_in(wire_d33_42),.data_out(wire_d33_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403344(.data_in(wire_d33_43),.data_out(wire_d33_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403345(.data_in(wire_d33_44),.data_out(wire_d33_45),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403346(.data_in(wire_d33_45),.data_out(wire_d33_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403347(.data_in(wire_d33_46),.data_out(wire_d33_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3403348(.data_in(wire_d33_47),.data_out(wire_d33_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3403349(.data_in(wire_d33_48),.data_out(wire_d33_49),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403350(.data_in(wire_d33_49),.data_out(wire_d33_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3403351(.data_in(wire_d33_50),.data_out(wire_d33_51),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403352(.data_in(wire_d33_51),.data_out(wire_d33_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403353(.data_in(wire_d33_52),.data_out(wire_d33_53),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403354(.data_in(wire_d33_53),.data_out(wire_d33_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3403355(.data_in(wire_d33_54),.data_out(wire_d33_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3403356(.data_in(wire_d33_55),.data_out(wire_d33_56),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403357(.data_in(wire_d33_56),.data_out(wire_d33_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403358(.data_in(wire_d33_57),.data_out(wire_d33_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3403359(.data_in(wire_d33_58),.data_out(wire_d33_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403360(.data_in(wire_d33_59),.data_out(wire_d33_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403361(.data_in(wire_d33_60),.data_out(wire_d33_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403362(.data_in(wire_d33_61),.data_out(wire_d33_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403363(.data_in(wire_d33_62),.data_out(wire_d33_63),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403364(.data_in(wire_d33_63),.data_out(wire_d33_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403365(.data_in(wire_d33_64),.data_out(wire_d33_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403366(.data_in(wire_d33_65),.data_out(wire_d33_66),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3403367(.data_in(wire_d33_66),.data_out(wire_d33_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403368(.data_in(wire_d33_67),.data_out(wire_d33_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403369(.data_in(wire_d33_68),.data_out(wire_d33_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403370(.data_in(wire_d33_69),.data_out(wire_d33_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3403371(.data_in(wire_d33_70),.data_out(wire_d33_71),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403372(.data_in(wire_d33_71),.data_out(wire_d33_72),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403373(.data_in(wire_d33_72),.data_out(wire_d33_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3403374(.data_in(wire_d33_73),.data_out(wire_d33_74),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3403375(.data_in(wire_d33_74),.data_out(wire_d33_75),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403376(.data_in(wire_d33_75),.data_out(wire_d33_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3403377(.data_in(wire_d33_76),.data_out(wire_d33_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403378(.data_in(wire_d33_77),.data_out(wire_d33_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3403379(.data_in(wire_d33_78),.data_out(d_out33),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance350340(.data_in(d_in34),.data_out(wire_d34_0),.clk(clk),.rst(rst));            //channel 35
	large_mux #(.WIDTH(WIDTH)) large_mux_instance350341(.data_in(wire_d34_0),.data_out(wire_d34_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance350342(.data_in(wire_d34_1),.data_out(wire_d34_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance350343(.data_in(wire_d34_2),.data_out(wire_d34_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance350344(.data_in(wire_d34_3),.data_out(wire_d34_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance350345(.data_in(wire_d34_4),.data_out(wire_d34_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance350346(.data_in(wire_d34_5),.data_out(wire_d34_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance350347(.data_in(wire_d34_6),.data_out(wire_d34_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance350348(.data_in(wire_d34_7),.data_out(wire_d34_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance350349(.data_in(wire_d34_8),.data_out(wire_d34_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503410(.data_in(wire_d34_9),.data_out(wire_d34_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503411(.data_in(wire_d34_10),.data_out(wire_d34_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503412(.data_in(wire_d34_11),.data_out(wire_d34_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503413(.data_in(wire_d34_12),.data_out(wire_d34_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503414(.data_in(wire_d34_13),.data_out(wire_d34_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503415(.data_in(wire_d34_14),.data_out(wire_d34_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503416(.data_in(wire_d34_15),.data_out(wire_d34_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503417(.data_in(wire_d34_16),.data_out(wire_d34_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503418(.data_in(wire_d34_17),.data_out(wire_d34_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503419(.data_in(wire_d34_18),.data_out(wire_d34_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503420(.data_in(wire_d34_19),.data_out(wire_d34_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503421(.data_in(wire_d34_20),.data_out(wire_d34_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503422(.data_in(wire_d34_21),.data_out(wire_d34_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503423(.data_in(wire_d34_22),.data_out(wire_d34_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503424(.data_in(wire_d34_23),.data_out(wire_d34_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503425(.data_in(wire_d34_24),.data_out(wire_d34_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503426(.data_in(wire_d34_25),.data_out(wire_d34_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503427(.data_in(wire_d34_26),.data_out(wire_d34_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503428(.data_in(wire_d34_27),.data_out(wire_d34_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503429(.data_in(wire_d34_28),.data_out(wire_d34_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3503430(.data_in(wire_d34_29),.data_out(wire_d34_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503431(.data_in(wire_d34_30),.data_out(wire_d34_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503432(.data_in(wire_d34_31),.data_out(wire_d34_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503433(.data_in(wire_d34_32),.data_out(wire_d34_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503434(.data_in(wire_d34_33),.data_out(wire_d34_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503435(.data_in(wire_d34_34),.data_out(wire_d34_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503436(.data_in(wire_d34_35),.data_out(wire_d34_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503437(.data_in(wire_d34_36),.data_out(wire_d34_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3503438(.data_in(wire_d34_37),.data_out(wire_d34_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503439(.data_in(wire_d34_38),.data_out(wire_d34_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503440(.data_in(wire_d34_39),.data_out(wire_d34_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503441(.data_in(wire_d34_40),.data_out(wire_d34_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503442(.data_in(wire_d34_41),.data_out(wire_d34_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3503443(.data_in(wire_d34_42),.data_out(wire_d34_43),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503444(.data_in(wire_d34_43),.data_out(wire_d34_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503445(.data_in(wire_d34_44),.data_out(wire_d34_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503446(.data_in(wire_d34_45),.data_out(wire_d34_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503447(.data_in(wire_d34_46),.data_out(wire_d34_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503448(.data_in(wire_d34_47),.data_out(wire_d34_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503449(.data_in(wire_d34_48),.data_out(wire_d34_49),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503450(.data_in(wire_d34_49),.data_out(wire_d34_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503451(.data_in(wire_d34_50),.data_out(wire_d34_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3503452(.data_in(wire_d34_51),.data_out(wire_d34_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3503453(.data_in(wire_d34_52),.data_out(wire_d34_53),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503454(.data_in(wire_d34_53),.data_out(wire_d34_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503455(.data_in(wire_d34_54),.data_out(wire_d34_55),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503456(.data_in(wire_d34_55),.data_out(wire_d34_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503457(.data_in(wire_d34_56),.data_out(wire_d34_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503458(.data_in(wire_d34_57),.data_out(wire_d34_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503459(.data_in(wire_d34_58),.data_out(wire_d34_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503460(.data_in(wire_d34_59),.data_out(wire_d34_60),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503461(.data_in(wire_d34_60),.data_out(wire_d34_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503462(.data_in(wire_d34_61),.data_out(wire_d34_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503463(.data_in(wire_d34_62),.data_out(wire_d34_63),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503464(.data_in(wire_d34_63),.data_out(wire_d34_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503465(.data_in(wire_d34_64),.data_out(wire_d34_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3503466(.data_in(wire_d34_65),.data_out(wire_d34_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503467(.data_in(wire_d34_66),.data_out(wire_d34_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3503468(.data_in(wire_d34_67),.data_out(wire_d34_68),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503469(.data_in(wire_d34_68),.data_out(wire_d34_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503470(.data_in(wire_d34_69),.data_out(wire_d34_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503471(.data_in(wire_d34_70),.data_out(wire_d34_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503472(.data_in(wire_d34_71),.data_out(wire_d34_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503473(.data_in(wire_d34_72),.data_out(wire_d34_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503474(.data_in(wire_d34_73),.data_out(wire_d34_74),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503475(.data_in(wire_d34_74),.data_out(wire_d34_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503476(.data_in(wire_d34_75),.data_out(wire_d34_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503477(.data_in(wire_d34_76),.data_out(wire_d34_77),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503478(.data_in(wire_d34_77),.data_out(wire_d34_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503479(.data_in(wire_d34_78),.data_out(d_out34),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance360350(.data_in(d_in35),.data_out(wire_d35_0),.clk(clk),.rst(rst));            //channel 36
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance360351(.data_in(wire_d35_0),.data_out(wire_d35_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance360352(.data_in(wire_d35_1),.data_out(wire_d35_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance360353(.data_in(wire_d35_2),.data_out(wire_d35_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance360354(.data_in(wire_d35_3),.data_out(wire_d35_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance360355(.data_in(wire_d35_4),.data_out(wire_d35_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance360356(.data_in(wire_d35_5),.data_out(wire_d35_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance360357(.data_in(wire_d35_6),.data_out(wire_d35_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance360358(.data_in(wire_d35_7),.data_out(wire_d35_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance360359(.data_in(wire_d35_8),.data_out(wire_d35_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603510(.data_in(wire_d35_9),.data_out(wire_d35_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603511(.data_in(wire_d35_10),.data_out(wire_d35_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603512(.data_in(wire_d35_11),.data_out(wire_d35_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603513(.data_in(wire_d35_12),.data_out(wire_d35_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603514(.data_in(wire_d35_13),.data_out(wire_d35_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603515(.data_in(wire_d35_14),.data_out(wire_d35_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603516(.data_in(wire_d35_15),.data_out(wire_d35_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603517(.data_in(wire_d35_16),.data_out(wire_d35_17),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603518(.data_in(wire_d35_17),.data_out(wire_d35_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603519(.data_in(wire_d35_18),.data_out(wire_d35_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603520(.data_in(wire_d35_19),.data_out(wire_d35_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603521(.data_in(wire_d35_20),.data_out(wire_d35_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603522(.data_in(wire_d35_21),.data_out(wire_d35_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603523(.data_in(wire_d35_22),.data_out(wire_d35_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603524(.data_in(wire_d35_23),.data_out(wire_d35_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603525(.data_in(wire_d35_24),.data_out(wire_d35_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603526(.data_in(wire_d35_25),.data_out(wire_d35_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603527(.data_in(wire_d35_26),.data_out(wire_d35_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603528(.data_in(wire_d35_27),.data_out(wire_d35_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603529(.data_in(wire_d35_28),.data_out(wire_d35_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603530(.data_in(wire_d35_29),.data_out(wire_d35_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603531(.data_in(wire_d35_30),.data_out(wire_d35_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603532(.data_in(wire_d35_31),.data_out(wire_d35_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603533(.data_in(wire_d35_32),.data_out(wire_d35_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603534(.data_in(wire_d35_33),.data_out(wire_d35_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603535(.data_in(wire_d35_34),.data_out(wire_d35_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603536(.data_in(wire_d35_35),.data_out(wire_d35_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603537(.data_in(wire_d35_36),.data_out(wire_d35_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603538(.data_in(wire_d35_37),.data_out(wire_d35_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603539(.data_in(wire_d35_38),.data_out(wire_d35_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603540(.data_in(wire_d35_39),.data_out(wire_d35_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603541(.data_in(wire_d35_40),.data_out(wire_d35_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603542(.data_in(wire_d35_41),.data_out(wire_d35_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603543(.data_in(wire_d35_42),.data_out(wire_d35_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603544(.data_in(wire_d35_43),.data_out(wire_d35_44),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603545(.data_in(wire_d35_44),.data_out(wire_d35_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603546(.data_in(wire_d35_45),.data_out(wire_d35_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603547(.data_in(wire_d35_46),.data_out(wire_d35_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603548(.data_in(wire_d35_47),.data_out(wire_d35_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603549(.data_in(wire_d35_48),.data_out(wire_d35_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603550(.data_in(wire_d35_49),.data_out(wire_d35_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603551(.data_in(wire_d35_50),.data_out(wire_d35_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603552(.data_in(wire_d35_51),.data_out(wire_d35_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603553(.data_in(wire_d35_52),.data_out(wire_d35_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603554(.data_in(wire_d35_53),.data_out(wire_d35_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603555(.data_in(wire_d35_54),.data_out(wire_d35_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603556(.data_in(wire_d35_55),.data_out(wire_d35_56),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603557(.data_in(wire_d35_56),.data_out(wire_d35_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603558(.data_in(wire_d35_57),.data_out(wire_d35_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603559(.data_in(wire_d35_58),.data_out(wire_d35_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603560(.data_in(wire_d35_59),.data_out(wire_d35_60),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603561(.data_in(wire_d35_60),.data_out(wire_d35_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603562(.data_in(wire_d35_61),.data_out(wire_d35_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603563(.data_in(wire_d35_62),.data_out(wire_d35_63),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603564(.data_in(wire_d35_63),.data_out(wire_d35_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603565(.data_in(wire_d35_64),.data_out(wire_d35_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603566(.data_in(wire_d35_65),.data_out(wire_d35_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603567(.data_in(wire_d35_66),.data_out(wire_d35_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603568(.data_in(wire_d35_67),.data_out(wire_d35_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603569(.data_in(wire_d35_68),.data_out(wire_d35_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603570(.data_in(wire_d35_69),.data_out(wire_d35_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603571(.data_in(wire_d35_70),.data_out(wire_d35_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603572(.data_in(wire_d35_71),.data_out(wire_d35_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603573(.data_in(wire_d35_72),.data_out(wire_d35_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603574(.data_in(wire_d35_73),.data_out(wire_d35_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603575(.data_in(wire_d35_74),.data_out(wire_d35_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603576(.data_in(wire_d35_75),.data_out(wire_d35_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603577(.data_in(wire_d35_76),.data_out(wire_d35_77),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603578(.data_in(wire_d35_77),.data_out(wire_d35_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603579(.data_in(wire_d35_78),.data_out(d_out35),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance370360(.data_in(d_in36),.data_out(wire_d36_0),.clk(clk),.rst(rst));            //channel 37
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance370361(.data_in(wire_d36_0),.data_out(wire_d36_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance370362(.data_in(wire_d36_1),.data_out(wire_d36_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance370363(.data_in(wire_d36_2),.data_out(wire_d36_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance370364(.data_in(wire_d36_3),.data_out(wire_d36_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance370365(.data_in(wire_d36_4),.data_out(wire_d36_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance370366(.data_in(wire_d36_5),.data_out(wire_d36_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance370367(.data_in(wire_d36_6),.data_out(wire_d36_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance370368(.data_in(wire_d36_7),.data_out(wire_d36_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance370369(.data_in(wire_d36_8),.data_out(wire_d36_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703610(.data_in(wire_d36_9),.data_out(wire_d36_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703611(.data_in(wire_d36_10),.data_out(wire_d36_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703612(.data_in(wire_d36_11),.data_out(wire_d36_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703613(.data_in(wire_d36_12),.data_out(wire_d36_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703614(.data_in(wire_d36_13),.data_out(wire_d36_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3703615(.data_in(wire_d36_14),.data_out(wire_d36_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703616(.data_in(wire_d36_15),.data_out(wire_d36_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703617(.data_in(wire_d36_16),.data_out(wire_d36_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703618(.data_in(wire_d36_17),.data_out(wire_d36_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703619(.data_in(wire_d36_18),.data_out(wire_d36_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3703620(.data_in(wire_d36_19),.data_out(wire_d36_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703621(.data_in(wire_d36_20),.data_out(wire_d36_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703622(.data_in(wire_d36_21),.data_out(wire_d36_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703623(.data_in(wire_d36_22),.data_out(wire_d36_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703624(.data_in(wire_d36_23),.data_out(wire_d36_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3703625(.data_in(wire_d36_24),.data_out(wire_d36_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3703626(.data_in(wire_d36_25),.data_out(wire_d36_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703627(.data_in(wire_d36_26),.data_out(wire_d36_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703628(.data_in(wire_d36_27),.data_out(wire_d36_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3703629(.data_in(wire_d36_28),.data_out(wire_d36_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703630(.data_in(wire_d36_29),.data_out(wire_d36_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703631(.data_in(wire_d36_30),.data_out(wire_d36_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3703632(.data_in(wire_d36_31),.data_out(wire_d36_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703633(.data_in(wire_d36_32),.data_out(wire_d36_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703634(.data_in(wire_d36_33),.data_out(wire_d36_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703635(.data_in(wire_d36_34),.data_out(wire_d36_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3703636(.data_in(wire_d36_35),.data_out(wire_d36_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703637(.data_in(wire_d36_36),.data_out(wire_d36_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703638(.data_in(wire_d36_37),.data_out(wire_d36_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3703639(.data_in(wire_d36_38),.data_out(wire_d36_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703640(.data_in(wire_d36_39),.data_out(wire_d36_40),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703641(.data_in(wire_d36_40),.data_out(wire_d36_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3703642(.data_in(wire_d36_41),.data_out(wire_d36_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703643(.data_in(wire_d36_42),.data_out(wire_d36_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703644(.data_in(wire_d36_43),.data_out(wire_d36_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3703645(.data_in(wire_d36_44),.data_out(wire_d36_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703646(.data_in(wire_d36_45),.data_out(wire_d36_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703647(.data_in(wire_d36_46),.data_out(wire_d36_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703648(.data_in(wire_d36_47),.data_out(wire_d36_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3703649(.data_in(wire_d36_48),.data_out(wire_d36_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3703650(.data_in(wire_d36_49),.data_out(wire_d36_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703651(.data_in(wire_d36_50),.data_out(wire_d36_51),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703652(.data_in(wire_d36_51),.data_out(wire_d36_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703653(.data_in(wire_d36_52),.data_out(wire_d36_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703654(.data_in(wire_d36_53),.data_out(wire_d36_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703655(.data_in(wire_d36_54),.data_out(wire_d36_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703656(.data_in(wire_d36_55),.data_out(wire_d36_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703657(.data_in(wire_d36_56),.data_out(wire_d36_57),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3703658(.data_in(wire_d36_57),.data_out(wire_d36_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3703659(.data_in(wire_d36_58),.data_out(wire_d36_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3703660(.data_in(wire_d36_59),.data_out(wire_d36_60),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703661(.data_in(wire_d36_60),.data_out(wire_d36_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703662(.data_in(wire_d36_61),.data_out(wire_d36_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703663(.data_in(wire_d36_62),.data_out(wire_d36_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3703664(.data_in(wire_d36_63),.data_out(wire_d36_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703665(.data_in(wire_d36_64),.data_out(wire_d36_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703666(.data_in(wire_d36_65),.data_out(wire_d36_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3703667(.data_in(wire_d36_66),.data_out(wire_d36_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703668(.data_in(wire_d36_67),.data_out(wire_d36_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703669(.data_in(wire_d36_68),.data_out(wire_d36_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703670(.data_in(wire_d36_69),.data_out(wire_d36_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3703671(.data_in(wire_d36_70),.data_out(wire_d36_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3703672(.data_in(wire_d36_71),.data_out(wire_d36_72),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703673(.data_in(wire_d36_72),.data_out(wire_d36_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703674(.data_in(wire_d36_73),.data_out(wire_d36_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703675(.data_in(wire_d36_74),.data_out(wire_d36_75),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703676(.data_in(wire_d36_75),.data_out(wire_d36_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3703677(.data_in(wire_d36_76),.data_out(wire_d36_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3703678(.data_in(wire_d36_77),.data_out(wire_d36_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703679(.data_in(wire_d36_78),.data_out(d_out36),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance380370(.data_in(d_in37),.data_out(wire_d37_0),.clk(clk),.rst(rst));            //channel 38
	register #(.WIDTH(WIDTH)) register_instance380371(.data_in(wire_d37_0),.data_out(wire_d37_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance380372(.data_in(wire_d37_1),.data_out(wire_d37_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance380373(.data_in(wire_d37_2),.data_out(wire_d37_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance380374(.data_in(wire_d37_3),.data_out(wire_d37_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance380375(.data_in(wire_d37_4),.data_out(wire_d37_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance380376(.data_in(wire_d37_5),.data_out(wire_d37_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance380377(.data_in(wire_d37_6),.data_out(wire_d37_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance380378(.data_in(wire_d37_7),.data_out(wire_d37_8),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance380379(.data_in(wire_d37_8),.data_out(wire_d37_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803710(.data_in(wire_d37_9),.data_out(wire_d37_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803711(.data_in(wire_d37_10),.data_out(wire_d37_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803712(.data_in(wire_d37_11),.data_out(wire_d37_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3803713(.data_in(wire_d37_12),.data_out(wire_d37_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803714(.data_in(wire_d37_13),.data_out(wire_d37_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803715(.data_in(wire_d37_14),.data_out(wire_d37_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3803716(.data_in(wire_d37_15),.data_out(wire_d37_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803717(.data_in(wire_d37_16),.data_out(wire_d37_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803718(.data_in(wire_d37_17),.data_out(wire_d37_18),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803719(.data_in(wire_d37_18),.data_out(wire_d37_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803720(.data_in(wire_d37_19),.data_out(wire_d37_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3803721(.data_in(wire_d37_20),.data_out(wire_d37_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803722(.data_in(wire_d37_21),.data_out(wire_d37_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803723(.data_in(wire_d37_22),.data_out(wire_d37_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803724(.data_in(wire_d37_23),.data_out(wire_d37_24),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803725(.data_in(wire_d37_24),.data_out(wire_d37_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803726(.data_in(wire_d37_25),.data_out(wire_d37_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803727(.data_in(wire_d37_26),.data_out(wire_d37_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803728(.data_in(wire_d37_27),.data_out(wire_d37_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803729(.data_in(wire_d37_28),.data_out(wire_d37_29),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803730(.data_in(wire_d37_29),.data_out(wire_d37_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803731(.data_in(wire_d37_30),.data_out(wire_d37_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803732(.data_in(wire_d37_31),.data_out(wire_d37_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803733(.data_in(wire_d37_32),.data_out(wire_d37_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803734(.data_in(wire_d37_33),.data_out(wire_d37_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803735(.data_in(wire_d37_34),.data_out(wire_d37_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803736(.data_in(wire_d37_35),.data_out(wire_d37_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803737(.data_in(wire_d37_36),.data_out(wire_d37_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803738(.data_in(wire_d37_37),.data_out(wire_d37_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803739(.data_in(wire_d37_38),.data_out(wire_d37_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803740(.data_in(wire_d37_39),.data_out(wire_d37_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3803741(.data_in(wire_d37_40),.data_out(wire_d37_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803742(.data_in(wire_d37_41),.data_out(wire_d37_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803743(.data_in(wire_d37_42),.data_out(wire_d37_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803744(.data_in(wire_d37_43),.data_out(wire_d37_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803745(.data_in(wire_d37_44),.data_out(wire_d37_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803746(.data_in(wire_d37_45),.data_out(wire_d37_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803747(.data_in(wire_d37_46),.data_out(wire_d37_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803748(.data_in(wire_d37_47),.data_out(wire_d37_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803749(.data_in(wire_d37_48),.data_out(wire_d37_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3803750(.data_in(wire_d37_49),.data_out(wire_d37_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803751(.data_in(wire_d37_50),.data_out(wire_d37_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803752(.data_in(wire_d37_51),.data_out(wire_d37_52),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803753(.data_in(wire_d37_52),.data_out(wire_d37_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803754(.data_in(wire_d37_53),.data_out(wire_d37_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803755(.data_in(wire_d37_54),.data_out(wire_d37_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803756(.data_in(wire_d37_55),.data_out(wire_d37_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803757(.data_in(wire_d37_56),.data_out(wire_d37_57),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803758(.data_in(wire_d37_57),.data_out(wire_d37_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803759(.data_in(wire_d37_58),.data_out(wire_d37_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3803760(.data_in(wire_d37_59),.data_out(wire_d37_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803761(.data_in(wire_d37_60),.data_out(wire_d37_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803762(.data_in(wire_d37_61),.data_out(wire_d37_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803763(.data_in(wire_d37_62),.data_out(wire_d37_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3803764(.data_in(wire_d37_63),.data_out(wire_d37_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803765(.data_in(wire_d37_64),.data_out(wire_d37_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803766(.data_in(wire_d37_65),.data_out(wire_d37_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803767(.data_in(wire_d37_66),.data_out(wire_d37_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803768(.data_in(wire_d37_67),.data_out(wire_d37_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803769(.data_in(wire_d37_68),.data_out(wire_d37_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803770(.data_in(wire_d37_69),.data_out(wire_d37_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803771(.data_in(wire_d37_70),.data_out(wire_d37_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803772(.data_in(wire_d37_71),.data_out(wire_d37_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803773(.data_in(wire_d37_72),.data_out(wire_d37_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803774(.data_in(wire_d37_73),.data_out(wire_d37_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803775(.data_in(wire_d37_74),.data_out(wire_d37_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803776(.data_in(wire_d37_75),.data_out(wire_d37_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803777(.data_in(wire_d37_76),.data_out(wire_d37_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803778(.data_in(wire_d37_77),.data_out(wire_d37_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803779(.data_in(wire_d37_78),.data_out(d_out37),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance390380(.data_in(d_in38),.data_out(wire_d38_0),.clk(clk),.rst(rst));            //channel 39
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance390381(.data_in(wire_d38_0),.data_out(wire_d38_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance390382(.data_in(wire_d38_1),.data_out(wire_d38_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance390383(.data_in(wire_d38_2),.data_out(wire_d38_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance390384(.data_in(wire_d38_3),.data_out(wire_d38_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance390385(.data_in(wire_d38_4),.data_out(wire_d38_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance390386(.data_in(wire_d38_5),.data_out(wire_d38_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance390387(.data_in(wire_d38_6),.data_out(wire_d38_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance390388(.data_in(wire_d38_7),.data_out(wire_d38_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance390389(.data_in(wire_d38_8),.data_out(wire_d38_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903810(.data_in(wire_d38_9),.data_out(wire_d38_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903811(.data_in(wire_d38_10),.data_out(wire_d38_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903812(.data_in(wire_d38_11),.data_out(wire_d38_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903813(.data_in(wire_d38_12),.data_out(wire_d38_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3903814(.data_in(wire_d38_13),.data_out(wire_d38_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903815(.data_in(wire_d38_14),.data_out(wire_d38_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903816(.data_in(wire_d38_15),.data_out(wire_d38_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903817(.data_in(wire_d38_16),.data_out(wire_d38_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903818(.data_in(wire_d38_17),.data_out(wire_d38_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903819(.data_in(wire_d38_18),.data_out(wire_d38_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903820(.data_in(wire_d38_19),.data_out(wire_d38_20),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903821(.data_in(wire_d38_20),.data_out(wire_d38_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903822(.data_in(wire_d38_21),.data_out(wire_d38_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903823(.data_in(wire_d38_22),.data_out(wire_d38_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903824(.data_in(wire_d38_23),.data_out(wire_d38_24),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903825(.data_in(wire_d38_24),.data_out(wire_d38_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3903826(.data_in(wire_d38_25),.data_out(wire_d38_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3903827(.data_in(wire_d38_26),.data_out(wire_d38_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903828(.data_in(wire_d38_27),.data_out(wire_d38_28),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903829(.data_in(wire_d38_28),.data_out(wire_d38_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903830(.data_in(wire_d38_29),.data_out(wire_d38_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903831(.data_in(wire_d38_30),.data_out(wire_d38_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3903832(.data_in(wire_d38_31),.data_out(wire_d38_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903833(.data_in(wire_d38_32),.data_out(wire_d38_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3903834(.data_in(wire_d38_33),.data_out(wire_d38_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3903835(.data_in(wire_d38_34),.data_out(wire_d38_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3903836(.data_in(wire_d38_35),.data_out(wire_d38_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903837(.data_in(wire_d38_36),.data_out(wire_d38_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903838(.data_in(wire_d38_37),.data_out(wire_d38_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903839(.data_in(wire_d38_38),.data_out(wire_d38_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903840(.data_in(wire_d38_39),.data_out(wire_d38_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3903841(.data_in(wire_d38_40),.data_out(wire_d38_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903842(.data_in(wire_d38_41),.data_out(wire_d38_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903843(.data_in(wire_d38_42),.data_out(wire_d38_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3903844(.data_in(wire_d38_43),.data_out(wire_d38_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903845(.data_in(wire_d38_44),.data_out(wire_d38_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903846(.data_in(wire_d38_45),.data_out(wire_d38_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3903847(.data_in(wire_d38_46),.data_out(wire_d38_47),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903848(.data_in(wire_d38_47),.data_out(wire_d38_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903849(.data_in(wire_d38_48),.data_out(wire_d38_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903850(.data_in(wire_d38_49),.data_out(wire_d38_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3903851(.data_in(wire_d38_50),.data_out(wire_d38_51),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903852(.data_in(wire_d38_51),.data_out(wire_d38_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3903853(.data_in(wire_d38_52),.data_out(wire_d38_53),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903854(.data_in(wire_d38_53),.data_out(wire_d38_54),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3903855(.data_in(wire_d38_54),.data_out(wire_d38_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903856(.data_in(wire_d38_55),.data_out(wire_d38_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903857(.data_in(wire_d38_56),.data_out(wire_d38_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903858(.data_in(wire_d38_57),.data_out(wire_d38_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903859(.data_in(wire_d38_58),.data_out(wire_d38_59),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3903860(.data_in(wire_d38_59),.data_out(wire_d38_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903861(.data_in(wire_d38_60),.data_out(wire_d38_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903862(.data_in(wire_d38_61),.data_out(wire_d38_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903863(.data_in(wire_d38_62),.data_out(wire_d38_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903864(.data_in(wire_d38_63),.data_out(wire_d38_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903865(.data_in(wire_d38_64),.data_out(wire_d38_65),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903866(.data_in(wire_d38_65),.data_out(wire_d38_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903867(.data_in(wire_d38_66),.data_out(wire_d38_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903868(.data_in(wire_d38_67),.data_out(wire_d38_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903869(.data_in(wire_d38_68),.data_out(wire_d38_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903870(.data_in(wire_d38_69),.data_out(wire_d38_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903871(.data_in(wire_d38_70),.data_out(wire_d38_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903872(.data_in(wire_d38_71),.data_out(wire_d38_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3903873(.data_in(wire_d38_72),.data_out(wire_d38_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903874(.data_in(wire_d38_73),.data_out(wire_d38_74),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903875(.data_in(wire_d38_74),.data_out(wire_d38_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903876(.data_in(wire_d38_75),.data_out(wire_d38_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3903877(.data_in(wire_d38_76),.data_out(wire_d38_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3903878(.data_in(wire_d38_77),.data_out(wire_d38_78),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903879(.data_in(wire_d38_78),.data_out(d_out38),.clk(clk),.rst(rst));

	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance400390(.data_in(d_in39),.data_out(wire_d39_0),.clk(clk),.rst(rst));            //channel 40
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance400391(.data_in(wire_d39_0),.data_out(wire_d39_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance400392(.data_in(wire_d39_1),.data_out(wire_d39_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance400393(.data_in(wire_d39_2),.data_out(wire_d39_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance400394(.data_in(wire_d39_3),.data_out(wire_d39_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance400395(.data_in(wire_d39_4),.data_out(wire_d39_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance400396(.data_in(wire_d39_5),.data_out(wire_d39_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance400397(.data_in(wire_d39_6),.data_out(wire_d39_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance400398(.data_in(wire_d39_7),.data_out(wire_d39_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance400399(.data_in(wire_d39_8),.data_out(wire_d39_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003910(.data_in(wire_d39_9),.data_out(wire_d39_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4003911(.data_in(wire_d39_10),.data_out(wire_d39_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003912(.data_in(wire_d39_11),.data_out(wire_d39_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003913(.data_in(wire_d39_12),.data_out(wire_d39_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003914(.data_in(wire_d39_13),.data_out(wire_d39_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4003915(.data_in(wire_d39_14),.data_out(wire_d39_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003916(.data_in(wire_d39_15),.data_out(wire_d39_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4003917(.data_in(wire_d39_16),.data_out(wire_d39_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003918(.data_in(wire_d39_17),.data_out(wire_d39_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003919(.data_in(wire_d39_18),.data_out(wire_d39_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003920(.data_in(wire_d39_19),.data_out(wire_d39_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4003921(.data_in(wire_d39_20),.data_out(wire_d39_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003922(.data_in(wire_d39_21),.data_out(wire_d39_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003923(.data_in(wire_d39_22),.data_out(wire_d39_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003924(.data_in(wire_d39_23),.data_out(wire_d39_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003925(.data_in(wire_d39_24),.data_out(wire_d39_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003926(.data_in(wire_d39_25),.data_out(wire_d39_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003927(.data_in(wire_d39_26),.data_out(wire_d39_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003928(.data_in(wire_d39_27),.data_out(wire_d39_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003929(.data_in(wire_d39_28),.data_out(wire_d39_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003930(.data_in(wire_d39_29),.data_out(wire_d39_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003931(.data_in(wire_d39_30),.data_out(wire_d39_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4003932(.data_in(wire_d39_31),.data_out(wire_d39_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003933(.data_in(wire_d39_32),.data_out(wire_d39_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003934(.data_in(wire_d39_33),.data_out(wire_d39_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003935(.data_in(wire_d39_34),.data_out(wire_d39_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003936(.data_in(wire_d39_35),.data_out(wire_d39_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003937(.data_in(wire_d39_36),.data_out(wire_d39_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003938(.data_in(wire_d39_37),.data_out(wire_d39_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003939(.data_in(wire_d39_38),.data_out(wire_d39_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003940(.data_in(wire_d39_39),.data_out(wire_d39_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003941(.data_in(wire_d39_40),.data_out(wire_d39_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4003942(.data_in(wire_d39_41),.data_out(wire_d39_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4003943(.data_in(wire_d39_42),.data_out(wire_d39_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003944(.data_in(wire_d39_43),.data_out(wire_d39_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003945(.data_in(wire_d39_44),.data_out(wire_d39_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4003946(.data_in(wire_d39_45),.data_out(wire_d39_46),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003947(.data_in(wire_d39_46),.data_out(wire_d39_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003948(.data_in(wire_d39_47),.data_out(wire_d39_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003949(.data_in(wire_d39_48),.data_out(wire_d39_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003950(.data_in(wire_d39_49),.data_out(wire_d39_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4003951(.data_in(wire_d39_50),.data_out(wire_d39_51),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003952(.data_in(wire_d39_51),.data_out(wire_d39_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003953(.data_in(wire_d39_52),.data_out(wire_d39_53),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003954(.data_in(wire_d39_53),.data_out(wire_d39_54),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003955(.data_in(wire_d39_54),.data_out(wire_d39_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4003956(.data_in(wire_d39_55),.data_out(wire_d39_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003957(.data_in(wire_d39_56),.data_out(wire_d39_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003958(.data_in(wire_d39_57),.data_out(wire_d39_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003959(.data_in(wire_d39_58),.data_out(wire_d39_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003960(.data_in(wire_d39_59),.data_out(wire_d39_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4003961(.data_in(wire_d39_60),.data_out(wire_d39_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003962(.data_in(wire_d39_61),.data_out(wire_d39_62),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003963(.data_in(wire_d39_62),.data_out(wire_d39_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003964(.data_in(wire_d39_63),.data_out(wire_d39_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4003965(.data_in(wire_d39_64),.data_out(wire_d39_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003966(.data_in(wire_d39_65),.data_out(wire_d39_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003967(.data_in(wire_d39_66),.data_out(wire_d39_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003968(.data_in(wire_d39_67),.data_out(wire_d39_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4003969(.data_in(wire_d39_68),.data_out(wire_d39_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003970(.data_in(wire_d39_69),.data_out(wire_d39_70),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4003971(.data_in(wire_d39_70),.data_out(wire_d39_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003972(.data_in(wire_d39_71),.data_out(wire_d39_72),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003973(.data_in(wire_d39_72),.data_out(wire_d39_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003974(.data_in(wire_d39_73),.data_out(wire_d39_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003975(.data_in(wire_d39_74),.data_out(wire_d39_75),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003976(.data_in(wire_d39_75),.data_out(wire_d39_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003977(.data_in(wire_d39_76),.data_out(wire_d39_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003978(.data_in(wire_d39_77),.data_out(wire_d39_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003979(.data_in(wire_d39_78),.data_out(d_out39),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance410400(.data_in(d_in40),.data_out(wire_d40_0),.clk(clk),.rst(rst));            //channel 41
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance410401(.data_in(wire_d40_0),.data_out(wire_d40_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance410402(.data_in(wire_d40_1),.data_out(wire_d40_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance410403(.data_in(wire_d40_2),.data_out(wire_d40_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance410404(.data_in(wire_d40_3),.data_out(wire_d40_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance410405(.data_in(wire_d40_4),.data_out(wire_d40_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance410406(.data_in(wire_d40_5),.data_out(wire_d40_6),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance410407(.data_in(wire_d40_6),.data_out(wire_d40_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance410408(.data_in(wire_d40_7),.data_out(wire_d40_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance410409(.data_in(wire_d40_8),.data_out(wire_d40_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104010(.data_in(wire_d40_9),.data_out(wire_d40_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4104011(.data_in(wire_d40_10),.data_out(wire_d40_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4104012(.data_in(wire_d40_11),.data_out(wire_d40_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4104013(.data_in(wire_d40_12),.data_out(wire_d40_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4104014(.data_in(wire_d40_13),.data_out(wire_d40_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4104015(.data_in(wire_d40_14),.data_out(wire_d40_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104016(.data_in(wire_d40_15),.data_out(wire_d40_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104017(.data_in(wire_d40_16),.data_out(wire_d40_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104018(.data_in(wire_d40_17),.data_out(wire_d40_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4104019(.data_in(wire_d40_18),.data_out(wire_d40_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104020(.data_in(wire_d40_19),.data_out(wire_d40_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104021(.data_in(wire_d40_20),.data_out(wire_d40_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104022(.data_in(wire_d40_21),.data_out(wire_d40_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4104023(.data_in(wire_d40_22),.data_out(wire_d40_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104024(.data_in(wire_d40_23),.data_out(wire_d40_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104025(.data_in(wire_d40_24),.data_out(wire_d40_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104026(.data_in(wire_d40_25),.data_out(wire_d40_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104027(.data_in(wire_d40_26),.data_out(wire_d40_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4104028(.data_in(wire_d40_27),.data_out(wire_d40_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4104029(.data_in(wire_d40_28),.data_out(wire_d40_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4104030(.data_in(wire_d40_29),.data_out(wire_d40_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104031(.data_in(wire_d40_30),.data_out(wire_d40_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104032(.data_in(wire_d40_31),.data_out(wire_d40_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104033(.data_in(wire_d40_32),.data_out(wire_d40_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4104034(.data_in(wire_d40_33),.data_out(wire_d40_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104035(.data_in(wire_d40_34),.data_out(wire_d40_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4104036(.data_in(wire_d40_35),.data_out(wire_d40_36),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104037(.data_in(wire_d40_36),.data_out(wire_d40_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104038(.data_in(wire_d40_37),.data_out(wire_d40_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104039(.data_in(wire_d40_38),.data_out(wire_d40_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104040(.data_in(wire_d40_39),.data_out(wire_d40_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4104041(.data_in(wire_d40_40),.data_out(wire_d40_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104042(.data_in(wire_d40_41),.data_out(wire_d40_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104043(.data_in(wire_d40_42),.data_out(wire_d40_43),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4104044(.data_in(wire_d40_43),.data_out(wire_d40_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104045(.data_in(wire_d40_44),.data_out(wire_d40_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104046(.data_in(wire_d40_45),.data_out(wire_d40_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4104047(.data_in(wire_d40_46),.data_out(wire_d40_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104048(.data_in(wire_d40_47),.data_out(wire_d40_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104049(.data_in(wire_d40_48),.data_out(wire_d40_49),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4104050(.data_in(wire_d40_49),.data_out(wire_d40_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104051(.data_in(wire_d40_50),.data_out(wire_d40_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104052(.data_in(wire_d40_51),.data_out(wire_d40_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104053(.data_in(wire_d40_52),.data_out(wire_d40_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104054(.data_in(wire_d40_53),.data_out(wire_d40_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104055(.data_in(wire_d40_54),.data_out(wire_d40_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104056(.data_in(wire_d40_55),.data_out(wire_d40_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104057(.data_in(wire_d40_56),.data_out(wire_d40_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104058(.data_in(wire_d40_57),.data_out(wire_d40_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104059(.data_in(wire_d40_58),.data_out(wire_d40_59),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104060(.data_in(wire_d40_59),.data_out(wire_d40_60),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4104061(.data_in(wire_d40_60),.data_out(wire_d40_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104062(.data_in(wire_d40_61),.data_out(wire_d40_62),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4104063(.data_in(wire_d40_62),.data_out(wire_d40_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104064(.data_in(wire_d40_63),.data_out(wire_d40_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104065(.data_in(wire_d40_64),.data_out(wire_d40_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104066(.data_in(wire_d40_65),.data_out(wire_d40_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4104067(.data_in(wire_d40_66),.data_out(wire_d40_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104068(.data_in(wire_d40_67),.data_out(wire_d40_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104069(.data_in(wire_d40_68),.data_out(wire_d40_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104070(.data_in(wire_d40_69),.data_out(wire_d40_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4104071(.data_in(wire_d40_70),.data_out(wire_d40_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104072(.data_in(wire_d40_71),.data_out(wire_d40_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104073(.data_in(wire_d40_72),.data_out(wire_d40_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104074(.data_in(wire_d40_73),.data_out(wire_d40_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104075(.data_in(wire_d40_74),.data_out(wire_d40_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104076(.data_in(wire_d40_75),.data_out(wire_d40_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104077(.data_in(wire_d40_76),.data_out(wire_d40_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104078(.data_in(wire_d40_77),.data_out(wire_d40_78),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104079(.data_in(wire_d40_78),.data_out(d_out40),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance420410(.data_in(d_in41),.data_out(wire_d41_0),.clk(clk),.rst(rst));            //channel 42
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance420411(.data_in(wire_d41_0),.data_out(wire_d41_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance420412(.data_in(wire_d41_1),.data_out(wire_d41_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance420413(.data_in(wire_d41_2),.data_out(wire_d41_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance420414(.data_in(wire_d41_3),.data_out(wire_d41_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance420415(.data_in(wire_d41_4),.data_out(wire_d41_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance420416(.data_in(wire_d41_5),.data_out(wire_d41_6),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance420417(.data_in(wire_d41_6),.data_out(wire_d41_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance420418(.data_in(wire_d41_7),.data_out(wire_d41_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance420419(.data_in(wire_d41_8),.data_out(wire_d41_9),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204110(.data_in(wire_d41_9),.data_out(wire_d41_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204111(.data_in(wire_d41_10),.data_out(wire_d41_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204112(.data_in(wire_d41_11),.data_out(wire_d41_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4204113(.data_in(wire_d41_12),.data_out(wire_d41_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204114(.data_in(wire_d41_13),.data_out(wire_d41_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4204115(.data_in(wire_d41_14),.data_out(wire_d41_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204116(.data_in(wire_d41_15),.data_out(wire_d41_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204117(.data_in(wire_d41_16),.data_out(wire_d41_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204118(.data_in(wire_d41_17),.data_out(wire_d41_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204119(.data_in(wire_d41_18),.data_out(wire_d41_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204120(.data_in(wire_d41_19),.data_out(wire_d41_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204121(.data_in(wire_d41_20),.data_out(wire_d41_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204122(.data_in(wire_d41_21),.data_out(wire_d41_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204123(.data_in(wire_d41_22),.data_out(wire_d41_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204124(.data_in(wire_d41_23),.data_out(wire_d41_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204125(.data_in(wire_d41_24),.data_out(wire_d41_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204126(.data_in(wire_d41_25),.data_out(wire_d41_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204127(.data_in(wire_d41_26),.data_out(wire_d41_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204128(.data_in(wire_d41_27),.data_out(wire_d41_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4204129(.data_in(wire_d41_28),.data_out(wire_d41_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204130(.data_in(wire_d41_29),.data_out(wire_d41_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204131(.data_in(wire_d41_30),.data_out(wire_d41_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204132(.data_in(wire_d41_31),.data_out(wire_d41_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4204133(.data_in(wire_d41_32),.data_out(wire_d41_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204134(.data_in(wire_d41_33),.data_out(wire_d41_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204135(.data_in(wire_d41_34),.data_out(wire_d41_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204136(.data_in(wire_d41_35),.data_out(wire_d41_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204137(.data_in(wire_d41_36),.data_out(wire_d41_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204138(.data_in(wire_d41_37),.data_out(wire_d41_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204139(.data_in(wire_d41_38),.data_out(wire_d41_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4204140(.data_in(wire_d41_39),.data_out(wire_d41_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204141(.data_in(wire_d41_40),.data_out(wire_d41_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4204142(.data_in(wire_d41_41),.data_out(wire_d41_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204143(.data_in(wire_d41_42),.data_out(wire_d41_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204144(.data_in(wire_d41_43),.data_out(wire_d41_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4204145(.data_in(wire_d41_44),.data_out(wire_d41_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204146(.data_in(wire_d41_45),.data_out(wire_d41_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204147(.data_in(wire_d41_46),.data_out(wire_d41_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204148(.data_in(wire_d41_47),.data_out(wire_d41_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204149(.data_in(wire_d41_48),.data_out(wire_d41_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204150(.data_in(wire_d41_49),.data_out(wire_d41_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204151(.data_in(wire_d41_50),.data_out(wire_d41_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204152(.data_in(wire_d41_51),.data_out(wire_d41_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4204153(.data_in(wire_d41_52),.data_out(wire_d41_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204154(.data_in(wire_d41_53),.data_out(wire_d41_54),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204155(.data_in(wire_d41_54),.data_out(wire_d41_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4204156(.data_in(wire_d41_55),.data_out(wire_d41_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204157(.data_in(wire_d41_56),.data_out(wire_d41_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204158(.data_in(wire_d41_57),.data_out(wire_d41_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204159(.data_in(wire_d41_58),.data_out(wire_d41_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204160(.data_in(wire_d41_59),.data_out(wire_d41_60),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204161(.data_in(wire_d41_60),.data_out(wire_d41_61),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204162(.data_in(wire_d41_61),.data_out(wire_d41_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204163(.data_in(wire_d41_62),.data_out(wire_d41_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4204164(.data_in(wire_d41_63),.data_out(wire_d41_64),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4204165(.data_in(wire_d41_64),.data_out(wire_d41_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204166(.data_in(wire_d41_65),.data_out(wire_d41_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4204167(.data_in(wire_d41_66),.data_out(wire_d41_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204168(.data_in(wire_d41_67),.data_out(wire_d41_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204169(.data_in(wire_d41_68),.data_out(wire_d41_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204170(.data_in(wire_d41_69),.data_out(wire_d41_70),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204171(.data_in(wire_d41_70),.data_out(wire_d41_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204172(.data_in(wire_d41_71),.data_out(wire_d41_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204173(.data_in(wire_d41_72),.data_out(wire_d41_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204174(.data_in(wire_d41_73),.data_out(wire_d41_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204175(.data_in(wire_d41_74),.data_out(wire_d41_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204176(.data_in(wire_d41_75),.data_out(wire_d41_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204177(.data_in(wire_d41_76),.data_out(wire_d41_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204178(.data_in(wire_d41_77),.data_out(wire_d41_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204179(.data_in(wire_d41_78),.data_out(d_out41),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance430420(.data_in(d_in42),.data_out(wire_d42_0),.clk(clk),.rst(rst));            //channel 43
	decoder_top #(.WIDTH(WIDTH)) decoder_instance430421(.data_in(wire_d42_0),.data_out(wire_d42_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance430422(.data_in(wire_d42_1),.data_out(wire_d42_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance430423(.data_in(wire_d42_2),.data_out(wire_d42_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance430424(.data_in(wire_d42_3),.data_out(wire_d42_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance430425(.data_in(wire_d42_4),.data_out(wire_d42_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance430426(.data_in(wire_d42_5),.data_out(wire_d42_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance430427(.data_in(wire_d42_6),.data_out(wire_d42_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance430428(.data_in(wire_d42_7),.data_out(wire_d42_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance430429(.data_in(wire_d42_8),.data_out(wire_d42_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304210(.data_in(wire_d42_9),.data_out(wire_d42_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4304211(.data_in(wire_d42_10),.data_out(wire_d42_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304212(.data_in(wire_d42_11),.data_out(wire_d42_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304213(.data_in(wire_d42_12),.data_out(wire_d42_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304214(.data_in(wire_d42_13),.data_out(wire_d42_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304215(.data_in(wire_d42_14),.data_out(wire_d42_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304216(.data_in(wire_d42_15),.data_out(wire_d42_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304217(.data_in(wire_d42_16),.data_out(wire_d42_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304218(.data_in(wire_d42_17),.data_out(wire_d42_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304219(.data_in(wire_d42_18),.data_out(wire_d42_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304220(.data_in(wire_d42_19),.data_out(wire_d42_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304221(.data_in(wire_d42_20),.data_out(wire_d42_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304222(.data_in(wire_d42_21),.data_out(wire_d42_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304223(.data_in(wire_d42_22),.data_out(wire_d42_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304224(.data_in(wire_d42_23),.data_out(wire_d42_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304225(.data_in(wire_d42_24),.data_out(wire_d42_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304226(.data_in(wire_d42_25),.data_out(wire_d42_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304227(.data_in(wire_d42_26),.data_out(wire_d42_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304228(.data_in(wire_d42_27),.data_out(wire_d42_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4304229(.data_in(wire_d42_28),.data_out(wire_d42_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304230(.data_in(wire_d42_29),.data_out(wire_d42_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304231(.data_in(wire_d42_30),.data_out(wire_d42_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304232(.data_in(wire_d42_31),.data_out(wire_d42_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304233(.data_in(wire_d42_32),.data_out(wire_d42_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304234(.data_in(wire_d42_33),.data_out(wire_d42_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304235(.data_in(wire_d42_34),.data_out(wire_d42_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304236(.data_in(wire_d42_35),.data_out(wire_d42_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304237(.data_in(wire_d42_36),.data_out(wire_d42_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304238(.data_in(wire_d42_37),.data_out(wire_d42_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304239(.data_in(wire_d42_38),.data_out(wire_d42_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304240(.data_in(wire_d42_39),.data_out(wire_d42_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4304241(.data_in(wire_d42_40),.data_out(wire_d42_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304242(.data_in(wire_d42_41),.data_out(wire_d42_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304243(.data_in(wire_d42_42),.data_out(wire_d42_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304244(.data_in(wire_d42_43),.data_out(wire_d42_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304245(.data_in(wire_d42_44),.data_out(wire_d42_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304246(.data_in(wire_d42_45),.data_out(wire_d42_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304247(.data_in(wire_d42_46),.data_out(wire_d42_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304248(.data_in(wire_d42_47),.data_out(wire_d42_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4304249(.data_in(wire_d42_48),.data_out(wire_d42_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304250(.data_in(wire_d42_49),.data_out(wire_d42_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304251(.data_in(wire_d42_50),.data_out(wire_d42_51),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304252(.data_in(wire_d42_51),.data_out(wire_d42_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304253(.data_in(wire_d42_52),.data_out(wire_d42_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304254(.data_in(wire_d42_53),.data_out(wire_d42_54),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304255(.data_in(wire_d42_54),.data_out(wire_d42_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304256(.data_in(wire_d42_55),.data_out(wire_d42_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304257(.data_in(wire_d42_56),.data_out(wire_d42_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304258(.data_in(wire_d42_57),.data_out(wire_d42_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304259(.data_in(wire_d42_58),.data_out(wire_d42_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304260(.data_in(wire_d42_59),.data_out(wire_d42_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4304261(.data_in(wire_d42_60),.data_out(wire_d42_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304262(.data_in(wire_d42_61),.data_out(wire_d42_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304263(.data_in(wire_d42_62),.data_out(wire_d42_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304264(.data_in(wire_d42_63),.data_out(wire_d42_64),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304265(.data_in(wire_d42_64),.data_out(wire_d42_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304266(.data_in(wire_d42_65),.data_out(wire_d42_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304267(.data_in(wire_d42_66),.data_out(wire_d42_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304268(.data_in(wire_d42_67),.data_out(wire_d42_68),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304269(.data_in(wire_d42_68),.data_out(wire_d42_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304270(.data_in(wire_d42_69),.data_out(wire_d42_70),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304271(.data_in(wire_d42_70),.data_out(wire_d42_71),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304272(.data_in(wire_d42_71),.data_out(wire_d42_72),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304273(.data_in(wire_d42_72),.data_out(wire_d42_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304274(.data_in(wire_d42_73),.data_out(wire_d42_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304275(.data_in(wire_d42_74),.data_out(wire_d42_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304276(.data_in(wire_d42_75),.data_out(wire_d42_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304277(.data_in(wire_d42_76),.data_out(wire_d42_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304278(.data_in(wire_d42_77),.data_out(wire_d42_78),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304279(.data_in(wire_d42_78),.data_out(d_out42),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance440430(.data_in(d_in43),.data_out(wire_d43_0),.clk(clk),.rst(rst));            //channel 44
	large_mux #(.WIDTH(WIDTH)) large_mux_instance440431(.data_in(wire_d43_0),.data_out(wire_d43_1),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance440432(.data_in(wire_d43_1),.data_out(wire_d43_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance440433(.data_in(wire_d43_2),.data_out(wire_d43_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance440434(.data_in(wire_d43_3),.data_out(wire_d43_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance440435(.data_in(wire_d43_4),.data_out(wire_d43_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance440436(.data_in(wire_d43_5),.data_out(wire_d43_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance440437(.data_in(wire_d43_6),.data_out(wire_d43_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance440438(.data_in(wire_d43_7),.data_out(wire_d43_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance440439(.data_in(wire_d43_8),.data_out(wire_d43_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404310(.data_in(wire_d43_9),.data_out(wire_d43_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4404311(.data_in(wire_d43_10),.data_out(wire_d43_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404312(.data_in(wire_d43_11),.data_out(wire_d43_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4404313(.data_in(wire_d43_12),.data_out(wire_d43_13),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404314(.data_in(wire_d43_13),.data_out(wire_d43_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404315(.data_in(wire_d43_14),.data_out(wire_d43_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4404316(.data_in(wire_d43_15),.data_out(wire_d43_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404317(.data_in(wire_d43_16),.data_out(wire_d43_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404318(.data_in(wire_d43_17),.data_out(wire_d43_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404319(.data_in(wire_d43_18),.data_out(wire_d43_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404320(.data_in(wire_d43_19),.data_out(wire_d43_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404321(.data_in(wire_d43_20),.data_out(wire_d43_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4404322(.data_in(wire_d43_21),.data_out(wire_d43_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4404323(.data_in(wire_d43_22),.data_out(wire_d43_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4404324(.data_in(wire_d43_23),.data_out(wire_d43_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404325(.data_in(wire_d43_24),.data_out(wire_d43_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404326(.data_in(wire_d43_25),.data_out(wire_d43_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4404327(.data_in(wire_d43_26),.data_out(wire_d43_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404328(.data_in(wire_d43_27),.data_out(wire_d43_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404329(.data_in(wire_d43_28),.data_out(wire_d43_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404330(.data_in(wire_d43_29),.data_out(wire_d43_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4404331(.data_in(wire_d43_30),.data_out(wire_d43_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404332(.data_in(wire_d43_31),.data_out(wire_d43_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404333(.data_in(wire_d43_32),.data_out(wire_d43_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404334(.data_in(wire_d43_33),.data_out(wire_d43_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404335(.data_in(wire_d43_34),.data_out(wire_d43_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404336(.data_in(wire_d43_35),.data_out(wire_d43_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404337(.data_in(wire_d43_36),.data_out(wire_d43_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404338(.data_in(wire_d43_37),.data_out(wire_d43_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404339(.data_in(wire_d43_38),.data_out(wire_d43_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4404340(.data_in(wire_d43_39),.data_out(wire_d43_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404341(.data_in(wire_d43_40),.data_out(wire_d43_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404342(.data_in(wire_d43_41),.data_out(wire_d43_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404343(.data_in(wire_d43_42),.data_out(wire_d43_43),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404344(.data_in(wire_d43_43),.data_out(wire_d43_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4404345(.data_in(wire_d43_44),.data_out(wire_d43_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404346(.data_in(wire_d43_45),.data_out(wire_d43_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404347(.data_in(wire_d43_46),.data_out(wire_d43_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404348(.data_in(wire_d43_47),.data_out(wire_d43_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4404349(.data_in(wire_d43_48),.data_out(wire_d43_49),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4404350(.data_in(wire_d43_49),.data_out(wire_d43_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404351(.data_in(wire_d43_50),.data_out(wire_d43_51),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404352(.data_in(wire_d43_51),.data_out(wire_d43_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4404353(.data_in(wire_d43_52),.data_out(wire_d43_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404354(.data_in(wire_d43_53),.data_out(wire_d43_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404355(.data_in(wire_d43_54),.data_out(wire_d43_55),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404356(.data_in(wire_d43_55),.data_out(wire_d43_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404357(.data_in(wire_d43_56),.data_out(wire_d43_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404358(.data_in(wire_d43_57),.data_out(wire_d43_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404359(.data_in(wire_d43_58),.data_out(wire_d43_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404360(.data_in(wire_d43_59),.data_out(wire_d43_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404361(.data_in(wire_d43_60),.data_out(wire_d43_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4404362(.data_in(wire_d43_61),.data_out(wire_d43_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404363(.data_in(wire_d43_62),.data_out(wire_d43_63),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404364(.data_in(wire_d43_63),.data_out(wire_d43_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404365(.data_in(wire_d43_64),.data_out(wire_d43_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404366(.data_in(wire_d43_65),.data_out(wire_d43_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404367(.data_in(wire_d43_66),.data_out(wire_d43_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404368(.data_in(wire_d43_67),.data_out(wire_d43_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404369(.data_in(wire_d43_68),.data_out(wire_d43_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404370(.data_in(wire_d43_69),.data_out(wire_d43_70),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404371(.data_in(wire_d43_70),.data_out(wire_d43_71),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404372(.data_in(wire_d43_71),.data_out(wire_d43_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404373(.data_in(wire_d43_72),.data_out(wire_d43_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404374(.data_in(wire_d43_73),.data_out(wire_d43_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404375(.data_in(wire_d43_74),.data_out(wire_d43_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404376(.data_in(wire_d43_75),.data_out(wire_d43_76),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404377(.data_in(wire_d43_76),.data_out(wire_d43_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404378(.data_in(wire_d43_77),.data_out(wire_d43_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404379(.data_in(wire_d43_78),.data_out(d_out43),.clk(clk),.rst(rst));

	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance450440(.data_in(d_in44),.data_out(wire_d44_0),.clk(clk),.rst(rst));            //channel 45
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance450441(.data_in(wire_d44_0),.data_out(wire_d44_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance450442(.data_in(wire_d44_1),.data_out(wire_d44_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance450443(.data_in(wire_d44_2),.data_out(wire_d44_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance450444(.data_in(wire_d44_3),.data_out(wire_d44_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance450445(.data_in(wire_d44_4),.data_out(wire_d44_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance450446(.data_in(wire_d44_5),.data_out(wire_d44_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance450447(.data_in(wire_d44_6),.data_out(wire_d44_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance450448(.data_in(wire_d44_7),.data_out(wire_d44_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance450449(.data_in(wire_d44_8),.data_out(wire_d44_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504410(.data_in(wire_d44_9),.data_out(wire_d44_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504411(.data_in(wire_d44_10),.data_out(wire_d44_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504412(.data_in(wire_d44_11),.data_out(wire_d44_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504413(.data_in(wire_d44_12),.data_out(wire_d44_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504414(.data_in(wire_d44_13),.data_out(wire_d44_14),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504415(.data_in(wire_d44_14),.data_out(wire_d44_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504416(.data_in(wire_d44_15),.data_out(wire_d44_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4504417(.data_in(wire_d44_16),.data_out(wire_d44_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504418(.data_in(wire_d44_17),.data_out(wire_d44_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504419(.data_in(wire_d44_18),.data_out(wire_d44_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504420(.data_in(wire_d44_19),.data_out(wire_d44_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504421(.data_in(wire_d44_20),.data_out(wire_d44_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4504422(.data_in(wire_d44_21),.data_out(wire_d44_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504423(.data_in(wire_d44_22),.data_out(wire_d44_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4504424(.data_in(wire_d44_23),.data_out(wire_d44_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504425(.data_in(wire_d44_24),.data_out(wire_d44_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504426(.data_in(wire_d44_25),.data_out(wire_d44_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4504427(.data_in(wire_d44_26),.data_out(wire_d44_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504428(.data_in(wire_d44_27),.data_out(wire_d44_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4504429(.data_in(wire_d44_28),.data_out(wire_d44_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4504430(.data_in(wire_d44_29),.data_out(wire_d44_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4504431(.data_in(wire_d44_30),.data_out(wire_d44_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4504432(.data_in(wire_d44_31),.data_out(wire_d44_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504433(.data_in(wire_d44_32),.data_out(wire_d44_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504434(.data_in(wire_d44_33),.data_out(wire_d44_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4504435(.data_in(wire_d44_34),.data_out(wire_d44_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504436(.data_in(wire_d44_35),.data_out(wire_d44_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504437(.data_in(wire_d44_36),.data_out(wire_d44_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504438(.data_in(wire_d44_37),.data_out(wire_d44_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504439(.data_in(wire_d44_38),.data_out(wire_d44_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504440(.data_in(wire_d44_39),.data_out(wire_d44_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504441(.data_in(wire_d44_40),.data_out(wire_d44_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4504442(.data_in(wire_d44_41),.data_out(wire_d44_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504443(.data_in(wire_d44_42),.data_out(wire_d44_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504444(.data_in(wire_d44_43),.data_out(wire_d44_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4504445(.data_in(wire_d44_44),.data_out(wire_d44_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504446(.data_in(wire_d44_45),.data_out(wire_d44_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504447(.data_in(wire_d44_46),.data_out(wire_d44_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4504448(.data_in(wire_d44_47),.data_out(wire_d44_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504449(.data_in(wire_d44_48),.data_out(wire_d44_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504450(.data_in(wire_d44_49),.data_out(wire_d44_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4504451(.data_in(wire_d44_50),.data_out(wire_d44_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4504452(.data_in(wire_d44_51),.data_out(wire_d44_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504453(.data_in(wire_d44_52),.data_out(wire_d44_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504454(.data_in(wire_d44_53),.data_out(wire_d44_54),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504455(.data_in(wire_d44_54),.data_out(wire_d44_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504456(.data_in(wire_d44_55),.data_out(wire_d44_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504457(.data_in(wire_d44_56),.data_out(wire_d44_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504458(.data_in(wire_d44_57),.data_out(wire_d44_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504459(.data_in(wire_d44_58),.data_out(wire_d44_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504460(.data_in(wire_d44_59),.data_out(wire_d44_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4504461(.data_in(wire_d44_60),.data_out(wire_d44_61),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504462(.data_in(wire_d44_61),.data_out(wire_d44_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4504463(.data_in(wire_d44_62),.data_out(wire_d44_63),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4504464(.data_in(wire_d44_63),.data_out(wire_d44_64),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504465(.data_in(wire_d44_64),.data_out(wire_d44_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504466(.data_in(wire_d44_65),.data_out(wire_d44_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4504467(.data_in(wire_d44_66),.data_out(wire_d44_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4504468(.data_in(wire_d44_67),.data_out(wire_d44_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504469(.data_in(wire_d44_68),.data_out(wire_d44_69),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504470(.data_in(wire_d44_69),.data_out(wire_d44_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504471(.data_in(wire_d44_70),.data_out(wire_d44_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504472(.data_in(wire_d44_71),.data_out(wire_d44_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4504473(.data_in(wire_d44_72),.data_out(wire_d44_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4504474(.data_in(wire_d44_73),.data_out(wire_d44_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504475(.data_in(wire_d44_74),.data_out(wire_d44_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504476(.data_in(wire_d44_75),.data_out(wire_d44_76),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504477(.data_in(wire_d44_76),.data_out(wire_d44_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4504478(.data_in(wire_d44_77),.data_out(wire_d44_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504479(.data_in(wire_d44_78),.data_out(d_out44),.clk(clk),.rst(rst));

	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance460450(.data_in(d_in45),.data_out(wire_d45_0),.clk(clk),.rst(rst));            //channel 46
	register #(.WIDTH(WIDTH)) register_instance460451(.data_in(wire_d45_0),.data_out(wire_d45_1),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance460452(.data_in(wire_d45_1),.data_out(wire_d45_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance460453(.data_in(wire_d45_2),.data_out(wire_d45_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance460454(.data_in(wire_d45_3),.data_out(wire_d45_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance460455(.data_in(wire_d45_4),.data_out(wire_d45_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance460456(.data_in(wire_d45_5),.data_out(wire_d45_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance460457(.data_in(wire_d45_6),.data_out(wire_d45_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance460458(.data_in(wire_d45_7),.data_out(wire_d45_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance460459(.data_in(wire_d45_8),.data_out(wire_d45_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604510(.data_in(wire_d45_9),.data_out(wire_d45_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4604511(.data_in(wire_d45_10),.data_out(wire_d45_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4604512(.data_in(wire_d45_11),.data_out(wire_d45_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604513(.data_in(wire_d45_12),.data_out(wire_d45_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604514(.data_in(wire_d45_13),.data_out(wire_d45_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604515(.data_in(wire_d45_14),.data_out(wire_d45_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604516(.data_in(wire_d45_15),.data_out(wire_d45_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604517(.data_in(wire_d45_16),.data_out(wire_d45_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4604518(.data_in(wire_d45_17),.data_out(wire_d45_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4604519(.data_in(wire_d45_18),.data_out(wire_d45_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604520(.data_in(wire_d45_19),.data_out(wire_d45_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604521(.data_in(wire_d45_20),.data_out(wire_d45_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4604522(.data_in(wire_d45_21),.data_out(wire_d45_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604523(.data_in(wire_d45_22),.data_out(wire_d45_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604524(.data_in(wire_d45_23),.data_out(wire_d45_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604525(.data_in(wire_d45_24),.data_out(wire_d45_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604526(.data_in(wire_d45_25),.data_out(wire_d45_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604527(.data_in(wire_d45_26),.data_out(wire_d45_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4604528(.data_in(wire_d45_27),.data_out(wire_d45_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4604529(.data_in(wire_d45_28),.data_out(wire_d45_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4604530(.data_in(wire_d45_29),.data_out(wire_d45_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604531(.data_in(wire_d45_30),.data_out(wire_d45_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604532(.data_in(wire_d45_31),.data_out(wire_d45_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604533(.data_in(wire_d45_32),.data_out(wire_d45_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4604534(.data_in(wire_d45_33),.data_out(wire_d45_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604535(.data_in(wire_d45_34),.data_out(wire_d45_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604536(.data_in(wire_d45_35),.data_out(wire_d45_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604537(.data_in(wire_d45_36),.data_out(wire_d45_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604538(.data_in(wire_d45_37),.data_out(wire_d45_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4604539(.data_in(wire_d45_38),.data_out(wire_d45_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604540(.data_in(wire_d45_39),.data_out(wire_d45_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604541(.data_in(wire_d45_40),.data_out(wire_d45_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4604542(.data_in(wire_d45_41),.data_out(wire_d45_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604543(.data_in(wire_d45_42),.data_out(wire_d45_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4604544(.data_in(wire_d45_43),.data_out(wire_d45_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604545(.data_in(wire_d45_44),.data_out(wire_d45_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4604546(.data_in(wire_d45_45),.data_out(wire_d45_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4604547(.data_in(wire_d45_46),.data_out(wire_d45_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604548(.data_in(wire_d45_47),.data_out(wire_d45_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604549(.data_in(wire_d45_48),.data_out(wire_d45_49),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604550(.data_in(wire_d45_49),.data_out(wire_d45_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4604551(.data_in(wire_d45_50),.data_out(wire_d45_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604552(.data_in(wire_d45_51),.data_out(wire_d45_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4604553(.data_in(wire_d45_52),.data_out(wire_d45_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4604554(.data_in(wire_d45_53),.data_out(wire_d45_54),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604555(.data_in(wire_d45_54),.data_out(wire_d45_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604556(.data_in(wire_d45_55),.data_out(wire_d45_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4604557(.data_in(wire_d45_56),.data_out(wire_d45_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4604558(.data_in(wire_d45_57),.data_out(wire_d45_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604559(.data_in(wire_d45_58),.data_out(wire_d45_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4604560(.data_in(wire_d45_59),.data_out(wire_d45_60),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4604561(.data_in(wire_d45_60),.data_out(wire_d45_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4604562(.data_in(wire_d45_61),.data_out(wire_d45_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604563(.data_in(wire_d45_62),.data_out(wire_d45_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604564(.data_in(wire_d45_63),.data_out(wire_d45_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4604565(.data_in(wire_d45_64),.data_out(wire_d45_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604566(.data_in(wire_d45_65),.data_out(wire_d45_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604567(.data_in(wire_d45_66),.data_out(wire_d45_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4604568(.data_in(wire_d45_67),.data_out(wire_d45_68),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604569(.data_in(wire_d45_68),.data_out(wire_d45_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604570(.data_in(wire_d45_69),.data_out(wire_d45_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604571(.data_in(wire_d45_70),.data_out(wire_d45_71),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604572(.data_in(wire_d45_71),.data_out(wire_d45_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4604573(.data_in(wire_d45_72),.data_out(wire_d45_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604574(.data_in(wire_d45_73),.data_out(wire_d45_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4604575(.data_in(wire_d45_74),.data_out(wire_d45_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604576(.data_in(wire_d45_75),.data_out(wire_d45_76),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604577(.data_in(wire_d45_76),.data_out(wire_d45_77),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604578(.data_in(wire_d45_77),.data_out(wire_d45_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4604579(.data_in(wire_d45_78),.data_out(d_out45),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance470460(.data_in(d_in46),.data_out(wire_d46_0),.clk(clk),.rst(rst));            //channel 47
	large_mux #(.WIDTH(WIDTH)) large_mux_instance470461(.data_in(wire_d46_0),.data_out(wire_d46_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance470462(.data_in(wire_d46_1),.data_out(wire_d46_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance470463(.data_in(wire_d46_2),.data_out(wire_d46_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance470464(.data_in(wire_d46_3),.data_out(wire_d46_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance470465(.data_in(wire_d46_4),.data_out(wire_d46_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance470466(.data_in(wire_d46_5),.data_out(wire_d46_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance470467(.data_in(wire_d46_6),.data_out(wire_d46_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance470468(.data_in(wire_d46_7),.data_out(wire_d46_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance470469(.data_in(wire_d46_8),.data_out(wire_d46_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704610(.data_in(wire_d46_9),.data_out(wire_d46_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4704611(.data_in(wire_d46_10),.data_out(wire_d46_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4704612(.data_in(wire_d46_11),.data_out(wire_d46_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4704613(.data_in(wire_d46_12),.data_out(wire_d46_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704614(.data_in(wire_d46_13),.data_out(wire_d46_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704615(.data_in(wire_d46_14),.data_out(wire_d46_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704616(.data_in(wire_d46_15),.data_out(wire_d46_16),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704617(.data_in(wire_d46_16),.data_out(wire_d46_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704618(.data_in(wire_d46_17),.data_out(wire_d46_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704619(.data_in(wire_d46_18),.data_out(wire_d46_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704620(.data_in(wire_d46_19),.data_out(wire_d46_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704621(.data_in(wire_d46_20),.data_out(wire_d46_21),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704622(.data_in(wire_d46_21),.data_out(wire_d46_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704623(.data_in(wire_d46_22),.data_out(wire_d46_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4704624(.data_in(wire_d46_23),.data_out(wire_d46_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704625(.data_in(wire_d46_24),.data_out(wire_d46_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704626(.data_in(wire_d46_25),.data_out(wire_d46_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704627(.data_in(wire_d46_26),.data_out(wire_d46_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704628(.data_in(wire_d46_27),.data_out(wire_d46_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704629(.data_in(wire_d46_28),.data_out(wire_d46_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704630(.data_in(wire_d46_29),.data_out(wire_d46_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704631(.data_in(wire_d46_30),.data_out(wire_d46_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704632(.data_in(wire_d46_31),.data_out(wire_d46_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704633(.data_in(wire_d46_32),.data_out(wire_d46_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4704634(.data_in(wire_d46_33),.data_out(wire_d46_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4704635(.data_in(wire_d46_34),.data_out(wire_d46_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704636(.data_in(wire_d46_35),.data_out(wire_d46_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704637(.data_in(wire_d46_36),.data_out(wire_d46_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704638(.data_in(wire_d46_37),.data_out(wire_d46_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704639(.data_in(wire_d46_38),.data_out(wire_d46_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704640(.data_in(wire_d46_39),.data_out(wire_d46_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704641(.data_in(wire_d46_40),.data_out(wire_d46_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704642(.data_in(wire_d46_41),.data_out(wire_d46_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704643(.data_in(wire_d46_42),.data_out(wire_d46_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704644(.data_in(wire_d46_43),.data_out(wire_d46_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704645(.data_in(wire_d46_44),.data_out(wire_d46_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704646(.data_in(wire_d46_45),.data_out(wire_d46_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704647(.data_in(wire_d46_46),.data_out(wire_d46_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704648(.data_in(wire_d46_47),.data_out(wire_d46_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704649(.data_in(wire_d46_48),.data_out(wire_d46_49),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704650(.data_in(wire_d46_49),.data_out(wire_d46_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704651(.data_in(wire_d46_50),.data_out(wire_d46_51),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704652(.data_in(wire_d46_51),.data_out(wire_d46_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704653(.data_in(wire_d46_52),.data_out(wire_d46_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704654(.data_in(wire_d46_53),.data_out(wire_d46_54),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704655(.data_in(wire_d46_54),.data_out(wire_d46_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704656(.data_in(wire_d46_55),.data_out(wire_d46_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4704657(.data_in(wire_d46_56),.data_out(wire_d46_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704658(.data_in(wire_d46_57),.data_out(wire_d46_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704659(.data_in(wire_d46_58),.data_out(wire_d46_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704660(.data_in(wire_d46_59),.data_out(wire_d46_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4704661(.data_in(wire_d46_60),.data_out(wire_d46_61),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704662(.data_in(wire_d46_61),.data_out(wire_d46_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4704663(.data_in(wire_d46_62),.data_out(wire_d46_63),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704664(.data_in(wire_d46_63),.data_out(wire_d46_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4704665(.data_in(wire_d46_64),.data_out(wire_d46_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704666(.data_in(wire_d46_65),.data_out(wire_d46_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704667(.data_in(wire_d46_66),.data_out(wire_d46_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4704668(.data_in(wire_d46_67),.data_out(wire_d46_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704669(.data_in(wire_d46_68),.data_out(wire_d46_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704670(.data_in(wire_d46_69),.data_out(wire_d46_70),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704671(.data_in(wire_d46_70),.data_out(wire_d46_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704672(.data_in(wire_d46_71),.data_out(wire_d46_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704673(.data_in(wire_d46_72),.data_out(wire_d46_73),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704674(.data_in(wire_d46_73),.data_out(wire_d46_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4704675(.data_in(wire_d46_74),.data_out(wire_d46_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4704676(.data_in(wire_d46_75),.data_out(wire_d46_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704677(.data_in(wire_d46_76),.data_out(wire_d46_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704678(.data_in(wire_d46_77),.data_out(wire_d46_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704679(.data_in(wire_d46_78),.data_out(d_out46),.clk(clk),.rst(rst));

	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance480470(.data_in(d_in47),.data_out(wire_d47_0),.clk(clk),.rst(rst));            //channel 48
	register #(.WIDTH(WIDTH)) register_instance480471(.data_in(wire_d47_0),.data_out(wire_d47_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance480472(.data_in(wire_d47_1),.data_out(wire_d47_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance480473(.data_in(wire_d47_2),.data_out(wire_d47_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance480474(.data_in(wire_d47_3),.data_out(wire_d47_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance480475(.data_in(wire_d47_4),.data_out(wire_d47_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance480476(.data_in(wire_d47_5),.data_out(wire_d47_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance480477(.data_in(wire_d47_6),.data_out(wire_d47_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance480478(.data_in(wire_d47_7),.data_out(wire_d47_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance480479(.data_in(wire_d47_8),.data_out(wire_d47_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804710(.data_in(wire_d47_9),.data_out(wire_d47_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804711(.data_in(wire_d47_10),.data_out(wire_d47_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804712(.data_in(wire_d47_11),.data_out(wire_d47_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804713(.data_in(wire_d47_12),.data_out(wire_d47_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804714(.data_in(wire_d47_13),.data_out(wire_d47_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804715(.data_in(wire_d47_14),.data_out(wire_d47_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4804716(.data_in(wire_d47_15),.data_out(wire_d47_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804717(.data_in(wire_d47_16),.data_out(wire_d47_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4804718(.data_in(wire_d47_17),.data_out(wire_d47_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804719(.data_in(wire_d47_18),.data_out(wire_d47_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4804720(.data_in(wire_d47_19),.data_out(wire_d47_20),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804721(.data_in(wire_d47_20),.data_out(wire_d47_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804722(.data_in(wire_d47_21),.data_out(wire_d47_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804723(.data_in(wire_d47_22),.data_out(wire_d47_23),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804724(.data_in(wire_d47_23),.data_out(wire_d47_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804725(.data_in(wire_d47_24),.data_out(wire_d47_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4804726(.data_in(wire_d47_25),.data_out(wire_d47_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804727(.data_in(wire_d47_26),.data_out(wire_d47_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804728(.data_in(wire_d47_27),.data_out(wire_d47_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804729(.data_in(wire_d47_28),.data_out(wire_d47_29),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804730(.data_in(wire_d47_29),.data_out(wire_d47_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804731(.data_in(wire_d47_30),.data_out(wire_d47_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804732(.data_in(wire_d47_31),.data_out(wire_d47_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804733(.data_in(wire_d47_32),.data_out(wire_d47_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804734(.data_in(wire_d47_33),.data_out(wire_d47_34),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804735(.data_in(wire_d47_34),.data_out(wire_d47_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804736(.data_in(wire_d47_35),.data_out(wire_d47_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4804737(.data_in(wire_d47_36),.data_out(wire_d47_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4804738(.data_in(wire_d47_37),.data_out(wire_d47_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804739(.data_in(wire_d47_38),.data_out(wire_d47_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804740(.data_in(wire_d47_39),.data_out(wire_d47_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804741(.data_in(wire_d47_40),.data_out(wire_d47_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804742(.data_in(wire_d47_41),.data_out(wire_d47_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804743(.data_in(wire_d47_42),.data_out(wire_d47_43),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804744(.data_in(wire_d47_43),.data_out(wire_d47_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804745(.data_in(wire_d47_44),.data_out(wire_d47_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804746(.data_in(wire_d47_45),.data_out(wire_d47_46),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4804747(.data_in(wire_d47_46),.data_out(wire_d47_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804748(.data_in(wire_d47_47),.data_out(wire_d47_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4804749(.data_in(wire_d47_48),.data_out(wire_d47_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804750(.data_in(wire_d47_49),.data_out(wire_d47_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804751(.data_in(wire_d47_50),.data_out(wire_d47_51),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804752(.data_in(wire_d47_51),.data_out(wire_d47_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804753(.data_in(wire_d47_52),.data_out(wire_d47_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804754(.data_in(wire_d47_53),.data_out(wire_d47_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804755(.data_in(wire_d47_54),.data_out(wire_d47_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4804756(.data_in(wire_d47_55),.data_out(wire_d47_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804757(.data_in(wire_d47_56),.data_out(wire_d47_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4804758(.data_in(wire_d47_57),.data_out(wire_d47_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804759(.data_in(wire_d47_58),.data_out(wire_d47_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804760(.data_in(wire_d47_59),.data_out(wire_d47_60),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804761(.data_in(wire_d47_60),.data_out(wire_d47_61),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804762(.data_in(wire_d47_61),.data_out(wire_d47_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804763(.data_in(wire_d47_62),.data_out(wire_d47_63),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4804764(.data_in(wire_d47_63),.data_out(wire_d47_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804765(.data_in(wire_d47_64),.data_out(wire_d47_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804766(.data_in(wire_d47_65),.data_out(wire_d47_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804767(.data_in(wire_d47_66),.data_out(wire_d47_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804768(.data_in(wire_d47_67),.data_out(wire_d47_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804769(.data_in(wire_d47_68),.data_out(wire_d47_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804770(.data_in(wire_d47_69),.data_out(wire_d47_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804771(.data_in(wire_d47_70),.data_out(wire_d47_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4804772(.data_in(wire_d47_71),.data_out(wire_d47_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804773(.data_in(wire_d47_72),.data_out(wire_d47_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804774(.data_in(wire_d47_73),.data_out(wire_d47_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4804775(.data_in(wire_d47_74),.data_out(wire_d47_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804776(.data_in(wire_d47_75),.data_out(wire_d47_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4804777(.data_in(wire_d47_76),.data_out(wire_d47_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804778(.data_in(wire_d47_77),.data_out(wire_d47_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804779(.data_in(wire_d47_78),.data_out(d_out47),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance490480(.data_in(d_in48),.data_out(wire_d48_0),.clk(clk),.rst(rst));            //channel 49
	register #(.WIDTH(WIDTH)) register_instance490481(.data_in(wire_d48_0),.data_out(wire_d48_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance490482(.data_in(wire_d48_1),.data_out(wire_d48_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance490483(.data_in(wire_d48_2),.data_out(wire_d48_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance490484(.data_in(wire_d48_3),.data_out(wire_d48_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance490485(.data_in(wire_d48_4),.data_out(wire_d48_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance490486(.data_in(wire_d48_5),.data_out(wire_d48_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance490487(.data_in(wire_d48_6),.data_out(wire_d48_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance490488(.data_in(wire_d48_7),.data_out(wire_d48_8),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance490489(.data_in(wire_d48_8),.data_out(wire_d48_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904810(.data_in(wire_d48_9),.data_out(wire_d48_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904811(.data_in(wire_d48_10),.data_out(wire_d48_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904812(.data_in(wire_d48_11),.data_out(wire_d48_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904813(.data_in(wire_d48_12),.data_out(wire_d48_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904814(.data_in(wire_d48_13),.data_out(wire_d48_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904815(.data_in(wire_d48_14),.data_out(wire_d48_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4904816(.data_in(wire_d48_15),.data_out(wire_d48_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904817(.data_in(wire_d48_16),.data_out(wire_d48_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904818(.data_in(wire_d48_17),.data_out(wire_d48_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904819(.data_in(wire_d48_18),.data_out(wire_d48_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904820(.data_in(wire_d48_19),.data_out(wire_d48_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904821(.data_in(wire_d48_20),.data_out(wire_d48_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904822(.data_in(wire_d48_21),.data_out(wire_d48_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904823(.data_in(wire_d48_22),.data_out(wire_d48_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904824(.data_in(wire_d48_23),.data_out(wire_d48_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904825(.data_in(wire_d48_24),.data_out(wire_d48_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4904826(.data_in(wire_d48_25),.data_out(wire_d48_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4904827(.data_in(wire_d48_26),.data_out(wire_d48_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904828(.data_in(wire_d48_27),.data_out(wire_d48_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904829(.data_in(wire_d48_28),.data_out(wire_d48_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4904830(.data_in(wire_d48_29),.data_out(wire_d48_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904831(.data_in(wire_d48_30),.data_out(wire_d48_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4904832(.data_in(wire_d48_31),.data_out(wire_d48_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904833(.data_in(wire_d48_32),.data_out(wire_d48_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904834(.data_in(wire_d48_33),.data_out(wire_d48_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904835(.data_in(wire_d48_34),.data_out(wire_d48_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4904836(.data_in(wire_d48_35),.data_out(wire_d48_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4904837(.data_in(wire_d48_36),.data_out(wire_d48_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904838(.data_in(wire_d48_37),.data_out(wire_d48_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904839(.data_in(wire_d48_38),.data_out(wire_d48_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904840(.data_in(wire_d48_39),.data_out(wire_d48_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4904841(.data_in(wire_d48_40),.data_out(wire_d48_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904842(.data_in(wire_d48_41),.data_out(wire_d48_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904843(.data_in(wire_d48_42),.data_out(wire_d48_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904844(.data_in(wire_d48_43),.data_out(wire_d48_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904845(.data_in(wire_d48_44),.data_out(wire_d48_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904846(.data_in(wire_d48_45),.data_out(wire_d48_46),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904847(.data_in(wire_d48_46),.data_out(wire_d48_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904848(.data_in(wire_d48_47),.data_out(wire_d48_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4904849(.data_in(wire_d48_48),.data_out(wire_d48_49),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904850(.data_in(wire_d48_49),.data_out(wire_d48_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904851(.data_in(wire_d48_50),.data_out(wire_d48_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904852(.data_in(wire_d48_51),.data_out(wire_d48_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904853(.data_in(wire_d48_52),.data_out(wire_d48_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904854(.data_in(wire_d48_53),.data_out(wire_d48_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904855(.data_in(wire_d48_54),.data_out(wire_d48_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904856(.data_in(wire_d48_55),.data_out(wire_d48_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904857(.data_in(wire_d48_56),.data_out(wire_d48_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904858(.data_in(wire_d48_57),.data_out(wire_d48_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4904859(.data_in(wire_d48_58),.data_out(wire_d48_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904860(.data_in(wire_d48_59),.data_out(wire_d48_60),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904861(.data_in(wire_d48_60),.data_out(wire_d48_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904862(.data_in(wire_d48_61),.data_out(wire_d48_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904863(.data_in(wire_d48_62),.data_out(wire_d48_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904864(.data_in(wire_d48_63),.data_out(wire_d48_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904865(.data_in(wire_d48_64),.data_out(wire_d48_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904866(.data_in(wire_d48_65),.data_out(wire_d48_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904867(.data_in(wire_d48_66),.data_out(wire_d48_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904868(.data_in(wire_d48_67),.data_out(wire_d48_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904869(.data_in(wire_d48_68),.data_out(wire_d48_69),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904870(.data_in(wire_d48_69),.data_out(wire_d48_70),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904871(.data_in(wire_d48_70),.data_out(wire_d48_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4904872(.data_in(wire_d48_71),.data_out(wire_d48_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904873(.data_in(wire_d48_72),.data_out(wire_d48_73),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904874(.data_in(wire_d48_73),.data_out(wire_d48_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904875(.data_in(wire_d48_74),.data_out(wire_d48_75),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904876(.data_in(wire_d48_75),.data_out(wire_d48_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904877(.data_in(wire_d48_76),.data_out(wire_d48_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904878(.data_in(wire_d48_77),.data_out(wire_d48_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4904879(.data_in(wire_d48_78),.data_out(d_out48),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance500490(.data_in(d_in49),.data_out(wire_d49_0),.clk(clk),.rst(rst));            //channel 50
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance500491(.data_in(wire_d49_0),.data_out(wire_d49_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance500492(.data_in(wire_d49_1),.data_out(wire_d49_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance500493(.data_in(wire_d49_2),.data_out(wire_d49_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance500494(.data_in(wire_d49_3),.data_out(wire_d49_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance500495(.data_in(wire_d49_4),.data_out(wire_d49_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance500496(.data_in(wire_d49_5),.data_out(wire_d49_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance500497(.data_in(wire_d49_6),.data_out(wire_d49_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance500498(.data_in(wire_d49_7),.data_out(wire_d49_8),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance500499(.data_in(wire_d49_8),.data_out(wire_d49_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004910(.data_in(wire_d49_9),.data_out(wire_d49_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004911(.data_in(wire_d49_10),.data_out(wire_d49_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004912(.data_in(wire_d49_11),.data_out(wire_d49_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004913(.data_in(wire_d49_12),.data_out(wire_d49_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004914(.data_in(wire_d49_13),.data_out(wire_d49_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004915(.data_in(wire_d49_14),.data_out(wire_d49_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004916(.data_in(wire_d49_15),.data_out(wire_d49_16),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004917(.data_in(wire_d49_16),.data_out(wire_d49_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004918(.data_in(wire_d49_17),.data_out(wire_d49_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004919(.data_in(wire_d49_18),.data_out(wire_d49_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004920(.data_in(wire_d49_19),.data_out(wire_d49_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004921(.data_in(wire_d49_20),.data_out(wire_d49_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004922(.data_in(wire_d49_21),.data_out(wire_d49_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004923(.data_in(wire_d49_22),.data_out(wire_d49_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004924(.data_in(wire_d49_23),.data_out(wire_d49_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004925(.data_in(wire_d49_24),.data_out(wire_d49_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004926(.data_in(wire_d49_25),.data_out(wire_d49_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004927(.data_in(wire_d49_26),.data_out(wire_d49_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004928(.data_in(wire_d49_27),.data_out(wire_d49_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004929(.data_in(wire_d49_28),.data_out(wire_d49_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004930(.data_in(wire_d49_29),.data_out(wire_d49_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004931(.data_in(wire_d49_30),.data_out(wire_d49_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004932(.data_in(wire_d49_31),.data_out(wire_d49_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004933(.data_in(wire_d49_32),.data_out(wire_d49_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004934(.data_in(wire_d49_33),.data_out(wire_d49_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004935(.data_in(wire_d49_34),.data_out(wire_d49_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5004936(.data_in(wire_d49_35),.data_out(wire_d49_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004937(.data_in(wire_d49_36),.data_out(wire_d49_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004938(.data_in(wire_d49_37),.data_out(wire_d49_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004939(.data_in(wire_d49_38),.data_out(wire_d49_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5004940(.data_in(wire_d49_39),.data_out(wire_d49_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004941(.data_in(wire_d49_40),.data_out(wire_d49_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004942(.data_in(wire_d49_41),.data_out(wire_d49_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004943(.data_in(wire_d49_42),.data_out(wire_d49_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004944(.data_in(wire_d49_43),.data_out(wire_d49_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004945(.data_in(wire_d49_44),.data_out(wire_d49_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004946(.data_in(wire_d49_45),.data_out(wire_d49_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004947(.data_in(wire_d49_46),.data_out(wire_d49_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004948(.data_in(wire_d49_47),.data_out(wire_d49_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004949(.data_in(wire_d49_48),.data_out(wire_d49_49),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004950(.data_in(wire_d49_49),.data_out(wire_d49_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004951(.data_in(wire_d49_50),.data_out(wire_d49_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5004952(.data_in(wire_d49_51),.data_out(wire_d49_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004953(.data_in(wire_d49_52),.data_out(wire_d49_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004954(.data_in(wire_d49_53),.data_out(wire_d49_54),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004955(.data_in(wire_d49_54),.data_out(wire_d49_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004956(.data_in(wire_d49_55),.data_out(wire_d49_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004957(.data_in(wire_d49_56),.data_out(wire_d49_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004958(.data_in(wire_d49_57),.data_out(wire_d49_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004959(.data_in(wire_d49_58),.data_out(wire_d49_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004960(.data_in(wire_d49_59),.data_out(wire_d49_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004961(.data_in(wire_d49_60),.data_out(wire_d49_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004962(.data_in(wire_d49_61),.data_out(wire_d49_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004963(.data_in(wire_d49_62),.data_out(wire_d49_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004964(.data_in(wire_d49_63),.data_out(wire_d49_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004965(.data_in(wire_d49_64),.data_out(wire_d49_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004966(.data_in(wire_d49_65),.data_out(wire_d49_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004967(.data_in(wire_d49_66),.data_out(wire_d49_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004968(.data_in(wire_d49_67),.data_out(wire_d49_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004969(.data_in(wire_d49_68),.data_out(wire_d49_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5004970(.data_in(wire_d49_69),.data_out(wire_d49_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004971(.data_in(wire_d49_70),.data_out(wire_d49_71),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004972(.data_in(wire_d49_71),.data_out(wire_d49_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004973(.data_in(wire_d49_72),.data_out(wire_d49_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004974(.data_in(wire_d49_73),.data_out(wire_d49_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004975(.data_in(wire_d49_74),.data_out(wire_d49_75),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004976(.data_in(wire_d49_75),.data_out(wire_d49_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004977(.data_in(wire_d49_76),.data_out(wire_d49_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004978(.data_in(wire_d49_77),.data_out(wire_d49_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004979(.data_in(wire_d49_78),.data_out(d_out49),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance510500(.data_in(d_in50),.data_out(wire_d50_0),.clk(clk),.rst(rst));            //channel 51
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance510501(.data_in(wire_d50_0),.data_out(wire_d50_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance510502(.data_in(wire_d50_1),.data_out(wire_d50_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance510503(.data_in(wire_d50_2),.data_out(wire_d50_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance510504(.data_in(wire_d50_3),.data_out(wire_d50_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance510505(.data_in(wire_d50_4),.data_out(wire_d50_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance510506(.data_in(wire_d50_5),.data_out(wire_d50_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance510507(.data_in(wire_d50_6),.data_out(wire_d50_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance510508(.data_in(wire_d50_7),.data_out(wire_d50_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance510509(.data_in(wire_d50_8),.data_out(wire_d50_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105010(.data_in(wire_d50_9),.data_out(wire_d50_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105011(.data_in(wire_d50_10),.data_out(wire_d50_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5105012(.data_in(wire_d50_11),.data_out(wire_d50_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5105013(.data_in(wire_d50_12),.data_out(wire_d50_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105014(.data_in(wire_d50_13),.data_out(wire_d50_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105015(.data_in(wire_d50_14),.data_out(wire_d50_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105016(.data_in(wire_d50_15),.data_out(wire_d50_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5105017(.data_in(wire_d50_16),.data_out(wire_d50_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5105018(.data_in(wire_d50_17),.data_out(wire_d50_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5105019(.data_in(wire_d50_18),.data_out(wire_d50_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105020(.data_in(wire_d50_19),.data_out(wire_d50_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105021(.data_in(wire_d50_20),.data_out(wire_d50_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5105022(.data_in(wire_d50_21),.data_out(wire_d50_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5105023(.data_in(wire_d50_22),.data_out(wire_d50_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5105024(.data_in(wire_d50_23),.data_out(wire_d50_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5105025(.data_in(wire_d50_24),.data_out(wire_d50_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105026(.data_in(wire_d50_25),.data_out(wire_d50_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105027(.data_in(wire_d50_26),.data_out(wire_d50_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105028(.data_in(wire_d50_27),.data_out(wire_d50_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5105029(.data_in(wire_d50_28),.data_out(wire_d50_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105030(.data_in(wire_d50_29),.data_out(wire_d50_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105031(.data_in(wire_d50_30),.data_out(wire_d50_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105032(.data_in(wire_d50_31),.data_out(wire_d50_32),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105033(.data_in(wire_d50_32),.data_out(wire_d50_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105034(.data_in(wire_d50_33),.data_out(wire_d50_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105035(.data_in(wire_d50_34),.data_out(wire_d50_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105036(.data_in(wire_d50_35),.data_out(wire_d50_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5105037(.data_in(wire_d50_36),.data_out(wire_d50_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105038(.data_in(wire_d50_37),.data_out(wire_d50_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105039(.data_in(wire_d50_38),.data_out(wire_d50_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105040(.data_in(wire_d50_39),.data_out(wire_d50_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105041(.data_in(wire_d50_40),.data_out(wire_d50_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5105042(.data_in(wire_d50_41),.data_out(wire_d50_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105043(.data_in(wire_d50_42),.data_out(wire_d50_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5105044(.data_in(wire_d50_43),.data_out(wire_d50_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105045(.data_in(wire_d50_44),.data_out(wire_d50_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105046(.data_in(wire_d50_45),.data_out(wire_d50_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105047(.data_in(wire_d50_46),.data_out(wire_d50_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5105048(.data_in(wire_d50_47),.data_out(wire_d50_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105049(.data_in(wire_d50_48),.data_out(wire_d50_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5105050(.data_in(wire_d50_49),.data_out(wire_d50_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5105051(.data_in(wire_d50_50),.data_out(wire_d50_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105052(.data_in(wire_d50_51),.data_out(wire_d50_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5105053(.data_in(wire_d50_52),.data_out(wire_d50_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5105054(.data_in(wire_d50_53),.data_out(wire_d50_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105055(.data_in(wire_d50_54),.data_out(wire_d50_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5105056(.data_in(wire_d50_55),.data_out(wire_d50_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5105057(.data_in(wire_d50_56),.data_out(wire_d50_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5105058(.data_in(wire_d50_57),.data_out(wire_d50_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5105059(.data_in(wire_d50_58),.data_out(wire_d50_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105060(.data_in(wire_d50_59),.data_out(wire_d50_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105061(.data_in(wire_d50_60),.data_out(wire_d50_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105062(.data_in(wire_d50_61),.data_out(wire_d50_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5105063(.data_in(wire_d50_62),.data_out(wire_d50_63),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5105064(.data_in(wire_d50_63),.data_out(wire_d50_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105065(.data_in(wire_d50_64),.data_out(wire_d50_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105066(.data_in(wire_d50_65),.data_out(wire_d50_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5105067(.data_in(wire_d50_66),.data_out(wire_d50_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105068(.data_in(wire_d50_67),.data_out(wire_d50_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5105069(.data_in(wire_d50_68),.data_out(wire_d50_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105070(.data_in(wire_d50_69),.data_out(wire_d50_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105071(.data_in(wire_d50_70),.data_out(wire_d50_71),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5105072(.data_in(wire_d50_71),.data_out(wire_d50_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105073(.data_in(wire_d50_72),.data_out(wire_d50_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105074(.data_in(wire_d50_73),.data_out(wire_d50_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5105075(.data_in(wire_d50_74),.data_out(wire_d50_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105076(.data_in(wire_d50_75),.data_out(wire_d50_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105077(.data_in(wire_d50_76),.data_out(wire_d50_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105078(.data_in(wire_d50_77),.data_out(wire_d50_78),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5105079(.data_in(wire_d50_78),.data_out(d_out50),.clk(clk),.rst(rst));

	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance520510(.data_in(d_in51),.data_out(wire_d51_0),.clk(clk),.rst(rst));            //channel 52
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance520511(.data_in(wire_d51_0),.data_out(wire_d51_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance520512(.data_in(wire_d51_1),.data_out(wire_d51_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance520513(.data_in(wire_d51_2),.data_out(wire_d51_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance520514(.data_in(wire_d51_3),.data_out(wire_d51_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance520515(.data_in(wire_d51_4),.data_out(wire_d51_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance520516(.data_in(wire_d51_5),.data_out(wire_d51_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance520517(.data_in(wire_d51_6),.data_out(wire_d51_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance520518(.data_in(wire_d51_7),.data_out(wire_d51_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance520519(.data_in(wire_d51_8),.data_out(wire_d51_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205110(.data_in(wire_d51_9),.data_out(wire_d51_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5205111(.data_in(wire_d51_10),.data_out(wire_d51_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205112(.data_in(wire_d51_11),.data_out(wire_d51_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205113(.data_in(wire_d51_12),.data_out(wire_d51_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205114(.data_in(wire_d51_13),.data_out(wire_d51_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5205115(.data_in(wire_d51_14),.data_out(wire_d51_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205116(.data_in(wire_d51_15),.data_out(wire_d51_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205117(.data_in(wire_d51_16),.data_out(wire_d51_17),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205118(.data_in(wire_d51_17),.data_out(wire_d51_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205119(.data_in(wire_d51_18),.data_out(wire_d51_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5205120(.data_in(wire_d51_19),.data_out(wire_d51_20),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205121(.data_in(wire_d51_20),.data_out(wire_d51_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205122(.data_in(wire_d51_21),.data_out(wire_d51_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205123(.data_in(wire_d51_22),.data_out(wire_d51_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205124(.data_in(wire_d51_23),.data_out(wire_d51_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205125(.data_in(wire_d51_24),.data_out(wire_d51_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205126(.data_in(wire_d51_25),.data_out(wire_d51_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5205127(.data_in(wire_d51_26),.data_out(wire_d51_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205128(.data_in(wire_d51_27),.data_out(wire_d51_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5205129(.data_in(wire_d51_28),.data_out(wire_d51_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205130(.data_in(wire_d51_29),.data_out(wire_d51_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205131(.data_in(wire_d51_30),.data_out(wire_d51_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205132(.data_in(wire_d51_31),.data_out(wire_d51_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205133(.data_in(wire_d51_32),.data_out(wire_d51_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5205134(.data_in(wire_d51_33),.data_out(wire_d51_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5205135(.data_in(wire_d51_34),.data_out(wire_d51_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205136(.data_in(wire_d51_35),.data_out(wire_d51_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5205137(.data_in(wire_d51_36),.data_out(wire_d51_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5205138(.data_in(wire_d51_37),.data_out(wire_d51_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205139(.data_in(wire_d51_38),.data_out(wire_d51_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205140(.data_in(wire_d51_39),.data_out(wire_d51_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5205141(.data_in(wire_d51_40),.data_out(wire_d51_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205142(.data_in(wire_d51_41),.data_out(wire_d51_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205143(.data_in(wire_d51_42),.data_out(wire_d51_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5205144(.data_in(wire_d51_43),.data_out(wire_d51_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205145(.data_in(wire_d51_44),.data_out(wire_d51_45),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5205146(.data_in(wire_d51_45),.data_out(wire_d51_46),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205147(.data_in(wire_d51_46),.data_out(wire_d51_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205148(.data_in(wire_d51_47),.data_out(wire_d51_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205149(.data_in(wire_d51_48),.data_out(wire_d51_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205150(.data_in(wire_d51_49),.data_out(wire_d51_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205151(.data_in(wire_d51_50),.data_out(wire_d51_51),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205152(.data_in(wire_d51_51),.data_out(wire_d51_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205153(.data_in(wire_d51_52),.data_out(wire_d51_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5205154(.data_in(wire_d51_53),.data_out(wire_d51_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5205155(.data_in(wire_d51_54),.data_out(wire_d51_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205156(.data_in(wire_d51_55),.data_out(wire_d51_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205157(.data_in(wire_d51_56),.data_out(wire_d51_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5205158(.data_in(wire_d51_57),.data_out(wire_d51_58),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5205159(.data_in(wire_d51_58),.data_out(wire_d51_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205160(.data_in(wire_d51_59),.data_out(wire_d51_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205161(.data_in(wire_d51_60),.data_out(wire_d51_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205162(.data_in(wire_d51_61),.data_out(wire_d51_62),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205163(.data_in(wire_d51_62),.data_out(wire_d51_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5205164(.data_in(wire_d51_63),.data_out(wire_d51_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205165(.data_in(wire_d51_64),.data_out(wire_d51_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205166(.data_in(wire_d51_65),.data_out(wire_d51_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205167(.data_in(wire_d51_66),.data_out(wire_d51_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5205168(.data_in(wire_d51_67),.data_out(wire_d51_68),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205169(.data_in(wire_d51_68),.data_out(wire_d51_69),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205170(.data_in(wire_d51_69),.data_out(wire_d51_70),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5205171(.data_in(wire_d51_70),.data_out(wire_d51_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205172(.data_in(wire_d51_71),.data_out(wire_d51_72),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5205173(.data_in(wire_d51_72),.data_out(wire_d51_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205174(.data_in(wire_d51_73),.data_out(wire_d51_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205175(.data_in(wire_d51_74),.data_out(wire_d51_75),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205176(.data_in(wire_d51_75),.data_out(wire_d51_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205177(.data_in(wire_d51_76),.data_out(wire_d51_77),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205178(.data_in(wire_d51_77),.data_out(wire_d51_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205179(.data_in(wire_d51_78),.data_out(d_out51),.clk(clk),.rst(rst));

	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance530520(.data_in(d_in52),.data_out(wire_d52_0),.clk(clk),.rst(rst));            //channel 53
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance530521(.data_in(wire_d52_0),.data_out(wire_d52_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance530522(.data_in(wire_d52_1),.data_out(wire_d52_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance530523(.data_in(wire_d52_2),.data_out(wire_d52_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance530524(.data_in(wire_d52_3),.data_out(wire_d52_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance530525(.data_in(wire_d52_4),.data_out(wire_d52_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance530526(.data_in(wire_d52_5),.data_out(wire_d52_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance530527(.data_in(wire_d52_6),.data_out(wire_d52_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance530528(.data_in(wire_d52_7),.data_out(wire_d52_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance530529(.data_in(wire_d52_8),.data_out(wire_d52_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305210(.data_in(wire_d52_9),.data_out(wire_d52_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305211(.data_in(wire_d52_10),.data_out(wire_d52_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305212(.data_in(wire_d52_11),.data_out(wire_d52_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305213(.data_in(wire_d52_12),.data_out(wire_d52_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305214(.data_in(wire_d52_13),.data_out(wire_d52_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305215(.data_in(wire_d52_14),.data_out(wire_d52_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305216(.data_in(wire_d52_15),.data_out(wire_d52_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305217(.data_in(wire_d52_16),.data_out(wire_d52_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305218(.data_in(wire_d52_17),.data_out(wire_d52_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305219(.data_in(wire_d52_18),.data_out(wire_d52_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305220(.data_in(wire_d52_19),.data_out(wire_d52_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305221(.data_in(wire_d52_20),.data_out(wire_d52_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305222(.data_in(wire_d52_21),.data_out(wire_d52_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5305223(.data_in(wire_d52_22),.data_out(wire_d52_23),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305224(.data_in(wire_d52_23),.data_out(wire_d52_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305225(.data_in(wire_d52_24),.data_out(wire_d52_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5305226(.data_in(wire_d52_25),.data_out(wire_d52_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305227(.data_in(wire_d52_26),.data_out(wire_d52_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5305228(.data_in(wire_d52_27),.data_out(wire_d52_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305229(.data_in(wire_d52_28),.data_out(wire_d52_29),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5305230(.data_in(wire_d52_29),.data_out(wire_d52_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305231(.data_in(wire_d52_30),.data_out(wire_d52_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305232(.data_in(wire_d52_31),.data_out(wire_d52_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305233(.data_in(wire_d52_32),.data_out(wire_d52_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305234(.data_in(wire_d52_33),.data_out(wire_d52_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305235(.data_in(wire_d52_34),.data_out(wire_d52_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305236(.data_in(wire_d52_35),.data_out(wire_d52_36),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305237(.data_in(wire_d52_36),.data_out(wire_d52_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305238(.data_in(wire_d52_37),.data_out(wire_d52_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305239(.data_in(wire_d52_38),.data_out(wire_d52_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305240(.data_in(wire_d52_39),.data_out(wire_d52_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305241(.data_in(wire_d52_40),.data_out(wire_d52_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305242(.data_in(wire_d52_41),.data_out(wire_d52_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305243(.data_in(wire_d52_42),.data_out(wire_d52_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305244(.data_in(wire_d52_43),.data_out(wire_d52_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305245(.data_in(wire_d52_44),.data_out(wire_d52_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305246(.data_in(wire_d52_45),.data_out(wire_d52_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305247(.data_in(wire_d52_46),.data_out(wire_d52_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305248(.data_in(wire_d52_47),.data_out(wire_d52_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305249(.data_in(wire_d52_48),.data_out(wire_d52_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305250(.data_in(wire_d52_49),.data_out(wire_d52_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305251(.data_in(wire_d52_50),.data_out(wire_d52_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305252(.data_in(wire_d52_51),.data_out(wire_d52_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305253(.data_in(wire_d52_52),.data_out(wire_d52_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305254(.data_in(wire_d52_53),.data_out(wire_d52_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305255(.data_in(wire_d52_54),.data_out(wire_d52_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305256(.data_in(wire_d52_55),.data_out(wire_d52_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305257(.data_in(wire_d52_56),.data_out(wire_d52_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305258(.data_in(wire_d52_57),.data_out(wire_d52_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305259(.data_in(wire_d52_58),.data_out(wire_d52_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305260(.data_in(wire_d52_59),.data_out(wire_d52_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305261(.data_in(wire_d52_60),.data_out(wire_d52_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305262(.data_in(wire_d52_61),.data_out(wire_d52_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305263(.data_in(wire_d52_62),.data_out(wire_d52_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305264(.data_in(wire_d52_63),.data_out(wire_d52_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305265(.data_in(wire_d52_64),.data_out(wire_d52_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305266(.data_in(wire_d52_65),.data_out(wire_d52_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5305267(.data_in(wire_d52_66),.data_out(wire_d52_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305268(.data_in(wire_d52_67),.data_out(wire_d52_68),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305269(.data_in(wire_d52_68),.data_out(wire_d52_69),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305270(.data_in(wire_d52_69),.data_out(wire_d52_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305271(.data_in(wire_d52_70),.data_out(wire_d52_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305272(.data_in(wire_d52_71),.data_out(wire_d52_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305273(.data_in(wire_d52_72),.data_out(wire_d52_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305274(.data_in(wire_d52_73),.data_out(wire_d52_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305275(.data_in(wire_d52_74),.data_out(wire_d52_75),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305276(.data_in(wire_d52_75),.data_out(wire_d52_76),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305277(.data_in(wire_d52_76),.data_out(wire_d52_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305278(.data_in(wire_d52_77),.data_out(wire_d52_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305279(.data_in(wire_d52_78),.data_out(d_out52),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance540530(.data_in(d_in53),.data_out(wire_d53_0),.clk(clk),.rst(rst));            //channel 54
	register #(.WIDTH(WIDTH)) register_instance540531(.data_in(wire_d53_0),.data_out(wire_d53_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance540532(.data_in(wire_d53_1),.data_out(wire_d53_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance540533(.data_in(wire_d53_2),.data_out(wire_d53_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance540534(.data_in(wire_d53_3),.data_out(wire_d53_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance540535(.data_in(wire_d53_4),.data_out(wire_d53_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance540536(.data_in(wire_d53_5),.data_out(wire_d53_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance540537(.data_in(wire_d53_6),.data_out(wire_d53_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance540538(.data_in(wire_d53_7),.data_out(wire_d53_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance540539(.data_in(wire_d53_8),.data_out(wire_d53_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5405310(.data_in(wire_d53_9),.data_out(wire_d53_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405311(.data_in(wire_d53_10),.data_out(wire_d53_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5405312(.data_in(wire_d53_11),.data_out(wire_d53_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5405313(.data_in(wire_d53_12),.data_out(wire_d53_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405314(.data_in(wire_d53_13),.data_out(wire_d53_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405315(.data_in(wire_d53_14),.data_out(wire_d53_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405316(.data_in(wire_d53_15),.data_out(wire_d53_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405317(.data_in(wire_d53_16),.data_out(wire_d53_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5405318(.data_in(wire_d53_17),.data_out(wire_d53_18),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405319(.data_in(wire_d53_18),.data_out(wire_d53_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405320(.data_in(wire_d53_19),.data_out(wire_d53_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405321(.data_in(wire_d53_20),.data_out(wire_d53_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405322(.data_in(wire_d53_21),.data_out(wire_d53_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405323(.data_in(wire_d53_22),.data_out(wire_d53_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405324(.data_in(wire_d53_23),.data_out(wire_d53_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5405325(.data_in(wire_d53_24),.data_out(wire_d53_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405326(.data_in(wire_d53_25),.data_out(wire_d53_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405327(.data_in(wire_d53_26),.data_out(wire_d53_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405328(.data_in(wire_d53_27),.data_out(wire_d53_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5405329(.data_in(wire_d53_28),.data_out(wire_d53_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405330(.data_in(wire_d53_29),.data_out(wire_d53_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405331(.data_in(wire_d53_30),.data_out(wire_d53_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5405332(.data_in(wire_d53_31),.data_out(wire_d53_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405333(.data_in(wire_d53_32),.data_out(wire_d53_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405334(.data_in(wire_d53_33),.data_out(wire_d53_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405335(.data_in(wire_d53_34),.data_out(wire_d53_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5405336(.data_in(wire_d53_35),.data_out(wire_d53_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405337(.data_in(wire_d53_36),.data_out(wire_d53_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5405338(.data_in(wire_d53_37),.data_out(wire_d53_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405339(.data_in(wire_d53_38),.data_out(wire_d53_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405340(.data_in(wire_d53_39),.data_out(wire_d53_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405341(.data_in(wire_d53_40),.data_out(wire_d53_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405342(.data_in(wire_d53_41),.data_out(wire_d53_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5405343(.data_in(wire_d53_42),.data_out(wire_d53_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5405344(.data_in(wire_d53_43),.data_out(wire_d53_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5405345(.data_in(wire_d53_44),.data_out(wire_d53_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405346(.data_in(wire_d53_45),.data_out(wire_d53_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5405347(.data_in(wire_d53_46),.data_out(wire_d53_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405348(.data_in(wire_d53_47),.data_out(wire_d53_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405349(.data_in(wire_d53_48),.data_out(wire_d53_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405350(.data_in(wire_d53_49),.data_out(wire_d53_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5405351(.data_in(wire_d53_50),.data_out(wire_d53_51),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5405352(.data_in(wire_d53_51),.data_out(wire_d53_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405353(.data_in(wire_d53_52),.data_out(wire_d53_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405354(.data_in(wire_d53_53),.data_out(wire_d53_54),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5405355(.data_in(wire_d53_54),.data_out(wire_d53_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405356(.data_in(wire_d53_55),.data_out(wire_d53_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405357(.data_in(wire_d53_56),.data_out(wire_d53_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5405358(.data_in(wire_d53_57),.data_out(wire_d53_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5405359(.data_in(wire_d53_58),.data_out(wire_d53_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405360(.data_in(wire_d53_59),.data_out(wire_d53_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405361(.data_in(wire_d53_60),.data_out(wire_d53_61),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405362(.data_in(wire_d53_61),.data_out(wire_d53_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405363(.data_in(wire_d53_62),.data_out(wire_d53_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405364(.data_in(wire_d53_63),.data_out(wire_d53_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405365(.data_in(wire_d53_64),.data_out(wire_d53_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405366(.data_in(wire_d53_65),.data_out(wire_d53_66),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405367(.data_in(wire_d53_66),.data_out(wire_d53_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5405368(.data_in(wire_d53_67),.data_out(wire_d53_68),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405369(.data_in(wire_d53_68),.data_out(wire_d53_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5405370(.data_in(wire_d53_69),.data_out(wire_d53_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405371(.data_in(wire_d53_70),.data_out(wire_d53_71),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405372(.data_in(wire_d53_71),.data_out(wire_d53_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405373(.data_in(wire_d53_72),.data_out(wire_d53_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405374(.data_in(wire_d53_73),.data_out(wire_d53_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5405375(.data_in(wire_d53_74),.data_out(wire_d53_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5405376(.data_in(wire_d53_75),.data_out(wire_d53_76),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405377(.data_in(wire_d53_76),.data_out(wire_d53_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405378(.data_in(wire_d53_77),.data_out(wire_d53_78),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405379(.data_in(wire_d53_78),.data_out(d_out53),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance550540(.data_in(d_in54),.data_out(wire_d54_0),.clk(clk),.rst(rst));            //channel 55
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance550541(.data_in(wire_d54_0),.data_out(wire_d54_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance550542(.data_in(wire_d54_1),.data_out(wire_d54_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance550543(.data_in(wire_d54_2),.data_out(wire_d54_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance550544(.data_in(wire_d54_3),.data_out(wire_d54_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance550545(.data_in(wire_d54_4),.data_out(wire_d54_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance550546(.data_in(wire_d54_5),.data_out(wire_d54_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance550547(.data_in(wire_d54_6),.data_out(wire_d54_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance550548(.data_in(wire_d54_7),.data_out(wire_d54_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance550549(.data_in(wire_d54_8),.data_out(wire_d54_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505410(.data_in(wire_d54_9),.data_out(wire_d54_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505411(.data_in(wire_d54_10),.data_out(wire_d54_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505412(.data_in(wire_d54_11),.data_out(wire_d54_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505413(.data_in(wire_d54_12),.data_out(wire_d54_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505414(.data_in(wire_d54_13),.data_out(wire_d54_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505415(.data_in(wire_d54_14),.data_out(wire_d54_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5505416(.data_in(wire_d54_15),.data_out(wire_d54_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505417(.data_in(wire_d54_16),.data_out(wire_d54_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5505418(.data_in(wire_d54_17),.data_out(wire_d54_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505419(.data_in(wire_d54_18),.data_out(wire_d54_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505420(.data_in(wire_d54_19),.data_out(wire_d54_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505421(.data_in(wire_d54_20),.data_out(wire_d54_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505422(.data_in(wire_d54_21),.data_out(wire_d54_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505423(.data_in(wire_d54_22),.data_out(wire_d54_23),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505424(.data_in(wire_d54_23),.data_out(wire_d54_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5505425(.data_in(wire_d54_24),.data_out(wire_d54_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505426(.data_in(wire_d54_25),.data_out(wire_d54_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5505427(.data_in(wire_d54_26),.data_out(wire_d54_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505428(.data_in(wire_d54_27),.data_out(wire_d54_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505429(.data_in(wire_d54_28),.data_out(wire_d54_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5505430(.data_in(wire_d54_29),.data_out(wire_d54_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505431(.data_in(wire_d54_30),.data_out(wire_d54_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505432(.data_in(wire_d54_31),.data_out(wire_d54_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5505433(.data_in(wire_d54_32),.data_out(wire_d54_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505434(.data_in(wire_d54_33),.data_out(wire_d54_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505435(.data_in(wire_d54_34),.data_out(wire_d54_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505436(.data_in(wire_d54_35),.data_out(wire_d54_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505437(.data_in(wire_d54_36),.data_out(wire_d54_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505438(.data_in(wire_d54_37),.data_out(wire_d54_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505439(.data_in(wire_d54_38),.data_out(wire_d54_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505440(.data_in(wire_d54_39),.data_out(wire_d54_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5505441(.data_in(wire_d54_40),.data_out(wire_d54_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5505442(.data_in(wire_d54_41),.data_out(wire_d54_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505443(.data_in(wire_d54_42),.data_out(wire_d54_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505444(.data_in(wire_d54_43),.data_out(wire_d54_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505445(.data_in(wire_d54_44),.data_out(wire_d54_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505446(.data_in(wire_d54_45),.data_out(wire_d54_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505447(.data_in(wire_d54_46),.data_out(wire_d54_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5505448(.data_in(wire_d54_47),.data_out(wire_d54_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505449(.data_in(wire_d54_48),.data_out(wire_d54_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505450(.data_in(wire_d54_49),.data_out(wire_d54_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505451(.data_in(wire_d54_50),.data_out(wire_d54_51),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505452(.data_in(wire_d54_51),.data_out(wire_d54_52),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505453(.data_in(wire_d54_52),.data_out(wire_d54_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5505454(.data_in(wire_d54_53),.data_out(wire_d54_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505455(.data_in(wire_d54_54),.data_out(wire_d54_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505456(.data_in(wire_d54_55),.data_out(wire_d54_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505457(.data_in(wire_d54_56),.data_out(wire_d54_57),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505458(.data_in(wire_d54_57),.data_out(wire_d54_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5505459(.data_in(wire_d54_58),.data_out(wire_d54_59),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505460(.data_in(wire_d54_59),.data_out(wire_d54_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5505461(.data_in(wire_d54_60),.data_out(wire_d54_61),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505462(.data_in(wire_d54_61),.data_out(wire_d54_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505463(.data_in(wire_d54_62),.data_out(wire_d54_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505464(.data_in(wire_d54_63),.data_out(wire_d54_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505465(.data_in(wire_d54_64),.data_out(wire_d54_65),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505466(.data_in(wire_d54_65),.data_out(wire_d54_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505467(.data_in(wire_d54_66),.data_out(wire_d54_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505468(.data_in(wire_d54_67),.data_out(wire_d54_68),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505469(.data_in(wire_d54_68),.data_out(wire_d54_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505470(.data_in(wire_d54_69),.data_out(wire_d54_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5505471(.data_in(wire_d54_70),.data_out(wire_d54_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505472(.data_in(wire_d54_71),.data_out(wire_d54_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505473(.data_in(wire_d54_72),.data_out(wire_d54_73),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5505474(.data_in(wire_d54_73),.data_out(wire_d54_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505475(.data_in(wire_d54_74),.data_out(wire_d54_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505476(.data_in(wire_d54_75),.data_out(wire_d54_76),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505477(.data_in(wire_d54_76),.data_out(wire_d54_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505478(.data_in(wire_d54_77),.data_out(wire_d54_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505479(.data_in(wire_d54_78),.data_out(d_out54),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance560550(.data_in(d_in55),.data_out(wire_d55_0),.clk(clk),.rst(rst));            //channel 56
	register #(.WIDTH(WIDTH)) register_instance560551(.data_in(wire_d55_0),.data_out(wire_d55_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance560552(.data_in(wire_d55_1),.data_out(wire_d55_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance560553(.data_in(wire_d55_2),.data_out(wire_d55_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance560554(.data_in(wire_d55_3),.data_out(wire_d55_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance560555(.data_in(wire_d55_4),.data_out(wire_d55_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance560556(.data_in(wire_d55_5),.data_out(wire_d55_6),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance560557(.data_in(wire_d55_6),.data_out(wire_d55_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance560558(.data_in(wire_d55_7),.data_out(wire_d55_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance560559(.data_in(wire_d55_8),.data_out(wire_d55_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5605510(.data_in(wire_d55_9),.data_out(wire_d55_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5605511(.data_in(wire_d55_10),.data_out(wire_d55_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5605512(.data_in(wire_d55_11),.data_out(wire_d55_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605513(.data_in(wire_d55_12),.data_out(wire_d55_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605514(.data_in(wire_d55_13),.data_out(wire_d55_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5605515(.data_in(wire_d55_14),.data_out(wire_d55_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5605516(.data_in(wire_d55_15),.data_out(wire_d55_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605517(.data_in(wire_d55_16),.data_out(wire_d55_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5605518(.data_in(wire_d55_17),.data_out(wire_d55_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605519(.data_in(wire_d55_18),.data_out(wire_d55_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605520(.data_in(wire_d55_19),.data_out(wire_d55_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5605521(.data_in(wire_d55_20),.data_out(wire_d55_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5605522(.data_in(wire_d55_21),.data_out(wire_d55_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5605523(.data_in(wire_d55_22),.data_out(wire_d55_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5605524(.data_in(wire_d55_23),.data_out(wire_d55_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5605525(.data_in(wire_d55_24),.data_out(wire_d55_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5605526(.data_in(wire_d55_25),.data_out(wire_d55_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5605527(.data_in(wire_d55_26),.data_out(wire_d55_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5605528(.data_in(wire_d55_27),.data_out(wire_d55_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5605529(.data_in(wire_d55_28),.data_out(wire_d55_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5605530(.data_in(wire_d55_29),.data_out(wire_d55_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605531(.data_in(wire_d55_30),.data_out(wire_d55_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5605532(.data_in(wire_d55_31),.data_out(wire_d55_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605533(.data_in(wire_d55_32),.data_out(wire_d55_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605534(.data_in(wire_d55_33),.data_out(wire_d55_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605535(.data_in(wire_d55_34),.data_out(wire_d55_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5605536(.data_in(wire_d55_35),.data_out(wire_d55_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605537(.data_in(wire_d55_36),.data_out(wire_d55_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5605538(.data_in(wire_d55_37),.data_out(wire_d55_38),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5605539(.data_in(wire_d55_38),.data_out(wire_d55_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605540(.data_in(wire_d55_39),.data_out(wire_d55_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605541(.data_in(wire_d55_40),.data_out(wire_d55_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605542(.data_in(wire_d55_41),.data_out(wire_d55_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5605543(.data_in(wire_d55_42),.data_out(wire_d55_43),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605544(.data_in(wire_d55_43),.data_out(wire_d55_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5605545(.data_in(wire_d55_44),.data_out(wire_d55_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5605546(.data_in(wire_d55_45),.data_out(wire_d55_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5605547(.data_in(wire_d55_46),.data_out(wire_d55_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605548(.data_in(wire_d55_47),.data_out(wire_d55_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605549(.data_in(wire_d55_48),.data_out(wire_d55_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5605550(.data_in(wire_d55_49),.data_out(wire_d55_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605551(.data_in(wire_d55_50),.data_out(wire_d55_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605552(.data_in(wire_d55_51),.data_out(wire_d55_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5605553(.data_in(wire_d55_52),.data_out(wire_d55_53),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5605554(.data_in(wire_d55_53),.data_out(wire_d55_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5605555(.data_in(wire_d55_54),.data_out(wire_d55_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5605556(.data_in(wire_d55_55),.data_out(wire_d55_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605557(.data_in(wire_d55_56),.data_out(wire_d55_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5605558(.data_in(wire_d55_57),.data_out(wire_d55_58),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5605559(.data_in(wire_d55_58),.data_out(wire_d55_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5605560(.data_in(wire_d55_59),.data_out(wire_d55_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605561(.data_in(wire_d55_60),.data_out(wire_d55_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5605562(.data_in(wire_d55_61),.data_out(wire_d55_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5605563(.data_in(wire_d55_62),.data_out(wire_d55_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605564(.data_in(wire_d55_63),.data_out(wire_d55_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5605565(.data_in(wire_d55_64),.data_out(wire_d55_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5605566(.data_in(wire_d55_65),.data_out(wire_d55_66),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5605567(.data_in(wire_d55_66),.data_out(wire_d55_67),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5605568(.data_in(wire_d55_67),.data_out(wire_d55_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605569(.data_in(wire_d55_68),.data_out(wire_d55_69),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5605570(.data_in(wire_d55_69),.data_out(wire_d55_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5605571(.data_in(wire_d55_70),.data_out(wire_d55_71),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605572(.data_in(wire_d55_71),.data_out(wire_d55_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605573(.data_in(wire_d55_72),.data_out(wire_d55_73),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5605574(.data_in(wire_d55_73),.data_out(wire_d55_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605575(.data_in(wire_d55_74),.data_out(wire_d55_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5605576(.data_in(wire_d55_75),.data_out(wire_d55_76),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5605577(.data_in(wire_d55_76),.data_out(wire_d55_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605578(.data_in(wire_d55_77),.data_out(wire_d55_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605579(.data_in(wire_d55_78),.data_out(d_out55),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance570560(.data_in(d_in56),.data_out(wire_d56_0),.clk(clk),.rst(rst));            //channel 57
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance570561(.data_in(wire_d56_0),.data_out(wire_d56_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance570562(.data_in(wire_d56_1),.data_out(wire_d56_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance570563(.data_in(wire_d56_2),.data_out(wire_d56_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance570564(.data_in(wire_d56_3),.data_out(wire_d56_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance570565(.data_in(wire_d56_4),.data_out(wire_d56_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance570566(.data_in(wire_d56_5),.data_out(wire_d56_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance570567(.data_in(wire_d56_6),.data_out(wire_d56_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance570568(.data_in(wire_d56_7),.data_out(wire_d56_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance570569(.data_in(wire_d56_8),.data_out(wire_d56_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5705610(.data_in(wire_d56_9),.data_out(wire_d56_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5705611(.data_in(wire_d56_10),.data_out(wire_d56_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5705612(.data_in(wire_d56_11),.data_out(wire_d56_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5705613(.data_in(wire_d56_12),.data_out(wire_d56_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5705614(.data_in(wire_d56_13),.data_out(wire_d56_14),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5705615(.data_in(wire_d56_14),.data_out(wire_d56_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705616(.data_in(wire_d56_15),.data_out(wire_d56_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705617(.data_in(wire_d56_16),.data_out(wire_d56_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705618(.data_in(wire_d56_17),.data_out(wire_d56_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5705619(.data_in(wire_d56_18),.data_out(wire_d56_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5705620(.data_in(wire_d56_19),.data_out(wire_d56_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705621(.data_in(wire_d56_20),.data_out(wire_d56_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5705622(.data_in(wire_d56_21),.data_out(wire_d56_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5705623(.data_in(wire_d56_22),.data_out(wire_d56_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5705624(.data_in(wire_d56_23),.data_out(wire_d56_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705625(.data_in(wire_d56_24),.data_out(wire_d56_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705626(.data_in(wire_d56_25),.data_out(wire_d56_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5705627(.data_in(wire_d56_26),.data_out(wire_d56_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5705628(.data_in(wire_d56_27),.data_out(wire_d56_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705629(.data_in(wire_d56_28),.data_out(wire_d56_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705630(.data_in(wire_d56_29),.data_out(wire_d56_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705631(.data_in(wire_d56_30),.data_out(wire_d56_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705632(.data_in(wire_d56_31),.data_out(wire_d56_32),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5705633(.data_in(wire_d56_32),.data_out(wire_d56_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5705634(.data_in(wire_d56_33),.data_out(wire_d56_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5705635(.data_in(wire_d56_34),.data_out(wire_d56_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5705636(.data_in(wire_d56_35),.data_out(wire_d56_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5705637(.data_in(wire_d56_36),.data_out(wire_d56_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5705638(.data_in(wire_d56_37),.data_out(wire_d56_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705639(.data_in(wire_d56_38),.data_out(wire_d56_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5705640(.data_in(wire_d56_39),.data_out(wire_d56_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5705641(.data_in(wire_d56_40),.data_out(wire_d56_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705642(.data_in(wire_d56_41),.data_out(wire_d56_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5705643(.data_in(wire_d56_42),.data_out(wire_d56_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5705644(.data_in(wire_d56_43),.data_out(wire_d56_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5705645(.data_in(wire_d56_44),.data_out(wire_d56_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5705646(.data_in(wire_d56_45),.data_out(wire_d56_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5705647(.data_in(wire_d56_46),.data_out(wire_d56_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705648(.data_in(wire_d56_47),.data_out(wire_d56_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5705649(.data_in(wire_d56_48),.data_out(wire_d56_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5705650(.data_in(wire_d56_49),.data_out(wire_d56_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705651(.data_in(wire_d56_50),.data_out(wire_d56_51),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5705652(.data_in(wire_d56_51),.data_out(wire_d56_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5705653(.data_in(wire_d56_52),.data_out(wire_d56_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5705654(.data_in(wire_d56_53),.data_out(wire_d56_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5705655(.data_in(wire_d56_54),.data_out(wire_d56_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705656(.data_in(wire_d56_55),.data_out(wire_d56_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5705657(.data_in(wire_d56_56),.data_out(wire_d56_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5705658(.data_in(wire_d56_57),.data_out(wire_d56_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5705659(.data_in(wire_d56_58),.data_out(wire_d56_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5705660(.data_in(wire_d56_59),.data_out(wire_d56_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705661(.data_in(wire_d56_60),.data_out(wire_d56_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5705662(.data_in(wire_d56_61),.data_out(wire_d56_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5705663(.data_in(wire_d56_62),.data_out(wire_d56_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705664(.data_in(wire_d56_63),.data_out(wire_d56_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5705665(.data_in(wire_d56_64),.data_out(wire_d56_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705666(.data_in(wire_d56_65),.data_out(wire_d56_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5705667(.data_in(wire_d56_66),.data_out(wire_d56_67),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5705668(.data_in(wire_d56_67),.data_out(wire_d56_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5705669(.data_in(wire_d56_68),.data_out(wire_d56_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5705670(.data_in(wire_d56_69),.data_out(wire_d56_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5705671(.data_in(wire_d56_70),.data_out(wire_d56_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705672(.data_in(wire_d56_71),.data_out(wire_d56_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5705673(.data_in(wire_d56_72),.data_out(wire_d56_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705674(.data_in(wire_d56_73),.data_out(wire_d56_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5705675(.data_in(wire_d56_74),.data_out(wire_d56_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705676(.data_in(wire_d56_75),.data_out(wire_d56_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705677(.data_in(wire_d56_76),.data_out(wire_d56_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705678(.data_in(wire_d56_77),.data_out(wire_d56_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5705679(.data_in(wire_d56_78),.data_out(d_out56),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance580570(.data_in(d_in57),.data_out(wire_d57_0),.clk(clk),.rst(rst));            //channel 58
	decoder_top #(.WIDTH(WIDTH)) decoder_instance580571(.data_in(wire_d57_0),.data_out(wire_d57_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance580572(.data_in(wire_d57_1),.data_out(wire_d57_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance580573(.data_in(wire_d57_2),.data_out(wire_d57_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance580574(.data_in(wire_d57_3),.data_out(wire_d57_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance580575(.data_in(wire_d57_4),.data_out(wire_d57_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance580576(.data_in(wire_d57_5),.data_out(wire_d57_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance580577(.data_in(wire_d57_6),.data_out(wire_d57_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance580578(.data_in(wire_d57_7),.data_out(wire_d57_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance580579(.data_in(wire_d57_8),.data_out(wire_d57_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805710(.data_in(wire_d57_9),.data_out(wire_d57_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5805711(.data_in(wire_d57_10),.data_out(wire_d57_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5805712(.data_in(wire_d57_11),.data_out(wire_d57_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805713(.data_in(wire_d57_12),.data_out(wire_d57_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5805714(.data_in(wire_d57_13),.data_out(wire_d57_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5805715(.data_in(wire_d57_14),.data_out(wire_d57_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805716(.data_in(wire_d57_15),.data_out(wire_d57_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805717(.data_in(wire_d57_16),.data_out(wire_d57_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5805718(.data_in(wire_d57_17),.data_out(wire_d57_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5805719(.data_in(wire_d57_18),.data_out(wire_d57_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805720(.data_in(wire_d57_19),.data_out(wire_d57_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805721(.data_in(wire_d57_20),.data_out(wire_d57_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5805722(.data_in(wire_d57_21),.data_out(wire_d57_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5805723(.data_in(wire_d57_22),.data_out(wire_d57_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805724(.data_in(wire_d57_23),.data_out(wire_d57_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5805725(.data_in(wire_d57_24),.data_out(wire_d57_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5805726(.data_in(wire_d57_25),.data_out(wire_d57_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805727(.data_in(wire_d57_26),.data_out(wire_d57_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805728(.data_in(wire_d57_27),.data_out(wire_d57_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5805729(.data_in(wire_d57_28),.data_out(wire_d57_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805730(.data_in(wire_d57_29),.data_out(wire_d57_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5805731(.data_in(wire_d57_30),.data_out(wire_d57_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805732(.data_in(wire_d57_31),.data_out(wire_d57_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805733(.data_in(wire_d57_32),.data_out(wire_d57_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805734(.data_in(wire_d57_33),.data_out(wire_d57_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5805735(.data_in(wire_d57_34),.data_out(wire_d57_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5805736(.data_in(wire_d57_35),.data_out(wire_d57_36),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5805737(.data_in(wire_d57_36),.data_out(wire_d57_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805738(.data_in(wire_d57_37),.data_out(wire_d57_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805739(.data_in(wire_d57_38),.data_out(wire_d57_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805740(.data_in(wire_d57_39),.data_out(wire_d57_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805741(.data_in(wire_d57_40),.data_out(wire_d57_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805742(.data_in(wire_d57_41),.data_out(wire_d57_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805743(.data_in(wire_d57_42),.data_out(wire_d57_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5805744(.data_in(wire_d57_43),.data_out(wire_d57_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5805745(.data_in(wire_d57_44),.data_out(wire_d57_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805746(.data_in(wire_d57_45),.data_out(wire_d57_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5805747(.data_in(wire_d57_46),.data_out(wire_d57_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805748(.data_in(wire_d57_47),.data_out(wire_d57_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805749(.data_in(wire_d57_48),.data_out(wire_d57_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5805750(.data_in(wire_d57_49),.data_out(wire_d57_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5805751(.data_in(wire_d57_50),.data_out(wire_d57_51),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5805752(.data_in(wire_d57_51),.data_out(wire_d57_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805753(.data_in(wire_d57_52),.data_out(wire_d57_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5805754(.data_in(wire_d57_53),.data_out(wire_d57_54),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805755(.data_in(wire_d57_54),.data_out(wire_d57_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805756(.data_in(wire_d57_55),.data_out(wire_d57_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5805757(.data_in(wire_d57_56),.data_out(wire_d57_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805758(.data_in(wire_d57_57),.data_out(wire_d57_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805759(.data_in(wire_d57_58),.data_out(wire_d57_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805760(.data_in(wire_d57_59),.data_out(wire_d57_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805761(.data_in(wire_d57_60),.data_out(wire_d57_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5805762(.data_in(wire_d57_61),.data_out(wire_d57_62),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805763(.data_in(wire_d57_62),.data_out(wire_d57_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5805764(.data_in(wire_d57_63),.data_out(wire_d57_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5805765(.data_in(wire_d57_64),.data_out(wire_d57_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5805766(.data_in(wire_d57_65),.data_out(wire_d57_66),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5805767(.data_in(wire_d57_66),.data_out(wire_d57_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5805768(.data_in(wire_d57_67),.data_out(wire_d57_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5805769(.data_in(wire_d57_68),.data_out(wire_d57_69),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5805770(.data_in(wire_d57_69),.data_out(wire_d57_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805771(.data_in(wire_d57_70),.data_out(wire_d57_71),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5805772(.data_in(wire_d57_71),.data_out(wire_d57_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5805773(.data_in(wire_d57_72),.data_out(wire_d57_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805774(.data_in(wire_d57_73),.data_out(wire_d57_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5805775(.data_in(wire_d57_74),.data_out(wire_d57_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5805776(.data_in(wire_d57_75),.data_out(wire_d57_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805777(.data_in(wire_d57_76),.data_out(wire_d57_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805778(.data_in(wire_d57_77),.data_out(wire_d57_78),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805779(.data_in(wire_d57_78),.data_out(d_out57),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance590580(.data_in(d_in58),.data_out(wire_d58_0),.clk(clk),.rst(rst));            //channel 59
	large_mux #(.WIDTH(WIDTH)) large_mux_instance590581(.data_in(wire_d58_0),.data_out(wire_d58_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance590582(.data_in(wire_d58_1),.data_out(wire_d58_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance590583(.data_in(wire_d58_2),.data_out(wire_d58_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance590584(.data_in(wire_d58_3),.data_out(wire_d58_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance590585(.data_in(wire_d58_4),.data_out(wire_d58_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance590586(.data_in(wire_d58_5),.data_out(wire_d58_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance590587(.data_in(wire_d58_6),.data_out(wire_d58_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance590588(.data_in(wire_d58_7),.data_out(wire_d58_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance590589(.data_in(wire_d58_8),.data_out(wire_d58_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5905810(.data_in(wire_d58_9),.data_out(wire_d58_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5905811(.data_in(wire_d58_10),.data_out(wire_d58_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5905812(.data_in(wire_d58_11),.data_out(wire_d58_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905813(.data_in(wire_d58_12),.data_out(wire_d58_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5905814(.data_in(wire_d58_13),.data_out(wire_d58_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5905815(.data_in(wire_d58_14),.data_out(wire_d58_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5905816(.data_in(wire_d58_15),.data_out(wire_d58_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5905817(.data_in(wire_d58_16),.data_out(wire_d58_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905818(.data_in(wire_d58_17),.data_out(wire_d58_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905819(.data_in(wire_d58_18),.data_out(wire_d58_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5905820(.data_in(wire_d58_19),.data_out(wire_d58_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5905821(.data_in(wire_d58_20),.data_out(wire_d58_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5905822(.data_in(wire_d58_21),.data_out(wire_d58_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5905823(.data_in(wire_d58_22),.data_out(wire_d58_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905824(.data_in(wire_d58_23),.data_out(wire_d58_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5905825(.data_in(wire_d58_24),.data_out(wire_d58_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5905826(.data_in(wire_d58_25),.data_out(wire_d58_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5905827(.data_in(wire_d58_26),.data_out(wire_d58_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905828(.data_in(wire_d58_27),.data_out(wire_d58_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5905829(.data_in(wire_d58_28),.data_out(wire_d58_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905830(.data_in(wire_d58_29),.data_out(wire_d58_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5905831(.data_in(wire_d58_30),.data_out(wire_d58_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905832(.data_in(wire_d58_31),.data_out(wire_d58_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5905833(.data_in(wire_d58_32),.data_out(wire_d58_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5905834(.data_in(wire_d58_33),.data_out(wire_d58_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5905835(.data_in(wire_d58_34),.data_out(wire_d58_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5905836(.data_in(wire_d58_35),.data_out(wire_d58_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5905837(.data_in(wire_d58_36),.data_out(wire_d58_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5905838(.data_in(wire_d58_37),.data_out(wire_d58_38),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5905839(.data_in(wire_d58_38),.data_out(wire_d58_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5905840(.data_in(wire_d58_39),.data_out(wire_d58_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5905841(.data_in(wire_d58_40),.data_out(wire_d58_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5905842(.data_in(wire_d58_41),.data_out(wire_d58_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5905843(.data_in(wire_d58_42),.data_out(wire_d58_43),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5905844(.data_in(wire_d58_43),.data_out(wire_d58_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5905845(.data_in(wire_d58_44),.data_out(wire_d58_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5905846(.data_in(wire_d58_45),.data_out(wire_d58_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5905847(.data_in(wire_d58_46),.data_out(wire_d58_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5905848(.data_in(wire_d58_47),.data_out(wire_d58_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5905849(.data_in(wire_d58_48),.data_out(wire_d58_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5905850(.data_in(wire_d58_49),.data_out(wire_d58_50),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5905851(.data_in(wire_d58_50),.data_out(wire_d58_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5905852(.data_in(wire_d58_51),.data_out(wire_d58_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905853(.data_in(wire_d58_52),.data_out(wire_d58_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5905854(.data_in(wire_d58_53),.data_out(wire_d58_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5905855(.data_in(wire_d58_54),.data_out(wire_d58_55),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5905856(.data_in(wire_d58_55),.data_out(wire_d58_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905857(.data_in(wire_d58_56),.data_out(wire_d58_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5905858(.data_in(wire_d58_57),.data_out(wire_d58_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5905859(.data_in(wire_d58_58),.data_out(wire_d58_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905860(.data_in(wire_d58_59),.data_out(wire_d58_60),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905861(.data_in(wire_d58_60),.data_out(wire_d58_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5905862(.data_in(wire_d58_61),.data_out(wire_d58_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905863(.data_in(wire_d58_62),.data_out(wire_d58_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5905864(.data_in(wire_d58_63),.data_out(wire_d58_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5905865(.data_in(wire_d58_64),.data_out(wire_d58_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905866(.data_in(wire_d58_65),.data_out(wire_d58_66),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905867(.data_in(wire_d58_66),.data_out(wire_d58_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5905868(.data_in(wire_d58_67),.data_out(wire_d58_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5905869(.data_in(wire_d58_68),.data_out(wire_d58_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5905870(.data_in(wire_d58_69),.data_out(wire_d58_70),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5905871(.data_in(wire_d58_70),.data_out(wire_d58_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5905872(.data_in(wire_d58_71),.data_out(wire_d58_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5905873(.data_in(wire_d58_72),.data_out(wire_d58_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905874(.data_in(wire_d58_73),.data_out(wire_d58_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5905875(.data_in(wire_d58_74),.data_out(wire_d58_75),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905876(.data_in(wire_d58_75),.data_out(wire_d58_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5905877(.data_in(wire_d58_76),.data_out(wire_d58_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905878(.data_in(wire_d58_77),.data_out(wire_d58_78),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905879(.data_in(wire_d58_78),.data_out(d_out58),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance600590(.data_in(d_in59),.data_out(wire_d59_0),.clk(clk),.rst(rst));            //channel 60
	decoder_top #(.WIDTH(WIDTH)) decoder_instance600591(.data_in(wire_d59_0),.data_out(wire_d59_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance600592(.data_in(wire_d59_1),.data_out(wire_d59_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance600593(.data_in(wire_d59_2),.data_out(wire_d59_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance600594(.data_in(wire_d59_3),.data_out(wire_d59_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance600595(.data_in(wire_d59_4),.data_out(wire_d59_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance600596(.data_in(wire_d59_5),.data_out(wire_d59_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance600597(.data_in(wire_d59_6),.data_out(wire_d59_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance600598(.data_in(wire_d59_7),.data_out(wire_d59_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance600599(.data_in(wire_d59_8),.data_out(wire_d59_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6005910(.data_in(wire_d59_9),.data_out(wire_d59_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005911(.data_in(wire_d59_10),.data_out(wire_d59_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6005912(.data_in(wire_d59_11),.data_out(wire_d59_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005913(.data_in(wire_d59_12),.data_out(wire_d59_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6005914(.data_in(wire_d59_13),.data_out(wire_d59_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005915(.data_in(wire_d59_14),.data_out(wire_d59_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6005916(.data_in(wire_d59_15),.data_out(wire_d59_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005917(.data_in(wire_d59_16),.data_out(wire_d59_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6005918(.data_in(wire_d59_17),.data_out(wire_d59_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005919(.data_in(wire_d59_18),.data_out(wire_d59_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005920(.data_in(wire_d59_19),.data_out(wire_d59_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6005921(.data_in(wire_d59_20),.data_out(wire_d59_21),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005922(.data_in(wire_d59_21),.data_out(wire_d59_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005923(.data_in(wire_d59_22),.data_out(wire_d59_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005924(.data_in(wire_d59_23),.data_out(wire_d59_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6005925(.data_in(wire_d59_24),.data_out(wire_d59_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005926(.data_in(wire_d59_25),.data_out(wire_d59_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005927(.data_in(wire_d59_26),.data_out(wire_d59_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6005928(.data_in(wire_d59_27),.data_out(wire_d59_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005929(.data_in(wire_d59_28),.data_out(wire_d59_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6005930(.data_in(wire_d59_29),.data_out(wire_d59_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005931(.data_in(wire_d59_30),.data_out(wire_d59_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6005932(.data_in(wire_d59_31),.data_out(wire_d59_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6005933(.data_in(wire_d59_32),.data_out(wire_d59_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6005934(.data_in(wire_d59_33),.data_out(wire_d59_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005935(.data_in(wire_d59_34),.data_out(wire_d59_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005936(.data_in(wire_d59_35),.data_out(wire_d59_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005937(.data_in(wire_d59_36),.data_out(wire_d59_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005938(.data_in(wire_d59_37),.data_out(wire_d59_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6005939(.data_in(wire_d59_38),.data_out(wire_d59_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005940(.data_in(wire_d59_39),.data_out(wire_d59_40),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6005941(.data_in(wire_d59_40),.data_out(wire_d59_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005942(.data_in(wire_d59_41),.data_out(wire_d59_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6005943(.data_in(wire_d59_42),.data_out(wire_d59_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6005944(.data_in(wire_d59_43),.data_out(wire_d59_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6005945(.data_in(wire_d59_44),.data_out(wire_d59_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6005946(.data_in(wire_d59_45),.data_out(wire_d59_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6005947(.data_in(wire_d59_46),.data_out(wire_d59_47),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005948(.data_in(wire_d59_47),.data_out(wire_d59_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005949(.data_in(wire_d59_48),.data_out(wire_d59_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6005950(.data_in(wire_d59_49),.data_out(wire_d59_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005951(.data_in(wire_d59_50),.data_out(wire_d59_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6005952(.data_in(wire_d59_51),.data_out(wire_d59_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005953(.data_in(wire_d59_52),.data_out(wire_d59_53),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6005954(.data_in(wire_d59_53),.data_out(wire_d59_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6005955(.data_in(wire_d59_54),.data_out(wire_d59_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005956(.data_in(wire_d59_55),.data_out(wire_d59_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005957(.data_in(wire_d59_56),.data_out(wire_d59_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005958(.data_in(wire_d59_57),.data_out(wire_d59_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6005959(.data_in(wire_d59_58),.data_out(wire_d59_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6005960(.data_in(wire_d59_59),.data_out(wire_d59_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6005961(.data_in(wire_d59_60),.data_out(wire_d59_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6005962(.data_in(wire_d59_61),.data_out(wire_d59_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6005963(.data_in(wire_d59_62),.data_out(wire_d59_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6005964(.data_in(wire_d59_63),.data_out(wire_d59_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005965(.data_in(wire_d59_64),.data_out(wire_d59_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005966(.data_in(wire_d59_65),.data_out(wire_d59_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005967(.data_in(wire_d59_66),.data_out(wire_d59_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6005968(.data_in(wire_d59_67),.data_out(wire_d59_68),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6005969(.data_in(wire_d59_68),.data_out(wire_d59_69),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6005970(.data_in(wire_d59_69),.data_out(wire_d59_70),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6005971(.data_in(wire_d59_70),.data_out(wire_d59_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005972(.data_in(wire_d59_71),.data_out(wire_d59_72),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6005973(.data_in(wire_d59_72),.data_out(wire_d59_73),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6005974(.data_in(wire_d59_73),.data_out(wire_d59_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005975(.data_in(wire_d59_74),.data_out(wire_d59_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005976(.data_in(wire_d59_75),.data_out(wire_d59_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005977(.data_in(wire_d59_76),.data_out(wire_d59_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005978(.data_in(wire_d59_77),.data_out(wire_d59_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6005979(.data_in(wire_d59_78),.data_out(d_out59),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance610600(.data_in(d_in60),.data_out(wire_d60_0),.clk(clk),.rst(rst));            //channel 61
	large_mux #(.WIDTH(WIDTH)) large_mux_instance610601(.data_in(wire_d60_0),.data_out(wire_d60_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance610602(.data_in(wire_d60_1),.data_out(wire_d60_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance610603(.data_in(wire_d60_2),.data_out(wire_d60_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance610604(.data_in(wire_d60_3),.data_out(wire_d60_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance610605(.data_in(wire_d60_4),.data_out(wire_d60_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance610606(.data_in(wire_d60_5),.data_out(wire_d60_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance610607(.data_in(wire_d60_6),.data_out(wire_d60_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance610608(.data_in(wire_d60_7),.data_out(wire_d60_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance610609(.data_in(wire_d60_8),.data_out(wire_d60_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6106010(.data_in(wire_d60_9),.data_out(wire_d60_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6106011(.data_in(wire_d60_10),.data_out(wire_d60_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6106012(.data_in(wire_d60_11),.data_out(wire_d60_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6106013(.data_in(wire_d60_12),.data_out(wire_d60_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6106014(.data_in(wire_d60_13),.data_out(wire_d60_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6106015(.data_in(wire_d60_14),.data_out(wire_d60_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6106016(.data_in(wire_d60_15),.data_out(wire_d60_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6106017(.data_in(wire_d60_16),.data_out(wire_d60_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6106018(.data_in(wire_d60_17),.data_out(wire_d60_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6106019(.data_in(wire_d60_18),.data_out(wire_d60_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6106020(.data_in(wire_d60_19),.data_out(wire_d60_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6106021(.data_in(wire_d60_20),.data_out(wire_d60_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6106022(.data_in(wire_d60_21),.data_out(wire_d60_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6106023(.data_in(wire_d60_22),.data_out(wire_d60_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6106024(.data_in(wire_d60_23),.data_out(wire_d60_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6106025(.data_in(wire_d60_24),.data_out(wire_d60_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6106026(.data_in(wire_d60_25),.data_out(wire_d60_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6106027(.data_in(wire_d60_26),.data_out(wire_d60_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6106028(.data_in(wire_d60_27),.data_out(wire_d60_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6106029(.data_in(wire_d60_28),.data_out(wire_d60_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6106030(.data_in(wire_d60_29),.data_out(wire_d60_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6106031(.data_in(wire_d60_30),.data_out(wire_d60_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6106032(.data_in(wire_d60_31),.data_out(wire_d60_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6106033(.data_in(wire_d60_32),.data_out(wire_d60_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6106034(.data_in(wire_d60_33),.data_out(wire_d60_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6106035(.data_in(wire_d60_34),.data_out(wire_d60_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6106036(.data_in(wire_d60_35),.data_out(wire_d60_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6106037(.data_in(wire_d60_36),.data_out(wire_d60_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6106038(.data_in(wire_d60_37),.data_out(wire_d60_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6106039(.data_in(wire_d60_38),.data_out(wire_d60_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6106040(.data_in(wire_d60_39),.data_out(wire_d60_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6106041(.data_in(wire_d60_40),.data_out(wire_d60_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6106042(.data_in(wire_d60_41),.data_out(wire_d60_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6106043(.data_in(wire_d60_42),.data_out(wire_d60_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6106044(.data_in(wire_d60_43),.data_out(wire_d60_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6106045(.data_in(wire_d60_44),.data_out(wire_d60_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6106046(.data_in(wire_d60_45),.data_out(wire_d60_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6106047(.data_in(wire_d60_46),.data_out(wire_d60_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6106048(.data_in(wire_d60_47),.data_out(wire_d60_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6106049(.data_in(wire_d60_48),.data_out(wire_d60_49),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6106050(.data_in(wire_d60_49),.data_out(wire_d60_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6106051(.data_in(wire_d60_50),.data_out(wire_d60_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6106052(.data_in(wire_d60_51),.data_out(wire_d60_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6106053(.data_in(wire_d60_52),.data_out(wire_d60_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6106054(.data_in(wire_d60_53),.data_out(wire_d60_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6106055(.data_in(wire_d60_54),.data_out(wire_d60_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6106056(.data_in(wire_d60_55),.data_out(wire_d60_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6106057(.data_in(wire_d60_56),.data_out(wire_d60_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6106058(.data_in(wire_d60_57),.data_out(wire_d60_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6106059(.data_in(wire_d60_58),.data_out(wire_d60_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6106060(.data_in(wire_d60_59),.data_out(wire_d60_60),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6106061(.data_in(wire_d60_60),.data_out(wire_d60_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6106062(.data_in(wire_d60_61),.data_out(wire_d60_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6106063(.data_in(wire_d60_62),.data_out(wire_d60_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6106064(.data_in(wire_d60_63),.data_out(wire_d60_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6106065(.data_in(wire_d60_64),.data_out(wire_d60_65),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6106066(.data_in(wire_d60_65),.data_out(wire_d60_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6106067(.data_in(wire_d60_66),.data_out(wire_d60_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6106068(.data_in(wire_d60_67),.data_out(wire_d60_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6106069(.data_in(wire_d60_68),.data_out(wire_d60_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6106070(.data_in(wire_d60_69),.data_out(wire_d60_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6106071(.data_in(wire_d60_70),.data_out(wire_d60_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6106072(.data_in(wire_d60_71),.data_out(wire_d60_72),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6106073(.data_in(wire_d60_72),.data_out(wire_d60_73),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6106074(.data_in(wire_d60_73),.data_out(wire_d60_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6106075(.data_in(wire_d60_74),.data_out(wire_d60_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6106076(.data_in(wire_d60_75),.data_out(wire_d60_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6106077(.data_in(wire_d60_76),.data_out(wire_d60_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6106078(.data_in(wire_d60_77),.data_out(wire_d60_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6106079(.data_in(wire_d60_78),.data_out(d_out60),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance620610(.data_in(d_in61),.data_out(wire_d61_0),.clk(clk),.rst(rst));            //channel 62
	decoder_top #(.WIDTH(WIDTH)) decoder_instance620611(.data_in(wire_d61_0),.data_out(wire_d61_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance620612(.data_in(wire_d61_1),.data_out(wire_d61_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance620613(.data_in(wire_d61_2),.data_out(wire_d61_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance620614(.data_in(wire_d61_3),.data_out(wire_d61_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance620615(.data_in(wire_d61_4),.data_out(wire_d61_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance620616(.data_in(wire_d61_5),.data_out(wire_d61_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance620617(.data_in(wire_d61_6),.data_out(wire_d61_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance620618(.data_in(wire_d61_7),.data_out(wire_d61_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance620619(.data_in(wire_d61_8),.data_out(wire_d61_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6206110(.data_in(wire_d61_9),.data_out(wire_d61_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6206111(.data_in(wire_d61_10),.data_out(wire_d61_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6206112(.data_in(wire_d61_11),.data_out(wire_d61_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6206113(.data_in(wire_d61_12),.data_out(wire_d61_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6206114(.data_in(wire_d61_13),.data_out(wire_d61_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6206115(.data_in(wire_d61_14),.data_out(wire_d61_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6206116(.data_in(wire_d61_15),.data_out(wire_d61_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6206117(.data_in(wire_d61_16),.data_out(wire_d61_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6206118(.data_in(wire_d61_17),.data_out(wire_d61_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6206119(.data_in(wire_d61_18),.data_out(wire_d61_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6206120(.data_in(wire_d61_19),.data_out(wire_d61_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6206121(.data_in(wire_d61_20),.data_out(wire_d61_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6206122(.data_in(wire_d61_21),.data_out(wire_d61_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6206123(.data_in(wire_d61_22),.data_out(wire_d61_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6206124(.data_in(wire_d61_23),.data_out(wire_d61_24),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6206125(.data_in(wire_d61_24),.data_out(wire_d61_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6206126(.data_in(wire_d61_25),.data_out(wire_d61_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6206127(.data_in(wire_d61_26),.data_out(wire_d61_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6206128(.data_in(wire_d61_27),.data_out(wire_d61_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6206129(.data_in(wire_d61_28),.data_out(wire_d61_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6206130(.data_in(wire_d61_29),.data_out(wire_d61_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6206131(.data_in(wire_d61_30),.data_out(wire_d61_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6206132(.data_in(wire_d61_31),.data_out(wire_d61_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6206133(.data_in(wire_d61_32),.data_out(wire_d61_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6206134(.data_in(wire_d61_33),.data_out(wire_d61_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6206135(.data_in(wire_d61_34),.data_out(wire_d61_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6206136(.data_in(wire_d61_35),.data_out(wire_d61_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6206137(.data_in(wire_d61_36),.data_out(wire_d61_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6206138(.data_in(wire_d61_37),.data_out(wire_d61_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6206139(.data_in(wire_d61_38),.data_out(wire_d61_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6206140(.data_in(wire_d61_39),.data_out(wire_d61_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6206141(.data_in(wire_d61_40),.data_out(wire_d61_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6206142(.data_in(wire_d61_41),.data_out(wire_d61_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6206143(.data_in(wire_d61_42),.data_out(wire_d61_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6206144(.data_in(wire_d61_43),.data_out(wire_d61_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6206145(.data_in(wire_d61_44),.data_out(wire_d61_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6206146(.data_in(wire_d61_45),.data_out(wire_d61_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6206147(.data_in(wire_d61_46),.data_out(wire_d61_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6206148(.data_in(wire_d61_47),.data_out(wire_d61_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6206149(.data_in(wire_d61_48),.data_out(wire_d61_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6206150(.data_in(wire_d61_49),.data_out(wire_d61_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6206151(.data_in(wire_d61_50),.data_out(wire_d61_51),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6206152(.data_in(wire_d61_51),.data_out(wire_d61_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6206153(.data_in(wire_d61_52),.data_out(wire_d61_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6206154(.data_in(wire_d61_53),.data_out(wire_d61_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6206155(.data_in(wire_d61_54),.data_out(wire_d61_55),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6206156(.data_in(wire_d61_55),.data_out(wire_d61_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6206157(.data_in(wire_d61_56),.data_out(wire_d61_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6206158(.data_in(wire_d61_57),.data_out(wire_d61_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6206159(.data_in(wire_d61_58),.data_out(wire_d61_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6206160(.data_in(wire_d61_59),.data_out(wire_d61_60),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6206161(.data_in(wire_d61_60),.data_out(wire_d61_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6206162(.data_in(wire_d61_61),.data_out(wire_d61_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6206163(.data_in(wire_d61_62),.data_out(wire_d61_63),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6206164(.data_in(wire_d61_63),.data_out(wire_d61_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6206165(.data_in(wire_d61_64),.data_out(wire_d61_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6206166(.data_in(wire_d61_65),.data_out(wire_d61_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6206167(.data_in(wire_d61_66),.data_out(wire_d61_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6206168(.data_in(wire_d61_67),.data_out(wire_d61_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6206169(.data_in(wire_d61_68),.data_out(wire_d61_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6206170(.data_in(wire_d61_69),.data_out(wire_d61_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6206171(.data_in(wire_d61_70),.data_out(wire_d61_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6206172(.data_in(wire_d61_71),.data_out(wire_d61_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6206173(.data_in(wire_d61_72),.data_out(wire_d61_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6206174(.data_in(wire_d61_73),.data_out(wire_d61_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6206175(.data_in(wire_d61_74),.data_out(wire_d61_75),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6206176(.data_in(wire_d61_75),.data_out(wire_d61_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6206177(.data_in(wire_d61_76),.data_out(wire_d61_77),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6206178(.data_in(wire_d61_77),.data_out(wire_d61_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6206179(.data_in(wire_d61_78),.data_out(d_out61),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance630620(.data_in(d_in62),.data_out(wire_d62_0),.clk(clk),.rst(rst));            //channel 63
	large_mux #(.WIDTH(WIDTH)) large_mux_instance630621(.data_in(wire_d62_0),.data_out(wire_d62_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance630622(.data_in(wire_d62_1),.data_out(wire_d62_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance630623(.data_in(wire_d62_2),.data_out(wire_d62_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance630624(.data_in(wire_d62_3),.data_out(wire_d62_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance630625(.data_in(wire_d62_4),.data_out(wire_d62_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance630626(.data_in(wire_d62_5),.data_out(wire_d62_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance630627(.data_in(wire_d62_6),.data_out(wire_d62_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance630628(.data_in(wire_d62_7),.data_out(wire_d62_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance630629(.data_in(wire_d62_8),.data_out(wire_d62_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6306210(.data_in(wire_d62_9),.data_out(wire_d62_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6306211(.data_in(wire_d62_10),.data_out(wire_d62_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6306212(.data_in(wire_d62_11),.data_out(wire_d62_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6306213(.data_in(wire_d62_12),.data_out(wire_d62_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6306214(.data_in(wire_d62_13),.data_out(wire_d62_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6306215(.data_in(wire_d62_14),.data_out(wire_d62_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6306216(.data_in(wire_d62_15),.data_out(wire_d62_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6306217(.data_in(wire_d62_16),.data_out(wire_d62_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6306218(.data_in(wire_d62_17),.data_out(wire_d62_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6306219(.data_in(wire_d62_18),.data_out(wire_d62_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6306220(.data_in(wire_d62_19),.data_out(wire_d62_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6306221(.data_in(wire_d62_20),.data_out(wire_d62_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6306222(.data_in(wire_d62_21),.data_out(wire_d62_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6306223(.data_in(wire_d62_22),.data_out(wire_d62_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6306224(.data_in(wire_d62_23),.data_out(wire_d62_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6306225(.data_in(wire_d62_24),.data_out(wire_d62_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6306226(.data_in(wire_d62_25),.data_out(wire_d62_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6306227(.data_in(wire_d62_26),.data_out(wire_d62_27),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6306228(.data_in(wire_d62_27),.data_out(wire_d62_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6306229(.data_in(wire_d62_28),.data_out(wire_d62_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6306230(.data_in(wire_d62_29),.data_out(wire_d62_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6306231(.data_in(wire_d62_30),.data_out(wire_d62_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6306232(.data_in(wire_d62_31),.data_out(wire_d62_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6306233(.data_in(wire_d62_32),.data_out(wire_d62_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6306234(.data_in(wire_d62_33),.data_out(wire_d62_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6306235(.data_in(wire_d62_34),.data_out(wire_d62_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6306236(.data_in(wire_d62_35),.data_out(wire_d62_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6306237(.data_in(wire_d62_36),.data_out(wire_d62_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6306238(.data_in(wire_d62_37),.data_out(wire_d62_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6306239(.data_in(wire_d62_38),.data_out(wire_d62_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6306240(.data_in(wire_d62_39),.data_out(wire_d62_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6306241(.data_in(wire_d62_40),.data_out(wire_d62_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6306242(.data_in(wire_d62_41),.data_out(wire_d62_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6306243(.data_in(wire_d62_42),.data_out(wire_d62_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6306244(.data_in(wire_d62_43),.data_out(wire_d62_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6306245(.data_in(wire_d62_44),.data_out(wire_d62_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6306246(.data_in(wire_d62_45),.data_out(wire_d62_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6306247(.data_in(wire_d62_46),.data_out(wire_d62_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6306248(.data_in(wire_d62_47),.data_out(wire_d62_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6306249(.data_in(wire_d62_48),.data_out(wire_d62_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6306250(.data_in(wire_d62_49),.data_out(wire_d62_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6306251(.data_in(wire_d62_50),.data_out(wire_d62_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6306252(.data_in(wire_d62_51),.data_out(wire_d62_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6306253(.data_in(wire_d62_52),.data_out(wire_d62_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6306254(.data_in(wire_d62_53),.data_out(wire_d62_54),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6306255(.data_in(wire_d62_54),.data_out(wire_d62_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6306256(.data_in(wire_d62_55),.data_out(wire_d62_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6306257(.data_in(wire_d62_56),.data_out(wire_d62_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6306258(.data_in(wire_d62_57),.data_out(wire_d62_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6306259(.data_in(wire_d62_58),.data_out(wire_d62_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6306260(.data_in(wire_d62_59),.data_out(wire_d62_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6306261(.data_in(wire_d62_60),.data_out(wire_d62_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6306262(.data_in(wire_d62_61),.data_out(wire_d62_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6306263(.data_in(wire_d62_62),.data_out(wire_d62_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6306264(.data_in(wire_d62_63),.data_out(wire_d62_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6306265(.data_in(wire_d62_64),.data_out(wire_d62_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6306266(.data_in(wire_d62_65),.data_out(wire_d62_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6306267(.data_in(wire_d62_66),.data_out(wire_d62_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6306268(.data_in(wire_d62_67),.data_out(wire_d62_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6306269(.data_in(wire_d62_68),.data_out(wire_d62_69),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6306270(.data_in(wire_d62_69),.data_out(wire_d62_70),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6306271(.data_in(wire_d62_70),.data_out(wire_d62_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6306272(.data_in(wire_d62_71),.data_out(wire_d62_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6306273(.data_in(wire_d62_72),.data_out(wire_d62_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6306274(.data_in(wire_d62_73),.data_out(wire_d62_74),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6306275(.data_in(wire_d62_74),.data_out(wire_d62_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6306276(.data_in(wire_d62_75),.data_out(wire_d62_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6306277(.data_in(wire_d62_76),.data_out(wire_d62_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6306278(.data_in(wire_d62_77),.data_out(wire_d62_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6306279(.data_in(wire_d62_78),.data_out(d_out62),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance640630(.data_in(d_in63),.data_out(wire_d63_0),.clk(clk),.rst(rst));            //channel 64
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance640631(.data_in(wire_d63_0),.data_out(wire_d63_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance640632(.data_in(wire_d63_1),.data_out(wire_d63_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance640633(.data_in(wire_d63_2),.data_out(wire_d63_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance640634(.data_in(wire_d63_3),.data_out(wire_d63_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance640635(.data_in(wire_d63_4),.data_out(wire_d63_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance640636(.data_in(wire_d63_5),.data_out(wire_d63_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance640637(.data_in(wire_d63_6),.data_out(wire_d63_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance640638(.data_in(wire_d63_7),.data_out(wire_d63_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance640639(.data_in(wire_d63_8),.data_out(wire_d63_9),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6406310(.data_in(wire_d63_9),.data_out(wire_d63_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6406311(.data_in(wire_d63_10),.data_out(wire_d63_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6406312(.data_in(wire_d63_11),.data_out(wire_d63_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6406313(.data_in(wire_d63_12),.data_out(wire_d63_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6406314(.data_in(wire_d63_13),.data_out(wire_d63_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6406315(.data_in(wire_d63_14),.data_out(wire_d63_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6406316(.data_in(wire_d63_15),.data_out(wire_d63_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6406317(.data_in(wire_d63_16),.data_out(wire_d63_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6406318(.data_in(wire_d63_17),.data_out(wire_d63_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6406319(.data_in(wire_d63_18),.data_out(wire_d63_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6406320(.data_in(wire_d63_19),.data_out(wire_d63_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6406321(.data_in(wire_d63_20),.data_out(wire_d63_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6406322(.data_in(wire_d63_21),.data_out(wire_d63_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6406323(.data_in(wire_d63_22),.data_out(wire_d63_23),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6406324(.data_in(wire_d63_23),.data_out(wire_d63_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6406325(.data_in(wire_d63_24),.data_out(wire_d63_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6406326(.data_in(wire_d63_25),.data_out(wire_d63_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6406327(.data_in(wire_d63_26),.data_out(wire_d63_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6406328(.data_in(wire_d63_27),.data_out(wire_d63_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6406329(.data_in(wire_d63_28),.data_out(wire_d63_29),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6406330(.data_in(wire_d63_29),.data_out(wire_d63_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6406331(.data_in(wire_d63_30),.data_out(wire_d63_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6406332(.data_in(wire_d63_31),.data_out(wire_d63_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6406333(.data_in(wire_d63_32),.data_out(wire_d63_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6406334(.data_in(wire_d63_33),.data_out(wire_d63_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6406335(.data_in(wire_d63_34),.data_out(wire_d63_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6406336(.data_in(wire_d63_35),.data_out(wire_d63_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6406337(.data_in(wire_d63_36),.data_out(wire_d63_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6406338(.data_in(wire_d63_37),.data_out(wire_d63_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6406339(.data_in(wire_d63_38),.data_out(wire_d63_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6406340(.data_in(wire_d63_39),.data_out(wire_d63_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6406341(.data_in(wire_d63_40),.data_out(wire_d63_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6406342(.data_in(wire_d63_41),.data_out(wire_d63_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6406343(.data_in(wire_d63_42),.data_out(wire_d63_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6406344(.data_in(wire_d63_43),.data_out(wire_d63_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6406345(.data_in(wire_d63_44),.data_out(wire_d63_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6406346(.data_in(wire_d63_45),.data_out(wire_d63_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6406347(.data_in(wire_d63_46),.data_out(wire_d63_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6406348(.data_in(wire_d63_47),.data_out(wire_d63_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6406349(.data_in(wire_d63_48),.data_out(wire_d63_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6406350(.data_in(wire_d63_49),.data_out(wire_d63_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6406351(.data_in(wire_d63_50),.data_out(wire_d63_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6406352(.data_in(wire_d63_51),.data_out(wire_d63_52),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6406353(.data_in(wire_d63_52),.data_out(wire_d63_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6406354(.data_in(wire_d63_53),.data_out(wire_d63_54),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6406355(.data_in(wire_d63_54),.data_out(wire_d63_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6406356(.data_in(wire_d63_55),.data_out(wire_d63_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6406357(.data_in(wire_d63_56),.data_out(wire_d63_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6406358(.data_in(wire_d63_57),.data_out(wire_d63_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6406359(.data_in(wire_d63_58),.data_out(wire_d63_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6406360(.data_in(wire_d63_59),.data_out(wire_d63_60),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6406361(.data_in(wire_d63_60),.data_out(wire_d63_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6406362(.data_in(wire_d63_61),.data_out(wire_d63_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6406363(.data_in(wire_d63_62),.data_out(wire_d63_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6406364(.data_in(wire_d63_63),.data_out(wire_d63_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6406365(.data_in(wire_d63_64),.data_out(wire_d63_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6406366(.data_in(wire_d63_65),.data_out(wire_d63_66),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6406367(.data_in(wire_d63_66),.data_out(wire_d63_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6406368(.data_in(wire_d63_67),.data_out(wire_d63_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6406369(.data_in(wire_d63_68),.data_out(wire_d63_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6406370(.data_in(wire_d63_69),.data_out(wire_d63_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6406371(.data_in(wire_d63_70),.data_out(wire_d63_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6406372(.data_in(wire_d63_71),.data_out(wire_d63_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6406373(.data_in(wire_d63_72),.data_out(wire_d63_73),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6406374(.data_in(wire_d63_73),.data_out(wire_d63_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6406375(.data_in(wire_d63_74),.data_out(wire_d63_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6406376(.data_in(wire_d63_75),.data_out(wire_d63_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6406377(.data_in(wire_d63_76),.data_out(wire_d63_77),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6406378(.data_in(wire_d63_77),.data_out(wire_d63_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6406379(.data_in(wire_d63_78),.data_out(d_out63),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance650640(.data_in(d_in64),.data_out(wire_d64_0),.clk(clk),.rst(rst));            //channel 65
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance650641(.data_in(wire_d64_0),.data_out(wire_d64_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance650642(.data_in(wire_d64_1),.data_out(wire_d64_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance650643(.data_in(wire_d64_2),.data_out(wire_d64_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance650644(.data_in(wire_d64_3),.data_out(wire_d64_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance650645(.data_in(wire_d64_4),.data_out(wire_d64_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance650646(.data_in(wire_d64_5),.data_out(wire_d64_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance650647(.data_in(wire_d64_6),.data_out(wire_d64_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance650648(.data_in(wire_d64_7),.data_out(wire_d64_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance650649(.data_in(wire_d64_8),.data_out(wire_d64_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6506410(.data_in(wire_d64_9),.data_out(wire_d64_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6506411(.data_in(wire_d64_10),.data_out(wire_d64_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6506412(.data_in(wire_d64_11),.data_out(wire_d64_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6506413(.data_in(wire_d64_12),.data_out(wire_d64_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6506414(.data_in(wire_d64_13),.data_out(wire_d64_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6506415(.data_in(wire_d64_14),.data_out(wire_d64_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6506416(.data_in(wire_d64_15),.data_out(wire_d64_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6506417(.data_in(wire_d64_16),.data_out(wire_d64_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6506418(.data_in(wire_d64_17),.data_out(wire_d64_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6506419(.data_in(wire_d64_18),.data_out(wire_d64_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6506420(.data_in(wire_d64_19),.data_out(wire_d64_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6506421(.data_in(wire_d64_20),.data_out(wire_d64_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6506422(.data_in(wire_d64_21),.data_out(wire_d64_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6506423(.data_in(wire_d64_22),.data_out(wire_d64_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6506424(.data_in(wire_d64_23),.data_out(wire_d64_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6506425(.data_in(wire_d64_24),.data_out(wire_d64_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6506426(.data_in(wire_d64_25),.data_out(wire_d64_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6506427(.data_in(wire_d64_26),.data_out(wire_d64_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6506428(.data_in(wire_d64_27),.data_out(wire_d64_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6506429(.data_in(wire_d64_28),.data_out(wire_d64_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6506430(.data_in(wire_d64_29),.data_out(wire_d64_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6506431(.data_in(wire_d64_30),.data_out(wire_d64_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6506432(.data_in(wire_d64_31),.data_out(wire_d64_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6506433(.data_in(wire_d64_32),.data_out(wire_d64_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6506434(.data_in(wire_d64_33),.data_out(wire_d64_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6506435(.data_in(wire_d64_34),.data_out(wire_d64_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6506436(.data_in(wire_d64_35),.data_out(wire_d64_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6506437(.data_in(wire_d64_36),.data_out(wire_d64_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6506438(.data_in(wire_d64_37),.data_out(wire_d64_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6506439(.data_in(wire_d64_38),.data_out(wire_d64_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6506440(.data_in(wire_d64_39),.data_out(wire_d64_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6506441(.data_in(wire_d64_40),.data_out(wire_d64_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6506442(.data_in(wire_d64_41),.data_out(wire_d64_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6506443(.data_in(wire_d64_42),.data_out(wire_d64_43),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6506444(.data_in(wire_d64_43),.data_out(wire_d64_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6506445(.data_in(wire_d64_44),.data_out(wire_d64_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6506446(.data_in(wire_d64_45),.data_out(wire_d64_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6506447(.data_in(wire_d64_46),.data_out(wire_d64_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6506448(.data_in(wire_d64_47),.data_out(wire_d64_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6506449(.data_in(wire_d64_48),.data_out(wire_d64_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6506450(.data_in(wire_d64_49),.data_out(wire_d64_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6506451(.data_in(wire_d64_50),.data_out(wire_d64_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6506452(.data_in(wire_d64_51),.data_out(wire_d64_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6506453(.data_in(wire_d64_52),.data_out(wire_d64_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6506454(.data_in(wire_d64_53),.data_out(wire_d64_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6506455(.data_in(wire_d64_54),.data_out(wire_d64_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6506456(.data_in(wire_d64_55),.data_out(wire_d64_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6506457(.data_in(wire_d64_56),.data_out(wire_d64_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6506458(.data_in(wire_d64_57),.data_out(wire_d64_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6506459(.data_in(wire_d64_58),.data_out(wire_d64_59),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6506460(.data_in(wire_d64_59),.data_out(wire_d64_60),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6506461(.data_in(wire_d64_60),.data_out(wire_d64_61),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6506462(.data_in(wire_d64_61),.data_out(wire_d64_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6506463(.data_in(wire_d64_62),.data_out(wire_d64_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6506464(.data_in(wire_d64_63),.data_out(wire_d64_64),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6506465(.data_in(wire_d64_64),.data_out(wire_d64_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6506466(.data_in(wire_d64_65),.data_out(wire_d64_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6506467(.data_in(wire_d64_66),.data_out(wire_d64_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6506468(.data_in(wire_d64_67),.data_out(wire_d64_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6506469(.data_in(wire_d64_68),.data_out(wire_d64_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6506470(.data_in(wire_d64_69),.data_out(wire_d64_70),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6506471(.data_in(wire_d64_70),.data_out(wire_d64_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6506472(.data_in(wire_d64_71),.data_out(wire_d64_72),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6506473(.data_in(wire_d64_72),.data_out(wire_d64_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6506474(.data_in(wire_d64_73),.data_out(wire_d64_74),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6506475(.data_in(wire_d64_74),.data_out(wire_d64_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6506476(.data_in(wire_d64_75),.data_out(wire_d64_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6506477(.data_in(wire_d64_76),.data_out(wire_d64_77),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6506478(.data_in(wire_d64_77),.data_out(wire_d64_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6506479(.data_in(wire_d64_78),.data_out(d_out64),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance660650(.data_in(d_in65),.data_out(wire_d65_0),.clk(clk),.rst(rst));            //channel 66
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance660651(.data_in(wire_d65_0),.data_out(wire_d65_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance660652(.data_in(wire_d65_1),.data_out(wire_d65_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance660653(.data_in(wire_d65_2),.data_out(wire_d65_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance660654(.data_in(wire_d65_3),.data_out(wire_d65_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance660655(.data_in(wire_d65_4),.data_out(wire_d65_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance660656(.data_in(wire_d65_5),.data_out(wire_d65_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance660657(.data_in(wire_d65_6),.data_out(wire_d65_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance660658(.data_in(wire_d65_7),.data_out(wire_d65_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance660659(.data_in(wire_d65_8),.data_out(wire_d65_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6606510(.data_in(wire_d65_9),.data_out(wire_d65_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6606511(.data_in(wire_d65_10),.data_out(wire_d65_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6606512(.data_in(wire_d65_11),.data_out(wire_d65_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6606513(.data_in(wire_d65_12),.data_out(wire_d65_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6606514(.data_in(wire_d65_13),.data_out(wire_d65_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6606515(.data_in(wire_d65_14),.data_out(wire_d65_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6606516(.data_in(wire_d65_15),.data_out(wire_d65_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6606517(.data_in(wire_d65_16),.data_out(wire_d65_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6606518(.data_in(wire_d65_17),.data_out(wire_d65_18),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6606519(.data_in(wire_d65_18),.data_out(wire_d65_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6606520(.data_in(wire_d65_19),.data_out(wire_d65_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6606521(.data_in(wire_d65_20),.data_out(wire_d65_21),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6606522(.data_in(wire_d65_21),.data_out(wire_d65_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6606523(.data_in(wire_d65_22),.data_out(wire_d65_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6606524(.data_in(wire_d65_23),.data_out(wire_d65_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6606525(.data_in(wire_d65_24),.data_out(wire_d65_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6606526(.data_in(wire_d65_25),.data_out(wire_d65_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6606527(.data_in(wire_d65_26),.data_out(wire_d65_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6606528(.data_in(wire_d65_27),.data_out(wire_d65_28),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6606529(.data_in(wire_d65_28),.data_out(wire_d65_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6606530(.data_in(wire_d65_29),.data_out(wire_d65_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6606531(.data_in(wire_d65_30),.data_out(wire_d65_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6606532(.data_in(wire_d65_31),.data_out(wire_d65_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6606533(.data_in(wire_d65_32),.data_out(wire_d65_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6606534(.data_in(wire_d65_33),.data_out(wire_d65_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6606535(.data_in(wire_d65_34),.data_out(wire_d65_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6606536(.data_in(wire_d65_35),.data_out(wire_d65_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6606537(.data_in(wire_d65_36),.data_out(wire_d65_37),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6606538(.data_in(wire_d65_37),.data_out(wire_d65_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6606539(.data_in(wire_d65_38),.data_out(wire_d65_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6606540(.data_in(wire_d65_39),.data_out(wire_d65_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6606541(.data_in(wire_d65_40),.data_out(wire_d65_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6606542(.data_in(wire_d65_41),.data_out(wire_d65_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6606543(.data_in(wire_d65_42),.data_out(wire_d65_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6606544(.data_in(wire_d65_43),.data_out(wire_d65_44),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6606545(.data_in(wire_d65_44),.data_out(wire_d65_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6606546(.data_in(wire_d65_45),.data_out(wire_d65_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6606547(.data_in(wire_d65_46),.data_out(wire_d65_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6606548(.data_in(wire_d65_47),.data_out(wire_d65_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6606549(.data_in(wire_d65_48),.data_out(wire_d65_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6606550(.data_in(wire_d65_49),.data_out(wire_d65_50),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6606551(.data_in(wire_d65_50),.data_out(wire_d65_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6606552(.data_in(wire_d65_51),.data_out(wire_d65_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6606553(.data_in(wire_d65_52),.data_out(wire_d65_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6606554(.data_in(wire_d65_53),.data_out(wire_d65_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6606555(.data_in(wire_d65_54),.data_out(wire_d65_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6606556(.data_in(wire_d65_55),.data_out(wire_d65_56),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6606557(.data_in(wire_d65_56),.data_out(wire_d65_57),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6606558(.data_in(wire_d65_57),.data_out(wire_d65_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6606559(.data_in(wire_d65_58),.data_out(wire_d65_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6606560(.data_in(wire_d65_59),.data_out(wire_d65_60),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6606561(.data_in(wire_d65_60),.data_out(wire_d65_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6606562(.data_in(wire_d65_61),.data_out(wire_d65_62),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6606563(.data_in(wire_d65_62),.data_out(wire_d65_63),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6606564(.data_in(wire_d65_63),.data_out(wire_d65_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6606565(.data_in(wire_d65_64),.data_out(wire_d65_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6606566(.data_in(wire_d65_65),.data_out(wire_d65_66),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6606567(.data_in(wire_d65_66),.data_out(wire_d65_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6606568(.data_in(wire_d65_67),.data_out(wire_d65_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6606569(.data_in(wire_d65_68),.data_out(wire_d65_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6606570(.data_in(wire_d65_69),.data_out(wire_d65_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6606571(.data_in(wire_d65_70),.data_out(wire_d65_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6606572(.data_in(wire_d65_71),.data_out(wire_d65_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6606573(.data_in(wire_d65_72),.data_out(wire_d65_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6606574(.data_in(wire_d65_73),.data_out(wire_d65_74),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6606575(.data_in(wire_d65_74),.data_out(wire_d65_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6606576(.data_in(wire_d65_75),.data_out(wire_d65_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6606577(.data_in(wire_d65_76),.data_out(wire_d65_77),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6606578(.data_in(wire_d65_77),.data_out(wire_d65_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6606579(.data_in(wire_d65_78),.data_out(d_out65),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance670660(.data_in(d_in66),.data_out(wire_d66_0),.clk(clk),.rst(rst));            //channel 67
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance670661(.data_in(wire_d66_0),.data_out(wire_d66_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance670662(.data_in(wire_d66_1),.data_out(wire_d66_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance670663(.data_in(wire_d66_2),.data_out(wire_d66_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance670664(.data_in(wire_d66_3),.data_out(wire_d66_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance670665(.data_in(wire_d66_4),.data_out(wire_d66_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance670666(.data_in(wire_d66_5),.data_out(wire_d66_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance670667(.data_in(wire_d66_6),.data_out(wire_d66_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance670668(.data_in(wire_d66_7),.data_out(wire_d66_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance670669(.data_in(wire_d66_8),.data_out(wire_d66_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6706610(.data_in(wire_d66_9),.data_out(wire_d66_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6706611(.data_in(wire_d66_10),.data_out(wire_d66_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6706612(.data_in(wire_d66_11),.data_out(wire_d66_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6706613(.data_in(wire_d66_12),.data_out(wire_d66_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6706614(.data_in(wire_d66_13),.data_out(wire_d66_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6706615(.data_in(wire_d66_14),.data_out(wire_d66_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6706616(.data_in(wire_d66_15),.data_out(wire_d66_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6706617(.data_in(wire_d66_16),.data_out(wire_d66_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6706618(.data_in(wire_d66_17),.data_out(wire_d66_18),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6706619(.data_in(wire_d66_18),.data_out(wire_d66_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6706620(.data_in(wire_d66_19),.data_out(wire_d66_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6706621(.data_in(wire_d66_20),.data_out(wire_d66_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6706622(.data_in(wire_d66_21),.data_out(wire_d66_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6706623(.data_in(wire_d66_22),.data_out(wire_d66_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6706624(.data_in(wire_d66_23),.data_out(wire_d66_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6706625(.data_in(wire_d66_24),.data_out(wire_d66_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6706626(.data_in(wire_d66_25),.data_out(wire_d66_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6706627(.data_in(wire_d66_26),.data_out(wire_d66_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6706628(.data_in(wire_d66_27),.data_out(wire_d66_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6706629(.data_in(wire_d66_28),.data_out(wire_d66_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6706630(.data_in(wire_d66_29),.data_out(wire_d66_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6706631(.data_in(wire_d66_30),.data_out(wire_d66_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6706632(.data_in(wire_d66_31),.data_out(wire_d66_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6706633(.data_in(wire_d66_32),.data_out(wire_d66_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6706634(.data_in(wire_d66_33),.data_out(wire_d66_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6706635(.data_in(wire_d66_34),.data_out(wire_d66_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6706636(.data_in(wire_d66_35),.data_out(wire_d66_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6706637(.data_in(wire_d66_36),.data_out(wire_d66_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6706638(.data_in(wire_d66_37),.data_out(wire_d66_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6706639(.data_in(wire_d66_38),.data_out(wire_d66_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6706640(.data_in(wire_d66_39),.data_out(wire_d66_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6706641(.data_in(wire_d66_40),.data_out(wire_d66_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6706642(.data_in(wire_d66_41),.data_out(wire_d66_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6706643(.data_in(wire_d66_42),.data_out(wire_d66_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6706644(.data_in(wire_d66_43),.data_out(wire_d66_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6706645(.data_in(wire_d66_44),.data_out(wire_d66_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6706646(.data_in(wire_d66_45),.data_out(wire_d66_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6706647(.data_in(wire_d66_46),.data_out(wire_d66_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6706648(.data_in(wire_d66_47),.data_out(wire_d66_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6706649(.data_in(wire_d66_48),.data_out(wire_d66_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6706650(.data_in(wire_d66_49),.data_out(wire_d66_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6706651(.data_in(wire_d66_50),.data_out(wire_d66_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6706652(.data_in(wire_d66_51),.data_out(wire_d66_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6706653(.data_in(wire_d66_52),.data_out(wire_d66_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6706654(.data_in(wire_d66_53),.data_out(wire_d66_54),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6706655(.data_in(wire_d66_54),.data_out(wire_d66_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6706656(.data_in(wire_d66_55),.data_out(wire_d66_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6706657(.data_in(wire_d66_56),.data_out(wire_d66_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6706658(.data_in(wire_d66_57),.data_out(wire_d66_58),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6706659(.data_in(wire_d66_58),.data_out(wire_d66_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6706660(.data_in(wire_d66_59),.data_out(wire_d66_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6706661(.data_in(wire_d66_60),.data_out(wire_d66_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6706662(.data_in(wire_d66_61),.data_out(wire_d66_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6706663(.data_in(wire_d66_62),.data_out(wire_d66_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6706664(.data_in(wire_d66_63),.data_out(wire_d66_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6706665(.data_in(wire_d66_64),.data_out(wire_d66_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6706666(.data_in(wire_d66_65),.data_out(wire_d66_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6706667(.data_in(wire_d66_66),.data_out(wire_d66_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6706668(.data_in(wire_d66_67),.data_out(wire_d66_68),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6706669(.data_in(wire_d66_68),.data_out(wire_d66_69),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6706670(.data_in(wire_d66_69),.data_out(wire_d66_70),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6706671(.data_in(wire_d66_70),.data_out(wire_d66_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6706672(.data_in(wire_d66_71),.data_out(wire_d66_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6706673(.data_in(wire_d66_72),.data_out(wire_d66_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6706674(.data_in(wire_d66_73),.data_out(wire_d66_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6706675(.data_in(wire_d66_74),.data_out(wire_d66_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6706676(.data_in(wire_d66_75),.data_out(wire_d66_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6706677(.data_in(wire_d66_76),.data_out(wire_d66_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6706678(.data_in(wire_d66_77),.data_out(wire_d66_78),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6706679(.data_in(wire_d66_78),.data_out(d_out66),.clk(clk),.rst(rst));

	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance680670(.data_in(d_in67),.data_out(wire_d67_0),.clk(clk),.rst(rst));            //channel 68
	register #(.WIDTH(WIDTH)) register_instance680671(.data_in(wire_d67_0),.data_out(wire_d67_1),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance680672(.data_in(wire_d67_1),.data_out(wire_d67_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance680673(.data_in(wire_d67_2),.data_out(wire_d67_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance680674(.data_in(wire_d67_3),.data_out(wire_d67_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance680675(.data_in(wire_d67_4),.data_out(wire_d67_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance680676(.data_in(wire_d67_5),.data_out(wire_d67_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance680677(.data_in(wire_d67_6),.data_out(wire_d67_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance680678(.data_in(wire_d67_7),.data_out(wire_d67_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance680679(.data_in(wire_d67_8),.data_out(wire_d67_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6806710(.data_in(wire_d67_9),.data_out(wire_d67_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6806711(.data_in(wire_d67_10),.data_out(wire_d67_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6806712(.data_in(wire_d67_11),.data_out(wire_d67_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6806713(.data_in(wire_d67_12),.data_out(wire_d67_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6806714(.data_in(wire_d67_13),.data_out(wire_d67_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6806715(.data_in(wire_d67_14),.data_out(wire_d67_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6806716(.data_in(wire_d67_15),.data_out(wire_d67_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6806717(.data_in(wire_d67_16),.data_out(wire_d67_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6806718(.data_in(wire_d67_17),.data_out(wire_d67_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6806719(.data_in(wire_d67_18),.data_out(wire_d67_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6806720(.data_in(wire_d67_19),.data_out(wire_d67_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6806721(.data_in(wire_d67_20),.data_out(wire_d67_21),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6806722(.data_in(wire_d67_21),.data_out(wire_d67_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6806723(.data_in(wire_d67_22),.data_out(wire_d67_23),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6806724(.data_in(wire_d67_23),.data_out(wire_d67_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6806725(.data_in(wire_d67_24),.data_out(wire_d67_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6806726(.data_in(wire_d67_25),.data_out(wire_d67_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6806727(.data_in(wire_d67_26),.data_out(wire_d67_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6806728(.data_in(wire_d67_27),.data_out(wire_d67_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6806729(.data_in(wire_d67_28),.data_out(wire_d67_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6806730(.data_in(wire_d67_29),.data_out(wire_d67_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6806731(.data_in(wire_d67_30),.data_out(wire_d67_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6806732(.data_in(wire_d67_31),.data_out(wire_d67_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6806733(.data_in(wire_d67_32),.data_out(wire_d67_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6806734(.data_in(wire_d67_33),.data_out(wire_d67_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6806735(.data_in(wire_d67_34),.data_out(wire_d67_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6806736(.data_in(wire_d67_35),.data_out(wire_d67_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6806737(.data_in(wire_d67_36),.data_out(wire_d67_37),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6806738(.data_in(wire_d67_37),.data_out(wire_d67_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6806739(.data_in(wire_d67_38),.data_out(wire_d67_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6806740(.data_in(wire_d67_39),.data_out(wire_d67_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6806741(.data_in(wire_d67_40),.data_out(wire_d67_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6806742(.data_in(wire_d67_41),.data_out(wire_d67_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6806743(.data_in(wire_d67_42),.data_out(wire_d67_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6806744(.data_in(wire_d67_43),.data_out(wire_d67_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6806745(.data_in(wire_d67_44),.data_out(wire_d67_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6806746(.data_in(wire_d67_45),.data_out(wire_d67_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6806747(.data_in(wire_d67_46),.data_out(wire_d67_47),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6806748(.data_in(wire_d67_47),.data_out(wire_d67_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6806749(.data_in(wire_d67_48),.data_out(wire_d67_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6806750(.data_in(wire_d67_49),.data_out(wire_d67_50),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6806751(.data_in(wire_d67_50),.data_out(wire_d67_51),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6806752(.data_in(wire_d67_51),.data_out(wire_d67_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6806753(.data_in(wire_d67_52),.data_out(wire_d67_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6806754(.data_in(wire_d67_53),.data_out(wire_d67_54),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6806755(.data_in(wire_d67_54),.data_out(wire_d67_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6806756(.data_in(wire_d67_55),.data_out(wire_d67_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6806757(.data_in(wire_d67_56),.data_out(wire_d67_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6806758(.data_in(wire_d67_57),.data_out(wire_d67_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6806759(.data_in(wire_d67_58),.data_out(wire_d67_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6806760(.data_in(wire_d67_59),.data_out(wire_d67_60),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6806761(.data_in(wire_d67_60),.data_out(wire_d67_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6806762(.data_in(wire_d67_61),.data_out(wire_d67_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6806763(.data_in(wire_d67_62),.data_out(wire_d67_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6806764(.data_in(wire_d67_63),.data_out(wire_d67_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6806765(.data_in(wire_d67_64),.data_out(wire_d67_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6806766(.data_in(wire_d67_65),.data_out(wire_d67_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6806767(.data_in(wire_d67_66),.data_out(wire_d67_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6806768(.data_in(wire_d67_67),.data_out(wire_d67_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6806769(.data_in(wire_d67_68),.data_out(wire_d67_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6806770(.data_in(wire_d67_69),.data_out(wire_d67_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6806771(.data_in(wire_d67_70),.data_out(wire_d67_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6806772(.data_in(wire_d67_71),.data_out(wire_d67_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6806773(.data_in(wire_d67_72),.data_out(wire_d67_73),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6806774(.data_in(wire_d67_73),.data_out(wire_d67_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6806775(.data_in(wire_d67_74),.data_out(wire_d67_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6806776(.data_in(wire_d67_75),.data_out(wire_d67_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6806777(.data_in(wire_d67_76),.data_out(wire_d67_77),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6806778(.data_in(wire_d67_77),.data_out(wire_d67_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6806779(.data_in(wire_d67_78),.data_out(d_out67),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance690680(.data_in(d_in68),.data_out(wire_d68_0),.clk(clk),.rst(rst));            //channel 69
	decoder_top #(.WIDTH(WIDTH)) decoder_instance690681(.data_in(wire_d68_0),.data_out(wire_d68_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance690682(.data_in(wire_d68_1),.data_out(wire_d68_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance690683(.data_in(wire_d68_2),.data_out(wire_d68_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance690684(.data_in(wire_d68_3),.data_out(wire_d68_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance690685(.data_in(wire_d68_4),.data_out(wire_d68_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance690686(.data_in(wire_d68_5),.data_out(wire_d68_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance690687(.data_in(wire_d68_6),.data_out(wire_d68_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance690688(.data_in(wire_d68_7),.data_out(wire_d68_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance690689(.data_in(wire_d68_8),.data_out(wire_d68_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6906810(.data_in(wire_d68_9),.data_out(wire_d68_10),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6906811(.data_in(wire_d68_10),.data_out(wire_d68_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6906812(.data_in(wire_d68_11),.data_out(wire_d68_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6906813(.data_in(wire_d68_12),.data_out(wire_d68_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6906814(.data_in(wire_d68_13),.data_out(wire_d68_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6906815(.data_in(wire_d68_14),.data_out(wire_d68_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6906816(.data_in(wire_d68_15),.data_out(wire_d68_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6906817(.data_in(wire_d68_16),.data_out(wire_d68_17),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6906818(.data_in(wire_d68_17),.data_out(wire_d68_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6906819(.data_in(wire_d68_18),.data_out(wire_d68_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6906820(.data_in(wire_d68_19),.data_out(wire_d68_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6906821(.data_in(wire_d68_20),.data_out(wire_d68_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6906822(.data_in(wire_d68_21),.data_out(wire_d68_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6906823(.data_in(wire_d68_22),.data_out(wire_d68_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6906824(.data_in(wire_d68_23),.data_out(wire_d68_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6906825(.data_in(wire_d68_24),.data_out(wire_d68_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6906826(.data_in(wire_d68_25),.data_out(wire_d68_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6906827(.data_in(wire_d68_26),.data_out(wire_d68_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6906828(.data_in(wire_d68_27),.data_out(wire_d68_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6906829(.data_in(wire_d68_28),.data_out(wire_d68_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6906830(.data_in(wire_d68_29),.data_out(wire_d68_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6906831(.data_in(wire_d68_30),.data_out(wire_d68_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6906832(.data_in(wire_d68_31),.data_out(wire_d68_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6906833(.data_in(wire_d68_32),.data_out(wire_d68_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6906834(.data_in(wire_d68_33),.data_out(wire_d68_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6906835(.data_in(wire_d68_34),.data_out(wire_d68_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6906836(.data_in(wire_d68_35),.data_out(wire_d68_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6906837(.data_in(wire_d68_36),.data_out(wire_d68_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6906838(.data_in(wire_d68_37),.data_out(wire_d68_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6906839(.data_in(wire_d68_38),.data_out(wire_d68_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6906840(.data_in(wire_d68_39),.data_out(wire_d68_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6906841(.data_in(wire_d68_40),.data_out(wire_d68_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6906842(.data_in(wire_d68_41),.data_out(wire_d68_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6906843(.data_in(wire_d68_42),.data_out(wire_d68_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6906844(.data_in(wire_d68_43),.data_out(wire_d68_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6906845(.data_in(wire_d68_44),.data_out(wire_d68_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6906846(.data_in(wire_d68_45),.data_out(wire_d68_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6906847(.data_in(wire_d68_46),.data_out(wire_d68_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6906848(.data_in(wire_d68_47),.data_out(wire_d68_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6906849(.data_in(wire_d68_48),.data_out(wire_d68_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6906850(.data_in(wire_d68_49),.data_out(wire_d68_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6906851(.data_in(wire_d68_50),.data_out(wire_d68_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6906852(.data_in(wire_d68_51),.data_out(wire_d68_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6906853(.data_in(wire_d68_52),.data_out(wire_d68_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6906854(.data_in(wire_d68_53),.data_out(wire_d68_54),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6906855(.data_in(wire_d68_54),.data_out(wire_d68_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6906856(.data_in(wire_d68_55),.data_out(wire_d68_56),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6906857(.data_in(wire_d68_56),.data_out(wire_d68_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6906858(.data_in(wire_d68_57),.data_out(wire_d68_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6906859(.data_in(wire_d68_58),.data_out(wire_d68_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6906860(.data_in(wire_d68_59),.data_out(wire_d68_60),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6906861(.data_in(wire_d68_60),.data_out(wire_d68_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6906862(.data_in(wire_d68_61),.data_out(wire_d68_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6906863(.data_in(wire_d68_62),.data_out(wire_d68_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6906864(.data_in(wire_d68_63),.data_out(wire_d68_64),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6906865(.data_in(wire_d68_64),.data_out(wire_d68_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6906866(.data_in(wire_d68_65),.data_out(wire_d68_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6906867(.data_in(wire_d68_66),.data_out(wire_d68_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6906868(.data_in(wire_d68_67),.data_out(wire_d68_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6906869(.data_in(wire_d68_68),.data_out(wire_d68_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6906870(.data_in(wire_d68_69),.data_out(wire_d68_70),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6906871(.data_in(wire_d68_70),.data_out(wire_d68_71),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6906872(.data_in(wire_d68_71),.data_out(wire_d68_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6906873(.data_in(wire_d68_72),.data_out(wire_d68_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6906874(.data_in(wire_d68_73),.data_out(wire_d68_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6906875(.data_in(wire_d68_74),.data_out(wire_d68_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6906876(.data_in(wire_d68_75),.data_out(wire_d68_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6906877(.data_in(wire_d68_76),.data_out(wire_d68_77),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6906878(.data_in(wire_d68_77),.data_out(wire_d68_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6906879(.data_in(wire_d68_78),.data_out(d_out68),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance700690(.data_in(d_in69),.data_out(wire_d69_0),.clk(clk),.rst(rst));            //channel 70
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance700691(.data_in(wire_d69_0),.data_out(wire_d69_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance700692(.data_in(wire_d69_1),.data_out(wire_d69_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance700693(.data_in(wire_d69_2),.data_out(wire_d69_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance700694(.data_in(wire_d69_3),.data_out(wire_d69_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance700695(.data_in(wire_d69_4),.data_out(wire_d69_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance700696(.data_in(wire_d69_5),.data_out(wire_d69_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance700697(.data_in(wire_d69_6),.data_out(wire_d69_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance700698(.data_in(wire_d69_7),.data_out(wire_d69_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance700699(.data_in(wire_d69_8),.data_out(wire_d69_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7006910(.data_in(wire_d69_9),.data_out(wire_d69_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7006911(.data_in(wire_d69_10),.data_out(wire_d69_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7006912(.data_in(wire_d69_11),.data_out(wire_d69_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7006913(.data_in(wire_d69_12),.data_out(wire_d69_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7006914(.data_in(wire_d69_13),.data_out(wire_d69_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7006915(.data_in(wire_d69_14),.data_out(wire_d69_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7006916(.data_in(wire_d69_15),.data_out(wire_d69_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7006917(.data_in(wire_d69_16),.data_out(wire_d69_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7006918(.data_in(wire_d69_17),.data_out(wire_d69_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7006919(.data_in(wire_d69_18),.data_out(wire_d69_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7006920(.data_in(wire_d69_19),.data_out(wire_d69_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7006921(.data_in(wire_d69_20),.data_out(wire_d69_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7006922(.data_in(wire_d69_21),.data_out(wire_d69_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7006923(.data_in(wire_d69_22),.data_out(wire_d69_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7006924(.data_in(wire_d69_23),.data_out(wire_d69_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7006925(.data_in(wire_d69_24),.data_out(wire_d69_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7006926(.data_in(wire_d69_25),.data_out(wire_d69_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7006927(.data_in(wire_d69_26),.data_out(wire_d69_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7006928(.data_in(wire_d69_27),.data_out(wire_d69_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7006929(.data_in(wire_d69_28),.data_out(wire_d69_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7006930(.data_in(wire_d69_29),.data_out(wire_d69_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7006931(.data_in(wire_d69_30),.data_out(wire_d69_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7006932(.data_in(wire_d69_31),.data_out(wire_d69_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7006933(.data_in(wire_d69_32),.data_out(wire_d69_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7006934(.data_in(wire_d69_33),.data_out(wire_d69_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7006935(.data_in(wire_d69_34),.data_out(wire_d69_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7006936(.data_in(wire_d69_35),.data_out(wire_d69_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7006937(.data_in(wire_d69_36),.data_out(wire_d69_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7006938(.data_in(wire_d69_37),.data_out(wire_d69_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7006939(.data_in(wire_d69_38),.data_out(wire_d69_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7006940(.data_in(wire_d69_39),.data_out(wire_d69_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7006941(.data_in(wire_d69_40),.data_out(wire_d69_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7006942(.data_in(wire_d69_41),.data_out(wire_d69_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7006943(.data_in(wire_d69_42),.data_out(wire_d69_43),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7006944(.data_in(wire_d69_43),.data_out(wire_d69_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7006945(.data_in(wire_d69_44),.data_out(wire_d69_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7006946(.data_in(wire_d69_45),.data_out(wire_d69_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7006947(.data_in(wire_d69_46),.data_out(wire_d69_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7006948(.data_in(wire_d69_47),.data_out(wire_d69_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7006949(.data_in(wire_d69_48),.data_out(wire_d69_49),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7006950(.data_in(wire_d69_49),.data_out(wire_d69_50),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7006951(.data_in(wire_d69_50),.data_out(wire_d69_51),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7006952(.data_in(wire_d69_51),.data_out(wire_d69_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7006953(.data_in(wire_d69_52),.data_out(wire_d69_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7006954(.data_in(wire_d69_53),.data_out(wire_d69_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7006955(.data_in(wire_d69_54),.data_out(wire_d69_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7006956(.data_in(wire_d69_55),.data_out(wire_d69_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7006957(.data_in(wire_d69_56),.data_out(wire_d69_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7006958(.data_in(wire_d69_57),.data_out(wire_d69_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7006959(.data_in(wire_d69_58),.data_out(wire_d69_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7006960(.data_in(wire_d69_59),.data_out(wire_d69_60),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7006961(.data_in(wire_d69_60),.data_out(wire_d69_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7006962(.data_in(wire_d69_61),.data_out(wire_d69_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7006963(.data_in(wire_d69_62),.data_out(wire_d69_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7006964(.data_in(wire_d69_63),.data_out(wire_d69_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7006965(.data_in(wire_d69_64),.data_out(wire_d69_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7006966(.data_in(wire_d69_65),.data_out(wire_d69_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7006967(.data_in(wire_d69_66),.data_out(wire_d69_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7006968(.data_in(wire_d69_67),.data_out(wire_d69_68),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7006969(.data_in(wire_d69_68),.data_out(wire_d69_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7006970(.data_in(wire_d69_69),.data_out(wire_d69_70),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7006971(.data_in(wire_d69_70),.data_out(wire_d69_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7006972(.data_in(wire_d69_71),.data_out(wire_d69_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7006973(.data_in(wire_d69_72),.data_out(wire_d69_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7006974(.data_in(wire_d69_73),.data_out(wire_d69_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7006975(.data_in(wire_d69_74),.data_out(wire_d69_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7006976(.data_in(wire_d69_75),.data_out(wire_d69_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7006977(.data_in(wire_d69_76),.data_out(wire_d69_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7006978(.data_in(wire_d69_77),.data_out(wire_d69_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7006979(.data_in(wire_d69_78),.data_out(d_out69),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance710700(.data_in(d_in70),.data_out(wire_d70_0),.clk(clk),.rst(rst));            //channel 71
	large_mux #(.WIDTH(WIDTH)) large_mux_instance710701(.data_in(wire_d70_0),.data_out(wire_d70_1),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance710702(.data_in(wire_d70_1),.data_out(wire_d70_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance710703(.data_in(wire_d70_2),.data_out(wire_d70_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance710704(.data_in(wire_d70_3),.data_out(wire_d70_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance710705(.data_in(wire_d70_4),.data_out(wire_d70_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance710706(.data_in(wire_d70_5),.data_out(wire_d70_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance710707(.data_in(wire_d70_6),.data_out(wire_d70_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance710708(.data_in(wire_d70_7),.data_out(wire_d70_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance710709(.data_in(wire_d70_8),.data_out(wire_d70_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7107010(.data_in(wire_d70_9),.data_out(wire_d70_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7107011(.data_in(wire_d70_10),.data_out(wire_d70_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7107012(.data_in(wire_d70_11),.data_out(wire_d70_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7107013(.data_in(wire_d70_12),.data_out(wire_d70_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7107014(.data_in(wire_d70_13),.data_out(wire_d70_14),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7107015(.data_in(wire_d70_14),.data_out(wire_d70_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7107016(.data_in(wire_d70_15),.data_out(wire_d70_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7107017(.data_in(wire_d70_16),.data_out(wire_d70_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7107018(.data_in(wire_d70_17),.data_out(wire_d70_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7107019(.data_in(wire_d70_18),.data_out(wire_d70_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7107020(.data_in(wire_d70_19),.data_out(wire_d70_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7107021(.data_in(wire_d70_20),.data_out(wire_d70_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7107022(.data_in(wire_d70_21),.data_out(wire_d70_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7107023(.data_in(wire_d70_22),.data_out(wire_d70_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7107024(.data_in(wire_d70_23),.data_out(wire_d70_24),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7107025(.data_in(wire_d70_24),.data_out(wire_d70_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7107026(.data_in(wire_d70_25),.data_out(wire_d70_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7107027(.data_in(wire_d70_26),.data_out(wire_d70_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7107028(.data_in(wire_d70_27),.data_out(wire_d70_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7107029(.data_in(wire_d70_28),.data_out(wire_d70_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7107030(.data_in(wire_d70_29),.data_out(wire_d70_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7107031(.data_in(wire_d70_30),.data_out(wire_d70_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7107032(.data_in(wire_d70_31),.data_out(wire_d70_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7107033(.data_in(wire_d70_32),.data_out(wire_d70_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7107034(.data_in(wire_d70_33),.data_out(wire_d70_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7107035(.data_in(wire_d70_34),.data_out(wire_d70_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7107036(.data_in(wire_d70_35),.data_out(wire_d70_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7107037(.data_in(wire_d70_36),.data_out(wire_d70_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7107038(.data_in(wire_d70_37),.data_out(wire_d70_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7107039(.data_in(wire_d70_38),.data_out(wire_d70_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7107040(.data_in(wire_d70_39),.data_out(wire_d70_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7107041(.data_in(wire_d70_40),.data_out(wire_d70_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7107042(.data_in(wire_d70_41),.data_out(wire_d70_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7107043(.data_in(wire_d70_42),.data_out(wire_d70_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7107044(.data_in(wire_d70_43),.data_out(wire_d70_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7107045(.data_in(wire_d70_44),.data_out(wire_d70_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7107046(.data_in(wire_d70_45),.data_out(wire_d70_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7107047(.data_in(wire_d70_46),.data_out(wire_d70_47),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7107048(.data_in(wire_d70_47),.data_out(wire_d70_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7107049(.data_in(wire_d70_48),.data_out(wire_d70_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7107050(.data_in(wire_d70_49),.data_out(wire_d70_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7107051(.data_in(wire_d70_50),.data_out(wire_d70_51),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7107052(.data_in(wire_d70_51),.data_out(wire_d70_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7107053(.data_in(wire_d70_52),.data_out(wire_d70_53),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7107054(.data_in(wire_d70_53),.data_out(wire_d70_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7107055(.data_in(wire_d70_54),.data_out(wire_d70_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7107056(.data_in(wire_d70_55),.data_out(wire_d70_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7107057(.data_in(wire_d70_56),.data_out(wire_d70_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7107058(.data_in(wire_d70_57),.data_out(wire_d70_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7107059(.data_in(wire_d70_58),.data_out(wire_d70_59),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7107060(.data_in(wire_d70_59),.data_out(wire_d70_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7107061(.data_in(wire_d70_60),.data_out(wire_d70_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7107062(.data_in(wire_d70_61),.data_out(wire_d70_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7107063(.data_in(wire_d70_62),.data_out(wire_d70_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7107064(.data_in(wire_d70_63),.data_out(wire_d70_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7107065(.data_in(wire_d70_64),.data_out(wire_d70_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7107066(.data_in(wire_d70_65),.data_out(wire_d70_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7107067(.data_in(wire_d70_66),.data_out(wire_d70_67),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7107068(.data_in(wire_d70_67),.data_out(wire_d70_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7107069(.data_in(wire_d70_68),.data_out(wire_d70_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7107070(.data_in(wire_d70_69),.data_out(wire_d70_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7107071(.data_in(wire_d70_70),.data_out(wire_d70_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7107072(.data_in(wire_d70_71),.data_out(wire_d70_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7107073(.data_in(wire_d70_72),.data_out(wire_d70_73),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7107074(.data_in(wire_d70_73),.data_out(wire_d70_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7107075(.data_in(wire_d70_74),.data_out(wire_d70_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7107076(.data_in(wire_d70_75),.data_out(wire_d70_76),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7107077(.data_in(wire_d70_76),.data_out(wire_d70_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7107078(.data_in(wire_d70_77),.data_out(wire_d70_78),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7107079(.data_in(wire_d70_78),.data_out(d_out70),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance720710(.data_in(d_in71),.data_out(wire_d71_0),.clk(clk),.rst(rst));            //channel 72
	decoder_top #(.WIDTH(WIDTH)) decoder_instance720711(.data_in(wire_d71_0),.data_out(wire_d71_1),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance720712(.data_in(wire_d71_1),.data_out(wire_d71_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance720713(.data_in(wire_d71_2),.data_out(wire_d71_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance720714(.data_in(wire_d71_3),.data_out(wire_d71_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance720715(.data_in(wire_d71_4),.data_out(wire_d71_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance720716(.data_in(wire_d71_5),.data_out(wire_d71_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance720717(.data_in(wire_d71_6),.data_out(wire_d71_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance720718(.data_in(wire_d71_7),.data_out(wire_d71_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance720719(.data_in(wire_d71_8),.data_out(wire_d71_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7207110(.data_in(wire_d71_9),.data_out(wire_d71_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7207111(.data_in(wire_d71_10),.data_out(wire_d71_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7207112(.data_in(wire_d71_11),.data_out(wire_d71_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7207113(.data_in(wire_d71_12),.data_out(wire_d71_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7207114(.data_in(wire_d71_13),.data_out(wire_d71_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7207115(.data_in(wire_d71_14),.data_out(wire_d71_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7207116(.data_in(wire_d71_15),.data_out(wire_d71_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7207117(.data_in(wire_d71_16),.data_out(wire_d71_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7207118(.data_in(wire_d71_17),.data_out(wire_d71_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7207119(.data_in(wire_d71_18),.data_out(wire_d71_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7207120(.data_in(wire_d71_19),.data_out(wire_d71_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7207121(.data_in(wire_d71_20),.data_out(wire_d71_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7207122(.data_in(wire_d71_21),.data_out(wire_d71_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7207123(.data_in(wire_d71_22),.data_out(wire_d71_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7207124(.data_in(wire_d71_23),.data_out(wire_d71_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7207125(.data_in(wire_d71_24),.data_out(wire_d71_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7207126(.data_in(wire_d71_25),.data_out(wire_d71_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7207127(.data_in(wire_d71_26),.data_out(wire_d71_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7207128(.data_in(wire_d71_27),.data_out(wire_d71_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7207129(.data_in(wire_d71_28),.data_out(wire_d71_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7207130(.data_in(wire_d71_29),.data_out(wire_d71_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7207131(.data_in(wire_d71_30),.data_out(wire_d71_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7207132(.data_in(wire_d71_31),.data_out(wire_d71_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7207133(.data_in(wire_d71_32),.data_out(wire_d71_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7207134(.data_in(wire_d71_33),.data_out(wire_d71_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7207135(.data_in(wire_d71_34),.data_out(wire_d71_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7207136(.data_in(wire_d71_35),.data_out(wire_d71_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7207137(.data_in(wire_d71_36),.data_out(wire_d71_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7207138(.data_in(wire_d71_37),.data_out(wire_d71_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7207139(.data_in(wire_d71_38),.data_out(wire_d71_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7207140(.data_in(wire_d71_39),.data_out(wire_d71_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7207141(.data_in(wire_d71_40),.data_out(wire_d71_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7207142(.data_in(wire_d71_41),.data_out(wire_d71_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7207143(.data_in(wire_d71_42),.data_out(wire_d71_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7207144(.data_in(wire_d71_43),.data_out(wire_d71_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7207145(.data_in(wire_d71_44),.data_out(wire_d71_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7207146(.data_in(wire_d71_45),.data_out(wire_d71_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7207147(.data_in(wire_d71_46),.data_out(wire_d71_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7207148(.data_in(wire_d71_47),.data_out(wire_d71_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7207149(.data_in(wire_d71_48),.data_out(wire_d71_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7207150(.data_in(wire_d71_49),.data_out(wire_d71_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7207151(.data_in(wire_d71_50),.data_out(wire_d71_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7207152(.data_in(wire_d71_51),.data_out(wire_d71_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7207153(.data_in(wire_d71_52),.data_out(wire_d71_53),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7207154(.data_in(wire_d71_53),.data_out(wire_d71_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7207155(.data_in(wire_d71_54),.data_out(wire_d71_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7207156(.data_in(wire_d71_55),.data_out(wire_d71_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7207157(.data_in(wire_d71_56),.data_out(wire_d71_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7207158(.data_in(wire_d71_57),.data_out(wire_d71_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7207159(.data_in(wire_d71_58),.data_out(wire_d71_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7207160(.data_in(wire_d71_59),.data_out(wire_d71_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7207161(.data_in(wire_d71_60),.data_out(wire_d71_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7207162(.data_in(wire_d71_61),.data_out(wire_d71_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7207163(.data_in(wire_d71_62),.data_out(wire_d71_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7207164(.data_in(wire_d71_63),.data_out(wire_d71_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7207165(.data_in(wire_d71_64),.data_out(wire_d71_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7207166(.data_in(wire_d71_65),.data_out(wire_d71_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7207167(.data_in(wire_d71_66),.data_out(wire_d71_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7207168(.data_in(wire_d71_67),.data_out(wire_d71_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7207169(.data_in(wire_d71_68),.data_out(wire_d71_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7207170(.data_in(wire_d71_69),.data_out(wire_d71_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7207171(.data_in(wire_d71_70),.data_out(wire_d71_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7207172(.data_in(wire_d71_71),.data_out(wire_d71_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7207173(.data_in(wire_d71_72),.data_out(wire_d71_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7207174(.data_in(wire_d71_73),.data_out(wire_d71_74),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7207175(.data_in(wire_d71_74),.data_out(wire_d71_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7207176(.data_in(wire_d71_75),.data_out(wire_d71_76),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7207177(.data_in(wire_d71_76),.data_out(wire_d71_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7207178(.data_in(wire_d71_77),.data_out(wire_d71_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7207179(.data_in(wire_d71_78),.data_out(d_out71),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance730720(.data_in(d_in72),.data_out(wire_d72_0),.clk(clk),.rst(rst));            //channel 73
	register #(.WIDTH(WIDTH)) register_instance730721(.data_in(wire_d72_0),.data_out(wire_d72_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance730722(.data_in(wire_d72_1),.data_out(wire_d72_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance730723(.data_in(wire_d72_2),.data_out(wire_d72_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance730724(.data_in(wire_d72_3),.data_out(wire_d72_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance730725(.data_in(wire_d72_4),.data_out(wire_d72_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance730726(.data_in(wire_d72_5),.data_out(wire_d72_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance730727(.data_in(wire_d72_6),.data_out(wire_d72_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance730728(.data_in(wire_d72_7),.data_out(wire_d72_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance730729(.data_in(wire_d72_8),.data_out(wire_d72_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7307210(.data_in(wire_d72_9),.data_out(wire_d72_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7307211(.data_in(wire_d72_10),.data_out(wire_d72_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7307212(.data_in(wire_d72_11),.data_out(wire_d72_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7307213(.data_in(wire_d72_12),.data_out(wire_d72_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7307214(.data_in(wire_d72_13),.data_out(wire_d72_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7307215(.data_in(wire_d72_14),.data_out(wire_d72_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7307216(.data_in(wire_d72_15),.data_out(wire_d72_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7307217(.data_in(wire_d72_16),.data_out(wire_d72_17),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7307218(.data_in(wire_d72_17),.data_out(wire_d72_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7307219(.data_in(wire_d72_18),.data_out(wire_d72_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7307220(.data_in(wire_d72_19),.data_out(wire_d72_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7307221(.data_in(wire_d72_20),.data_out(wire_d72_21),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7307222(.data_in(wire_d72_21),.data_out(wire_d72_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7307223(.data_in(wire_d72_22),.data_out(wire_d72_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7307224(.data_in(wire_d72_23),.data_out(wire_d72_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7307225(.data_in(wire_d72_24),.data_out(wire_d72_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7307226(.data_in(wire_d72_25),.data_out(wire_d72_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7307227(.data_in(wire_d72_26),.data_out(wire_d72_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7307228(.data_in(wire_d72_27),.data_out(wire_d72_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7307229(.data_in(wire_d72_28),.data_out(wire_d72_29),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7307230(.data_in(wire_d72_29),.data_out(wire_d72_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7307231(.data_in(wire_d72_30),.data_out(wire_d72_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7307232(.data_in(wire_d72_31),.data_out(wire_d72_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7307233(.data_in(wire_d72_32),.data_out(wire_d72_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7307234(.data_in(wire_d72_33),.data_out(wire_d72_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7307235(.data_in(wire_d72_34),.data_out(wire_d72_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7307236(.data_in(wire_d72_35),.data_out(wire_d72_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7307237(.data_in(wire_d72_36),.data_out(wire_d72_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7307238(.data_in(wire_d72_37),.data_out(wire_d72_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7307239(.data_in(wire_d72_38),.data_out(wire_d72_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7307240(.data_in(wire_d72_39),.data_out(wire_d72_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7307241(.data_in(wire_d72_40),.data_out(wire_d72_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7307242(.data_in(wire_d72_41),.data_out(wire_d72_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7307243(.data_in(wire_d72_42),.data_out(wire_d72_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7307244(.data_in(wire_d72_43),.data_out(wire_d72_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7307245(.data_in(wire_d72_44),.data_out(wire_d72_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7307246(.data_in(wire_d72_45),.data_out(wire_d72_46),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7307247(.data_in(wire_d72_46),.data_out(wire_d72_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7307248(.data_in(wire_d72_47),.data_out(wire_d72_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7307249(.data_in(wire_d72_48),.data_out(wire_d72_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7307250(.data_in(wire_d72_49),.data_out(wire_d72_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7307251(.data_in(wire_d72_50),.data_out(wire_d72_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7307252(.data_in(wire_d72_51),.data_out(wire_d72_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7307253(.data_in(wire_d72_52),.data_out(wire_d72_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7307254(.data_in(wire_d72_53),.data_out(wire_d72_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7307255(.data_in(wire_d72_54),.data_out(wire_d72_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7307256(.data_in(wire_d72_55),.data_out(wire_d72_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7307257(.data_in(wire_d72_56),.data_out(wire_d72_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7307258(.data_in(wire_d72_57),.data_out(wire_d72_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7307259(.data_in(wire_d72_58),.data_out(wire_d72_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7307260(.data_in(wire_d72_59),.data_out(wire_d72_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7307261(.data_in(wire_d72_60),.data_out(wire_d72_61),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7307262(.data_in(wire_d72_61),.data_out(wire_d72_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7307263(.data_in(wire_d72_62),.data_out(wire_d72_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7307264(.data_in(wire_d72_63),.data_out(wire_d72_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7307265(.data_in(wire_d72_64),.data_out(wire_d72_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7307266(.data_in(wire_d72_65),.data_out(wire_d72_66),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7307267(.data_in(wire_d72_66),.data_out(wire_d72_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7307268(.data_in(wire_d72_67),.data_out(wire_d72_68),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7307269(.data_in(wire_d72_68),.data_out(wire_d72_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7307270(.data_in(wire_d72_69),.data_out(wire_d72_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7307271(.data_in(wire_d72_70),.data_out(wire_d72_71),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7307272(.data_in(wire_d72_71),.data_out(wire_d72_72),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7307273(.data_in(wire_d72_72),.data_out(wire_d72_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7307274(.data_in(wire_d72_73),.data_out(wire_d72_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7307275(.data_in(wire_d72_74),.data_out(wire_d72_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7307276(.data_in(wire_d72_75),.data_out(wire_d72_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7307277(.data_in(wire_d72_76),.data_out(wire_d72_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7307278(.data_in(wire_d72_77),.data_out(wire_d72_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7307279(.data_in(wire_d72_78),.data_out(d_out72),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance740730(.data_in(d_in73),.data_out(wire_d73_0),.clk(clk),.rst(rst));            //channel 74
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance740731(.data_in(wire_d73_0),.data_out(wire_d73_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance740732(.data_in(wire_d73_1),.data_out(wire_d73_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance740733(.data_in(wire_d73_2),.data_out(wire_d73_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance740734(.data_in(wire_d73_3),.data_out(wire_d73_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance740735(.data_in(wire_d73_4),.data_out(wire_d73_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance740736(.data_in(wire_d73_5),.data_out(wire_d73_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance740737(.data_in(wire_d73_6),.data_out(wire_d73_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance740738(.data_in(wire_d73_7),.data_out(wire_d73_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance740739(.data_in(wire_d73_8),.data_out(wire_d73_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7407310(.data_in(wire_d73_9),.data_out(wire_d73_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7407311(.data_in(wire_d73_10),.data_out(wire_d73_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7407312(.data_in(wire_d73_11),.data_out(wire_d73_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7407313(.data_in(wire_d73_12),.data_out(wire_d73_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7407314(.data_in(wire_d73_13),.data_out(wire_d73_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7407315(.data_in(wire_d73_14),.data_out(wire_d73_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7407316(.data_in(wire_d73_15),.data_out(wire_d73_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7407317(.data_in(wire_d73_16),.data_out(wire_d73_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7407318(.data_in(wire_d73_17),.data_out(wire_d73_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7407319(.data_in(wire_d73_18),.data_out(wire_d73_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7407320(.data_in(wire_d73_19),.data_out(wire_d73_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7407321(.data_in(wire_d73_20),.data_out(wire_d73_21),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7407322(.data_in(wire_d73_21),.data_out(wire_d73_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7407323(.data_in(wire_d73_22),.data_out(wire_d73_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7407324(.data_in(wire_d73_23),.data_out(wire_d73_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7407325(.data_in(wire_d73_24),.data_out(wire_d73_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7407326(.data_in(wire_d73_25),.data_out(wire_d73_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7407327(.data_in(wire_d73_26),.data_out(wire_d73_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7407328(.data_in(wire_d73_27),.data_out(wire_d73_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7407329(.data_in(wire_d73_28),.data_out(wire_d73_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7407330(.data_in(wire_d73_29),.data_out(wire_d73_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7407331(.data_in(wire_d73_30),.data_out(wire_d73_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7407332(.data_in(wire_d73_31),.data_out(wire_d73_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7407333(.data_in(wire_d73_32),.data_out(wire_d73_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7407334(.data_in(wire_d73_33),.data_out(wire_d73_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7407335(.data_in(wire_d73_34),.data_out(wire_d73_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7407336(.data_in(wire_d73_35),.data_out(wire_d73_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7407337(.data_in(wire_d73_36),.data_out(wire_d73_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7407338(.data_in(wire_d73_37),.data_out(wire_d73_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7407339(.data_in(wire_d73_38),.data_out(wire_d73_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7407340(.data_in(wire_d73_39),.data_out(wire_d73_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7407341(.data_in(wire_d73_40),.data_out(wire_d73_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7407342(.data_in(wire_d73_41),.data_out(wire_d73_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7407343(.data_in(wire_d73_42),.data_out(wire_d73_43),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7407344(.data_in(wire_d73_43),.data_out(wire_d73_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7407345(.data_in(wire_d73_44),.data_out(wire_d73_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7407346(.data_in(wire_d73_45),.data_out(wire_d73_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7407347(.data_in(wire_d73_46),.data_out(wire_d73_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7407348(.data_in(wire_d73_47),.data_out(wire_d73_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7407349(.data_in(wire_d73_48),.data_out(wire_d73_49),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7407350(.data_in(wire_d73_49),.data_out(wire_d73_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7407351(.data_in(wire_d73_50),.data_out(wire_d73_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7407352(.data_in(wire_d73_51),.data_out(wire_d73_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7407353(.data_in(wire_d73_52),.data_out(wire_d73_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7407354(.data_in(wire_d73_53),.data_out(wire_d73_54),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7407355(.data_in(wire_d73_54),.data_out(wire_d73_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7407356(.data_in(wire_d73_55),.data_out(wire_d73_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7407357(.data_in(wire_d73_56),.data_out(wire_d73_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7407358(.data_in(wire_d73_57),.data_out(wire_d73_58),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7407359(.data_in(wire_d73_58),.data_out(wire_d73_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7407360(.data_in(wire_d73_59),.data_out(wire_d73_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7407361(.data_in(wire_d73_60),.data_out(wire_d73_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7407362(.data_in(wire_d73_61),.data_out(wire_d73_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7407363(.data_in(wire_d73_62),.data_out(wire_d73_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7407364(.data_in(wire_d73_63),.data_out(wire_d73_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7407365(.data_in(wire_d73_64),.data_out(wire_d73_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7407366(.data_in(wire_d73_65),.data_out(wire_d73_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7407367(.data_in(wire_d73_66),.data_out(wire_d73_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7407368(.data_in(wire_d73_67),.data_out(wire_d73_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7407369(.data_in(wire_d73_68),.data_out(wire_d73_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7407370(.data_in(wire_d73_69),.data_out(wire_d73_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7407371(.data_in(wire_d73_70),.data_out(wire_d73_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7407372(.data_in(wire_d73_71),.data_out(wire_d73_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7407373(.data_in(wire_d73_72),.data_out(wire_d73_73),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7407374(.data_in(wire_d73_73),.data_out(wire_d73_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7407375(.data_in(wire_d73_74),.data_out(wire_d73_75),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7407376(.data_in(wire_d73_75),.data_out(wire_d73_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7407377(.data_in(wire_d73_76),.data_out(wire_d73_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7407378(.data_in(wire_d73_77),.data_out(wire_d73_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7407379(.data_in(wire_d73_78),.data_out(d_out73),.clk(clk),.rst(rst));

	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance750740(.data_in(d_in74),.data_out(wire_d74_0),.clk(clk),.rst(rst));            //channel 75
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance750741(.data_in(wire_d74_0),.data_out(wire_d74_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance750742(.data_in(wire_d74_1),.data_out(wire_d74_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance750743(.data_in(wire_d74_2),.data_out(wire_d74_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance750744(.data_in(wire_d74_3),.data_out(wire_d74_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance750745(.data_in(wire_d74_4),.data_out(wire_d74_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance750746(.data_in(wire_d74_5),.data_out(wire_d74_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance750747(.data_in(wire_d74_6),.data_out(wire_d74_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance750748(.data_in(wire_d74_7),.data_out(wire_d74_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance750749(.data_in(wire_d74_8),.data_out(wire_d74_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7507410(.data_in(wire_d74_9),.data_out(wire_d74_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7507411(.data_in(wire_d74_10),.data_out(wire_d74_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7507412(.data_in(wire_d74_11),.data_out(wire_d74_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7507413(.data_in(wire_d74_12),.data_out(wire_d74_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7507414(.data_in(wire_d74_13),.data_out(wire_d74_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7507415(.data_in(wire_d74_14),.data_out(wire_d74_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7507416(.data_in(wire_d74_15),.data_out(wire_d74_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7507417(.data_in(wire_d74_16),.data_out(wire_d74_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7507418(.data_in(wire_d74_17),.data_out(wire_d74_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7507419(.data_in(wire_d74_18),.data_out(wire_d74_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7507420(.data_in(wire_d74_19),.data_out(wire_d74_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7507421(.data_in(wire_d74_20),.data_out(wire_d74_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7507422(.data_in(wire_d74_21),.data_out(wire_d74_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7507423(.data_in(wire_d74_22),.data_out(wire_d74_23),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7507424(.data_in(wire_d74_23),.data_out(wire_d74_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7507425(.data_in(wire_d74_24),.data_out(wire_d74_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7507426(.data_in(wire_d74_25),.data_out(wire_d74_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7507427(.data_in(wire_d74_26),.data_out(wire_d74_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7507428(.data_in(wire_d74_27),.data_out(wire_d74_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7507429(.data_in(wire_d74_28),.data_out(wire_d74_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7507430(.data_in(wire_d74_29),.data_out(wire_d74_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7507431(.data_in(wire_d74_30),.data_out(wire_d74_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7507432(.data_in(wire_d74_31),.data_out(wire_d74_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7507433(.data_in(wire_d74_32),.data_out(wire_d74_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7507434(.data_in(wire_d74_33),.data_out(wire_d74_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7507435(.data_in(wire_d74_34),.data_out(wire_d74_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7507436(.data_in(wire_d74_35),.data_out(wire_d74_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7507437(.data_in(wire_d74_36),.data_out(wire_d74_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7507438(.data_in(wire_d74_37),.data_out(wire_d74_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7507439(.data_in(wire_d74_38),.data_out(wire_d74_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7507440(.data_in(wire_d74_39),.data_out(wire_d74_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7507441(.data_in(wire_d74_40),.data_out(wire_d74_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7507442(.data_in(wire_d74_41),.data_out(wire_d74_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7507443(.data_in(wire_d74_42),.data_out(wire_d74_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7507444(.data_in(wire_d74_43),.data_out(wire_d74_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7507445(.data_in(wire_d74_44),.data_out(wire_d74_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7507446(.data_in(wire_d74_45),.data_out(wire_d74_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7507447(.data_in(wire_d74_46),.data_out(wire_d74_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7507448(.data_in(wire_d74_47),.data_out(wire_d74_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7507449(.data_in(wire_d74_48),.data_out(wire_d74_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7507450(.data_in(wire_d74_49),.data_out(wire_d74_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7507451(.data_in(wire_d74_50),.data_out(wire_d74_51),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7507452(.data_in(wire_d74_51),.data_out(wire_d74_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7507453(.data_in(wire_d74_52),.data_out(wire_d74_53),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7507454(.data_in(wire_d74_53),.data_out(wire_d74_54),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7507455(.data_in(wire_d74_54),.data_out(wire_d74_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7507456(.data_in(wire_d74_55),.data_out(wire_d74_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7507457(.data_in(wire_d74_56),.data_out(wire_d74_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7507458(.data_in(wire_d74_57),.data_out(wire_d74_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7507459(.data_in(wire_d74_58),.data_out(wire_d74_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7507460(.data_in(wire_d74_59),.data_out(wire_d74_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7507461(.data_in(wire_d74_60),.data_out(wire_d74_61),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7507462(.data_in(wire_d74_61),.data_out(wire_d74_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7507463(.data_in(wire_d74_62),.data_out(wire_d74_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7507464(.data_in(wire_d74_63),.data_out(wire_d74_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7507465(.data_in(wire_d74_64),.data_out(wire_d74_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7507466(.data_in(wire_d74_65),.data_out(wire_d74_66),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7507467(.data_in(wire_d74_66),.data_out(wire_d74_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7507468(.data_in(wire_d74_67),.data_out(wire_d74_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7507469(.data_in(wire_d74_68),.data_out(wire_d74_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7507470(.data_in(wire_d74_69),.data_out(wire_d74_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7507471(.data_in(wire_d74_70),.data_out(wire_d74_71),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7507472(.data_in(wire_d74_71),.data_out(wire_d74_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7507473(.data_in(wire_d74_72),.data_out(wire_d74_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7507474(.data_in(wire_d74_73),.data_out(wire_d74_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7507475(.data_in(wire_d74_74),.data_out(wire_d74_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7507476(.data_in(wire_d74_75),.data_out(wire_d74_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7507477(.data_in(wire_d74_76),.data_out(wire_d74_77),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7507478(.data_in(wire_d74_77),.data_out(wire_d74_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7507479(.data_in(wire_d74_78),.data_out(d_out74),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance760750(.data_in(d_in75),.data_out(wire_d75_0),.clk(clk),.rst(rst));            //channel 76
	decoder_top #(.WIDTH(WIDTH)) decoder_instance760751(.data_in(wire_d75_0),.data_out(wire_d75_1),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance760752(.data_in(wire_d75_1),.data_out(wire_d75_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance760753(.data_in(wire_d75_2),.data_out(wire_d75_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance760754(.data_in(wire_d75_3),.data_out(wire_d75_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance760755(.data_in(wire_d75_4),.data_out(wire_d75_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance760756(.data_in(wire_d75_5),.data_out(wire_d75_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance760757(.data_in(wire_d75_6),.data_out(wire_d75_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance760758(.data_in(wire_d75_7),.data_out(wire_d75_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance760759(.data_in(wire_d75_8),.data_out(wire_d75_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7607510(.data_in(wire_d75_9),.data_out(wire_d75_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7607511(.data_in(wire_d75_10),.data_out(wire_d75_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7607512(.data_in(wire_d75_11),.data_out(wire_d75_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7607513(.data_in(wire_d75_12),.data_out(wire_d75_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7607514(.data_in(wire_d75_13),.data_out(wire_d75_14),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7607515(.data_in(wire_d75_14),.data_out(wire_d75_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7607516(.data_in(wire_d75_15),.data_out(wire_d75_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7607517(.data_in(wire_d75_16),.data_out(wire_d75_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7607518(.data_in(wire_d75_17),.data_out(wire_d75_18),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7607519(.data_in(wire_d75_18),.data_out(wire_d75_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7607520(.data_in(wire_d75_19),.data_out(wire_d75_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7607521(.data_in(wire_d75_20),.data_out(wire_d75_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7607522(.data_in(wire_d75_21),.data_out(wire_d75_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7607523(.data_in(wire_d75_22),.data_out(wire_d75_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7607524(.data_in(wire_d75_23),.data_out(wire_d75_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7607525(.data_in(wire_d75_24),.data_out(wire_d75_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7607526(.data_in(wire_d75_25),.data_out(wire_d75_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7607527(.data_in(wire_d75_26),.data_out(wire_d75_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7607528(.data_in(wire_d75_27),.data_out(wire_d75_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7607529(.data_in(wire_d75_28),.data_out(wire_d75_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7607530(.data_in(wire_d75_29),.data_out(wire_d75_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7607531(.data_in(wire_d75_30),.data_out(wire_d75_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7607532(.data_in(wire_d75_31),.data_out(wire_d75_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7607533(.data_in(wire_d75_32),.data_out(wire_d75_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7607534(.data_in(wire_d75_33),.data_out(wire_d75_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7607535(.data_in(wire_d75_34),.data_out(wire_d75_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7607536(.data_in(wire_d75_35),.data_out(wire_d75_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7607537(.data_in(wire_d75_36),.data_out(wire_d75_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7607538(.data_in(wire_d75_37),.data_out(wire_d75_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7607539(.data_in(wire_d75_38),.data_out(wire_d75_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7607540(.data_in(wire_d75_39),.data_out(wire_d75_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7607541(.data_in(wire_d75_40),.data_out(wire_d75_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7607542(.data_in(wire_d75_41),.data_out(wire_d75_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7607543(.data_in(wire_d75_42),.data_out(wire_d75_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7607544(.data_in(wire_d75_43),.data_out(wire_d75_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7607545(.data_in(wire_d75_44),.data_out(wire_d75_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7607546(.data_in(wire_d75_45),.data_out(wire_d75_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7607547(.data_in(wire_d75_46),.data_out(wire_d75_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7607548(.data_in(wire_d75_47),.data_out(wire_d75_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7607549(.data_in(wire_d75_48),.data_out(wire_d75_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7607550(.data_in(wire_d75_49),.data_out(wire_d75_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7607551(.data_in(wire_d75_50),.data_out(wire_d75_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7607552(.data_in(wire_d75_51),.data_out(wire_d75_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7607553(.data_in(wire_d75_52),.data_out(wire_d75_53),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7607554(.data_in(wire_d75_53),.data_out(wire_d75_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7607555(.data_in(wire_d75_54),.data_out(wire_d75_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7607556(.data_in(wire_d75_55),.data_out(wire_d75_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7607557(.data_in(wire_d75_56),.data_out(wire_d75_57),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7607558(.data_in(wire_d75_57),.data_out(wire_d75_58),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7607559(.data_in(wire_d75_58),.data_out(wire_d75_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7607560(.data_in(wire_d75_59),.data_out(wire_d75_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7607561(.data_in(wire_d75_60),.data_out(wire_d75_61),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7607562(.data_in(wire_d75_61),.data_out(wire_d75_62),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7607563(.data_in(wire_d75_62),.data_out(wire_d75_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7607564(.data_in(wire_d75_63),.data_out(wire_d75_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7607565(.data_in(wire_d75_64),.data_out(wire_d75_65),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7607566(.data_in(wire_d75_65),.data_out(wire_d75_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7607567(.data_in(wire_d75_66),.data_out(wire_d75_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7607568(.data_in(wire_d75_67),.data_out(wire_d75_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7607569(.data_in(wire_d75_68),.data_out(wire_d75_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7607570(.data_in(wire_d75_69),.data_out(wire_d75_70),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7607571(.data_in(wire_d75_70),.data_out(wire_d75_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7607572(.data_in(wire_d75_71),.data_out(wire_d75_72),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7607573(.data_in(wire_d75_72),.data_out(wire_d75_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7607574(.data_in(wire_d75_73),.data_out(wire_d75_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7607575(.data_in(wire_d75_74),.data_out(wire_d75_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7607576(.data_in(wire_d75_75),.data_out(wire_d75_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7607577(.data_in(wire_d75_76),.data_out(wire_d75_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7607578(.data_in(wire_d75_77),.data_out(wire_d75_78),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7607579(.data_in(wire_d75_78),.data_out(d_out75),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance770760(.data_in(d_in76),.data_out(wire_d76_0),.clk(clk),.rst(rst));            //channel 77
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance770761(.data_in(wire_d76_0),.data_out(wire_d76_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance770762(.data_in(wire_d76_1),.data_out(wire_d76_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance770763(.data_in(wire_d76_2),.data_out(wire_d76_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance770764(.data_in(wire_d76_3),.data_out(wire_d76_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance770765(.data_in(wire_d76_4),.data_out(wire_d76_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance770766(.data_in(wire_d76_5),.data_out(wire_d76_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance770767(.data_in(wire_d76_6),.data_out(wire_d76_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance770768(.data_in(wire_d76_7),.data_out(wire_d76_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance770769(.data_in(wire_d76_8),.data_out(wire_d76_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7707610(.data_in(wire_d76_9),.data_out(wire_d76_10),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7707611(.data_in(wire_d76_10),.data_out(wire_d76_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7707612(.data_in(wire_d76_11),.data_out(wire_d76_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7707613(.data_in(wire_d76_12),.data_out(wire_d76_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7707614(.data_in(wire_d76_13),.data_out(wire_d76_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7707615(.data_in(wire_d76_14),.data_out(wire_d76_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7707616(.data_in(wire_d76_15),.data_out(wire_d76_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7707617(.data_in(wire_d76_16),.data_out(wire_d76_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7707618(.data_in(wire_d76_17),.data_out(wire_d76_18),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7707619(.data_in(wire_d76_18),.data_out(wire_d76_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7707620(.data_in(wire_d76_19),.data_out(wire_d76_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7707621(.data_in(wire_d76_20),.data_out(wire_d76_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7707622(.data_in(wire_d76_21),.data_out(wire_d76_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7707623(.data_in(wire_d76_22),.data_out(wire_d76_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7707624(.data_in(wire_d76_23),.data_out(wire_d76_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7707625(.data_in(wire_d76_24),.data_out(wire_d76_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7707626(.data_in(wire_d76_25),.data_out(wire_d76_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7707627(.data_in(wire_d76_26),.data_out(wire_d76_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7707628(.data_in(wire_d76_27),.data_out(wire_d76_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7707629(.data_in(wire_d76_28),.data_out(wire_d76_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7707630(.data_in(wire_d76_29),.data_out(wire_d76_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7707631(.data_in(wire_d76_30),.data_out(wire_d76_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7707632(.data_in(wire_d76_31),.data_out(wire_d76_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7707633(.data_in(wire_d76_32),.data_out(wire_d76_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7707634(.data_in(wire_d76_33),.data_out(wire_d76_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7707635(.data_in(wire_d76_34),.data_out(wire_d76_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7707636(.data_in(wire_d76_35),.data_out(wire_d76_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7707637(.data_in(wire_d76_36),.data_out(wire_d76_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7707638(.data_in(wire_d76_37),.data_out(wire_d76_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7707639(.data_in(wire_d76_38),.data_out(wire_d76_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7707640(.data_in(wire_d76_39),.data_out(wire_d76_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7707641(.data_in(wire_d76_40),.data_out(wire_d76_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7707642(.data_in(wire_d76_41),.data_out(wire_d76_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7707643(.data_in(wire_d76_42),.data_out(wire_d76_43),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7707644(.data_in(wire_d76_43),.data_out(wire_d76_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7707645(.data_in(wire_d76_44),.data_out(wire_d76_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7707646(.data_in(wire_d76_45),.data_out(wire_d76_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7707647(.data_in(wire_d76_46),.data_out(wire_d76_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7707648(.data_in(wire_d76_47),.data_out(wire_d76_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7707649(.data_in(wire_d76_48),.data_out(wire_d76_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7707650(.data_in(wire_d76_49),.data_out(wire_d76_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7707651(.data_in(wire_d76_50),.data_out(wire_d76_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7707652(.data_in(wire_d76_51),.data_out(wire_d76_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7707653(.data_in(wire_d76_52),.data_out(wire_d76_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7707654(.data_in(wire_d76_53),.data_out(wire_d76_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7707655(.data_in(wire_d76_54),.data_out(wire_d76_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7707656(.data_in(wire_d76_55),.data_out(wire_d76_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7707657(.data_in(wire_d76_56),.data_out(wire_d76_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7707658(.data_in(wire_d76_57),.data_out(wire_d76_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7707659(.data_in(wire_d76_58),.data_out(wire_d76_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7707660(.data_in(wire_d76_59),.data_out(wire_d76_60),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7707661(.data_in(wire_d76_60),.data_out(wire_d76_61),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7707662(.data_in(wire_d76_61),.data_out(wire_d76_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7707663(.data_in(wire_d76_62),.data_out(wire_d76_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7707664(.data_in(wire_d76_63),.data_out(wire_d76_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7707665(.data_in(wire_d76_64),.data_out(wire_d76_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7707666(.data_in(wire_d76_65),.data_out(wire_d76_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7707667(.data_in(wire_d76_66),.data_out(wire_d76_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7707668(.data_in(wire_d76_67),.data_out(wire_d76_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7707669(.data_in(wire_d76_68),.data_out(wire_d76_69),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7707670(.data_in(wire_d76_69),.data_out(wire_d76_70),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7707671(.data_in(wire_d76_70),.data_out(wire_d76_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7707672(.data_in(wire_d76_71),.data_out(wire_d76_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7707673(.data_in(wire_d76_72),.data_out(wire_d76_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7707674(.data_in(wire_d76_73),.data_out(wire_d76_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7707675(.data_in(wire_d76_74),.data_out(wire_d76_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7707676(.data_in(wire_d76_75),.data_out(wire_d76_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7707677(.data_in(wire_d76_76),.data_out(wire_d76_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7707678(.data_in(wire_d76_77),.data_out(wire_d76_78),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7707679(.data_in(wire_d76_78),.data_out(d_out76),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance780770(.data_in(d_in77),.data_out(wire_d77_0),.clk(clk),.rst(rst));            //channel 78
	decoder_top #(.WIDTH(WIDTH)) decoder_instance780771(.data_in(wire_d77_0),.data_out(wire_d77_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance780772(.data_in(wire_d77_1),.data_out(wire_d77_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance780773(.data_in(wire_d77_2),.data_out(wire_d77_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance780774(.data_in(wire_d77_3),.data_out(wire_d77_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance780775(.data_in(wire_d77_4),.data_out(wire_d77_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance780776(.data_in(wire_d77_5),.data_out(wire_d77_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance780777(.data_in(wire_d77_6),.data_out(wire_d77_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance780778(.data_in(wire_d77_7),.data_out(wire_d77_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance780779(.data_in(wire_d77_8),.data_out(wire_d77_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7807710(.data_in(wire_d77_9),.data_out(wire_d77_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7807711(.data_in(wire_d77_10),.data_out(wire_d77_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7807712(.data_in(wire_d77_11),.data_out(wire_d77_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7807713(.data_in(wire_d77_12),.data_out(wire_d77_13),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7807714(.data_in(wire_d77_13),.data_out(wire_d77_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7807715(.data_in(wire_d77_14),.data_out(wire_d77_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7807716(.data_in(wire_d77_15),.data_out(wire_d77_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7807717(.data_in(wire_d77_16),.data_out(wire_d77_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7807718(.data_in(wire_d77_17),.data_out(wire_d77_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7807719(.data_in(wire_d77_18),.data_out(wire_d77_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7807720(.data_in(wire_d77_19),.data_out(wire_d77_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7807721(.data_in(wire_d77_20),.data_out(wire_d77_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7807722(.data_in(wire_d77_21),.data_out(wire_d77_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7807723(.data_in(wire_d77_22),.data_out(wire_d77_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7807724(.data_in(wire_d77_23),.data_out(wire_d77_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7807725(.data_in(wire_d77_24),.data_out(wire_d77_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7807726(.data_in(wire_d77_25),.data_out(wire_d77_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7807727(.data_in(wire_d77_26),.data_out(wire_d77_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7807728(.data_in(wire_d77_27),.data_out(wire_d77_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7807729(.data_in(wire_d77_28),.data_out(wire_d77_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7807730(.data_in(wire_d77_29),.data_out(wire_d77_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7807731(.data_in(wire_d77_30),.data_out(wire_d77_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7807732(.data_in(wire_d77_31),.data_out(wire_d77_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7807733(.data_in(wire_d77_32),.data_out(wire_d77_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7807734(.data_in(wire_d77_33),.data_out(wire_d77_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7807735(.data_in(wire_d77_34),.data_out(wire_d77_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7807736(.data_in(wire_d77_35),.data_out(wire_d77_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7807737(.data_in(wire_d77_36),.data_out(wire_d77_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7807738(.data_in(wire_d77_37),.data_out(wire_d77_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7807739(.data_in(wire_d77_38),.data_out(wire_d77_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7807740(.data_in(wire_d77_39),.data_out(wire_d77_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7807741(.data_in(wire_d77_40),.data_out(wire_d77_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7807742(.data_in(wire_d77_41),.data_out(wire_d77_42),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7807743(.data_in(wire_d77_42),.data_out(wire_d77_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7807744(.data_in(wire_d77_43),.data_out(wire_d77_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7807745(.data_in(wire_d77_44),.data_out(wire_d77_45),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7807746(.data_in(wire_d77_45),.data_out(wire_d77_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7807747(.data_in(wire_d77_46),.data_out(wire_d77_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7807748(.data_in(wire_d77_47),.data_out(wire_d77_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7807749(.data_in(wire_d77_48),.data_out(wire_d77_49),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7807750(.data_in(wire_d77_49),.data_out(wire_d77_50),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7807751(.data_in(wire_d77_50),.data_out(wire_d77_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7807752(.data_in(wire_d77_51),.data_out(wire_d77_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7807753(.data_in(wire_d77_52),.data_out(wire_d77_53),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7807754(.data_in(wire_d77_53),.data_out(wire_d77_54),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7807755(.data_in(wire_d77_54),.data_out(wire_d77_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7807756(.data_in(wire_d77_55),.data_out(wire_d77_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7807757(.data_in(wire_d77_56),.data_out(wire_d77_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7807758(.data_in(wire_d77_57),.data_out(wire_d77_58),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7807759(.data_in(wire_d77_58),.data_out(wire_d77_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7807760(.data_in(wire_d77_59),.data_out(wire_d77_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7807761(.data_in(wire_d77_60),.data_out(wire_d77_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7807762(.data_in(wire_d77_61),.data_out(wire_d77_62),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7807763(.data_in(wire_d77_62),.data_out(wire_d77_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7807764(.data_in(wire_d77_63),.data_out(wire_d77_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7807765(.data_in(wire_d77_64),.data_out(wire_d77_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7807766(.data_in(wire_d77_65),.data_out(wire_d77_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7807767(.data_in(wire_d77_66),.data_out(wire_d77_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7807768(.data_in(wire_d77_67),.data_out(wire_d77_68),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7807769(.data_in(wire_d77_68),.data_out(wire_d77_69),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7807770(.data_in(wire_d77_69),.data_out(wire_d77_70),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7807771(.data_in(wire_d77_70),.data_out(wire_d77_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7807772(.data_in(wire_d77_71),.data_out(wire_d77_72),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7807773(.data_in(wire_d77_72),.data_out(wire_d77_73),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7807774(.data_in(wire_d77_73),.data_out(wire_d77_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7807775(.data_in(wire_d77_74),.data_out(wire_d77_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7807776(.data_in(wire_d77_75),.data_out(wire_d77_76),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7807777(.data_in(wire_d77_76),.data_out(wire_d77_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7807778(.data_in(wire_d77_77),.data_out(wire_d77_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7807779(.data_in(wire_d77_78),.data_out(d_out77),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance790780(.data_in(d_in78),.data_out(wire_d78_0),.clk(clk),.rst(rst));            //channel 79
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance790781(.data_in(wire_d78_0),.data_out(wire_d78_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance790782(.data_in(wire_d78_1),.data_out(wire_d78_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance790783(.data_in(wire_d78_2),.data_out(wire_d78_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance790784(.data_in(wire_d78_3),.data_out(wire_d78_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance790785(.data_in(wire_d78_4),.data_out(wire_d78_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance790786(.data_in(wire_d78_5),.data_out(wire_d78_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance790787(.data_in(wire_d78_6),.data_out(wire_d78_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance790788(.data_in(wire_d78_7),.data_out(wire_d78_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance790789(.data_in(wire_d78_8),.data_out(wire_d78_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7907810(.data_in(wire_d78_9),.data_out(wire_d78_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7907811(.data_in(wire_d78_10),.data_out(wire_d78_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7907812(.data_in(wire_d78_11),.data_out(wire_d78_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7907813(.data_in(wire_d78_12),.data_out(wire_d78_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7907814(.data_in(wire_d78_13),.data_out(wire_d78_14),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7907815(.data_in(wire_d78_14),.data_out(wire_d78_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7907816(.data_in(wire_d78_15),.data_out(wire_d78_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7907817(.data_in(wire_d78_16),.data_out(wire_d78_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7907818(.data_in(wire_d78_17),.data_out(wire_d78_18),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7907819(.data_in(wire_d78_18),.data_out(wire_d78_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7907820(.data_in(wire_d78_19),.data_out(wire_d78_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7907821(.data_in(wire_d78_20),.data_out(wire_d78_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7907822(.data_in(wire_d78_21),.data_out(wire_d78_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7907823(.data_in(wire_d78_22),.data_out(wire_d78_23),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7907824(.data_in(wire_d78_23),.data_out(wire_d78_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7907825(.data_in(wire_d78_24),.data_out(wire_d78_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7907826(.data_in(wire_d78_25),.data_out(wire_d78_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7907827(.data_in(wire_d78_26),.data_out(wire_d78_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7907828(.data_in(wire_d78_27),.data_out(wire_d78_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7907829(.data_in(wire_d78_28),.data_out(wire_d78_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7907830(.data_in(wire_d78_29),.data_out(wire_d78_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7907831(.data_in(wire_d78_30),.data_out(wire_d78_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7907832(.data_in(wire_d78_31),.data_out(wire_d78_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7907833(.data_in(wire_d78_32),.data_out(wire_d78_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7907834(.data_in(wire_d78_33),.data_out(wire_d78_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7907835(.data_in(wire_d78_34),.data_out(wire_d78_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7907836(.data_in(wire_d78_35),.data_out(wire_d78_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7907837(.data_in(wire_d78_36),.data_out(wire_d78_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7907838(.data_in(wire_d78_37),.data_out(wire_d78_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7907839(.data_in(wire_d78_38),.data_out(wire_d78_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7907840(.data_in(wire_d78_39),.data_out(wire_d78_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7907841(.data_in(wire_d78_40),.data_out(wire_d78_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7907842(.data_in(wire_d78_41),.data_out(wire_d78_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7907843(.data_in(wire_d78_42),.data_out(wire_d78_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7907844(.data_in(wire_d78_43),.data_out(wire_d78_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7907845(.data_in(wire_d78_44),.data_out(wire_d78_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7907846(.data_in(wire_d78_45),.data_out(wire_d78_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7907847(.data_in(wire_d78_46),.data_out(wire_d78_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7907848(.data_in(wire_d78_47),.data_out(wire_d78_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7907849(.data_in(wire_d78_48),.data_out(wire_d78_49),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7907850(.data_in(wire_d78_49),.data_out(wire_d78_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7907851(.data_in(wire_d78_50),.data_out(wire_d78_51),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7907852(.data_in(wire_d78_51),.data_out(wire_d78_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7907853(.data_in(wire_d78_52),.data_out(wire_d78_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7907854(.data_in(wire_d78_53),.data_out(wire_d78_54),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7907855(.data_in(wire_d78_54),.data_out(wire_d78_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7907856(.data_in(wire_d78_55),.data_out(wire_d78_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7907857(.data_in(wire_d78_56),.data_out(wire_d78_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7907858(.data_in(wire_d78_57),.data_out(wire_d78_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7907859(.data_in(wire_d78_58),.data_out(wire_d78_59),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7907860(.data_in(wire_d78_59),.data_out(wire_d78_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7907861(.data_in(wire_d78_60),.data_out(wire_d78_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7907862(.data_in(wire_d78_61),.data_out(wire_d78_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7907863(.data_in(wire_d78_62),.data_out(wire_d78_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7907864(.data_in(wire_d78_63),.data_out(wire_d78_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7907865(.data_in(wire_d78_64),.data_out(wire_d78_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7907866(.data_in(wire_d78_65),.data_out(wire_d78_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7907867(.data_in(wire_d78_66),.data_out(wire_d78_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7907868(.data_in(wire_d78_67),.data_out(wire_d78_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7907869(.data_in(wire_d78_68),.data_out(wire_d78_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7907870(.data_in(wire_d78_69),.data_out(wire_d78_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7907871(.data_in(wire_d78_70),.data_out(wire_d78_71),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7907872(.data_in(wire_d78_71),.data_out(wire_d78_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7907873(.data_in(wire_d78_72),.data_out(wire_d78_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7907874(.data_in(wire_d78_73),.data_out(wire_d78_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7907875(.data_in(wire_d78_74),.data_out(wire_d78_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7907876(.data_in(wire_d78_75),.data_out(wire_d78_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7907877(.data_in(wire_d78_76),.data_out(wire_d78_77),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7907878(.data_in(wire_d78_77),.data_out(wire_d78_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7907879(.data_in(wire_d78_78),.data_out(d_out78),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance800790(.data_in(d_in79),.data_out(wire_d79_0),.clk(clk),.rst(rst));            //channel 80
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance800791(.data_in(wire_d79_0),.data_out(wire_d79_1),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance800792(.data_in(wire_d79_1),.data_out(wire_d79_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance800793(.data_in(wire_d79_2),.data_out(wire_d79_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance800794(.data_in(wire_d79_3),.data_out(wire_d79_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance800795(.data_in(wire_d79_4),.data_out(wire_d79_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance800796(.data_in(wire_d79_5),.data_out(wire_d79_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance800797(.data_in(wire_d79_6),.data_out(wire_d79_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance800798(.data_in(wire_d79_7),.data_out(wire_d79_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance800799(.data_in(wire_d79_8),.data_out(wire_d79_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8007910(.data_in(wire_d79_9),.data_out(wire_d79_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8007911(.data_in(wire_d79_10),.data_out(wire_d79_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8007912(.data_in(wire_d79_11),.data_out(wire_d79_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8007913(.data_in(wire_d79_12),.data_out(wire_d79_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8007914(.data_in(wire_d79_13),.data_out(wire_d79_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8007915(.data_in(wire_d79_14),.data_out(wire_d79_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8007916(.data_in(wire_d79_15),.data_out(wire_d79_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8007917(.data_in(wire_d79_16),.data_out(wire_d79_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8007918(.data_in(wire_d79_17),.data_out(wire_d79_18),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8007919(.data_in(wire_d79_18),.data_out(wire_d79_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8007920(.data_in(wire_d79_19),.data_out(wire_d79_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8007921(.data_in(wire_d79_20),.data_out(wire_d79_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8007922(.data_in(wire_d79_21),.data_out(wire_d79_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8007923(.data_in(wire_d79_22),.data_out(wire_d79_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8007924(.data_in(wire_d79_23),.data_out(wire_d79_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8007925(.data_in(wire_d79_24),.data_out(wire_d79_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8007926(.data_in(wire_d79_25),.data_out(wire_d79_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8007927(.data_in(wire_d79_26),.data_out(wire_d79_27),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8007928(.data_in(wire_d79_27),.data_out(wire_d79_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8007929(.data_in(wire_d79_28),.data_out(wire_d79_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8007930(.data_in(wire_d79_29),.data_out(wire_d79_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8007931(.data_in(wire_d79_30),.data_out(wire_d79_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8007932(.data_in(wire_d79_31),.data_out(wire_d79_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8007933(.data_in(wire_d79_32),.data_out(wire_d79_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8007934(.data_in(wire_d79_33),.data_out(wire_d79_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8007935(.data_in(wire_d79_34),.data_out(wire_d79_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8007936(.data_in(wire_d79_35),.data_out(wire_d79_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8007937(.data_in(wire_d79_36),.data_out(wire_d79_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8007938(.data_in(wire_d79_37),.data_out(wire_d79_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8007939(.data_in(wire_d79_38),.data_out(wire_d79_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8007940(.data_in(wire_d79_39),.data_out(wire_d79_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8007941(.data_in(wire_d79_40),.data_out(wire_d79_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8007942(.data_in(wire_d79_41),.data_out(wire_d79_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8007943(.data_in(wire_d79_42),.data_out(wire_d79_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8007944(.data_in(wire_d79_43),.data_out(wire_d79_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8007945(.data_in(wire_d79_44),.data_out(wire_d79_45),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8007946(.data_in(wire_d79_45),.data_out(wire_d79_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8007947(.data_in(wire_d79_46),.data_out(wire_d79_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8007948(.data_in(wire_d79_47),.data_out(wire_d79_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8007949(.data_in(wire_d79_48),.data_out(wire_d79_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8007950(.data_in(wire_d79_49),.data_out(wire_d79_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8007951(.data_in(wire_d79_50),.data_out(wire_d79_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8007952(.data_in(wire_d79_51),.data_out(wire_d79_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8007953(.data_in(wire_d79_52),.data_out(wire_d79_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8007954(.data_in(wire_d79_53),.data_out(wire_d79_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8007955(.data_in(wire_d79_54),.data_out(wire_d79_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8007956(.data_in(wire_d79_55),.data_out(wire_d79_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8007957(.data_in(wire_d79_56),.data_out(wire_d79_57),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8007958(.data_in(wire_d79_57),.data_out(wire_d79_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8007959(.data_in(wire_d79_58),.data_out(wire_d79_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8007960(.data_in(wire_d79_59),.data_out(wire_d79_60),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8007961(.data_in(wire_d79_60),.data_out(wire_d79_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8007962(.data_in(wire_d79_61),.data_out(wire_d79_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8007963(.data_in(wire_d79_62),.data_out(wire_d79_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8007964(.data_in(wire_d79_63),.data_out(wire_d79_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8007965(.data_in(wire_d79_64),.data_out(wire_d79_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8007966(.data_in(wire_d79_65),.data_out(wire_d79_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8007967(.data_in(wire_d79_66),.data_out(wire_d79_67),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8007968(.data_in(wire_d79_67),.data_out(wire_d79_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8007969(.data_in(wire_d79_68),.data_out(wire_d79_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8007970(.data_in(wire_d79_69),.data_out(wire_d79_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8007971(.data_in(wire_d79_70),.data_out(wire_d79_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8007972(.data_in(wire_d79_71),.data_out(wire_d79_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8007973(.data_in(wire_d79_72),.data_out(wire_d79_73),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8007974(.data_in(wire_d79_73),.data_out(wire_d79_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8007975(.data_in(wire_d79_74),.data_out(wire_d79_75),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8007976(.data_in(wire_d79_75),.data_out(wire_d79_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8007977(.data_in(wire_d79_76),.data_out(wire_d79_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8007978(.data_in(wire_d79_77),.data_out(wire_d79_78),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8007979(.data_in(wire_d79_78),.data_out(d_out79),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance810800(.data_in(d_in80),.data_out(wire_d80_0),.clk(clk),.rst(rst));            //channel 81
	register #(.WIDTH(WIDTH)) register_instance810801(.data_in(wire_d80_0),.data_out(wire_d80_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance810802(.data_in(wire_d80_1),.data_out(wire_d80_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance810803(.data_in(wire_d80_2),.data_out(wire_d80_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance810804(.data_in(wire_d80_3),.data_out(wire_d80_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance810805(.data_in(wire_d80_4),.data_out(wire_d80_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance810806(.data_in(wire_d80_5),.data_out(wire_d80_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance810807(.data_in(wire_d80_6),.data_out(wire_d80_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance810808(.data_in(wire_d80_7),.data_out(wire_d80_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance810809(.data_in(wire_d80_8),.data_out(wire_d80_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8108010(.data_in(wire_d80_9),.data_out(wire_d80_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8108011(.data_in(wire_d80_10),.data_out(wire_d80_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8108012(.data_in(wire_d80_11),.data_out(wire_d80_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8108013(.data_in(wire_d80_12),.data_out(wire_d80_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8108014(.data_in(wire_d80_13),.data_out(wire_d80_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8108015(.data_in(wire_d80_14),.data_out(wire_d80_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8108016(.data_in(wire_d80_15),.data_out(wire_d80_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8108017(.data_in(wire_d80_16),.data_out(wire_d80_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8108018(.data_in(wire_d80_17),.data_out(wire_d80_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8108019(.data_in(wire_d80_18),.data_out(wire_d80_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8108020(.data_in(wire_d80_19),.data_out(wire_d80_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8108021(.data_in(wire_d80_20),.data_out(wire_d80_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8108022(.data_in(wire_d80_21),.data_out(wire_d80_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8108023(.data_in(wire_d80_22),.data_out(wire_d80_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8108024(.data_in(wire_d80_23),.data_out(wire_d80_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8108025(.data_in(wire_d80_24),.data_out(wire_d80_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8108026(.data_in(wire_d80_25),.data_out(wire_d80_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8108027(.data_in(wire_d80_26),.data_out(wire_d80_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8108028(.data_in(wire_d80_27),.data_out(wire_d80_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8108029(.data_in(wire_d80_28),.data_out(wire_d80_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8108030(.data_in(wire_d80_29),.data_out(wire_d80_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8108031(.data_in(wire_d80_30),.data_out(wire_d80_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8108032(.data_in(wire_d80_31),.data_out(wire_d80_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8108033(.data_in(wire_d80_32),.data_out(wire_d80_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8108034(.data_in(wire_d80_33),.data_out(wire_d80_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8108035(.data_in(wire_d80_34),.data_out(wire_d80_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8108036(.data_in(wire_d80_35),.data_out(wire_d80_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8108037(.data_in(wire_d80_36),.data_out(wire_d80_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8108038(.data_in(wire_d80_37),.data_out(wire_d80_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8108039(.data_in(wire_d80_38),.data_out(wire_d80_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8108040(.data_in(wire_d80_39),.data_out(wire_d80_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8108041(.data_in(wire_d80_40),.data_out(wire_d80_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8108042(.data_in(wire_d80_41),.data_out(wire_d80_42),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8108043(.data_in(wire_d80_42),.data_out(wire_d80_43),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8108044(.data_in(wire_d80_43),.data_out(wire_d80_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8108045(.data_in(wire_d80_44),.data_out(wire_d80_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8108046(.data_in(wire_d80_45),.data_out(wire_d80_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8108047(.data_in(wire_d80_46),.data_out(wire_d80_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8108048(.data_in(wire_d80_47),.data_out(wire_d80_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8108049(.data_in(wire_d80_48),.data_out(wire_d80_49),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8108050(.data_in(wire_d80_49),.data_out(wire_d80_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8108051(.data_in(wire_d80_50),.data_out(wire_d80_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8108052(.data_in(wire_d80_51),.data_out(wire_d80_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8108053(.data_in(wire_d80_52),.data_out(wire_d80_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8108054(.data_in(wire_d80_53),.data_out(wire_d80_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8108055(.data_in(wire_d80_54),.data_out(wire_d80_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8108056(.data_in(wire_d80_55),.data_out(wire_d80_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8108057(.data_in(wire_d80_56),.data_out(wire_d80_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8108058(.data_in(wire_d80_57),.data_out(wire_d80_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8108059(.data_in(wire_d80_58),.data_out(wire_d80_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8108060(.data_in(wire_d80_59),.data_out(wire_d80_60),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8108061(.data_in(wire_d80_60),.data_out(wire_d80_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8108062(.data_in(wire_d80_61),.data_out(wire_d80_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8108063(.data_in(wire_d80_62),.data_out(wire_d80_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8108064(.data_in(wire_d80_63),.data_out(wire_d80_64),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8108065(.data_in(wire_d80_64),.data_out(wire_d80_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8108066(.data_in(wire_d80_65),.data_out(wire_d80_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8108067(.data_in(wire_d80_66),.data_out(wire_d80_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8108068(.data_in(wire_d80_67),.data_out(wire_d80_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8108069(.data_in(wire_d80_68),.data_out(wire_d80_69),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8108070(.data_in(wire_d80_69),.data_out(wire_d80_70),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8108071(.data_in(wire_d80_70),.data_out(wire_d80_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8108072(.data_in(wire_d80_71),.data_out(wire_d80_72),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8108073(.data_in(wire_d80_72),.data_out(wire_d80_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8108074(.data_in(wire_d80_73),.data_out(wire_d80_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8108075(.data_in(wire_d80_74),.data_out(wire_d80_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8108076(.data_in(wire_d80_75),.data_out(wire_d80_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8108077(.data_in(wire_d80_76),.data_out(wire_d80_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8108078(.data_in(wire_d80_77),.data_out(wire_d80_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8108079(.data_in(wire_d80_78),.data_out(d_out80),.clk(clk),.rst(rst));

	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance820810(.data_in(d_in81),.data_out(wire_d81_0),.clk(clk),.rst(rst));            //channel 82
	large_mux #(.WIDTH(WIDTH)) large_mux_instance820811(.data_in(wire_d81_0),.data_out(wire_d81_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance820812(.data_in(wire_d81_1),.data_out(wire_d81_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance820813(.data_in(wire_d81_2),.data_out(wire_d81_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance820814(.data_in(wire_d81_3),.data_out(wire_d81_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance820815(.data_in(wire_d81_4),.data_out(wire_d81_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance820816(.data_in(wire_d81_5),.data_out(wire_d81_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance820817(.data_in(wire_d81_6),.data_out(wire_d81_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance820818(.data_in(wire_d81_7),.data_out(wire_d81_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance820819(.data_in(wire_d81_8),.data_out(wire_d81_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8208110(.data_in(wire_d81_9),.data_out(wire_d81_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8208111(.data_in(wire_d81_10),.data_out(wire_d81_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8208112(.data_in(wire_d81_11),.data_out(wire_d81_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8208113(.data_in(wire_d81_12),.data_out(wire_d81_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8208114(.data_in(wire_d81_13),.data_out(wire_d81_14),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8208115(.data_in(wire_d81_14),.data_out(wire_d81_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8208116(.data_in(wire_d81_15),.data_out(wire_d81_16),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8208117(.data_in(wire_d81_16),.data_out(wire_d81_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8208118(.data_in(wire_d81_17),.data_out(wire_d81_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8208119(.data_in(wire_d81_18),.data_out(wire_d81_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8208120(.data_in(wire_d81_19),.data_out(wire_d81_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8208121(.data_in(wire_d81_20),.data_out(wire_d81_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8208122(.data_in(wire_d81_21),.data_out(wire_d81_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8208123(.data_in(wire_d81_22),.data_out(wire_d81_23),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8208124(.data_in(wire_d81_23),.data_out(wire_d81_24),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8208125(.data_in(wire_d81_24),.data_out(wire_d81_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8208126(.data_in(wire_d81_25),.data_out(wire_d81_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8208127(.data_in(wire_d81_26),.data_out(wire_d81_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8208128(.data_in(wire_d81_27),.data_out(wire_d81_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8208129(.data_in(wire_d81_28),.data_out(wire_d81_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8208130(.data_in(wire_d81_29),.data_out(wire_d81_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8208131(.data_in(wire_d81_30),.data_out(wire_d81_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8208132(.data_in(wire_d81_31),.data_out(wire_d81_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8208133(.data_in(wire_d81_32),.data_out(wire_d81_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8208134(.data_in(wire_d81_33),.data_out(wire_d81_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8208135(.data_in(wire_d81_34),.data_out(wire_d81_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8208136(.data_in(wire_d81_35),.data_out(wire_d81_36),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8208137(.data_in(wire_d81_36),.data_out(wire_d81_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8208138(.data_in(wire_d81_37),.data_out(wire_d81_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8208139(.data_in(wire_d81_38),.data_out(wire_d81_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8208140(.data_in(wire_d81_39),.data_out(wire_d81_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8208141(.data_in(wire_d81_40),.data_out(wire_d81_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8208142(.data_in(wire_d81_41),.data_out(wire_d81_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8208143(.data_in(wire_d81_42),.data_out(wire_d81_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8208144(.data_in(wire_d81_43),.data_out(wire_d81_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8208145(.data_in(wire_d81_44),.data_out(wire_d81_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8208146(.data_in(wire_d81_45),.data_out(wire_d81_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8208147(.data_in(wire_d81_46),.data_out(wire_d81_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8208148(.data_in(wire_d81_47),.data_out(wire_d81_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8208149(.data_in(wire_d81_48),.data_out(wire_d81_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8208150(.data_in(wire_d81_49),.data_out(wire_d81_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8208151(.data_in(wire_d81_50),.data_out(wire_d81_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8208152(.data_in(wire_d81_51),.data_out(wire_d81_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8208153(.data_in(wire_d81_52),.data_out(wire_d81_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8208154(.data_in(wire_d81_53),.data_out(wire_d81_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8208155(.data_in(wire_d81_54),.data_out(wire_d81_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8208156(.data_in(wire_d81_55),.data_out(wire_d81_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8208157(.data_in(wire_d81_56),.data_out(wire_d81_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8208158(.data_in(wire_d81_57),.data_out(wire_d81_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8208159(.data_in(wire_d81_58),.data_out(wire_d81_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8208160(.data_in(wire_d81_59),.data_out(wire_d81_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8208161(.data_in(wire_d81_60),.data_out(wire_d81_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8208162(.data_in(wire_d81_61),.data_out(wire_d81_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8208163(.data_in(wire_d81_62),.data_out(wire_d81_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8208164(.data_in(wire_d81_63),.data_out(wire_d81_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8208165(.data_in(wire_d81_64),.data_out(wire_d81_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8208166(.data_in(wire_d81_65),.data_out(wire_d81_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8208167(.data_in(wire_d81_66),.data_out(wire_d81_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8208168(.data_in(wire_d81_67),.data_out(wire_d81_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8208169(.data_in(wire_d81_68),.data_out(wire_d81_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8208170(.data_in(wire_d81_69),.data_out(wire_d81_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8208171(.data_in(wire_d81_70),.data_out(wire_d81_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8208172(.data_in(wire_d81_71),.data_out(wire_d81_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8208173(.data_in(wire_d81_72),.data_out(wire_d81_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8208174(.data_in(wire_d81_73),.data_out(wire_d81_74),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8208175(.data_in(wire_d81_74),.data_out(wire_d81_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8208176(.data_in(wire_d81_75),.data_out(wire_d81_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8208177(.data_in(wire_d81_76),.data_out(wire_d81_77),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8208178(.data_in(wire_d81_77),.data_out(wire_d81_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8208179(.data_in(wire_d81_78),.data_out(d_out81),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance830820(.data_in(d_in82),.data_out(wire_d82_0),.clk(clk),.rst(rst));            //channel 83
	register #(.WIDTH(WIDTH)) register_instance830821(.data_in(wire_d82_0),.data_out(wire_d82_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance830822(.data_in(wire_d82_1),.data_out(wire_d82_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance830823(.data_in(wire_d82_2),.data_out(wire_d82_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance830824(.data_in(wire_d82_3),.data_out(wire_d82_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance830825(.data_in(wire_d82_4),.data_out(wire_d82_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance830826(.data_in(wire_d82_5),.data_out(wire_d82_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance830827(.data_in(wire_d82_6),.data_out(wire_d82_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance830828(.data_in(wire_d82_7),.data_out(wire_d82_8),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance830829(.data_in(wire_d82_8),.data_out(wire_d82_9),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8308210(.data_in(wire_d82_9),.data_out(wire_d82_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8308211(.data_in(wire_d82_10),.data_out(wire_d82_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8308212(.data_in(wire_d82_11),.data_out(wire_d82_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8308213(.data_in(wire_d82_12),.data_out(wire_d82_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8308214(.data_in(wire_d82_13),.data_out(wire_d82_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8308215(.data_in(wire_d82_14),.data_out(wire_d82_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8308216(.data_in(wire_d82_15),.data_out(wire_d82_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8308217(.data_in(wire_d82_16),.data_out(wire_d82_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8308218(.data_in(wire_d82_17),.data_out(wire_d82_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8308219(.data_in(wire_d82_18),.data_out(wire_d82_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8308220(.data_in(wire_d82_19),.data_out(wire_d82_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8308221(.data_in(wire_d82_20),.data_out(wire_d82_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8308222(.data_in(wire_d82_21),.data_out(wire_d82_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8308223(.data_in(wire_d82_22),.data_out(wire_d82_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8308224(.data_in(wire_d82_23),.data_out(wire_d82_24),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8308225(.data_in(wire_d82_24),.data_out(wire_d82_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8308226(.data_in(wire_d82_25),.data_out(wire_d82_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8308227(.data_in(wire_d82_26),.data_out(wire_d82_27),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8308228(.data_in(wire_d82_27),.data_out(wire_d82_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8308229(.data_in(wire_d82_28),.data_out(wire_d82_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8308230(.data_in(wire_d82_29),.data_out(wire_d82_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8308231(.data_in(wire_d82_30),.data_out(wire_d82_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8308232(.data_in(wire_d82_31),.data_out(wire_d82_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8308233(.data_in(wire_d82_32),.data_out(wire_d82_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8308234(.data_in(wire_d82_33),.data_out(wire_d82_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8308235(.data_in(wire_d82_34),.data_out(wire_d82_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8308236(.data_in(wire_d82_35),.data_out(wire_d82_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8308237(.data_in(wire_d82_36),.data_out(wire_d82_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8308238(.data_in(wire_d82_37),.data_out(wire_d82_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8308239(.data_in(wire_d82_38),.data_out(wire_d82_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8308240(.data_in(wire_d82_39),.data_out(wire_d82_40),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8308241(.data_in(wire_d82_40),.data_out(wire_d82_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8308242(.data_in(wire_d82_41),.data_out(wire_d82_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8308243(.data_in(wire_d82_42),.data_out(wire_d82_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8308244(.data_in(wire_d82_43),.data_out(wire_d82_44),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8308245(.data_in(wire_d82_44),.data_out(wire_d82_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8308246(.data_in(wire_d82_45),.data_out(wire_d82_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8308247(.data_in(wire_d82_46),.data_out(wire_d82_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8308248(.data_in(wire_d82_47),.data_out(wire_d82_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8308249(.data_in(wire_d82_48),.data_out(wire_d82_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8308250(.data_in(wire_d82_49),.data_out(wire_d82_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8308251(.data_in(wire_d82_50),.data_out(wire_d82_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8308252(.data_in(wire_d82_51),.data_out(wire_d82_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8308253(.data_in(wire_d82_52),.data_out(wire_d82_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8308254(.data_in(wire_d82_53),.data_out(wire_d82_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8308255(.data_in(wire_d82_54),.data_out(wire_d82_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8308256(.data_in(wire_d82_55),.data_out(wire_d82_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8308257(.data_in(wire_d82_56),.data_out(wire_d82_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8308258(.data_in(wire_d82_57),.data_out(wire_d82_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8308259(.data_in(wire_d82_58),.data_out(wire_d82_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8308260(.data_in(wire_d82_59),.data_out(wire_d82_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8308261(.data_in(wire_d82_60),.data_out(wire_d82_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8308262(.data_in(wire_d82_61),.data_out(wire_d82_62),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8308263(.data_in(wire_d82_62),.data_out(wire_d82_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8308264(.data_in(wire_d82_63),.data_out(wire_d82_64),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8308265(.data_in(wire_d82_64),.data_out(wire_d82_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8308266(.data_in(wire_d82_65),.data_out(wire_d82_66),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8308267(.data_in(wire_d82_66),.data_out(wire_d82_67),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8308268(.data_in(wire_d82_67),.data_out(wire_d82_68),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8308269(.data_in(wire_d82_68),.data_out(wire_d82_69),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8308270(.data_in(wire_d82_69),.data_out(wire_d82_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8308271(.data_in(wire_d82_70),.data_out(wire_d82_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8308272(.data_in(wire_d82_71),.data_out(wire_d82_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8308273(.data_in(wire_d82_72),.data_out(wire_d82_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8308274(.data_in(wire_d82_73),.data_out(wire_d82_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8308275(.data_in(wire_d82_74),.data_out(wire_d82_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8308276(.data_in(wire_d82_75),.data_out(wire_d82_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8308277(.data_in(wire_d82_76),.data_out(wire_d82_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8308278(.data_in(wire_d82_77),.data_out(wire_d82_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8308279(.data_in(wire_d82_78),.data_out(d_out82),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance840830(.data_in(d_in83),.data_out(wire_d83_0),.clk(clk),.rst(rst));            //channel 84
	register #(.WIDTH(WIDTH)) register_instance840831(.data_in(wire_d83_0),.data_out(wire_d83_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance840832(.data_in(wire_d83_1),.data_out(wire_d83_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance840833(.data_in(wire_d83_2),.data_out(wire_d83_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance840834(.data_in(wire_d83_3),.data_out(wire_d83_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance840835(.data_in(wire_d83_4),.data_out(wire_d83_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance840836(.data_in(wire_d83_5),.data_out(wire_d83_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance840837(.data_in(wire_d83_6),.data_out(wire_d83_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance840838(.data_in(wire_d83_7),.data_out(wire_d83_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance840839(.data_in(wire_d83_8),.data_out(wire_d83_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8408310(.data_in(wire_d83_9),.data_out(wire_d83_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8408311(.data_in(wire_d83_10),.data_out(wire_d83_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8408312(.data_in(wire_d83_11),.data_out(wire_d83_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8408313(.data_in(wire_d83_12),.data_out(wire_d83_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8408314(.data_in(wire_d83_13),.data_out(wire_d83_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8408315(.data_in(wire_d83_14),.data_out(wire_d83_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8408316(.data_in(wire_d83_15),.data_out(wire_d83_16),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8408317(.data_in(wire_d83_16),.data_out(wire_d83_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8408318(.data_in(wire_d83_17),.data_out(wire_d83_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8408319(.data_in(wire_d83_18),.data_out(wire_d83_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8408320(.data_in(wire_d83_19),.data_out(wire_d83_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8408321(.data_in(wire_d83_20),.data_out(wire_d83_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8408322(.data_in(wire_d83_21),.data_out(wire_d83_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8408323(.data_in(wire_d83_22),.data_out(wire_d83_23),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8408324(.data_in(wire_d83_23),.data_out(wire_d83_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8408325(.data_in(wire_d83_24),.data_out(wire_d83_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8408326(.data_in(wire_d83_25),.data_out(wire_d83_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8408327(.data_in(wire_d83_26),.data_out(wire_d83_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8408328(.data_in(wire_d83_27),.data_out(wire_d83_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8408329(.data_in(wire_d83_28),.data_out(wire_d83_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8408330(.data_in(wire_d83_29),.data_out(wire_d83_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8408331(.data_in(wire_d83_30),.data_out(wire_d83_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8408332(.data_in(wire_d83_31),.data_out(wire_d83_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8408333(.data_in(wire_d83_32),.data_out(wire_d83_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8408334(.data_in(wire_d83_33),.data_out(wire_d83_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8408335(.data_in(wire_d83_34),.data_out(wire_d83_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8408336(.data_in(wire_d83_35),.data_out(wire_d83_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8408337(.data_in(wire_d83_36),.data_out(wire_d83_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8408338(.data_in(wire_d83_37),.data_out(wire_d83_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8408339(.data_in(wire_d83_38),.data_out(wire_d83_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8408340(.data_in(wire_d83_39),.data_out(wire_d83_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8408341(.data_in(wire_d83_40),.data_out(wire_d83_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8408342(.data_in(wire_d83_41),.data_out(wire_d83_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8408343(.data_in(wire_d83_42),.data_out(wire_d83_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8408344(.data_in(wire_d83_43),.data_out(wire_d83_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8408345(.data_in(wire_d83_44),.data_out(wire_d83_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8408346(.data_in(wire_d83_45),.data_out(wire_d83_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8408347(.data_in(wire_d83_46),.data_out(wire_d83_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8408348(.data_in(wire_d83_47),.data_out(wire_d83_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8408349(.data_in(wire_d83_48),.data_out(wire_d83_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8408350(.data_in(wire_d83_49),.data_out(wire_d83_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8408351(.data_in(wire_d83_50),.data_out(wire_d83_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8408352(.data_in(wire_d83_51),.data_out(wire_d83_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8408353(.data_in(wire_d83_52),.data_out(wire_d83_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8408354(.data_in(wire_d83_53),.data_out(wire_d83_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8408355(.data_in(wire_d83_54),.data_out(wire_d83_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8408356(.data_in(wire_d83_55),.data_out(wire_d83_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8408357(.data_in(wire_d83_56),.data_out(wire_d83_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8408358(.data_in(wire_d83_57),.data_out(wire_d83_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8408359(.data_in(wire_d83_58),.data_out(wire_d83_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8408360(.data_in(wire_d83_59),.data_out(wire_d83_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8408361(.data_in(wire_d83_60),.data_out(wire_d83_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8408362(.data_in(wire_d83_61),.data_out(wire_d83_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8408363(.data_in(wire_d83_62),.data_out(wire_d83_63),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8408364(.data_in(wire_d83_63),.data_out(wire_d83_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8408365(.data_in(wire_d83_64),.data_out(wire_d83_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8408366(.data_in(wire_d83_65),.data_out(wire_d83_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8408367(.data_in(wire_d83_66),.data_out(wire_d83_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8408368(.data_in(wire_d83_67),.data_out(wire_d83_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8408369(.data_in(wire_d83_68),.data_out(wire_d83_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8408370(.data_in(wire_d83_69),.data_out(wire_d83_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8408371(.data_in(wire_d83_70),.data_out(wire_d83_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8408372(.data_in(wire_d83_71),.data_out(wire_d83_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8408373(.data_in(wire_d83_72),.data_out(wire_d83_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8408374(.data_in(wire_d83_73),.data_out(wire_d83_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8408375(.data_in(wire_d83_74),.data_out(wire_d83_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8408376(.data_in(wire_d83_75),.data_out(wire_d83_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8408377(.data_in(wire_d83_76),.data_out(wire_d83_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8408378(.data_in(wire_d83_77),.data_out(wire_d83_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8408379(.data_in(wire_d83_78),.data_out(d_out83),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance850840(.data_in(d_in84),.data_out(wire_d84_0),.clk(clk),.rst(rst));            //channel 85
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance850841(.data_in(wire_d84_0),.data_out(wire_d84_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance850842(.data_in(wire_d84_1),.data_out(wire_d84_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance850843(.data_in(wire_d84_2),.data_out(wire_d84_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance850844(.data_in(wire_d84_3),.data_out(wire_d84_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance850845(.data_in(wire_d84_4),.data_out(wire_d84_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance850846(.data_in(wire_d84_5),.data_out(wire_d84_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance850847(.data_in(wire_d84_6),.data_out(wire_d84_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance850848(.data_in(wire_d84_7),.data_out(wire_d84_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance850849(.data_in(wire_d84_8),.data_out(wire_d84_9),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8508410(.data_in(wire_d84_9),.data_out(wire_d84_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8508411(.data_in(wire_d84_10),.data_out(wire_d84_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8508412(.data_in(wire_d84_11),.data_out(wire_d84_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8508413(.data_in(wire_d84_12),.data_out(wire_d84_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8508414(.data_in(wire_d84_13),.data_out(wire_d84_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8508415(.data_in(wire_d84_14),.data_out(wire_d84_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8508416(.data_in(wire_d84_15),.data_out(wire_d84_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8508417(.data_in(wire_d84_16),.data_out(wire_d84_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8508418(.data_in(wire_d84_17),.data_out(wire_d84_18),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8508419(.data_in(wire_d84_18),.data_out(wire_d84_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8508420(.data_in(wire_d84_19),.data_out(wire_d84_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8508421(.data_in(wire_d84_20),.data_out(wire_d84_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8508422(.data_in(wire_d84_21),.data_out(wire_d84_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8508423(.data_in(wire_d84_22),.data_out(wire_d84_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8508424(.data_in(wire_d84_23),.data_out(wire_d84_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8508425(.data_in(wire_d84_24),.data_out(wire_d84_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8508426(.data_in(wire_d84_25),.data_out(wire_d84_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8508427(.data_in(wire_d84_26),.data_out(wire_d84_27),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8508428(.data_in(wire_d84_27),.data_out(wire_d84_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8508429(.data_in(wire_d84_28),.data_out(wire_d84_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8508430(.data_in(wire_d84_29),.data_out(wire_d84_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8508431(.data_in(wire_d84_30),.data_out(wire_d84_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8508432(.data_in(wire_d84_31),.data_out(wire_d84_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8508433(.data_in(wire_d84_32),.data_out(wire_d84_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8508434(.data_in(wire_d84_33),.data_out(wire_d84_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8508435(.data_in(wire_d84_34),.data_out(wire_d84_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8508436(.data_in(wire_d84_35),.data_out(wire_d84_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8508437(.data_in(wire_d84_36),.data_out(wire_d84_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8508438(.data_in(wire_d84_37),.data_out(wire_d84_38),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8508439(.data_in(wire_d84_38),.data_out(wire_d84_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8508440(.data_in(wire_d84_39),.data_out(wire_d84_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8508441(.data_in(wire_d84_40),.data_out(wire_d84_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8508442(.data_in(wire_d84_41),.data_out(wire_d84_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8508443(.data_in(wire_d84_42),.data_out(wire_d84_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8508444(.data_in(wire_d84_43),.data_out(wire_d84_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8508445(.data_in(wire_d84_44),.data_out(wire_d84_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8508446(.data_in(wire_d84_45),.data_out(wire_d84_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8508447(.data_in(wire_d84_46),.data_out(wire_d84_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8508448(.data_in(wire_d84_47),.data_out(wire_d84_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8508449(.data_in(wire_d84_48),.data_out(wire_d84_49),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8508450(.data_in(wire_d84_49),.data_out(wire_d84_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8508451(.data_in(wire_d84_50),.data_out(wire_d84_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8508452(.data_in(wire_d84_51),.data_out(wire_d84_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8508453(.data_in(wire_d84_52),.data_out(wire_d84_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8508454(.data_in(wire_d84_53),.data_out(wire_d84_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8508455(.data_in(wire_d84_54),.data_out(wire_d84_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8508456(.data_in(wire_d84_55),.data_out(wire_d84_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8508457(.data_in(wire_d84_56),.data_out(wire_d84_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8508458(.data_in(wire_d84_57),.data_out(wire_d84_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8508459(.data_in(wire_d84_58),.data_out(wire_d84_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8508460(.data_in(wire_d84_59),.data_out(wire_d84_60),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8508461(.data_in(wire_d84_60),.data_out(wire_d84_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8508462(.data_in(wire_d84_61),.data_out(wire_d84_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8508463(.data_in(wire_d84_62),.data_out(wire_d84_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8508464(.data_in(wire_d84_63),.data_out(wire_d84_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8508465(.data_in(wire_d84_64),.data_out(wire_d84_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8508466(.data_in(wire_d84_65),.data_out(wire_d84_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8508467(.data_in(wire_d84_66),.data_out(wire_d84_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8508468(.data_in(wire_d84_67),.data_out(wire_d84_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8508469(.data_in(wire_d84_68),.data_out(wire_d84_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8508470(.data_in(wire_d84_69),.data_out(wire_d84_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8508471(.data_in(wire_d84_70),.data_out(wire_d84_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8508472(.data_in(wire_d84_71),.data_out(wire_d84_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8508473(.data_in(wire_d84_72),.data_out(wire_d84_73),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8508474(.data_in(wire_d84_73),.data_out(wire_d84_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8508475(.data_in(wire_d84_74),.data_out(wire_d84_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8508476(.data_in(wire_d84_75),.data_out(wire_d84_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8508477(.data_in(wire_d84_76),.data_out(wire_d84_77),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8508478(.data_in(wire_d84_77),.data_out(wire_d84_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8508479(.data_in(wire_d84_78),.data_out(d_out84),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance860850(.data_in(d_in85),.data_out(wire_d85_0),.clk(clk),.rst(rst));            //channel 86
	register #(.WIDTH(WIDTH)) register_instance860851(.data_in(wire_d85_0),.data_out(wire_d85_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance860852(.data_in(wire_d85_1),.data_out(wire_d85_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance860853(.data_in(wire_d85_2),.data_out(wire_d85_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance860854(.data_in(wire_d85_3),.data_out(wire_d85_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance860855(.data_in(wire_d85_4),.data_out(wire_d85_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance860856(.data_in(wire_d85_5),.data_out(wire_d85_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance860857(.data_in(wire_d85_6),.data_out(wire_d85_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance860858(.data_in(wire_d85_7),.data_out(wire_d85_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance860859(.data_in(wire_d85_8),.data_out(wire_d85_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8608510(.data_in(wire_d85_9),.data_out(wire_d85_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8608511(.data_in(wire_d85_10),.data_out(wire_d85_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8608512(.data_in(wire_d85_11),.data_out(wire_d85_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8608513(.data_in(wire_d85_12),.data_out(wire_d85_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8608514(.data_in(wire_d85_13),.data_out(wire_d85_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8608515(.data_in(wire_d85_14),.data_out(wire_d85_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8608516(.data_in(wire_d85_15),.data_out(wire_d85_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8608517(.data_in(wire_d85_16),.data_out(wire_d85_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8608518(.data_in(wire_d85_17),.data_out(wire_d85_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8608519(.data_in(wire_d85_18),.data_out(wire_d85_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8608520(.data_in(wire_d85_19),.data_out(wire_d85_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8608521(.data_in(wire_d85_20),.data_out(wire_d85_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8608522(.data_in(wire_d85_21),.data_out(wire_d85_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8608523(.data_in(wire_d85_22),.data_out(wire_d85_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8608524(.data_in(wire_d85_23),.data_out(wire_d85_24),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8608525(.data_in(wire_d85_24),.data_out(wire_d85_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8608526(.data_in(wire_d85_25),.data_out(wire_d85_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8608527(.data_in(wire_d85_26),.data_out(wire_d85_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8608528(.data_in(wire_d85_27),.data_out(wire_d85_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8608529(.data_in(wire_d85_28),.data_out(wire_d85_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8608530(.data_in(wire_d85_29),.data_out(wire_d85_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8608531(.data_in(wire_d85_30),.data_out(wire_d85_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8608532(.data_in(wire_d85_31),.data_out(wire_d85_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8608533(.data_in(wire_d85_32),.data_out(wire_d85_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8608534(.data_in(wire_d85_33),.data_out(wire_d85_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8608535(.data_in(wire_d85_34),.data_out(wire_d85_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8608536(.data_in(wire_d85_35),.data_out(wire_d85_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8608537(.data_in(wire_d85_36),.data_out(wire_d85_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8608538(.data_in(wire_d85_37),.data_out(wire_d85_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8608539(.data_in(wire_d85_38),.data_out(wire_d85_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8608540(.data_in(wire_d85_39),.data_out(wire_d85_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8608541(.data_in(wire_d85_40),.data_out(wire_d85_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8608542(.data_in(wire_d85_41),.data_out(wire_d85_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8608543(.data_in(wire_d85_42),.data_out(wire_d85_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8608544(.data_in(wire_d85_43),.data_out(wire_d85_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8608545(.data_in(wire_d85_44),.data_out(wire_d85_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8608546(.data_in(wire_d85_45),.data_out(wire_d85_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8608547(.data_in(wire_d85_46),.data_out(wire_d85_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8608548(.data_in(wire_d85_47),.data_out(wire_d85_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8608549(.data_in(wire_d85_48),.data_out(wire_d85_49),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8608550(.data_in(wire_d85_49),.data_out(wire_d85_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8608551(.data_in(wire_d85_50),.data_out(wire_d85_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8608552(.data_in(wire_d85_51),.data_out(wire_d85_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8608553(.data_in(wire_d85_52),.data_out(wire_d85_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8608554(.data_in(wire_d85_53),.data_out(wire_d85_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8608555(.data_in(wire_d85_54),.data_out(wire_d85_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8608556(.data_in(wire_d85_55),.data_out(wire_d85_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8608557(.data_in(wire_d85_56),.data_out(wire_d85_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8608558(.data_in(wire_d85_57),.data_out(wire_d85_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8608559(.data_in(wire_d85_58),.data_out(wire_d85_59),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8608560(.data_in(wire_d85_59),.data_out(wire_d85_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8608561(.data_in(wire_d85_60),.data_out(wire_d85_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8608562(.data_in(wire_d85_61),.data_out(wire_d85_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8608563(.data_in(wire_d85_62),.data_out(wire_d85_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8608564(.data_in(wire_d85_63),.data_out(wire_d85_64),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8608565(.data_in(wire_d85_64),.data_out(wire_d85_65),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8608566(.data_in(wire_d85_65),.data_out(wire_d85_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8608567(.data_in(wire_d85_66),.data_out(wire_d85_67),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8608568(.data_in(wire_d85_67),.data_out(wire_d85_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8608569(.data_in(wire_d85_68),.data_out(wire_d85_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8608570(.data_in(wire_d85_69),.data_out(wire_d85_70),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8608571(.data_in(wire_d85_70),.data_out(wire_d85_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8608572(.data_in(wire_d85_71),.data_out(wire_d85_72),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8608573(.data_in(wire_d85_72),.data_out(wire_d85_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8608574(.data_in(wire_d85_73),.data_out(wire_d85_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8608575(.data_in(wire_d85_74),.data_out(wire_d85_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8608576(.data_in(wire_d85_75),.data_out(wire_d85_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8608577(.data_in(wire_d85_76),.data_out(wire_d85_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8608578(.data_in(wire_d85_77),.data_out(wire_d85_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8608579(.data_in(wire_d85_78),.data_out(d_out85),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance870860(.data_in(d_in86),.data_out(wire_d86_0),.clk(clk),.rst(rst));            //channel 87
	large_mux #(.WIDTH(WIDTH)) large_mux_instance870861(.data_in(wire_d86_0),.data_out(wire_d86_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance870862(.data_in(wire_d86_1),.data_out(wire_d86_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance870863(.data_in(wire_d86_2),.data_out(wire_d86_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance870864(.data_in(wire_d86_3),.data_out(wire_d86_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance870865(.data_in(wire_d86_4),.data_out(wire_d86_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance870866(.data_in(wire_d86_5),.data_out(wire_d86_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance870867(.data_in(wire_d86_6),.data_out(wire_d86_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance870868(.data_in(wire_d86_7),.data_out(wire_d86_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance870869(.data_in(wire_d86_8),.data_out(wire_d86_9),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8708610(.data_in(wire_d86_9),.data_out(wire_d86_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8708611(.data_in(wire_d86_10),.data_out(wire_d86_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8708612(.data_in(wire_d86_11),.data_out(wire_d86_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8708613(.data_in(wire_d86_12),.data_out(wire_d86_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8708614(.data_in(wire_d86_13),.data_out(wire_d86_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8708615(.data_in(wire_d86_14),.data_out(wire_d86_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8708616(.data_in(wire_d86_15),.data_out(wire_d86_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8708617(.data_in(wire_d86_16),.data_out(wire_d86_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8708618(.data_in(wire_d86_17),.data_out(wire_d86_18),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8708619(.data_in(wire_d86_18),.data_out(wire_d86_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8708620(.data_in(wire_d86_19),.data_out(wire_d86_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8708621(.data_in(wire_d86_20),.data_out(wire_d86_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8708622(.data_in(wire_d86_21),.data_out(wire_d86_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8708623(.data_in(wire_d86_22),.data_out(wire_d86_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8708624(.data_in(wire_d86_23),.data_out(wire_d86_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8708625(.data_in(wire_d86_24),.data_out(wire_d86_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8708626(.data_in(wire_d86_25),.data_out(wire_d86_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8708627(.data_in(wire_d86_26),.data_out(wire_d86_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8708628(.data_in(wire_d86_27),.data_out(wire_d86_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8708629(.data_in(wire_d86_28),.data_out(wire_d86_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8708630(.data_in(wire_d86_29),.data_out(wire_d86_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8708631(.data_in(wire_d86_30),.data_out(wire_d86_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8708632(.data_in(wire_d86_31),.data_out(wire_d86_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8708633(.data_in(wire_d86_32),.data_out(wire_d86_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8708634(.data_in(wire_d86_33),.data_out(wire_d86_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8708635(.data_in(wire_d86_34),.data_out(wire_d86_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8708636(.data_in(wire_d86_35),.data_out(wire_d86_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8708637(.data_in(wire_d86_36),.data_out(wire_d86_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8708638(.data_in(wire_d86_37),.data_out(wire_d86_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8708639(.data_in(wire_d86_38),.data_out(wire_d86_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8708640(.data_in(wire_d86_39),.data_out(wire_d86_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8708641(.data_in(wire_d86_40),.data_out(wire_d86_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8708642(.data_in(wire_d86_41),.data_out(wire_d86_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8708643(.data_in(wire_d86_42),.data_out(wire_d86_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8708644(.data_in(wire_d86_43),.data_out(wire_d86_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8708645(.data_in(wire_d86_44),.data_out(wire_d86_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8708646(.data_in(wire_d86_45),.data_out(wire_d86_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8708647(.data_in(wire_d86_46),.data_out(wire_d86_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8708648(.data_in(wire_d86_47),.data_out(wire_d86_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8708649(.data_in(wire_d86_48),.data_out(wire_d86_49),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8708650(.data_in(wire_d86_49),.data_out(wire_d86_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8708651(.data_in(wire_d86_50),.data_out(wire_d86_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8708652(.data_in(wire_d86_51),.data_out(wire_d86_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8708653(.data_in(wire_d86_52),.data_out(wire_d86_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8708654(.data_in(wire_d86_53),.data_out(wire_d86_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8708655(.data_in(wire_d86_54),.data_out(wire_d86_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8708656(.data_in(wire_d86_55),.data_out(wire_d86_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8708657(.data_in(wire_d86_56),.data_out(wire_d86_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8708658(.data_in(wire_d86_57),.data_out(wire_d86_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8708659(.data_in(wire_d86_58),.data_out(wire_d86_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8708660(.data_in(wire_d86_59),.data_out(wire_d86_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8708661(.data_in(wire_d86_60),.data_out(wire_d86_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8708662(.data_in(wire_d86_61),.data_out(wire_d86_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8708663(.data_in(wire_d86_62),.data_out(wire_d86_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8708664(.data_in(wire_d86_63),.data_out(wire_d86_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8708665(.data_in(wire_d86_64),.data_out(wire_d86_65),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8708666(.data_in(wire_d86_65),.data_out(wire_d86_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8708667(.data_in(wire_d86_66),.data_out(wire_d86_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8708668(.data_in(wire_d86_67),.data_out(wire_d86_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8708669(.data_in(wire_d86_68),.data_out(wire_d86_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8708670(.data_in(wire_d86_69),.data_out(wire_d86_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8708671(.data_in(wire_d86_70),.data_out(wire_d86_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8708672(.data_in(wire_d86_71),.data_out(wire_d86_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8708673(.data_in(wire_d86_72),.data_out(wire_d86_73),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8708674(.data_in(wire_d86_73),.data_out(wire_d86_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8708675(.data_in(wire_d86_74),.data_out(wire_d86_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8708676(.data_in(wire_d86_75),.data_out(wire_d86_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8708677(.data_in(wire_d86_76),.data_out(wire_d86_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8708678(.data_in(wire_d86_77),.data_out(wire_d86_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8708679(.data_in(wire_d86_78),.data_out(d_out86),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance880870(.data_in(d_in87),.data_out(wire_d87_0),.clk(clk),.rst(rst));            //channel 88
	large_mux #(.WIDTH(WIDTH)) large_mux_instance880871(.data_in(wire_d87_0),.data_out(wire_d87_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance880872(.data_in(wire_d87_1),.data_out(wire_d87_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance880873(.data_in(wire_d87_2),.data_out(wire_d87_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance880874(.data_in(wire_d87_3),.data_out(wire_d87_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance880875(.data_in(wire_d87_4),.data_out(wire_d87_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance880876(.data_in(wire_d87_5),.data_out(wire_d87_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance880877(.data_in(wire_d87_6),.data_out(wire_d87_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance880878(.data_in(wire_d87_7),.data_out(wire_d87_8),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance880879(.data_in(wire_d87_8),.data_out(wire_d87_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8808710(.data_in(wire_d87_9),.data_out(wire_d87_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8808711(.data_in(wire_d87_10),.data_out(wire_d87_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8808712(.data_in(wire_d87_11),.data_out(wire_d87_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8808713(.data_in(wire_d87_12),.data_out(wire_d87_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8808714(.data_in(wire_d87_13),.data_out(wire_d87_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8808715(.data_in(wire_d87_14),.data_out(wire_d87_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8808716(.data_in(wire_d87_15),.data_out(wire_d87_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8808717(.data_in(wire_d87_16),.data_out(wire_d87_17),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8808718(.data_in(wire_d87_17),.data_out(wire_d87_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8808719(.data_in(wire_d87_18),.data_out(wire_d87_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8808720(.data_in(wire_d87_19),.data_out(wire_d87_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8808721(.data_in(wire_d87_20),.data_out(wire_d87_21),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8808722(.data_in(wire_d87_21),.data_out(wire_d87_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8808723(.data_in(wire_d87_22),.data_out(wire_d87_23),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8808724(.data_in(wire_d87_23),.data_out(wire_d87_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8808725(.data_in(wire_d87_24),.data_out(wire_d87_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8808726(.data_in(wire_d87_25),.data_out(wire_d87_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8808727(.data_in(wire_d87_26),.data_out(wire_d87_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8808728(.data_in(wire_d87_27),.data_out(wire_d87_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8808729(.data_in(wire_d87_28),.data_out(wire_d87_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8808730(.data_in(wire_d87_29),.data_out(wire_d87_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8808731(.data_in(wire_d87_30),.data_out(wire_d87_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8808732(.data_in(wire_d87_31),.data_out(wire_d87_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8808733(.data_in(wire_d87_32),.data_out(wire_d87_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8808734(.data_in(wire_d87_33),.data_out(wire_d87_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8808735(.data_in(wire_d87_34),.data_out(wire_d87_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8808736(.data_in(wire_d87_35),.data_out(wire_d87_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8808737(.data_in(wire_d87_36),.data_out(wire_d87_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8808738(.data_in(wire_d87_37),.data_out(wire_d87_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8808739(.data_in(wire_d87_38),.data_out(wire_d87_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8808740(.data_in(wire_d87_39),.data_out(wire_d87_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8808741(.data_in(wire_d87_40),.data_out(wire_d87_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8808742(.data_in(wire_d87_41),.data_out(wire_d87_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8808743(.data_in(wire_d87_42),.data_out(wire_d87_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8808744(.data_in(wire_d87_43),.data_out(wire_d87_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8808745(.data_in(wire_d87_44),.data_out(wire_d87_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8808746(.data_in(wire_d87_45),.data_out(wire_d87_46),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8808747(.data_in(wire_d87_46),.data_out(wire_d87_47),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8808748(.data_in(wire_d87_47),.data_out(wire_d87_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8808749(.data_in(wire_d87_48),.data_out(wire_d87_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8808750(.data_in(wire_d87_49),.data_out(wire_d87_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8808751(.data_in(wire_d87_50),.data_out(wire_d87_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8808752(.data_in(wire_d87_51),.data_out(wire_d87_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8808753(.data_in(wire_d87_52),.data_out(wire_d87_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8808754(.data_in(wire_d87_53),.data_out(wire_d87_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8808755(.data_in(wire_d87_54),.data_out(wire_d87_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8808756(.data_in(wire_d87_55),.data_out(wire_d87_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8808757(.data_in(wire_d87_56),.data_out(wire_d87_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8808758(.data_in(wire_d87_57),.data_out(wire_d87_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8808759(.data_in(wire_d87_58),.data_out(wire_d87_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8808760(.data_in(wire_d87_59),.data_out(wire_d87_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8808761(.data_in(wire_d87_60),.data_out(wire_d87_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8808762(.data_in(wire_d87_61),.data_out(wire_d87_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8808763(.data_in(wire_d87_62),.data_out(wire_d87_63),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8808764(.data_in(wire_d87_63),.data_out(wire_d87_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8808765(.data_in(wire_d87_64),.data_out(wire_d87_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8808766(.data_in(wire_d87_65),.data_out(wire_d87_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8808767(.data_in(wire_d87_66),.data_out(wire_d87_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8808768(.data_in(wire_d87_67),.data_out(wire_d87_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8808769(.data_in(wire_d87_68),.data_out(wire_d87_69),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8808770(.data_in(wire_d87_69),.data_out(wire_d87_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8808771(.data_in(wire_d87_70),.data_out(wire_d87_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8808772(.data_in(wire_d87_71),.data_out(wire_d87_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8808773(.data_in(wire_d87_72),.data_out(wire_d87_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8808774(.data_in(wire_d87_73),.data_out(wire_d87_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8808775(.data_in(wire_d87_74),.data_out(wire_d87_75),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8808776(.data_in(wire_d87_75),.data_out(wire_d87_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8808777(.data_in(wire_d87_76),.data_out(wire_d87_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8808778(.data_in(wire_d87_77),.data_out(wire_d87_78),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8808779(.data_in(wire_d87_78),.data_out(d_out87),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance890880(.data_in(d_in88),.data_out(wire_d88_0),.clk(clk),.rst(rst));            //channel 89
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance890881(.data_in(wire_d88_0),.data_out(wire_d88_1),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance890882(.data_in(wire_d88_1),.data_out(wire_d88_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance890883(.data_in(wire_d88_2),.data_out(wire_d88_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance890884(.data_in(wire_d88_3),.data_out(wire_d88_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance890885(.data_in(wire_d88_4),.data_out(wire_d88_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance890886(.data_in(wire_d88_5),.data_out(wire_d88_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance890887(.data_in(wire_d88_6),.data_out(wire_d88_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance890888(.data_in(wire_d88_7),.data_out(wire_d88_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance890889(.data_in(wire_d88_8),.data_out(wire_d88_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8908810(.data_in(wire_d88_9),.data_out(wire_d88_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8908811(.data_in(wire_d88_10),.data_out(wire_d88_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8908812(.data_in(wire_d88_11),.data_out(wire_d88_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8908813(.data_in(wire_d88_12),.data_out(wire_d88_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8908814(.data_in(wire_d88_13),.data_out(wire_d88_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8908815(.data_in(wire_d88_14),.data_out(wire_d88_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8908816(.data_in(wire_d88_15),.data_out(wire_d88_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8908817(.data_in(wire_d88_16),.data_out(wire_d88_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8908818(.data_in(wire_d88_17),.data_out(wire_d88_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8908819(.data_in(wire_d88_18),.data_out(wire_d88_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8908820(.data_in(wire_d88_19),.data_out(wire_d88_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8908821(.data_in(wire_d88_20),.data_out(wire_d88_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8908822(.data_in(wire_d88_21),.data_out(wire_d88_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8908823(.data_in(wire_d88_22),.data_out(wire_d88_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8908824(.data_in(wire_d88_23),.data_out(wire_d88_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8908825(.data_in(wire_d88_24),.data_out(wire_d88_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8908826(.data_in(wire_d88_25),.data_out(wire_d88_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8908827(.data_in(wire_d88_26),.data_out(wire_d88_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8908828(.data_in(wire_d88_27),.data_out(wire_d88_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8908829(.data_in(wire_d88_28),.data_out(wire_d88_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8908830(.data_in(wire_d88_29),.data_out(wire_d88_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8908831(.data_in(wire_d88_30),.data_out(wire_d88_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8908832(.data_in(wire_d88_31),.data_out(wire_d88_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8908833(.data_in(wire_d88_32),.data_out(wire_d88_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8908834(.data_in(wire_d88_33),.data_out(wire_d88_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8908835(.data_in(wire_d88_34),.data_out(wire_d88_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8908836(.data_in(wire_d88_35),.data_out(wire_d88_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8908837(.data_in(wire_d88_36),.data_out(wire_d88_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8908838(.data_in(wire_d88_37),.data_out(wire_d88_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8908839(.data_in(wire_d88_38),.data_out(wire_d88_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8908840(.data_in(wire_d88_39),.data_out(wire_d88_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8908841(.data_in(wire_d88_40),.data_out(wire_d88_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8908842(.data_in(wire_d88_41),.data_out(wire_d88_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8908843(.data_in(wire_d88_42),.data_out(wire_d88_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8908844(.data_in(wire_d88_43),.data_out(wire_d88_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8908845(.data_in(wire_d88_44),.data_out(wire_d88_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8908846(.data_in(wire_d88_45),.data_out(wire_d88_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8908847(.data_in(wire_d88_46),.data_out(wire_d88_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8908848(.data_in(wire_d88_47),.data_out(wire_d88_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8908849(.data_in(wire_d88_48),.data_out(wire_d88_49),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8908850(.data_in(wire_d88_49),.data_out(wire_d88_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8908851(.data_in(wire_d88_50),.data_out(wire_d88_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8908852(.data_in(wire_d88_51),.data_out(wire_d88_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8908853(.data_in(wire_d88_52),.data_out(wire_d88_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8908854(.data_in(wire_d88_53),.data_out(wire_d88_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8908855(.data_in(wire_d88_54),.data_out(wire_d88_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8908856(.data_in(wire_d88_55),.data_out(wire_d88_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8908857(.data_in(wire_d88_56),.data_out(wire_d88_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8908858(.data_in(wire_d88_57),.data_out(wire_d88_58),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8908859(.data_in(wire_d88_58),.data_out(wire_d88_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8908860(.data_in(wire_d88_59),.data_out(wire_d88_60),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8908861(.data_in(wire_d88_60),.data_out(wire_d88_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8908862(.data_in(wire_d88_61),.data_out(wire_d88_62),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8908863(.data_in(wire_d88_62),.data_out(wire_d88_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8908864(.data_in(wire_d88_63),.data_out(wire_d88_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8908865(.data_in(wire_d88_64),.data_out(wire_d88_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8908866(.data_in(wire_d88_65),.data_out(wire_d88_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8908867(.data_in(wire_d88_66),.data_out(wire_d88_67),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8908868(.data_in(wire_d88_67),.data_out(wire_d88_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8908869(.data_in(wire_d88_68),.data_out(wire_d88_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8908870(.data_in(wire_d88_69),.data_out(wire_d88_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8908871(.data_in(wire_d88_70),.data_out(wire_d88_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8908872(.data_in(wire_d88_71),.data_out(wire_d88_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8908873(.data_in(wire_d88_72),.data_out(wire_d88_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8908874(.data_in(wire_d88_73),.data_out(wire_d88_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8908875(.data_in(wire_d88_74),.data_out(wire_d88_75),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8908876(.data_in(wire_d88_75),.data_out(wire_d88_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8908877(.data_in(wire_d88_76),.data_out(wire_d88_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8908878(.data_in(wire_d88_77),.data_out(wire_d88_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8908879(.data_in(wire_d88_78),.data_out(d_out88),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance900890(.data_in(d_in89),.data_out(wire_d89_0),.clk(clk),.rst(rst));            //channel 90
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance900891(.data_in(wire_d89_0),.data_out(wire_d89_1),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance900892(.data_in(wire_d89_1),.data_out(wire_d89_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance900893(.data_in(wire_d89_2),.data_out(wire_d89_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance900894(.data_in(wire_d89_3),.data_out(wire_d89_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance900895(.data_in(wire_d89_4),.data_out(wire_d89_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance900896(.data_in(wire_d89_5),.data_out(wire_d89_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance900897(.data_in(wire_d89_6),.data_out(wire_d89_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance900898(.data_in(wire_d89_7),.data_out(wire_d89_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance900899(.data_in(wire_d89_8),.data_out(wire_d89_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9008910(.data_in(wire_d89_9),.data_out(wire_d89_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9008911(.data_in(wire_d89_10),.data_out(wire_d89_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9008912(.data_in(wire_d89_11),.data_out(wire_d89_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9008913(.data_in(wire_d89_12),.data_out(wire_d89_13),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9008914(.data_in(wire_d89_13),.data_out(wire_d89_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9008915(.data_in(wire_d89_14),.data_out(wire_d89_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9008916(.data_in(wire_d89_15),.data_out(wire_d89_16),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9008917(.data_in(wire_d89_16),.data_out(wire_d89_17),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9008918(.data_in(wire_d89_17),.data_out(wire_d89_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9008919(.data_in(wire_d89_18),.data_out(wire_d89_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9008920(.data_in(wire_d89_19),.data_out(wire_d89_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9008921(.data_in(wire_d89_20),.data_out(wire_d89_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9008922(.data_in(wire_d89_21),.data_out(wire_d89_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9008923(.data_in(wire_d89_22),.data_out(wire_d89_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9008924(.data_in(wire_d89_23),.data_out(wire_d89_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9008925(.data_in(wire_d89_24),.data_out(wire_d89_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9008926(.data_in(wire_d89_25),.data_out(wire_d89_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9008927(.data_in(wire_d89_26),.data_out(wire_d89_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9008928(.data_in(wire_d89_27),.data_out(wire_d89_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9008929(.data_in(wire_d89_28),.data_out(wire_d89_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9008930(.data_in(wire_d89_29),.data_out(wire_d89_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9008931(.data_in(wire_d89_30),.data_out(wire_d89_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9008932(.data_in(wire_d89_31),.data_out(wire_d89_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9008933(.data_in(wire_d89_32),.data_out(wire_d89_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9008934(.data_in(wire_d89_33),.data_out(wire_d89_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9008935(.data_in(wire_d89_34),.data_out(wire_d89_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9008936(.data_in(wire_d89_35),.data_out(wire_d89_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9008937(.data_in(wire_d89_36),.data_out(wire_d89_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9008938(.data_in(wire_d89_37),.data_out(wire_d89_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9008939(.data_in(wire_d89_38),.data_out(wire_d89_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9008940(.data_in(wire_d89_39),.data_out(wire_d89_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9008941(.data_in(wire_d89_40),.data_out(wire_d89_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9008942(.data_in(wire_d89_41),.data_out(wire_d89_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9008943(.data_in(wire_d89_42),.data_out(wire_d89_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9008944(.data_in(wire_d89_43),.data_out(wire_d89_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9008945(.data_in(wire_d89_44),.data_out(wire_d89_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9008946(.data_in(wire_d89_45),.data_out(wire_d89_46),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9008947(.data_in(wire_d89_46),.data_out(wire_d89_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9008948(.data_in(wire_d89_47),.data_out(wire_d89_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9008949(.data_in(wire_d89_48),.data_out(wire_d89_49),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9008950(.data_in(wire_d89_49),.data_out(wire_d89_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9008951(.data_in(wire_d89_50),.data_out(wire_d89_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9008952(.data_in(wire_d89_51),.data_out(wire_d89_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9008953(.data_in(wire_d89_52),.data_out(wire_d89_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9008954(.data_in(wire_d89_53),.data_out(wire_d89_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9008955(.data_in(wire_d89_54),.data_out(wire_d89_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9008956(.data_in(wire_d89_55),.data_out(wire_d89_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9008957(.data_in(wire_d89_56),.data_out(wire_d89_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9008958(.data_in(wire_d89_57),.data_out(wire_d89_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9008959(.data_in(wire_d89_58),.data_out(wire_d89_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9008960(.data_in(wire_d89_59),.data_out(wire_d89_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9008961(.data_in(wire_d89_60),.data_out(wire_d89_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9008962(.data_in(wire_d89_61),.data_out(wire_d89_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9008963(.data_in(wire_d89_62),.data_out(wire_d89_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9008964(.data_in(wire_d89_63),.data_out(wire_d89_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9008965(.data_in(wire_d89_64),.data_out(wire_d89_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9008966(.data_in(wire_d89_65),.data_out(wire_d89_66),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9008967(.data_in(wire_d89_66),.data_out(wire_d89_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9008968(.data_in(wire_d89_67),.data_out(wire_d89_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9008969(.data_in(wire_d89_68),.data_out(wire_d89_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9008970(.data_in(wire_d89_69),.data_out(wire_d89_70),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9008971(.data_in(wire_d89_70),.data_out(wire_d89_71),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9008972(.data_in(wire_d89_71),.data_out(wire_d89_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9008973(.data_in(wire_d89_72),.data_out(wire_d89_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9008974(.data_in(wire_d89_73),.data_out(wire_d89_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9008975(.data_in(wire_d89_74),.data_out(wire_d89_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9008976(.data_in(wire_d89_75),.data_out(wire_d89_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9008977(.data_in(wire_d89_76),.data_out(wire_d89_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9008978(.data_in(wire_d89_77),.data_out(wire_d89_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9008979(.data_in(wire_d89_78),.data_out(d_out89),.clk(clk),.rst(rst));

	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance910900(.data_in(d_in90),.data_out(wire_d90_0),.clk(clk),.rst(rst));            //channel 91
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance910901(.data_in(wire_d90_0),.data_out(wire_d90_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance910902(.data_in(wire_d90_1),.data_out(wire_d90_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance910903(.data_in(wire_d90_2),.data_out(wire_d90_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance910904(.data_in(wire_d90_3),.data_out(wire_d90_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance910905(.data_in(wire_d90_4),.data_out(wire_d90_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance910906(.data_in(wire_d90_5),.data_out(wire_d90_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance910907(.data_in(wire_d90_6),.data_out(wire_d90_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance910908(.data_in(wire_d90_7),.data_out(wire_d90_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance910909(.data_in(wire_d90_8),.data_out(wire_d90_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9109010(.data_in(wire_d90_9),.data_out(wire_d90_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9109011(.data_in(wire_d90_10),.data_out(wire_d90_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9109012(.data_in(wire_d90_11),.data_out(wire_d90_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9109013(.data_in(wire_d90_12),.data_out(wire_d90_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9109014(.data_in(wire_d90_13),.data_out(wire_d90_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9109015(.data_in(wire_d90_14),.data_out(wire_d90_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9109016(.data_in(wire_d90_15),.data_out(wire_d90_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9109017(.data_in(wire_d90_16),.data_out(wire_d90_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9109018(.data_in(wire_d90_17),.data_out(wire_d90_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9109019(.data_in(wire_d90_18),.data_out(wire_d90_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9109020(.data_in(wire_d90_19),.data_out(wire_d90_20),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9109021(.data_in(wire_d90_20),.data_out(wire_d90_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9109022(.data_in(wire_d90_21),.data_out(wire_d90_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9109023(.data_in(wire_d90_22),.data_out(wire_d90_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9109024(.data_in(wire_d90_23),.data_out(wire_d90_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9109025(.data_in(wire_d90_24),.data_out(wire_d90_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9109026(.data_in(wire_d90_25),.data_out(wire_d90_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9109027(.data_in(wire_d90_26),.data_out(wire_d90_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9109028(.data_in(wire_d90_27),.data_out(wire_d90_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9109029(.data_in(wire_d90_28),.data_out(wire_d90_29),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9109030(.data_in(wire_d90_29),.data_out(wire_d90_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9109031(.data_in(wire_d90_30),.data_out(wire_d90_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9109032(.data_in(wire_d90_31),.data_out(wire_d90_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9109033(.data_in(wire_d90_32),.data_out(wire_d90_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9109034(.data_in(wire_d90_33),.data_out(wire_d90_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9109035(.data_in(wire_d90_34),.data_out(wire_d90_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9109036(.data_in(wire_d90_35),.data_out(wire_d90_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9109037(.data_in(wire_d90_36),.data_out(wire_d90_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9109038(.data_in(wire_d90_37),.data_out(wire_d90_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9109039(.data_in(wire_d90_38),.data_out(wire_d90_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9109040(.data_in(wire_d90_39),.data_out(wire_d90_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9109041(.data_in(wire_d90_40),.data_out(wire_d90_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9109042(.data_in(wire_d90_41),.data_out(wire_d90_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9109043(.data_in(wire_d90_42),.data_out(wire_d90_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9109044(.data_in(wire_d90_43),.data_out(wire_d90_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9109045(.data_in(wire_d90_44),.data_out(wire_d90_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9109046(.data_in(wire_d90_45),.data_out(wire_d90_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9109047(.data_in(wire_d90_46),.data_out(wire_d90_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9109048(.data_in(wire_d90_47),.data_out(wire_d90_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9109049(.data_in(wire_d90_48),.data_out(wire_d90_49),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9109050(.data_in(wire_d90_49),.data_out(wire_d90_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9109051(.data_in(wire_d90_50),.data_out(wire_d90_51),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9109052(.data_in(wire_d90_51),.data_out(wire_d90_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9109053(.data_in(wire_d90_52),.data_out(wire_d90_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9109054(.data_in(wire_d90_53),.data_out(wire_d90_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9109055(.data_in(wire_d90_54),.data_out(wire_d90_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9109056(.data_in(wire_d90_55),.data_out(wire_d90_56),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9109057(.data_in(wire_d90_56),.data_out(wire_d90_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9109058(.data_in(wire_d90_57),.data_out(wire_d90_58),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9109059(.data_in(wire_d90_58),.data_out(wire_d90_59),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9109060(.data_in(wire_d90_59),.data_out(wire_d90_60),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9109061(.data_in(wire_d90_60),.data_out(wire_d90_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9109062(.data_in(wire_d90_61),.data_out(wire_d90_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9109063(.data_in(wire_d90_62),.data_out(wire_d90_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9109064(.data_in(wire_d90_63),.data_out(wire_d90_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9109065(.data_in(wire_d90_64),.data_out(wire_d90_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9109066(.data_in(wire_d90_65),.data_out(wire_d90_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9109067(.data_in(wire_d90_66),.data_out(wire_d90_67),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9109068(.data_in(wire_d90_67),.data_out(wire_d90_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9109069(.data_in(wire_d90_68),.data_out(wire_d90_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9109070(.data_in(wire_d90_69),.data_out(wire_d90_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9109071(.data_in(wire_d90_70),.data_out(wire_d90_71),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9109072(.data_in(wire_d90_71),.data_out(wire_d90_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9109073(.data_in(wire_d90_72),.data_out(wire_d90_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9109074(.data_in(wire_d90_73),.data_out(wire_d90_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9109075(.data_in(wire_d90_74),.data_out(wire_d90_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9109076(.data_in(wire_d90_75),.data_out(wire_d90_76),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9109077(.data_in(wire_d90_76),.data_out(wire_d90_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9109078(.data_in(wire_d90_77),.data_out(wire_d90_78),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9109079(.data_in(wire_d90_78),.data_out(d_out90),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance920910(.data_in(d_in91),.data_out(wire_d91_0),.clk(clk),.rst(rst));            //channel 92
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance920911(.data_in(wire_d91_0),.data_out(wire_d91_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance920912(.data_in(wire_d91_1),.data_out(wire_d91_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance920913(.data_in(wire_d91_2),.data_out(wire_d91_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance920914(.data_in(wire_d91_3),.data_out(wire_d91_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance920915(.data_in(wire_d91_4),.data_out(wire_d91_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance920916(.data_in(wire_d91_5),.data_out(wire_d91_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance920917(.data_in(wire_d91_6),.data_out(wire_d91_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance920918(.data_in(wire_d91_7),.data_out(wire_d91_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance920919(.data_in(wire_d91_8),.data_out(wire_d91_9),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9209110(.data_in(wire_d91_9),.data_out(wire_d91_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9209111(.data_in(wire_d91_10),.data_out(wire_d91_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9209112(.data_in(wire_d91_11),.data_out(wire_d91_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9209113(.data_in(wire_d91_12),.data_out(wire_d91_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9209114(.data_in(wire_d91_13),.data_out(wire_d91_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9209115(.data_in(wire_d91_14),.data_out(wire_d91_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9209116(.data_in(wire_d91_15),.data_out(wire_d91_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9209117(.data_in(wire_d91_16),.data_out(wire_d91_17),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9209118(.data_in(wire_d91_17),.data_out(wire_d91_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9209119(.data_in(wire_d91_18),.data_out(wire_d91_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9209120(.data_in(wire_d91_19),.data_out(wire_d91_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9209121(.data_in(wire_d91_20),.data_out(wire_d91_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9209122(.data_in(wire_d91_21),.data_out(wire_d91_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9209123(.data_in(wire_d91_22),.data_out(wire_d91_23),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9209124(.data_in(wire_d91_23),.data_out(wire_d91_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9209125(.data_in(wire_d91_24),.data_out(wire_d91_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9209126(.data_in(wire_d91_25),.data_out(wire_d91_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9209127(.data_in(wire_d91_26),.data_out(wire_d91_27),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9209128(.data_in(wire_d91_27),.data_out(wire_d91_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9209129(.data_in(wire_d91_28),.data_out(wire_d91_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9209130(.data_in(wire_d91_29),.data_out(wire_d91_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9209131(.data_in(wire_d91_30),.data_out(wire_d91_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9209132(.data_in(wire_d91_31),.data_out(wire_d91_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9209133(.data_in(wire_d91_32),.data_out(wire_d91_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9209134(.data_in(wire_d91_33),.data_out(wire_d91_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9209135(.data_in(wire_d91_34),.data_out(wire_d91_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9209136(.data_in(wire_d91_35),.data_out(wire_d91_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9209137(.data_in(wire_d91_36),.data_out(wire_d91_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9209138(.data_in(wire_d91_37),.data_out(wire_d91_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9209139(.data_in(wire_d91_38),.data_out(wire_d91_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9209140(.data_in(wire_d91_39),.data_out(wire_d91_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9209141(.data_in(wire_d91_40),.data_out(wire_d91_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9209142(.data_in(wire_d91_41),.data_out(wire_d91_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9209143(.data_in(wire_d91_42),.data_out(wire_d91_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9209144(.data_in(wire_d91_43),.data_out(wire_d91_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9209145(.data_in(wire_d91_44),.data_out(wire_d91_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9209146(.data_in(wire_d91_45),.data_out(wire_d91_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9209147(.data_in(wire_d91_46),.data_out(wire_d91_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9209148(.data_in(wire_d91_47),.data_out(wire_d91_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9209149(.data_in(wire_d91_48),.data_out(wire_d91_49),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9209150(.data_in(wire_d91_49),.data_out(wire_d91_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9209151(.data_in(wire_d91_50),.data_out(wire_d91_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9209152(.data_in(wire_d91_51),.data_out(wire_d91_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9209153(.data_in(wire_d91_52),.data_out(wire_d91_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9209154(.data_in(wire_d91_53),.data_out(wire_d91_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9209155(.data_in(wire_d91_54),.data_out(wire_d91_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9209156(.data_in(wire_d91_55),.data_out(wire_d91_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9209157(.data_in(wire_d91_56),.data_out(wire_d91_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9209158(.data_in(wire_d91_57),.data_out(wire_d91_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9209159(.data_in(wire_d91_58),.data_out(wire_d91_59),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9209160(.data_in(wire_d91_59),.data_out(wire_d91_60),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9209161(.data_in(wire_d91_60),.data_out(wire_d91_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9209162(.data_in(wire_d91_61),.data_out(wire_d91_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9209163(.data_in(wire_d91_62),.data_out(wire_d91_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9209164(.data_in(wire_d91_63),.data_out(wire_d91_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9209165(.data_in(wire_d91_64),.data_out(wire_d91_65),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9209166(.data_in(wire_d91_65),.data_out(wire_d91_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9209167(.data_in(wire_d91_66),.data_out(wire_d91_67),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9209168(.data_in(wire_d91_67),.data_out(wire_d91_68),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9209169(.data_in(wire_d91_68),.data_out(wire_d91_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9209170(.data_in(wire_d91_69),.data_out(wire_d91_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9209171(.data_in(wire_d91_70),.data_out(wire_d91_71),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9209172(.data_in(wire_d91_71),.data_out(wire_d91_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9209173(.data_in(wire_d91_72),.data_out(wire_d91_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9209174(.data_in(wire_d91_73),.data_out(wire_d91_74),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9209175(.data_in(wire_d91_74),.data_out(wire_d91_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9209176(.data_in(wire_d91_75),.data_out(wire_d91_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9209177(.data_in(wire_d91_76),.data_out(wire_d91_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9209178(.data_in(wire_d91_77),.data_out(wire_d91_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9209179(.data_in(wire_d91_78),.data_out(d_out91),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance930920(.data_in(d_in92),.data_out(wire_d92_0),.clk(clk),.rst(rst));            //channel 93
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance930921(.data_in(wire_d92_0),.data_out(wire_d92_1),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance930922(.data_in(wire_d92_1),.data_out(wire_d92_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance930923(.data_in(wire_d92_2),.data_out(wire_d92_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance930924(.data_in(wire_d92_3),.data_out(wire_d92_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance930925(.data_in(wire_d92_4),.data_out(wire_d92_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance930926(.data_in(wire_d92_5),.data_out(wire_d92_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance930927(.data_in(wire_d92_6),.data_out(wire_d92_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance930928(.data_in(wire_d92_7),.data_out(wire_d92_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance930929(.data_in(wire_d92_8),.data_out(wire_d92_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9309210(.data_in(wire_d92_9),.data_out(wire_d92_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9309211(.data_in(wire_d92_10),.data_out(wire_d92_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9309212(.data_in(wire_d92_11),.data_out(wire_d92_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9309213(.data_in(wire_d92_12),.data_out(wire_d92_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9309214(.data_in(wire_d92_13),.data_out(wire_d92_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9309215(.data_in(wire_d92_14),.data_out(wire_d92_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9309216(.data_in(wire_d92_15),.data_out(wire_d92_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9309217(.data_in(wire_d92_16),.data_out(wire_d92_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9309218(.data_in(wire_d92_17),.data_out(wire_d92_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9309219(.data_in(wire_d92_18),.data_out(wire_d92_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9309220(.data_in(wire_d92_19),.data_out(wire_d92_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9309221(.data_in(wire_d92_20),.data_out(wire_d92_21),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9309222(.data_in(wire_d92_21),.data_out(wire_d92_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9309223(.data_in(wire_d92_22),.data_out(wire_d92_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9309224(.data_in(wire_d92_23),.data_out(wire_d92_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9309225(.data_in(wire_d92_24),.data_out(wire_d92_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9309226(.data_in(wire_d92_25),.data_out(wire_d92_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9309227(.data_in(wire_d92_26),.data_out(wire_d92_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9309228(.data_in(wire_d92_27),.data_out(wire_d92_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9309229(.data_in(wire_d92_28),.data_out(wire_d92_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9309230(.data_in(wire_d92_29),.data_out(wire_d92_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9309231(.data_in(wire_d92_30),.data_out(wire_d92_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9309232(.data_in(wire_d92_31),.data_out(wire_d92_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9309233(.data_in(wire_d92_32),.data_out(wire_d92_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9309234(.data_in(wire_d92_33),.data_out(wire_d92_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9309235(.data_in(wire_d92_34),.data_out(wire_d92_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9309236(.data_in(wire_d92_35),.data_out(wire_d92_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9309237(.data_in(wire_d92_36),.data_out(wire_d92_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9309238(.data_in(wire_d92_37),.data_out(wire_d92_38),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9309239(.data_in(wire_d92_38),.data_out(wire_d92_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9309240(.data_in(wire_d92_39),.data_out(wire_d92_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9309241(.data_in(wire_d92_40),.data_out(wire_d92_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9309242(.data_in(wire_d92_41),.data_out(wire_d92_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9309243(.data_in(wire_d92_42),.data_out(wire_d92_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9309244(.data_in(wire_d92_43),.data_out(wire_d92_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9309245(.data_in(wire_d92_44),.data_out(wire_d92_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9309246(.data_in(wire_d92_45),.data_out(wire_d92_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9309247(.data_in(wire_d92_46),.data_out(wire_d92_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9309248(.data_in(wire_d92_47),.data_out(wire_d92_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9309249(.data_in(wire_d92_48),.data_out(wire_d92_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9309250(.data_in(wire_d92_49),.data_out(wire_d92_50),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9309251(.data_in(wire_d92_50),.data_out(wire_d92_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9309252(.data_in(wire_d92_51),.data_out(wire_d92_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9309253(.data_in(wire_d92_52),.data_out(wire_d92_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9309254(.data_in(wire_d92_53),.data_out(wire_d92_54),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9309255(.data_in(wire_d92_54),.data_out(wire_d92_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9309256(.data_in(wire_d92_55),.data_out(wire_d92_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9309257(.data_in(wire_d92_56),.data_out(wire_d92_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9309258(.data_in(wire_d92_57),.data_out(wire_d92_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9309259(.data_in(wire_d92_58),.data_out(wire_d92_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9309260(.data_in(wire_d92_59),.data_out(wire_d92_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9309261(.data_in(wire_d92_60),.data_out(wire_d92_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9309262(.data_in(wire_d92_61),.data_out(wire_d92_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9309263(.data_in(wire_d92_62),.data_out(wire_d92_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9309264(.data_in(wire_d92_63),.data_out(wire_d92_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9309265(.data_in(wire_d92_64),.data_out(wire_d92_65),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9309266(.data_in(wire_d92_65),.data_out(wire_d92_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9309267(.data_in(wire_d92_66),.data_out(wire_d92_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9309268(.data_in(wire_d92_67),.data_out(wire_d92_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9309269(.data_in(wire_d92_68),.data_out(wire_d92_69),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9309270(.data_in(wire_d92_69),.data_out(wire_d92_70),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9309271(.data_in(wire_d92_70),.data_out(wire_d92_71),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9309272(.data_in(wire_d92_71),.data_out(wire_d92_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9309273(.data_in(wire_d92_72),.data_out(wire_d92_73),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9309274(.data_in(wire_d92_73),.data_out(wire_d92_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9309275(.data_in(wire_d92_74),.data_out(wire_d92_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9309276(.data_in(wire_d92_75),.data_out(wire_d92_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9309277(.data_in(wire_d92_76),.data_out(wire_d92_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9309278(.data_in(wire_d92_77),.data_out(wire_d92_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9309279(.data_in(wire_d92_78),.data_out(d_out92),.clk(clk),.rst(rst));

	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance940930(.data_in(d_in93),.data_out(wire_d93_0),.clk(clk),.rst(rst));            //channel 94
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance940931(.data_in(wire_d93_0),.data_out(wire_d93_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance940932(.data_in(wire_d93_1),.data_out(wire_d93_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance940933(.data_in(wire_d93_2),.data_out(wire_d93_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance940934(.data_in(wire_d93_3),.data_out(wire_d93_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance940935(.data_in(wire_d93_4),.data_out(wire_d93_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance940936(.data_in(wire_d93_5),.data_out(wire_d93_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance940937(.data_in(wire_d93_6),.data_out(wire_d93_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance940938(.data_in(wire_d93_7),.data_out(wire_d93_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance940939(.data_in(wire_d93_8),.data_out(wire_d93_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9409310(.data_in(wire_d93_9),.data_out(wire_d93_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9409311(.data_in(wire_d93_10),.data_out(wire_d93_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9409312(.data_in(wire_d93_11),.data_out(wire_d93_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9409313(.data_in(wire_d93_12),.data_out(wire_d93_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9409314(.data_in(wire_d93_13),.data_out(wire_d93_14),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9409315(.data_in(wire_d93_14),.data_out(wire_d93_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9409316(.data_in(wire_d93_15),.data_out(wire_d93_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9409317(.data_in(wire_d93_16),.data_out(wire_d93_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9409318(.data_in(wire_d93_17),.data_out(wire_d93_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9409319(.data_in(wire_d93_18),.data_out(wire_d93_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9409320(.data_in(wire_d93_19),.data_out(wire_d93_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9409321(.data_in(wire_d93_20),.data_out(wire_d93_21),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9409322(.data_in(wire_d93_21),.data_out(wire_d93_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9409323(.data_in(wire_d93_22),.data_out(wire_d93_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9409324(.data_in(wire_d93_23),.data_out(wire_d93_24),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9409325(.data_in(wire_d93_24),.data_out(wire_d93_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9409326(.data_in(wire_d93_25),.data_out(wire_d93_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9409327(.data_in(wire_d93_26),.data_out(wire_d93_27),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9409328(.data_in(wire_d93_27),.data_out(wire_d93_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9409329(.data_in(wire_d93_28),.data_out(wire_d93_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9409330(.data_in(wire_d93_29),.data_out(wire_d93_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9409331(.data_in(wire_d93_30),.data_out(wire_d93_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9409332(.data_in(wire_d93_31),.data_out(wire_d93_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9409333(.data_in(wire_d93_32),.data_out(wire_d93_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9409334(.data_in(wire_d93_33),.data_out(wire_d93_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9409335(.data_in(wire_d93_34),.data_out(wire_d93_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9409336(.data_in(wire_d93_35),.data_out(wire_d93_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9409337(.data_in(wire_d93_36),.data_out(wire_d93_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9409338(.data_in(wire_d93_37),.data_out(wire_d93_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9409339(.data_in(wire_d93_38),.data_out(wire_d93_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9409340(.data_in(wire_d93_39),.data_out(wire_d93_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9409341(.data_in(wire_d93_40),.data_out(wire_d93_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9409342(.data_in(wire_d93_41),.data_out(wire_d93_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9409343(.data_in(wire_d93_42),.data_out(wire_d93_43),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9409344(.data_in(wire_d93_43),.data_out(wire_d93_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9409345(.data_in(wire_d93_44),.data_out(wire_d93_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9409346(.data_in(wire_d93_45),.data_out(wire_d93_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9409347(.data_in(wire_d93_46),.data_out(wire_d93_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9409348(.data_in(wire_d93_47),.data_out(wire_d93_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9409349(.data_in(wire_d93_48),.data_out(wire_d93_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9409350(.data_in(wire_d93_49),.data_out(wire_d93_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9409351(.data_in(wire_d93_50),.data_out(wire_d93_51),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9409352(.data_in(wire_d93_51),.data_out(wire_d93_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9409353(.data_in(wire_d93_52),.data_out(wire_d93_53),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9409354(.data_in(wire_d93_53),.data_out(wire_d93_54),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9409355(.data_in(wire_d93_54),.data_out(wire_d93_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9409356(.data_in(wire_d93_55),.data_out(wire_d93_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9409357(.data_in(wire_d93_56),.data_out(wire_d93_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9409358(.data_in(wire_d93_57),.data_out(wire_d93_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9409359(.data_in(wire_d93_58),.data_out(wire_d93_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9409360(.data_in(wire_d93_59),.data_out(wire_d93_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9409361(.data_in(wire_d93_60),.data_out(wire_d93_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9409362(.data_in(wire_d93_61),.data_out(wire_d93_62),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9409363(.data_in(wire_d93_62),.data_out(wire_d93_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9409364(.data_in(wire_d93_63),.data_out(wire_d93_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9409365(.data_in(wire_d93_64),.data_out(wire_d93_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9409366(.data_in(wire_d93_65),.data_out(wire_d93_66),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9409367(.data_in(wire_d93_66),.data_out(wire_d93_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9409368(.data_in(wire_d93_67),.data_out(wire_d93_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9409369(.data_in(wire_d93_68),.data_out(wire_d93_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9409370(.data_in(wire_d93_69),.data_out(wire_d93_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9409371(.data_in(wire_d93_70),.data_out(wire_d93_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9409372(.data_in(wire_d93_71),.data_out(wire_d93_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9409373(.data_in(wire_d93_72),.data_out(wire_d93_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9409374(.data_in(wire_d93_73),.data_out(wire_d93_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9409375(.data_in(wire_d93_74),.data_out(wire_d93_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9409376(.data_in(wire_d93_75),.data_out(wire_d93_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9409377(.data_in(wire_d93_76),.data_out(wire_d93_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9409378(.data_in(wire_d93_77),.data_out(wire_d93_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9409379(.data_in(wire_d93_78),.data_out(d_out93),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance950940(.data_in(d_in94),.data_out(wire_d94_0),.clk(clk),.rst(rst));            //channel 95
	large_mux #(.WIDTH(WIDTH)) large_mux_instance950941(.data_in(wire_d94_0),.data_out(wire_d94_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance950942(.data_in(wire_d94_1),.data_out(wire_d94_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance950943(.data_in(wire_d94_2),.data_out(wire_d94_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance950944(.data_in(wire_d94_3),.data_out(wire_d94_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance950945(.data_in(wire_d94_4),.data_out(wire_d94_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance950946(.data_in(wire_d94_5),.data_out(wire_d94_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance950947(.data_in(wire_d94_6),.data_out(wire_d94_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance950948(.data_in(wire_d94_7),.data_out(wire_d94_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance950949(.data_in(wire_d94_8),.data_out(wire_d94_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9509410(.data_in(wire_d94_9),.data_out(wire_d94_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9509411(.data_in(wire_d94_10),.data_out(wire_d94_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9509412(.data_in(wire_d94_11),.data_out(wire_d94_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9509413(.data_in(wire_d94_12),.data_out(wire_d94_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9509414(.data_in(wire_d94_13),.data_out(wire_d94_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9509415(.data_in(wire_d94_14),.data_out(wire_d94_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9509416(.data_in(wire_d94_15),.data_out(wire_d94_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9509417(.data_in(wire_d94_16),.data_out(wire_d94_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9509418(.data_in(wire_d94_17),.data_out(wire_d94_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9509419(.data_in(wire_d94_18),.data_out(wire_d94_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9509420(.data_in(wire_d94_19),.data_out(wire_d94_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9509421(.data_in(wire_d94_20),.data_out(wire_d94_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9509422(.data_in(wire_d94_21),.data_out(wire_d94_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9509423(.data_in(wire_d94_22),.data_out(wire_d94_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9509424(.data_in(wire_d94_23),.data_out(wire_d94_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9509425(.data_in(wire_d94_24),.data_out(wire_d94_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9509426(.data_in(wire_d94_25),.data_out(wire_d94_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9509427(.data_in(wire_d94_26),.data_out(wire_d94_27),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9509428(.data_in(wire_d94_27),.data_out(wire_d94_28),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9509429(.data_in(wire_d94_28),.data_out(wire_d94_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9509430(.data_in(wire_d94_29),.data_out(wire_d94_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9509431(.data_in(wire_d94_30),.data_out(wire_d94_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9509432(.data_in(wire_d94_31),.data_out(wire_d94_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9509433(.data_in(wire_d94_32),.data_out(wire_d94_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9509434(.data_in(wire_d94_33),.data_out(wire_d94_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9509435(.data_in(wire_d94_34),.data_out(wire_d94_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9509436(.data_in(wire_d94_35),.data_out(wire_d94_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9509437(.data_in(wire_d94_36),.data_out(wire_d94_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9509438(.data_in(wire_d94_37),.data_out(wire_d94_38),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9509439(.data_in(wire_d94_38),.data_out(wire_d94_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9509440(.data_in(wire_d94_39),.data_out(wire_d94_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9509441(.data_in(wire_d94_40),.data_out(wire_d94_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9509442(.data_in(wire_d94_41),.data_out(wire_d94_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9509443(.data_in(wire_d94_42),.data_out(wire_d94_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9509444(.data_in(wire_d94_43),.data_out(wire_d94_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9509445(.data_in(wire_d94_44),.data_out(wire_d94_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9509446(.data_in(wire_d94_45),.data_out(wire_d94_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9509447(.data_in(wire_d94_46),.data_out(wire_d94_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9509448(.data_in(wire_d94_47),.data_out(wire_d94_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9509449(.data_in(wire_d94_48),.data_out(wire_d94_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9509450(.data_in(wire_d94_49),.data_out(wire_d94_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9509451(.data_in(wire_d94_50),.data_out(wire_d94_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9509452(.data_in(wire_d94_51),.data_out(wire_d94_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9509453(.data_in(wire_d94_52),.data_out(wire_d94_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9509454(.data_in(wire_d94_53),.data_out(wire_d94_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9509455(.data_in(wire_d94_54),.data_out(wire_d94_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9509456(.data_in(wire_d94_55),.data_out(wire_d94_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9509457(.data_in(wire_d94_56),.data_out(wire_d94_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9509458(.data_in(wire_d94_57),.data_out(wire_d94_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9509459(.data_in(wire_d94_58),.data_out(wire_d94_59),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9509460(.data_in(wire_d94_59),.data_out(wire_d94_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9509461(.data_in(wire_d94_60),.data_out(wire_d94_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9509462(.data_in(wire_d94_61),.data_out(wire_d94_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9509463(.data_in(wire_d94_62),.data_out(wire_d94_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9509464(.data_in(wire_d94_63),.data_out(wire_d94_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9509465(.data_in(wire_d94_64),.data_out(wire_d94_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9509466(.data_in(wire_d94_65),.data_out(wire_d94_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9509467(.data_in(wire_d94_66),.data_out(wire_d94_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9509468(.data_in(wire_d94_67),.data_out(wire_d94_68),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9509469(.data_in(wire_d94_68),.data_out(wire_d94_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9509470(.data_in(wire_d94_69),.data_out(wire_d94_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9509471(.data_in(wire_d94_70),.data_out(wire_d94_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9509472(.data_in(wire_d94_71),.data_out(wire_d94_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9509473(.data_in(wire_d94_72),.data_out(wire_d94_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9509474(.data_in(wire_d94_73),.data_out(wire_d94_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9509475(.data_in(wire_d94_74),.data_out(wire_d94_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9509476(.data_in(wire_d94_75),.data_out(wire_d94_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9509477(.data_in(wire_d94_76),.data_out(wire_d94_77),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9509478(.data_in(wire_d94_77),.data_out(wire_d94_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9509479(.data_in(wire_d94_78),.data_out(d_out94),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance960950(.data_in(d_in95),.data_out(wire_d95_0),.clk(clk),.rst(rst));            //channel 96
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance960951(.data_in(wire_d95_0),.data_out(wire_d95_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance960952(.data_in(wire_d95_1),.data_out(wire_d95_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance960953(.data_in(wire_d95_2),.data_out(wire_d95_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance960954(.data_in(wire_d95_3),.data_out(wire_d95_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance960955(.data_in(wire_d95_4),.data_out(wire_d95_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance960956(.data_in(wire_d95_5),.data_out(wire_d95_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance960957(.data_in(wire_d95_6),.data_out(wire_d95_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance960958(.data_in(wire_d95_7),.data_out(wire_d95_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance960959(.data_in(wire_d95_8),.data_out(wire_d95_9),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9609510(.data_in(wire_d95_9),.data_out(wire_d95_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9609511(.data_in(wire_d95_10),.data_out(wire_d95_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9609512(.data_in(wire_d95_11),.data_out(wire_d95_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9609513(.data_in(wire_d95_12),.data_out(wire_d95_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9609514(.data_in(wire_d95_13),.data_out(wire_d95_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9609515(.data_in(wire_d95_14),.data_out(wire_d95_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9609516(.data_in(wire_d95_15),.data_out(wire_d95_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9609517(.data_in(wire_d95_16),.data_out(wire_d95_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9609518(.data_in(wire_d95_17),.data_out(wire_d95_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9609519(.data_in(wire_d95_18),.data_out(wire_d95_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9609520(.data_in(wire_d95_19),.data_out(wire_d95_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9609521(.data_in(wire_d95_20),.data_out(wire_d95_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9609522(.data_in(wire_d95_21),.data_out(wire_d95_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9609523(.data_in(wire_d95_22),.data_out(wire_d95_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9609524(.data_in(wire_d95_23),.data_out(wire_d95_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9609525(.data_in(wire_d95_24),.data_out(wire_d95_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9609526(.data_in(wire_d95_25),.data_out(wire_d95_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9609527(.data_in(wire_d95_26),.data_out(wire_d95_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9609528(.data_in(wire_d95_27),.data_out(wire_d95_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9609529(.data_in(wire_d95_28),.data_out(wire_d95_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9609530(.data_in(wire_d95_29),.data_out(wire_d95_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9609531(.data_in(wire_d95_30),.data_out(wire_d95_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9609532(.data_in(wire_d95_31),.data_out(wire_d95_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9609533(.data_in(wire_d95_32),.data_out(wire_d95_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9609534(.data_in(wire_d95_33),.data_out(wire_d95_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9609535(.data_in(wire_d95_34),.data_out(wire_d95_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9609536(.data_in(wire_d95_35),.data_out(wire_d95_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9609537(.data_in(wire_d95_36),.data_out(wire_d95_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9609538(.data_in(wire_d95_37),.data_out(wire_d95_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9609539(.data_in(wire_d95_38),.data_out(wire_d95_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9609540(.data_in(wire_d95_39),.data_out(wire_d95_40),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9609541(.data_in(wire_d95_40),.data_out(wire_d95_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9609542(.data_in(wire_d95_41),.data_out(wire_d95_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9609543(.data_in(wire_d95_42),.data_out(wire_d95_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9609544(.data_in(wire_d95_43),.data_out(wire_d95_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9609545(.data_in(wire_d95_44),.data_out(wire_d95_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9609546(.data_in(wire_d95_45),.data_out(wire_d95_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9609547(.data_in(wire_d95_46),.data_out(wire_d95_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9609548(.data_in(wire_d95_47),.data_out(wire_d95_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9609549(.data_in(wire_d95_48),.data_out(wire_d95_49),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9609550(.data_in(wire_d95_49),.data_out(wire_d95_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9609551(.data_in(wire_d95_50),.data_out(wire_d95_51),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9609552(.data_in(wire_d95_51),.data_out(wire_d95_52),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9609553(.data_in(wire_d95_52),.data_out(wire_d95_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9609554(.data_in(wire_d95_53),.data_out(wire_d95_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9609555(.data_in(wire_d95_54),.data_out(wire_d95_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9609556(.data_in(wire_d95_55),.data_out(wire_d95_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9609557(.data_in(wire_d95_56),.data_out(wire_d95_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9609558(.data_in(wire_d95_57),.data_out(wire_d95_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9609559(.data_in(wire_d95_58),.data_out(wire_d95_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9609560(.data_in(wire_d95_59),.data_out(wire_d95_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9609561(.data_in(wire_d95_60),.data_out(wire_d95_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9609562(.data_in(wire_d95_61),.data_out(wire_d95_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9609563(.data_in(wire_d95_62),.data_out(wire_d95_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9609564(.data_in(wire_d95_63),.data_out(wire_d95_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9609565(.data_in(wire_d95_64),.data_out(wire_d95_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9609566(.data_in(wire_d95_65),.data_out(wire_d95_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9609567(.data_in(wire_d95_66),.data_out(wire_d95_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9609568(.data_in(wire_d95_67),.data_out(wire_d95_68),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9609569(.data_in(wire_d95_68),.data_out(wire_d95_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9609570(.data_in(wire_d95_69),.data_out(wire_d95_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9609571(.data_in(wire_d95_70),.data_out(wire_d95_71),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9609572(.data_in(wire_d95_71),.data_out(wire_d95_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9609573(.data_in(wire_d95_72),.data_out(wire_d95_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9609574(.data_in(wire_d95_73),.data_out(wire_d95_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9609575(.data_in(wire_d95_74),.data_out(wire_d95_75),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9609576(.data_in(wire_d95_75),.data_out(wire_d95_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9609577(.data_in(wire_d95_76),.data_out(wire_d95_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9609578(.data_in(wire_d95_77),.data_out(wire_d95_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9609579(.data_in(wire_d95_78),.data_out(d_out95),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance970960(.data_in(d_in96),.data_out(wire_d96_0),.clk(clk),.rst(rst));            //channel 97
	register #(.WIDTH(WIDTH)) register_instance970961(.data_in(wire_d96_0),.data_out(wire_d96_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance970962(.data_in(wire_d96_1),.data_out(wire_d96_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance970963(.data_in(wire_d96_2),.data_out(wire_d96_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance970964(.data_in(wire_d96_3),.data_out(wire_d96_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance970965(.data_in(wire_d96_4),.data_out(wire_d96_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance970966(.data_in(wire_d96_5),.data_out(wire_d96_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance970967(.data_in(wire_d96_6),.data_out(wire_d96_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance970968(.data_in(wire_d96_7),.data_out(wire_d96_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance970969(.data_in(wire_d96_8),.data_out(wire_d96_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9709610(.data_in(wire_d96_9),.data_out(wire_d96_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9709611(.data_in(wire_d96_10),.data_out(wire_d96_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9709612(.data_in(wire_d96_11),.data_out(wire_d96_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9709613(.data_in(wire_d96_12),.data_out(wire_d96_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9709614(.data_in(wire_d96_13),.data_out(wire_d96_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9709615(.data_in(wire_d96_14),.data_out(wire_d96_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9709616(.data_in(wire_d96_15),.data_out(wire_d96_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9709617(.data_in(wire_d96_16),.data_out(wire_d96_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9709618(.data_in(wire_d96_17),.data_out(wire_d96_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9709619(.data_in(wire_d96_18),.data_out(wire_d96_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9709620(.data_in(wire_d96_19),.data_out(wire_d96_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9709621(.data_in(wire_d96_20),.data_out(wire_d96_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9709622(.data_in(wire_d96_21),.data_out(wire_d96_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9709623(.data_in(wire_d96_22),.data_out(wire_d96_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9709624(.data_in(wire_d96_23),.data_out(wire_d96_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9709625(.data_in(wire_d96_24),.data_out(wire_d96_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9709626(.data_in(wire_d96_25),.data_out(wire_d96_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9709627(.data_in(wire_d96_26),.data_out(wire_d96_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9709628(.data_in(wire_d96_27),.data_out(wire_d96_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9709629(.data_in(wire_d96_28),.data_out(wire_d96_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9709630(.data_in(wire_d96_29),.data_out(wire_d96_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9709631(.data_in(wire_d96_30),.data_out(wire_d96_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9709632(.data_in(wire_d96_31),.data_out(wire_d96_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9709633(.data_in(wire_d96_32),.data_out(wire_d96_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9709634(.data_in(wire_d96_33),.data_out(wire_d96_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9709635(.data_in(wire_d96_34),.data_out(wire_d96_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9709636(.data_in(wire_d96_35),.data_out(wire_d96_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9709637(.data_in(wire_d96_36),.data_out(wire_d96_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9709638(.data_in(wire_d96_37),.data_out(wire_d96_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9709639(.data_in(wire_d96_38),.data_out(wire_d96_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9709640(.data_in(wire_d96_39),.data_out(wire_d96_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9709641(.data_in(wire_d96_40),.data_out(wire_d96_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9709642(.data_in(wire_d96_41),.data_out(wire_d96_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9709643(.data_in(wire_d96_42),.data_out(wire_d96_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9709644(.data_in(wire_d96_43),.data_out(wire_d96_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9709645(.data_in(wire_d96_44),.data_out(wire_d96_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9709646(.data_in(wire_d96_45),.data_out(wire_d96_46),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9709647(.data_in(wire_d96_46),.data_out(wire_d96_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9709648(.data_in(wire_d96_47),.data_out(wire_d96_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9709649(.data_in(wire_d96_48),.data_out(wire_d96_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9709650(.data_in(wire_d96_49),.data_out(wire_d96_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9709651(.data_in(wire_d96_50),.data_out(wire_d96_51),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9709652(.data_in(wire_d96_51),.data_out(wire_d96_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9709653(.data_in(wire_d96_52),.data_out(wire_d96_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9709654(.data_in(wire_d96_53),.data_out(wire_d96_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9709655(.data_in(wire_d96_54),.data_out(wire_d96_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9709656(.data_in(wire_d96_55),.data_out(wire_d96_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9709657(.data_in(wire_d96_56),.data_out(wire_d96_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9709658(.data_in(wire_d96_57),.data_out(wire_d96_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9709659(.data_in(wire_d96_58),.data_out(wire_d96_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9709660(.data_in(wire_d96_59),.data_out(wire_d96_60),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9709661(.data_in(wire_d96_60),.data_out(wire_d96_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9709662(.data_in(wire_d96_61),.data_out(wire_d96_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9709663(.data_in(wire_d96_62),.data_out(wire_d96_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9709664(.data_in(wire_d96_63),.data_out(wire_d96_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9709665(.data_in(wire_d96_64),.data_out(wire_d96_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9709666(.data_in(wire_d96_65),.data_out(wire_d96_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9709667(.data_in(wire_d96_66),.data_out(wire_d96_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9709668(.data_in(wire_d96_67),.data_out(wire_d96_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9709669(.data_in(wire_d96_68),.data_out(wire_d96_69),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9709670(.data_in(wire_d96_69),.data_out(wire_d96_70),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9709671(.data_in(wire_d96_70),.data_out(wire_d96_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9709672(.data_in(wire_d96_71),.data_out(wire_d96_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9709673(.data_in(wire_d96_72),.data_out(wire_d96_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9709674(.data_in(wire_d96_73),.data_out(wire_d96_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9709675(.data_in(wire_d96_74),.data_out(wire_d96_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9709676(.data_in(wire_d96_75),.data_out(wire_d96_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9709677(.data_in(wire_d96_76),.data_out(wire_d96_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9709678(.data_in(wire_d96_77),.data_out(wire_d96_78),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9709679(.data_in(wire_d96_78),.data_out(d_out96),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance980970(.data_in(d_in97),.data_out(wire_d97_0),.clk(clk),.rst(rst));            //channel 98
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance980971(.data_in(wire_d97_0),.data_out(wire_d97_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance980972(.data_in(wire_d97_1),.data_out(wire_d97_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance980973(.data_in(wire_d97_2),.data_out(wire_d97_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance980974(.data_in(wire_d97_3),.data_out(wire_d97_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance980975(.data_in(wire_d97_4),.data_out(wire_d97_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance980976(.data_in(wire_d97_5),.data_out(wire_d97_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance980977(.data_in(wire_d97_6),.data_out(wire_d97_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance980978(.data_in(wire_d97_7),.data_out(wire_d97_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance980979(.data_in(wire_d97_8),.data_out(wire_d97_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9809710(.data_in(wire_d97_9),.data_out(wire_d97_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9809711(.data_in(wire_d97_10),.data_out(wire_d97_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9809712(.data_in(wire_d97_11),.data_out(wire_d97_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9809713(.data_in(wire_d97_12),.data_out(wire_d97_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9809714(.data_in(wire_d97_13),.data_out(wire_d97_14),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9809715(.data_in(wire_d97_14),.data_out(wire_d97_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9809716(.data_in(wire_d97_15),.data_out(wire_d97_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9809717(.data_in(wire_d97_16),.data_out(wire_d97_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9809718(.data_in(wire_d97_17),.data_out(wire_d97_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9809719(.data_in(wire_d97_18),.data_out(wire_d97_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9809720(.data_in(wire_d97_19),.data_out(wire_d97_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9809721(.data_in(wire_d97_20),.data_out(wire_d97_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9809722(.data_in(wire_d97_21),.data_out(wire_d97_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9809723(.data_in(wire_d97_22),.data_out(wire_d97_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9809724(.data_in(wire_d97_23),.data_out(wire_d97_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9809725(.data_in(wire_d97_24),.data_out(wire_d97_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9809726(.data_in(wire_d97_25),.data_out(wire_d97_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9809727(.data_in(wire_d97_26),.data_out(wire_d97_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9809728(.data_in(wire_d97_27),.data_out(wire_d97_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9809729(.data_in(wire_d97_28),.data_out(wire_d97_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9809730(.data_in(wire_d97_29),.data_out(wire_d97_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9809731(.data_in(wire_d97_30),.data_out(wire_d97_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9809732(.data_in(wire_d97_31),.data_out(wire_d97_32),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9809733(.data_in(wire_d97_32),.data_out(wire_d97_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9809734(.data_in(wire_d97_33),.data_out(wire_d97_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9809735(.data_in(wire_d97_34),.data_out(wire_d97_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9809736(.data_in(wire_d97_35),.data_out(wire_d97_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9809737(.data_in(wire_d97_36),.data_out(wire_d97_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9809738(.data_in(wire_d97_37),.data_out(wire_d97_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9809739(.data_in(wire_d97_38),.data_out(wire_d97_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9809740(.data_in(wire_d97_39),.data_out(wire_d97_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9809741(.data_in(wire_d97_40),.data_out(wire_d97_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9809742(.data_in(wire_d97_41),.data_out(wire_d97_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9809743(.data_in(wire_d97_42),.data_out(wire_d97_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9809744(.data_in(wire_d97_43),.data_out(wire_d97_44),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9809745(.data_in(wire_d97_44),.data_out(wire_d97_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9809746(.data_in(wire_d97_45),.data_out(wire_d97_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9809747(.data_in(wire_d97_46),.data_out(wire_d97_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9809748(.data_in(wire_d97_47),.data_out(wire_d97_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9809749(.data_in(wire_d97_48),.data_out(wire_d97_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9809750(.data_in(wire_d97_49),.data_out(wire_d97_50),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9809751(.data_in(wire_d97_50),.data_out(wire_d97_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9809752(.data_in(wire_d97_51),.data_out(wire_d97_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9809753(.data_in(wire_d97_52),.data_out(wire_d97_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9809754(.data_in(wire_d97_53),.data_out(wire_d97_54),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9809755(.data_in(wire_d97_54),.data_out(wire_d97_55),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9809756(.data_in(wire_d97_55),.data_out(wire_d97_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9809757(.data_in(wire_d97_56),.data_out(wire_d97_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9809758(.data_in(wire_d97_57),.data_out(wire_d97_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9809759(.data_in(wire_d97_58),.data_out(wire_d97_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9809760(.data_in(wire_d97_59),.data_out(wire_d97_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9809761(.data_in(wire_d97_60),.data_out(wire_d97_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9809762(.data_in(wire_d97_61),.data_out(wire_d97_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9809763(.data_in(wire_d97_62),.data_out(wire_d97_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9809764(.data_in(wire_d97_63),.data_out(wire_d97_64),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9809765(.data_in(wire_d97_64),.data_out(wire_d97_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9809766(.data_in(wire_d97_65),.data_out(wire_d97_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9809767(.data_in(wire_d97_66),.data_out(wire_d97_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9809768(.data_in(wire_d97_67),.data_out(wire_d97_68),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9809769(.data_in(wire_d97_68),.data_out(wire_d97_69),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9809770(.data_in(wire_d97_69),.data_out(wire_d97_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9809771(.data_in(wire_d97_70),.data_out(wire_d97_71),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9809772(.data_in(wire_d97_71),.data_out(wire_d97_72),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9809773(.data_in(wire_d97_72),.data_out(wire_d97_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9809774(.data_in(wire_d97_73),.data_out(wire_d97_74),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9809775(.data_in(wire_d97_74),.data_out(wire_d97_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9809776(.data_in(wire_d97_75),.data_out(wire_d97_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9809777(.data_in(wire_d97_76),.data_out(wire_d97_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9809778(.data_in(wire_d97_77),.data_out(wire_d97_78),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9809779(.data_in(wire_d97_78),.data_out(d_out97),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance990980(.data_in(d_in98),.data_out(wire_d98_0),.clk(clk),.rst(rst));            //channel 99
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance990981(.data_in(wire_d98_0),.data_out(wire_d98_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance990982(.data_in(wire_d98_1),.data_out(wire_d98_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance990983(.data_in(wire_d98_2),.data_out(wire_d98_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance990984(.data_in(wire_d98_3),.data_out(wire_d98_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance990985(.data_in(wire_d98_4),.data_out(wire_d98_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance990986(.data_in(wire_d98_5),.data_out(wire_d98_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance990987(.data_in(wire_d98_6),.data_out(wire_d98_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance990988(.data_in(wire_d98_7),.data_out(wire_d98_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance990989(.data_in(wire_d98_8),.data_out(wire_d98_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9909810(.data_in(wire_d98_9),.data_out(wire_d98_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9909811(.data_in(wire_d98_10),.data_out(wire_d98_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9909812(.data_in(wire_d98_11),.data_out(wire_d98_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9909813(.data_in(wire_d98_12),.data_out(wire_d98_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9909814(.data_in(wire_d98_13),.data_out(wire_d98_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9909815(.data_in(wire_d98_14),.data_out(wire_d98_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9909816(.data_in(wire_d98_15),.data_out(wire_d98_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9909817(.data_in(wire_d98_16),.data_out(wire_d98_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9909818(.data_in(wire_d98_17),.data_out(wire_d98_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9909819(.data_in(wire_d98_18),.data_out(wire_d98_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9909820(.data_in(wire_d98_19),.data_out(wire_d98_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9909821(.data_in(wire_d98_20),.data_out(wire_d98_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9909822(.data_in(wire_d98_21),.data_out(wire_d98_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9909823(.data_in(wire_d98_22),.data_out(wire_d98_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9909824(.data_in(wire_d98_23),.data_out(wire_d98_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9909825(.data_in(wire_d98_24),.data_out(wire_d98_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9909826(.data_in(wire_d98_25),.data_out(wire_d98_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9909827(.data_in(wire_d98_26),.data_out(wire_d98_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9909828(.data_in(wire_d98_27),.data_out(wire_d98_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9909829(.data_in(wire_d98_28),.data_out(wire_d98_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9909830(.data_in(wire_d98_29),.data_out(wire_d98_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9909831(.data_in(wire_d98_30),.data_out(wire_d98_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9909832(.data_in(wire_d98_31),.data_out(wire_d98_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9909833(.data_in(wire_d98_32),.data_out(wire_d98_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9909834(.data_in(wire_d98_33),.data_out(wire_d98_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9909835(.data_in(wire_d98_34),.data_out(wire_d98_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9909836(.data_in(wire_d98_35),.data_out(wire_d98_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9909837(.data_in(wire_d98_36),.data_out(wire_d98_37),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9909838(.data_in(wire_d98_37),.data_out(wire_d98_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9909839(.data_in(wire_d98_38),.data_out(wire_d98_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9909840(.data_in(wire_d98_39),.data_out(wire_d98_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9909841(.data_in(wire_d98_40),.data_out(wire_d98_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9909842(.data_in(wire_d98_41),.data_out(wire_d98_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9909843(.data_in(wire_d98_42),.data_out(wire_d98_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9909844(.data_in(wire_d98_43),.data_out(wire_d98_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9909845(.data_in(wire_d98_44),.data_out(wire_d98_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9909846(.data_in(wire_d98_45),.data_out(wire_d98_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9909847(.data_in(wire_d98_46),.data_out(wire_d98_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9909848(.data_in(wire_d98_47),.data_out(wire_d98_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9909849(.data_in(wire_d98_48),.data_out(wire_d98_49),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9909850(.data_in(wire_d98_49),.data_out(wire_d98_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9909851(.data_in(wire_d98_50),.data_out(wire_d98_51),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9909852(.data_in(wire_d98_51),.data_out(wire_d98_52),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9909853(.data_in(wire_d98_52),.data_out(wire_d98_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9909854(.data_in(wire_d98_53),.data_out(wire_d98_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9909855(.data_in(wire_d98_54),.data_out(wire_d98_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9909856(.data_in(wire_d98_55),.data_out(wire_d98_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9909857(.data_in(wire_d98_56),.data_out(wire_d98_57),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9909858(.data_in(wire_d98_57),.data_out(wire_d98_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9909859(.data_in(wire_d98_58),.data_out(wire_d98_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9909860(.data_in(wire_d98_59),.data_out(wire_d98_60),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9909861(.data_in(wire_d98_60),.data_out(wire_d98_61),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9909862(.data_in(wire_d98_61),.data_out(wire_d98_62),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9909863(.data_in(wire_d98_62),.data_out(wire_d98_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9909864(.data_in(wire_d98_63),.data_out(wire_d98_64),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9909865(.data_in(wire_d98_64),.data_out(wire_d98_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9909866(.data_in(wire_d98_65),.data_out(wire_d98_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9909867(.data_in(wire_d98_66),.data_out(wire_d98_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9909868(.data_in(wire_d98_67),.data_out(wire_d98_68),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9909869(.data_in(wire_d98_68),.data_out(wire_d98_69),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9909870(.data_in(wire_d98_69),.data_out(wire_d98_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9909871(.data_in(wire_d98_70),.data_out(wire_d98_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9909872(.data_in(wire_d98_71),.data_out(wire_d98_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9909873(.data_in(wire_d98_72),.data_out(wire_d98_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9909874(.data_in(wire_d98_73),.data_out(wire_d98_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9909875(.data_in(wire_d98_74),.data_out(wire_d98_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9909876(.data_in(wire_d98_75),.data_out(wire_d98_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9909877(.data_in(wire_d98_76),.data_out(wire_d98_77),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9909878(.data_in(wire_d98_77),.data_out(wire_d98_78),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9909879(.data_in(wire_d98_78),.data_out(d_out98),.clk(clk),.rst(rst));

	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1000990(.data_in(d_in99),.data_out(wire_d99_0),.clk(clk),.rst(rst));            //channel 100
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1000991(.data_in(wire_d99_0),.data_out(wire_d99_1),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1000992(.data_in(wire_d99_1),.data_out(wire_d99_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1000993(.data_in(wire_d99_2),.data_out(wire_d99_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1000994(.data_in(wire_d99_3),.data_out(wire_d99_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1000995(.data_in(wire_d99_4),.data_out(wire_d99_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1000996(.data_in(wire_d99_5),.data_out(wire_d99_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1000997(.data_in(wire_d99_6),.data_out(wire_d99_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1000998(.data_in(wire_d99_7),.data_out(wire_d99_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1000999(.data_in(wire_d99_8),.data_out(wire_d99_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance10009910(.data_in(wire_d99_9),.data_out(wire_d99_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance10009911(.data_in(wire_d99_10),.data_out(wire_d99_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10009912(.data_in(wire_d99_11),.data_out(wire_d99_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10009913(.data_in(wire_d99_12),.data_out(wire_d99_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10009914(.data_in(wire_d99_13),.data_out(wire_d99_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance10009915(.data_in(wire_d99_14),.data_out(wire_d99_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance10009916(.data_in(wire_d99_15),.data_out(wire_d99_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10009917(.data_in(wire_d99_16),.data_out(wire_d99_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance10009918(.data_in(wire_d99_17),.data_out(wire_d99_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance10009919(.data_in(wire_d99_18),.data_out(wire_d99_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10009920(.data_in(wire_d99_19),.data_out(wire_d99_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10009921(.data_in(wire_d99_20),.data_out(wire_d99_21),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance10009922(.data_in(wire_d99_21),.data_out(wire_d99_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance10009923(.data_in(wire_d99_22),.data_out(wire_d99_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance10009924(.data_in(wire_d99_23),.data_out(wire_d99_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance10009925(.data_in(wire_d99_24),.data_out(wire_d99_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10009926(.data_in(wire_d99_25),.data_out(wire_d99_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance10009927(.data_in(wire_d99_26),.data_out(wire_d99_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance10009928(.data_in(wire_d99_27),.data_out(wire_d99_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10009929(.data_in(wire_d99_28),.data_out(wire_d99_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10009930(.data_in(wire_d99_29),.data_out(wire_d99_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance10009931(.data_in(wire_d99_30),.data_out(wire_d99_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10009932(.data_in(wire_d99_31),.data_out(wire_d99_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance10009933(.data_in(wire_d99_32),.data_out(wire_d99_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10009934(.data_in(wire_d99_33),.data_out(wire_d99_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance10009935(.data_in(wire_d99_34),.data_out(wire_d99_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance10009936(.data_in(wire_d99_35),.data_out(wire_d99_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance10009937(.data_in(wire_d99_36),.data_out(wire_d99_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance10009938(.data_in(wire_d99_37),.data_out(wire_d99_38),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance10009939(.data_in(wire_d99_38),.data_out(wire_d99_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10009940(.data_in(wire_d99_39),.data_out(wire_d99_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance10009941(.data_in(wire_d99_40),.data_out(wire_d99_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance10009942(.data_in(wire_d99_41),.data_out(wire_d99_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance10009943(.data_in(wire_d99_42),.data_out(wire_d99_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10009944(.data_in(wire_d99_43),.data_out(wire_d99_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance10009945(.data_in(wire_d99_44),.data_out(wire_d99_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10009946(.data_in(wire_d99_45),.data_out(wire_d99_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10009947(.data_in(wire_d99_46),.data_out(wire_d99_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance10009948(.data_in(wire_d99_47),.data_out(wire_d99_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance10009949(.data_in(wire_d99_48),.data_out(wire_d99_49),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10009950(.data_in(wire_d99_49),.data_out(wire_d99_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance10009951(.data_in(wire_d99_50),.data_out(wire_d99_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10009952(.data_in(wire_d99_51),.data_out(wire_d99_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance10009953(.data_in(wire_d99_52),.data_out(wire_d99_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance10009954(.data_in(wire_d99_53),.data_out(wire_d99_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance10009955(.data_in(wire_d99_54),.data_out(wire_d99_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance10009956(.data_in(wire_d99_55),.data_out(wire_d99_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance10009957(.data_in(wire_d99_56),.data_out(wire_d99_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance10009958(.data_in(wire_d99_57),.data_out(wire_d99_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance10009959(.data_in(wire_d99_58),.data_out(wire_d99_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance10009960(.data_in(wire_d99_59),.data_out(wire_d99_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance10009961(.data_in(wire_d99_60),.data_out(wire_d99_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10009962(.data_in(wire_d99_61),.data_out(wire_d99_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance10009963(.data_in(wire_d99_62),.data_out(wire_d99_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10009964(.data_in(wire_d99_63),.data_out(wire_d99_64),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance10009965(.data_in(wire_d99_64),.data_out(wire_d99_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10009966(.data_in(wire_d99_65),.data_out(wire_d99_66),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10009967(.data_in(wire_d99_66),.data_out(wire_d99_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance10009968(.data_in(wire_d99_67),.data_out(wire_d99_68),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance10009969(.data_in(wire_d99_68),.data_out(wire_d99_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10009970(.data_in(wire_d99_69),.data_out(wire_d99_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance10009971(.data_in(wire_d99_70),.data_out(wire_d99_71),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance10009972(.data_in(wire_d99_71),.data_out(wire_d99_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance10009973(.data_in(wire_d99_72),.data_out(wire_d99_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance10009974(.data_in(wire_d99_73),.data_out(wire_d99_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance10009975(.data_in(wire_d99_74),.data_out(wire_d99_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance10009976(.data_in(wire_d99_75),.data_out(wire_d99_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10009977(.data_in(wire_d99_76),.data_out(wire_d99_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance10009978(.data_in(wire_d99_77),.data_out(wire_d99_78),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance10009979(.data_in(wire_d99_78),.data_out(d_out99),.clk(clk),.rst(rst));


endmodule