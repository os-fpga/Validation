module LATCH_primitive_inst_old(D, G, Q);
  input D;
  input G;
  output Q;

LATCH inst (.*);

endmodule
