-----------------------------------------------------------------
--                                                             --
-----------------------------------------------------------------
--                                                             --
-- Copyright (C) 2013 Stefano Tonello                          --
--                                                             --
-- This source file may be used and distributed without        --
-- restriction provided that this copyright statement is not   --
-- removed from the file and that any derivative work contains --
-- the original copyright notice and the associated disclaimer.--
--                                                             --
-- THIS SOFTWARE IS PROVIDED ``AS IS'' AND WITHOUT ANY         --
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED   --
-- TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS   --
-- FOR A PARTICULAR PURPOSE. IN NO EVENT SHALL THE AUTHOR      --
-- OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT,         --
-- INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES    --
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE   --
-- GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR        --
-- BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF  --
-- LIABILITY, WHETHER IN  CONTRACT, STRICT LIABILITY, OR TORT  --
-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT  --
-- OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE         --
-- POSSIBILITY OF SUCH DAMAGE.                                 --
--                                                             --
-----------------------------------------------------------------

---------------------------------------------------------------
-- G.729a ASIP Instruction ROM content
---------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library WORK;
use work.G729A_ASIP_PKG.all;
use work.G729A_ASIP_CFG_PKG.all;

package G729A_ASIP_ROMI_PKG is

--WIDTH=48;
--DEPTH=4608;

--ADDRESS_RADIX=UNS;
--DATA_RADIX=HEX;

--CONTENT BEGIN

  subtype ROMI_WORD_T is std_logic_vector(ILEN*2-1 downto 0);

  type ROMI_DATA_T is array (0 to IMEM_SIZE/2-1) of ROMI_WORD_T;

  constant ROMI_INIT_DATA : ROMI_DATA_T := (

    X"80f11b3ff007", --    0
    X"80f33b80f22b", --    1
    X"81f07a80f44b", --    2
    X"83f05a82f06a", --    3
    X"c000eac000b9", --    4
    X"84100a00301e", --    5
    X"122001111001", --    6
    X"81f01a8f24fb", --    7
    X"83f03a82f02a", --    8
    X"1ff00784f04a", --    9
    X"3ff00a00e01a", --   10
    X"80f12b80f01b", --   11
    X"80f34b80f23b", --   12
    X"80f56b80f45b", --   13
    X"80000a80f0aa", --   14
    X"80100b81f07a", --   15
    X"c002a980f09a", --   16
    X"81f08ac0031a", --   17
    X"81f0aa00101e", --   18
    X"82f07a111001", --   19
    X"130000122001", --   20
    X"11100184100a", --   21
    X"04400904400b", --   22
    X"12200180240b", --   23
    X"00400904030b", --   24
    X"04400b84100a", --   25
    X"80240b044009", --   26
    X"81f02a80f01a", --   27
    X"83f04a82f03a", --   28
    X"85f06a84f05a", --   29
    X"00e01a1ff00a", --   30
    X"80f01b3ff00e", --   31
    X"80f23b80f12b", --   32
    X"80f45b80f34b", --   33
    X"80f67b80f56b", --   34
    X"80f89b80f78b", --   35
    X"80fabb80f9ab", --   36
    X"d10028d00000", --   37
    X"88f0ca82f0da", --   38
    X"86200a83f0ea", --   39
    X"13300187300a", --   40
    X"04670bc00589", --   41
    X"c0005bc005fa", --   42
    X"000024004023", --   43
    X"862ffa87300a", --   44
    X"8a2fea89301a", --   45
    X"322002133002", --   46
    X"049a13047613", --   47
    X"12200a100001", --   48
    X"044009844031", --   49
    X"122001188001", --   50
    X"8e01798f84fb", --   51
    X"81f02a80f01a", --   52
    X"83f04a82f03a", --   53
    X"85f06a84f05a", --   54
    X"87f08a86f07a", --   55
    X"89f0aa88f09a", --   56
    X"1ff00e8af0ba", --   57
    X"3ff07500e01a", --   58
    X"80f12b80f01b", --   59
    X"80f34b80f23b", --   60
    X"80f56b80f45b", --   61
    X"80f78b80f67b", --   62
    X"80f9ab80f89b", --   63
    X"80f71a80fabb", --   64
    X"c0086911f00c", --   65
    X"c000abc0089a", --   66
    X"10000182000a", --   67
    X"8f12fb111001", --   68
    X"84f72a80f74a", --   69
    X"11f00c040402", --   70
    X"81f75a15100a", --   71
    X"83100a82000a", --   72
    X"c009a9385001", --   73
    X"c00a1a06230b", --   74
    X"c0005b111001", --   75
    X"000024006023", --   76
    X"83100a82800a", --   77
    X"8a101a898ffa", --   78
    X"111002388002", --   79
    X"069a14062314", --   80
    X"066009866031", --   81
    X"80560b100001", --   82
    X"8e0489155001", --   83
    X"10000a10f00c", --   84
    X"c00af981f73a", --   85
    X"84f72ac00b2a", --   86
    X"83000a00401e", --   87
    X"111001100001", --   88
    X"80f70a8f13fb", --   89
    X"8001c8d10000", --   90
    X"00040280f73a", --   91
    X"81f71a30000a", --   92
    X"c00c0ac00bd9", --   93
    X"83000ac000ab", --   94
    X"111001100001", --   95
    X"80f01a8f13fb", --   96
    X"82f03a81f02a", --   97
    X"84f05a83f04a", --   98
    X"86f07a85f06a", --   99
    X"88f09a87f08a", --  100
    X"8af0ba89f0aa", --  101
    X"00e01a1ff075", --  102
    X"3ff00e00001d", --  103
    X"80f12b80f01b", --  104
    X"80f34b80f23b", --  105
    X"80f56b80f45b", --  106
    X"80f78b80f67b", --  107
    X"81f0ea80f89b", --  108
    X"d8000082f0da", --  109
    X"c02144c01154", --  110
    X"c00122001206", --  111
    X"d87fff801239", --  112
    X"641001c00f18", --  113
    X"662001844013", --  114
    X"c00eb9866013", --  115
    X"c000fbc00f0a", --  116
    X"888010844011", --  117
    X"c02035024607", --  118
    X"188001044607", --  119
    X"80f8cb844011", --  120
    X"81f02a80f01a", --  121
    X"83f04a82f03a", --  122
    X"85f06a84f05a", --  123
    X"87f08a86f07a", --  124
    X"1ff00e88f09a", --  125
    X"3ff02e00e01a", --  126
    X"80f12b80f01b", --  127
    X"80f34b80f23b", --  128
    X"80f56b80f45b", --  129
    X"80f78b80f67b", --  130
    X"80f9ab80f89b", --  131
    X"80fecb80fabb", --  132
    X"c0189ac010e9", --  133
    X"d60000c0002b", --  134
    X"80f00b80f2ea", --  135
    X"8ff0fb10f017", --  136
    X"d20004d01485", --  137
    X"02260c72200a", --  138
    X"8ff0eb000202", --  139
    X"8ff0dbd00303", --  140
    X"72600ad014e9", --  141
    X"8ff0cb000202", --  142
    X"10f017be01ce", --  143
    X"d00e4580f00b", --  144
    X"be02058ff0fb", --  145
    X"10f00d88ffea", --  146
    X"80080b000602", --  147
    X"80f00b10f017", --  148
    X"da0e4570800a", --  149
    X"8ff0fb000a02", --  150
    X"8ff0eb80f2da", --  151
    X"8ff0dbd01345", --  152
    X"87ffcabe023c", --  153
    X"00060210f00f", --  154
    X"10f02180070b", --  155
    X"da0e4571800a", --  156
    X"72700a011a02", --  157
    X"022a02da1345", --  158
    X"84100a170005", --  159
    X"03450285200a", --  160
    X"10000180030b", --  161
    X"122001111001", --  162
    X"10f0218f0799", --  163
    X"be028380f00b", --  164
    X"80f00b10f017", --  165
    X"da0e4570800a", --  166
    X"8ff0fb000a02", --  167
    X"8ff0eb80f2da", --  168
    X"8ff0dbd01345", --  169
    X"87ffcabe029f", --  170
    X"00060210f011", --  171
    X"10f02180070b", --  172
    X"71800a100005", --  173
    X"011a02da0e45", --  174
    X"72700a111005", --  175
    X"022a02da1345", --  176
    X"170005122005", --  177
    X"85200a84100a", --  178
    X"80030b034502", --  179
    X"111001100001", --  180
    X"8f0799122001", --  181
    X"80f00b10f021", --  182
    X"10f021be02e9", --  183
    X"d0000580f00b", --  184
    X"be03068ff0fb", --  185
    X"80f00b80f2da", --  186
    X"8ff0fb10f021", --  187
    X"8ff0cb10f017", --  188
    X"72600ad014d5", --  189
    X"8ff0bb000202", --  190
    X"87ffdabe0325", --  191
    X"72600210f013", --  192
    X"80070b000202", --  193
    X"10f01387ffea", --  194
    X"000202726002", --  195
    X"16600180071b", --  196
    X"10f013d60000", --  197
    X"83001a82000a", --  198
    X"85003a84002a", --  199
    X"c02027024207", --  200
    X"806070d60001", --  201
    X"01160211f00d", --  202
    X"00010281100a", --  203
    X"80200b82f2ba", --  204
    X"01160211f00f", --  205
    X"80105081100a", --  206
    X"01160211f011", --  207
    X"00010281100a", --  208
    X"80201b82f2ba", --  209
    X"00060210f00d", --  210
    X"80f00b80000a", --  211
    X"00060210f00f", --  212
    X"8ff0fb80000a", --  213
    X"00060210f011", --  214
    X"8ff0eb80000a", --  215
    X"d10004d01485", --  216
    X"01160c71100a", --  217
    X"8ff0db000102", --  218
    X"8ff0cbd00303", --  219
    X"8ff0bb80f2ca", --  220
    X"d1000ad014d5", --  221
    X"00010201160c", --  222
    X"be03548ff0ab", --  223
    X"81f02a80f01a", --  224
    X"83f04a82f03a", --  225
    X"85f06a84f05a", --  226
    X"87f08a86f07a", --  227
    X"89f0aa88f09a", --  228
    X"8ef0ca8af0ba", --  229
    X"00e01a1ff02e", --  230
    X"80f01b3ff00f", --  231
    X"80f23b80f12b", --  232
    X"80f45b80f34b", --  233
    X"80f67b80f56b", --  234
    X"80f89b80f78b", --  235
    X"d0000080f9ab", --  236
    X"03100281f0fa", --  237
    X"d2000083300a", --  238
    X"84f0ca002023", --  239
    X"d6000085f0da", --  240
    X"07700277600a", --  241
    X"88700a077402", --  242
    X"07700277600a", --  243
    X"89700a077502", --  244
    X"166001028914", --  245
    X"cf7f54376004", --  246
    X"07700287f0ba", --  247
    X"02370b87700a", --  248
    X"87f0ea822031", --  249
    X"80730b077002", --  250
    X"d7000a100001", --  251
    X"80f01a8e0739", --  252
    X"82f03a81f02a", --  253
    X"84f05a83f04a", --  254
    X"86f07a85f06a", --  255
    X"88f09a87f08a", --  256
    X"1ff00f89f0aa", --  257
    X"3ff00e00e01a", --  258
    X"80f12b80f01b", --  259
    X"80f34b80f23b", --  260
    X"80f56b80f45b", --  261
    X"80f78b80f67b", --  262
    X"80f9ab80f89b", --  263
    X"d8000080fabb", --  264
    X"d77fffd6ffff", --  265
    X"d9008082f0da", --  266
    X"d40000da0000", --  267
    X"004023d50000", --  268
    X"c0227ac021e9", --  269
    X"80f0eac0005b", --  270
    X"81200a83000a", --  271
    X"8c201a8b001a", --  272
    X"122002100002", --  273
    X"0bbc06013106", --  274
    X"04bb13041113", --  275
    X"c00037004607", --  276
    X"18a000264000", --  277
    X"8ea9a91aa001", --  278
    X"80f01a80f8cb", --  279
    X"82f03a81f02a", --  280
    X"84f05a83f04a", --  281
    X"86f07a85f06a", --  282
    X"88f09a87f08a", --  283
    X"8af0ba89f0aa", --  284
    X"00e01a1ff00e", --  285
    X"80f01b3ff01b", --  286
    X"80f23b80f12b", --  287
    X"80f45b80f34b", --  288
    X"80f67b80f56b", --  289
    X"80f89b80f78b", --  290
    X"80fabb80f9ab", --  291
    X"10f00d80fbcb", --  292
    X"82f1aa81f1ba", --  293
    X"84100a130005", --  294
    X"06450685200a", --  295
    X"10000180060b", --  296
    X"122001111001", --  297
    X"d6ffff8f0399", --  298
    X"82f18ad77fff", --  299
    X"d0002089f18a", --  300
    X"09900270000a", --  301
    X"c02659da0000", --  302
    X"10f00dc026da", --  303
    X"d4000088f19a", --  304
    X"004023d50000", --  305
    X"83000ac0005b", --  306
    X"8b800a81200a", --  307
    X"013106100001", --  308
    X"12200103b10a", --  309
    X"043113188001", --  310
    X"c00037004607", --  311
    X"81fa7b264000", --  312
    X"1220051aa001", --  313
    X"80f01a8e29b9", --  314
    X"82f03a81f02a", --  315
    X"84f05a83f04a", --  316
    X"86f07a85f06a", --  317
    X"88f09a87f08a", --  318
    X"8af0ba89f0aa", --  319
    X"1ff01b8bf0ca", --  320
    X"3ff00600e01a", --  321
    X"80f12b80f01b", --  322
    X"80f34b80f23b", --  323
    X"80f06a80f45b", --  324
    X"311001110005", --  325
    X"83001a82000a", --  326
    X"14400a042306", --  327
    X"c04050844012", --  328
    X"80020b022406", --  329
    X"80031b033402", --  330
    X"8f0159100001", --  331
    X"81f02a80f01a", --  332
    X"83f04a82f03a", --  333
    X"1ff00684f05a", --  334
    X"3ff01b00e01a", --  335
    X"80f12b80f01b", --  336
    X"80f34b80f23b", --  337
    X"80f56b80f45b", --  338
    X"80f78b80f67b", --  339
    X"80f9ab80f89b", --  340
    X"80fbcb80fabb", --  341
    X"10000510f00d", --  342
    X"11100581f1ba", --  343
    X"12200582f1aa", --  344
    X"84100a130005", --  345
    X"85200a111001", --  346
    X"064506122001", --  347
    X"10000180060b", --  348
    X"d6ffff8f0399", --  349
    X"82f18ad77fff", --  350
    X"d90020122005", --  351
    X"d40000da0000", --  352
    X"004023d50000", --  353
    X"c02d3ac02cb9", --  354
    X"10f00dc0005b", --  355
    X"88f19a100005", --  356
    X"83000a188005", --  357
    X"8b800a81200a", --  358
    X"013106100001", --  359
    X"188001122001", --  360
    X"04311303b10a", --  361
    X"c00037004607", --  362
    X"81fa7b264000", --  363
    X"1220051aa001", --  364
    X"80f01a8ea979", --  365
    X"82f03a81f02a", --  366
    X"84f05a83f04a", --  367
    X"86f07a85f06a", --  368
    X"88f09a87f08a", --  369
    X"8af0ba89f0aa", --  370
    X"1ff01b8bf0ca", --  371
    X"3ff00600e01a", --  372
    X"80f12b80f01b", --  373
    X"80f34b80f23b", --  374
    X"80f06a80f45b", --  375
    X"300001100005", --  376
    X"82000a110005", --  377
    X"04230683001a", --  378
    X"84401214400a", --  379
    X"022406c04050", --  380
    X"03340280020b", --  381
    X"10000180031b", --  382
    X"80f01a8f0159", --  383
    X"82f03a81f02a", --  384
    X"84f05a83f04a", --  385
    X"00e01a1ff006", --  386
    X"80f01b3ff008", --  387
    X"80f23b80f12b", --  388
    X"80f45b80f34b", --  389
    X"80f08a80f56b", --  390
    X"31100111000a", --  391
    X"82000a85f07a", --  392
    X"04230683001a", --  393
    X"844012044502", --  394
    X"022406c04050", --  395
    X"03340280020b", --  396
    X"10000180031b", --  397
    X"80f01a8f0159", --  398
    X"82f03a81f02a", --  399
    X"84f05a83f04a", --  400
    X"1ff00885f06a", --  401
    X"3ff01000e01a", --  402
    X"80f12b80f01b", --  403
    X"80f34b80f23b", --  404
    X"80f56b80f45b", --  405
    X"80f78b80f67b", --  406
    X"80f9ab80f89b", --  407
    X"d90000d80000", --  408
    X"81f0ca80f0fa", --  409
    X"83f10a82f0ba", --  410
    X"85000a14000a", --  411
    X"05560686100a", --  412
    X"05560a86200a", --  413
    X"06650b86300a", --  414
    X"06750b866041", --  415
    X"100001088603", --  416
    X"122001111001", --  417
    X"8f0429133001", --  418
    X"80f9eb80f8db", --  419
    X"81f02a80f01a", --  420
    X"83f04a82f03a", --  421
    X"85f06a84f05a", --  422
    X"87f08a86f07a", --  423
    X"89f0aa88f09a", --  424
    X"00e01a1ff010", --  425
    X"80f01b3ff01d", --  426
    X"80f23b80f12b", --  427
    X"80f45b80f34b", --  428
    X"80f67b80f56b", --  429
    X"80f89b80f78b", --  430
    X"80fabb80f9ab", --  431
    X"10f00d80fecb", --  432
    X"82f1da110005", --  433
    X"da0e4572200a", --  434
    X"83f1ca022a02", --  435
    X"da134573300a", --  436
    X"84200a033a02", --  437
    X"85300a122001", --  438
    X"044502133001", --  439
    X"10000180040b", --  440
    X"10f00d8f0199", --  441
    X"110005100005", --  442
    X"72200a82f1da", --  443
    X"022a02da0e45", --  444
    X"83f1ba122005", --  445
    X"da134573300a", --  446
    X"133005033a02", --  447
    X"12200184200a", --  448
    X"13300185300a", --  449
    X"80040b044502", --  450
    X"8f0199100001", --  451
    X"80f00b10f00d", --  452
    X"8ff0fbd0000a", --  453
    X"10f00dbe0306", --  454
    X"d0000580f00b", --  455
    X"be03068ff0fb", --  456
    X"80f00b10f00d", --  457
    X"8ff0fb80f18a", --  458
    X"8ff0eb80f1aa", --  459
    X"8ff0db80f19a", --  460
    X"8ff0cb80f17a", --  461
    X"10f00dbe03b3", --  462
    X"80f19a80f00b", --  463
    X"be03e98ff0fb", --  464
    X"80f00b80f18a", --  465
    X"80f01abe040c", --  466
    X"82f03a81f02a", --  467
    X"84f05a83f04a", --  468
    X"86f07a85f06a", --  469
    X"88f09a87f08a", --  470
    X"8af0ba89f0aa", --  471
    X"1ff01d8ef0ca", --  472
    X"3ff00f00e01a", --  473
    X"80f12b80f01b", --  474
    X"80f34b80f23b", --  475
    X"80f56b80f45b", --  476
    X"80f78b80f67b", --  477
    X"80f9ab80f89b", --  478
    X"80f0fa89f0ea", --  479
    X"82f0ba81f0ba", --  480
    X"d8000012200a", --  481
    X"10000183000a", --  482
    X"11100186100a", --  483
    X"00402304360b", --  484
    X"03380283f0ca", --  485
    X"06680286f0da", --  486
    X"d4000a87f0da", --  487
    X"077402744004", --  488
    X"84300a077802", --  489
    X"04451385600a", --  490
    X"16600a13300a", --  491
    X"80950b8f67b9", --  492
    X"188001199001", --  493
    X"80f01a8e1289", --  494
    X"82f03a81f02a", --  495
    X"84f05a83f04a", --  496
    X"86f07a85f06a", --  497
    X"88f09a87f08a", --  498
    X"1ff00f89f0aa", --  499
    X"3ff00500e01a", --  500
    X"80f12b80f01b", --  501
    X"80f04a80f23b", --  502
    X"71100ad10004", --  503
    X"000102311001", --  504
    X"31100a82f04a", --  505
    X"111001022102", --  506
    X"c03fcac03f99", --  507
    X"81200a00101e", --  508
    X"80010b322001", --  509
    X"c04039300001", --  510
    X"c000abc0406a", --  511
    X"12200a82f05a", --  512
    X"81200a322001", --  513
    X"80010b322001", --  514
    X"80f01a300001", --  515
    X"82f03a81f02a", --  516
    X"00e01a1ff005", --  517
    X"80f01b3ff007", --  518
    X"80f23b80f12b", --  519
    X"80f45b80f34b", --  520
    X"80f07a80f56b", --  521
    X"111fff11000a", --  522
    X"62200182000a", --  523
    X"84001a822013", --  524
    X"844013644001", --  525
    X"c06057064207", --  526
    X"84001a82000a", --  527
    X"80040b80021b", --  528
    X"8f0139100001", --  529
    X"81000a80f07a", --  530
    X"c01036311028", --  531
    X"80010bd10028", --  532
    X"111fff11000a", --  533
    X"62200182000a", --  534
    X"84001a822013", --  535
    X"844013644001", --  536
    X"466141064207", --  537
    X"82000ac06047", --  538
    X"80021b122141", --  539
    X"8f0139100001", --  540
    X"d2645181000a", --  541
    X"c01030011206", --  542
    X"80010bd16451", --  543
    X"81f02a80f01a", --  544
    X"83f04a82f03a", --  545
    X"85f06a84f05a", --  546
    X"00e01a1ff007", --  547
    X"80f01b3ff014", --  548
    X"80f23b80f12b", --  549
    X"80f45b80f34b", --  550
    X"80fe7b80f56b", --  551
    X"81f13a80f14a", --  552
    X"c0456912f008", --  553
    X"c000abc045ea", --  554
    X"10000183000a", --  555
    X"84100a833012", --  556
    X"844012111001", --  557
    X"80250b054302", --  558
    X"12f008122001", --  559
    X"80f12a80f20b", --  560
    X"be04748ff0fb", --  561
    X"80f00b80f13a", --  562
    X"10000a80f12a", --  563
    X"8ff0fb100001", --  564
    X"80f01abe0474", --  565
    X"82f03a81f02a", --  566
    X"84f05a83f04a", --  567
    X"8ef07a85f06a", --  568
    X"00e01a1ff014", --  569
    X"80f01b3ff025", --  570
    X"80f23b80f12b", --  571
    X"80f45b80f34b", --  572
    X"80f67b80f56b", --  573
    X"80f89b80f78b", --  574
    X"80febb80f9ab", --  575
    X"80f00b80f25a", --  576
    X"8ff0fb10f00c", --  577
    X"80f25abe04d6", --  578
    X"80f00b100001", --  579
    X"8ff0fb10f018", --  580
    X"c04939be04d6", --  581
    X"c0005bc04a2a", --  582
    X"11f00cd00005", --  583
    X"12f01811100a", --  584
    X"84100a12200a", --  585
    X"861fea85101a", --  586
    X"044603871ffa", --  587
    X"80151b80140b", --  588
    X"85201a84200a", --  589
    X"872ffa862fea", --  590
    X"80240b044607", --  591
    X"31100280251b", --  592
    X"d01000322002", --  593
    X"80100b81f24a", --  594
    X"c04c8ac04b19", --  595
    X"80f24ac0005b", --  596
    X"11f00c100001", --  597
    X"12f018111002", --  598
    X"83f24a122002", --  599
    X"84100a13300a", --  600
    X"86200a85101a", --  601
    X"08460387201a", --  602
    X"8ff8fb80f90b", --  603
    X"8ff9ebd9000d", --  604
    X"88ffcabe0528", --  605
    X"08460780080b", --  606
    X"8ff8fb80f90b", --  607
    X"8ff9ebd9000d", --  608
    X"88ffcabe0528", --  609
    X"10000180380b", --  610
    X"122002111002", --  611
    X"80f01a333001", --  612
    X"82f03a81f02a", --  613
    X"84f05a83f04a", --  614
    X"86f07a85f06a", --  615
    X"88f09a87f08a", --  616
    X"8ef0ba89f0aa", --  617
    X"00e01a1ff025", --  618
    X"80f01b3ff00c", --  619
    X"80f23b80f12b", --  620
    X"80f45b80f34b", --  621
    X"80f67b80f56b", --  622
    X"80f89b80f78b", --  623
    X"82f0ba80f9ab", --  624
    X"d10800d01000", --  625
    X"80200b00010b", --  626
    X"22200280211b", --  627
    X"d0000083f0ca", --  628
    X"000023d10000", --  629
    X"d1020080300a", --  630
    X"80200b000114", --  631
    X"12200280211b", --  632
    X"c04f79133002", --  633
    X"c0004bc051ba", --  634
    X"802fcad80002", --  635
    X"80200b812fda", --  636
    X"20000080211b", --  637
    X"802fead90001", --  638
    X"000008812ffa", --  639
    X"04061786300a", --  640
    X"80200a844011", --  641
    X"20000081201a", --  642
    X"872fda862fca", --  643
    X"000603266000", --  644
    X"80200b000407", --  645
    X"32200280211b", --  646
    X"8e98e9199001", --  647
    X"81201a80200a", --  648
    X"86300a000023", --  649
    X"006714d70200", --  650
    X"80211b80200b", --  651
    X"022802022802", --  652
    X"188001133002", --  653
    X"81f02a80f01a", --  654
    X"83f04a82f03a", --  655
    X"85f06a84f05a", --  656
    X"87f08a86f07a", --  657
    X"89f0aa88f09a", --  658
    X"00e01a1ff00c", --  659
    X"80f01b3ff00d", --  660
    X"80f23b80f12b", --  661
    X"80f45b80f34b", --  662
    X"80f67b80f56b", --  663
    X"80f0ba80f78b", --  664
    X"c0004430001f", --  665
    X"d10000d00000", --  666
    X"80f0cac05468", --  667
    X"82f0ba81f0da", --  668
    X"c020b0000210", --  669
    X"87f0da86f0ca", --  670
    X"d50000d40001", --  671
    X"04420e322001", --  672
    X"077518066418", --  673
    X"200001c06021", --  674
    X"80f1ab80f09b", --  675
    X"81f02a80f01a", --  676
    X"83f04a82f03a", --  677
    X"85f06a84f05a", --  678
    X"87f08a86f07a", --  679
    X"00e01a1ff00d", --  680
    X"80f01b3ff00f", --  681
    X"80f23b80f12b", --  682
    X"80f45b80f34b", --  683
    X"80f67b80f56b", --  684
    X"80f89b80f78b", --  685
    X"80fabb80f9ab", --  686
    X"81f0ea80fbcb", --  687
    X"00010680f0fa", --  688
    X"0bb0048bf0da", --  689
    X"1bb003c0b036", --  690
    X"89f0fa300001", --  691
    X"1aa0288af0fa", --  692
    X"100001110000", --  693
    X"120000d414fd", --  694
    X"d514fd044b02", --  695
    X"155003d60000", --  696
    X"055b06d70000", --  697
    X"c05789006023", --  698
    X"c000abc0581a", --  699
    X"87400a86100a", --  700
    X"88500a83200a", --  701
    X"122001066713", --  702
    X"155003144003", --  703
    X"311001063813", --  704
    X"80960b066009", --  705
    X"8e9a59199001", --  706
    X"81f02a80f01a", --  707
    X"83f04a82f03a", --  708
    X"85f06a84f05a", --  709
    X"87f08a86f07a", --  710
    X"89f0aa88f09a", --  711
    X"8bf0ca8af0ba", --  712
    X"00e01a1ff00f", --  713
    X"80f01b3ff00c", --  714
    X"80f23b80f12b", --  715
    X"80f45b80f34b", --  716
    X"80f67b80f56b", --  717
    X"80f89b80f78b", --  718
    X"80f0ca80f9ab", --  719
    X"11000a88f0ba", --  720
    X"d9517d82000a", --  721
    X"83208202290a", --  722
    X"042418d400ff", --  723
    X"c0502035303f", --  724
    X"d20dc5d3003f", --  725
    X"82200a022302", --  726
    X"8660d306240b", --  727
    X"022302d20d85", --  728
    X"05260282200a", --  729
    X"10000180850b", --  730
    X"8e01b9188001", --  731
    X"81f02a80f01a", --  732
    X"83f04a82f03a", --  733
    X"85f06a84f05a", --  734
    X"87f08a86f07a", --  735
    X"89f0aa88f09a", --  736
    X"00e01a1ff00c", --  737
    X"80f01b3ff00f", --  738
    X"80f23b80f12b", --  739
    X"80fe9b80f34b", --  740
    X"d10000d00000", --  741
    X"c05d19000023", --  742
    X"c0028bc05d3a", --  743
    X"80200a82f0ea", --  744
    X"000013122001", --  745
    X"8ff0fb80f10b", --  746
    X"80ffdabe05ff", --  747
    X"d29fac81ffea", --  748
    X"000023000217", --  749
    X"902020d27f4c", --  750
    X"0000238000a1", --  751
    X"c05e9ac05e59", --  752
    X"d2151cc0004b", --  753
    X"80200a83f0fa", --  754
    X"81300a122001", --  755
    X"000113133001", --  756
    X"d0153f80f1db", --  757
    X"80008300100b", --  758
    X"d2000e000008", --  759
    X"8ff0fb80f20b", --  760
    X"82ffdabe062f", --  761
    X"31100e80f2db", --  762
    X"80f1cb011004", --  763
    X"81f02a80f01a", --  764
    X"83f04a82f03a", --  765
    X"1ff00f8ef09a", --  766
    X"3ff00a00e01a", --  767
    X"80f12b80f01b", --  768
    X"80f34b80f23b", --  769
    X"80f56b80f45b", --  770
    X"81f0aa80f09a", --  771
    X"d00000c00053", --  772
    X"80f07b80f08b", --  773
    X"020012c06278", --  774
    X"32201e00020e", --  775
    X"80f28b022004", --  776
    X"121000800093", --  777
    X"130000800013", --  778
    X"033418d47fff", --  779
    X"d00000322020", --  780
    X"011202d115cc", --  781
    X"d415cc81100a", --  782
    X"84400a044202", --  783
    X"055202d515cc", --  784
    X"04450685501a", --  785
    X"004314000023", --  786
    X"80f01a80f17b", --  787
    X"82f03a81f02a", --  788
    X"84f05a83f04a", --  789
    X"1ff00a85f06a", --  790
    X"3ff00b00e01a", --  791
    X"80f12b80f01b", --  792
    X"80f34b80f23b", --  793
    X"80f56b80f45b", --  794
    X"80f0aa80fe7b", --  795
    X"121000600020", --  796
    X"130000800013", --  797
    X"033418d47fff", --  798
    X"d115abd00000", --  799
    X"81100a011202", --  800
    X"d515ab141000", --  801
    X"85501a055202", --  802
    X"000023044506", --  803
    X"84f0ba004314", --  804
    X"04400434401e", --  805
    X"8ff0fb80f10b", --  806
    X"be065d8ff4eb", --  807
    X"80ffca81ffda", --  808
    X"80f08b80f19b", --  809
    X"81f02a80f01a", --  810
    X"83f04a82f03a", --  811
    X"85f06a84f05a", --  812
    X"1ff00b8ef07a", --  813
    X"3ff00b00e01a", --  814
    X"80f12b80f01b", --  815
    X"80f34b80f23b", --  816
    X"80f56b80f45b", --  817
    X"11000080f09a", --  818
    X"c0104031101f", --  819
    X"d50000d40000", --  820
    X"82f0aac06758", --  821
    X"04201083f0ba", --  822
    X"300001c00070", --  823
    X"d10001022010", --  824
    X"c02020022118", --  825
    X"80f47b244001", --  826
    X"80f01a80f58b", --  827
    X"82f03a81f02a", --  828
    X"84f05a83f04a", --  829
    X"1ff00b85f06a", --  830
    X"3ff00800e01a", --  831
    X"80f12b80f01b", --  832
    X"80f34b80f23b", --  833
    X"80f08a80fe5b", --  834
    X"80013b81002a", --  835
    X"80012b81001a", --  836
    X"80011b81000a", --  837
    X"80f00b80f07a", --  838
    X"8ff0fb80f06a", --  839
    X"81ffeabe05ff", --  840
    X"31100d80ffda", --  841
    X"d20000131000", --  842
    X"920001002023", --  843
    X"d260548220d1", --  844
    X"80f08a03320a", --  845
    X"80f01a80030b", --  846
    X"82f03a81f02a", --  847
    X"8ef05a83f04a", --  848
    X"00e01a1ff008", --  849
    X"80f01b3ff00d", --  850
    X"80f23b80f12b", --  851
    X"80f45b80f34b", --  852
    X"80f67b80f56b", --  853
    X"80f89b80f78b", --  854
    X"80200a12f00c", --  855
    X"d47fff81201a", --  856
    X"c00215d53fff", --  857
    X"00020e020012", --  858
    X"02200432201e", --  859
    X"032318d30001", --  860
    X"800013c03022", --  861
    X"122001822012", --  862
    X"131000800093", --  863
    X"160000800013", --  864
    X"066018d07fff", --  865
    X"d015ed333010", --  866
    X"81000a000302", --  867
    X"d715edd00000", --  868
    X"177001077302", --  869
    X"07170687700a", --  870
    X"007614000023", --  871
    X"12f00a000210", --  872
    X"80211b80200b", --  873
    X"81f02a80f01a", --  874
    X"83f04a82f03a", --  875
    X"85f06a84f05a", --  876
    X"87f08a86f07a", --  877
    X"1ff00d88f09a", --  878
    X"3ff00200e01a", --  879
    X"80f12b80f01b", --  880
    X"d10000d0047c", --  881
    X"80011b80010b", --  882
    X"80013b80012b", --  883
    X"80015b80014b", --  884
    X"81f02a80f01a", --  885
    X"00e01a1ff002", --  886
    X"80f01b3ff00f", --  887
    X"80f23b80f12b", --  888
    X"80f45b80f34b", --  889
    X"80f67b80f56b", --  890
    X"80f89b80f78b", --  891
    X"80fabb80f9ab", --  892
    X"80fcdb80fbcb", --  893
    X"d6047c80fdeb", --  894
    X"81601a80600a", --  895
    X"83603a82602a", --  896
    X"85605a84604a", --  897
    X"c0708989f0fa", --  898
    X"c0050bc071da", --  899
    X"d83ddc86900a", --  900
    X"d8e20d0a2817", --  901
    X"0aac030c4817", --  902
    X"d81e1300a023", --  903
    X"d8c3da0a6813", --  904
    X"d81e130a0813", --  905
    X"8aa0210a1813", --  906
    X"106000110000", --  907
    X"06600986a011", --  908
    X"19900180960b", --  909
    X"02a008242000", --  910
    X"80600bd6047c", --  911
    X"80622b80611b", --  912
    X"80644b80633b", --  913
    X"80f01a80655b", --  914
    X"82f03a81f02a", --  915
    X"84f05a83f04a", --  916
    X"86f07a85f06a", --  917
    X"88f09a87f08a", --  918
    X"8af0ba89f0aa", --  919
    X"8cf0da8bf0ca", --  920
    X"1ff00f8df0ea", --  921
    X"3ff01400e01a", --  922
    X"80f12b80f01b", --  923
    X"80f34b80f23b", --  924
    X"80f56b80f45b", --  925
    X"80f78b80f67b", --  926
    X"80f9ab80f89b", --  927
    X"80fbcb80fabb", --  928
    X"80fdeb80fcdb", --  929
    X"80f12a80fefb", --  930
    X"01100681f13a", --  931
    X"d38000d20000", --  932
    X"84f11a150000", --  933
    X"d60000144001", --  934
    X"006023d70000", --  935
    X"19100088f13a", --  936
    X"c0759ac07559", --  937
    X"86800ac0028b", --  938
    X"18800187900a", --  939
    X"066713199001", --  940
    X"c0a0310a6207", --  941
    X"105000226000", --  942
    X"155001311001", --  943
    X"d600018e54d9", --  944
    X"006023d70000", --  945
    X"08800688f13a", --  946
    X"c076dac07699", --  947
    X"86800ac0014b", --  948
    X"1880028a801a", --  949
    X"06aa13066613", --  950
    X"db0000da0001", --  951
    X"88f13a00a023", --  952
    X"c0779ac07759", --  953
    X"8a800ac0014b", --  954
    X"18800284801a", --  955
    X"0a44130aaa13", --  956
    X"d20000c02037", --  957
    X"242000d30000", --  958
    X"c0c0210c6407", --  959
    X"0ca407246000", --  960
    X"24a000c0c021", --  961
    X"02290e094012", --  962
    X"06690e042009", --  963
    X"0aa90e056009", --  964
    X"0c440b09a009", --  965
    X"82201302590b", --  966
    X"c0c0b70cc207", --  967
    X"c0798ac07959", --  968
    X"88f14ac0028b", --  969
    X"80800a89f10a", --  970
    X"80900b188001", --  971
    X"c07bf8199001", --  972
    X"399001094506", --  973
    X"d65555c09044", --  974
    X"c07af8d72aab", --  975
    X"04480ad84000", --  976
    X"855012844012", --  977
    X"c09080094502", --  978
    X"8ff9fb80f40b", --  979
    X"87ffeabe00cf", --  980
    X"069706d97fff", --  981
    X"d70000c07af8", --  982
    X"c07b69d67fff", --  983
    X"c0028bc07bea", --  984
    X"88f14a85f14a", --  985
    X"89f10a088006", --  986
    X"1880018a800a", --  987
    X"8b500a0a7a0a", --  988
    X"0b6b0a155001", --  989
    X"809a0b0aab02", --  990
    X"80f01a199001", --  991
    X"82f03a81f02a", --  992
    X"84f05a83f04a", --  993
    X"86f07a85f06a", --  994
    X"88f09a87f08a", --  995
    X"8af0ba89f0aa", --  996
    X"8cf0da8bf0ca", --  997
    X"8ef0fa8df0ea", --  998
    X"00e01a1ff014", --  999
    X"80f01b3ff008", -- 1000
    X"80f23b80f12b", -- 1001
    X"80f45b80f34b", -- 1002
    X"81f08a80f56b", -- 1003
    X"311001111028", -- 1004
    X"80100a321001", -- 1005
    X"c07e8ac07e29", -- 1006
    X"333001d30028", -- 1007
    X"83f07a00301e", -- 1008
    X"32200184200a", -- 1009
    X"85100a04340a", -- 1010
    X"80140b045406", -- 1011
    X"d405f0311001", -- 1012
    X"04340a84400a", -- 1013
    X"04540685100a", -- 1014
    X"d405f080140b", -- 1015
    X"80f01a80400b", -- 1016
    X"82f03a81f02a", -- 1017
    X"84f05a83f04a", -- 1018
    X"1ff00885f06a", -- 1019
    X"3ff03900e01a", -- 1020
    X"80f12b80f01b", -- 1021
    X"80f34b80f23b", -- 1022
    X"80f56b80f45b", -- 1023
    X"80f78b80f67b", -- 1024
    X"80f9ab80f89b", -- 1025
    X"80fbcb80fabb", -- 1026
    X"80fdeb80fcdb", -- 1027
    X"c080e980fefb", -- 1028
    X"c0028bc0812a", -- 1029
    X"11f01080f38a", -- 1030
    X"10000182000a", -- 1031
    X"80120b822022", -- 1032
    X"d20000111001", -- 1033
    X"002023d30000", -- 1034
    X"c081cac081a9", -- 1035
    X"11f010c0028b", -- 1036
    X"11100182100a", -- 1037
    X"c02053022213", -- 1038
    X"d10000d005f1", -- 1039
    X"c0864880010b", -- 1040
    X"377001072012", -- 1041
    X"04200902270e", -- 1042
    X"c082fac082b9", -- 1043
    X"80f39ac0028b", -- 1044
    X"82000a11f010", -- 1045
    X"822022100001", -- 1046
    X"11100180120b", -- 1047
    X"d30000d20000", -- 1048
    X"c08379002023", -- 1049
    X"c0028bc0839a", -- 1050
    X"82100a11f010", -- 1051
    X"022213111001", -- 1052
    X"d60000c02033", -- 1053
    X"012012c08548", -- 1054
    X"05200902210e", -- 1055
    X"80f40b017106", -- 1056
    X"be00cf8ff5fb", -- 1057
    X"c0203682ffea", -- 1058
    X"c08498d38001", -- 1059
    X"822071d30000", -- 1060
    X"80f30b022110", -- 1061
    X"be06a48ff2fb", -- 1062
    X"82ffda83ffea", -- 1063
    X"012009822091", -- 1064
    X"06160ad60ccc", -- 1065
    X"85500ad505f1", -- 1066
    X"c0861ac085b9", -- 1067
    X"81f38ac0028b", -- 1068
    X"05570ad77333", -- 1069
    X"82100a055602", -- 1070
    X"82203102250b", -- 1071
    X"11100180130b", -- 1072
    X"80450bd405f1", -- 1073
    X"81f02a80f01a", -- 1074
    X"83f04a82f03a", -- 1075
    X"85f06a84f05a", -- 1076
    X"87f08a86f07a", -- 1077
    X"89f0aa88f09a", -- 1078
    X"8bf0ca8af0ba", -- 1079
    X"8df0ea8cf0da", -- 1080
    X"1ff0398ef0fa", -- 1081
    X"3ff00200e01a", -- 1082
    X"80f12b80f01b", -- 1083
    X"c087eac087d9", -- 1084
    X"d005f2c000ab", -- 1085
    X"80010bd10000", -- 1086
    X"c08859100001", -- 1087
    X"d0008fc0886a", -- 1088
    X"00001e100028", -- 1089
    X"80010bd00482", -- 1090
    X"c088d9100001", -- 1091
    X"d0008fc088ea", -- 1092
    X"00001e100028", -- 1093
    X"80010bd00539", -- 1094
    X"80f01a100001", -- 1095
    X"1ff00281f02a", -- 1096
    X"3ff0b000e01a", -- 1097
    X"80f12b80f01b", -- 1098
    X"80f34b80f23b", -- 1099
    X"80f56b80f45b", -- 1100
    X"80f78b80f67b", -- 1101
    X"11f0af80fe9b", -- 1102
    X"d1000080100a", -- 1103
    X"82300a13f0ae", -- 1104
    X"12200183200a", -- 1105
    X"143006333003", -- 1106
    X"c0503035408f", -- 1107
    X"334006d4008f", -- 1108
    X"d5466680f00b", -- 1109
    X"d5000a8ff5fb", -- 1110
    X"15f0828ff5eb", -- 1111
    X"be00158ff5db", -- 1112
    X"8ff5fbd5599a", -- 1113
    X"8ff5db15f08d", -- 1114
    X"15f082be0015", -- 1115
    X"15f0b080f50b", -- 1116
    X"05510285500a", -- 1117
    X"d505118ff5fb", -- 1118
    X"be003e8ff5eb", -- 1119
    X"c08c8ac08c49", -- 1120
    X"d605c8c0028b", -- 1121
    X"15500187500a", -- 1122
    X"80670b877022", -- 1123
    X"d50511166001", -- 1124
    X"d505c880f50b", -- 1125
    X"8ff3eb8ff5fb", -- 1126
    X"15f00a8ff4db", -- 1127
    X"be07358ff5cb", -- 1128
    X"80f50b15f082", -- 1129
    X"8ff5fb15f098", -- 1130
    X"155001d5000a", -- 1131
    X"be00008ff5eb", -- 1132
    X"c08e5ac08e49", -- 1133
    X"35500ad50016", -- 1134
    X"00501e355001", -- 1135
    X"15500a15f098", -- 1136
    X"d60000155001", -- 1137
    X"15500180560b", -- 1138
    X"80f50b15f08d", -- 1139
    X"8ff5fb15f098", -- 1140
    X"d500168ff5eb", -- 1141
    X"15f0988ff5db", -- 1142
    X"15500115500a", -- 1143
    X"d500008ff5cb", -- 1144
    X"be00758ff5bb", -- 1145
    X"84300a13f098", -- 1146
    X"04440b133001", -- 1147
    X"c08fe9004023", -- 1148
    X"d50016c0900a", -- 1149
    X"00501e355001", -- 1150
    X"13300184300a", -- 1151
    X"165000044413", -- 1152
    X"84300a13f098", -- 1153
    X"85300a133001", -- 1154
    X"00402304450b", -- 1155
    X"c0910ac090d9", -- 1156
    X"355002d50016", -- 1157
    X"84300a00501e", -- 1158
    X"13300185301a", -- 1159
    X"175000044513", -- 1160
    X"d70000c07022", -- 1161
    X"07750ad56666", -- 1162
    X"8ff6fb80f70b", -- 1163
    X"87ffeabe00cf", -- 1164
    X"80f50b15f00a", -- 1165
    X"be07d08ff7fb", -- 1166
    X"80f50b15f08d", -- 1167
    X"8ff5fb15f00a", -- 1168
    X"05510215f032", -- 1169
    X"d500288ff5eb", -- 1170
    X"d505f28ff5db", -- 1171
    X"d500018ff5cb", -- 1172
    X"be00758ff5bb", -- 1173
    X"85500a15f0b0", -- 1174
    X"80f50b055102", -- 1175
    X"05510215f032", -- 1176
    X"be07f98ff5fb", -- 1177
    X"155028d50511", -- 1178
    X"80f50b35508f", -- 1179
    X"35508fd50511", -- 1180
    X"d5008f8ff5fb", -- 1181
    X"be00008ff5eb", -- 1182
    X"155028d505c8", -- 1183
    X"80f50b35508f", -- 1184
    X"35508fd505c8", -- 1185
    X"d5008f8ff5fb", -- 1186
    X"be00008ff5eb", -- 1187
    X"10000110000a", -- 1188
    X"351050111028", -- 1189
    X"15f0b0cf5564", -- 1190
    X"15505085500a", -- 1191
    X"80f50b35500a", -- 1192
    X"85500a15f0b0", -- 1193
    X"8ff5fb35500a", -- 1194
    X"8ff5ebd5000a", -- 1195
    X"15f032be0000", -- 1196
    X"15f0b080f50b", -- 1197
    X"8ff5fb85500a", -- 1198
    X"8ff5ebd50050", -- 1199
    X"80f01abe0000", -- 1200
    X"82f03a81f02a", -- 1201
    X"84f05a83f04a", -- 1202
    X"86f07a85f06a", -- 1203
    X"8ef09a87f08a", -- 1204
    X"00e01a1ff0b0", -- 1205
    X"d00427df0bff", -- 1206
    X"80010bd17530", -- 1207
    X"80011bd16590", -- 1208
    X"80012bd15208", -- 1209
    X"80013bd13a98", -- 1210
    X"80014bd11f40", -- 1211
    X"80015bd10000", -- 1212
    X"80016bd1e0c0", -- 1213
    X"80017bd1c568", -- 1214
    X"80018bd1adf8", -- 1215
    X"80019bd19a70", -- 1216
    X"d10923d00467", -- 1217
    X"d1124780010b", -- 1218
    X"d11b6a80011b", -- 1219
    X"d1248e80012b", -- 1220
    X"d12db280013b", -- 1221
    X"d136d580014b", -- 1222
    X"d13ff980015b", -- 1223
    X"d1491d80016b", -- 1224
    X"d1524080017b", -- 1225
    X"d15b6480018b", -- 1226
    X"c099c980019b", -- 1227
    X"c000abc099da", -- 1228
    X"d10000d00601", -- 1229
    X"10000180010b", -- 1230
    X"d10000d0065b", -- 1231
    X"be0b5f80010b", -- 1232
    X"be06dfbe0875", -- 1233
    X"d10000d005f0", -- 1234
    X"d005f180010b", -- 1235
    X"80010bd11000", -- 1236
    X"d15555d005fc", -- 1237
    X"d005fd80010b", -- 1238
    X"80010bd1c800", -- 1239
    X"80012b80011b", -- 1240
    X"00001d80013b", -- 1241
    X"80f01b3ff015", -- 1242
    X"80f23b80f12b", -- 1243
    X"80f45b80f34b", -- 1244
    X"80f67b80f56b", -- 1245
    X"80f13a80fe8b", -- 1246
    X"830109d10000", -- 1247
    X"81000a80f15a", -- 1248
    X"d20001811072", -- 1249
    X"81000a031218", -- 1250
    X"322001d20080", -- 1251
    X"81001a041218", -- 1252
    X"d20020811052", -- 1253
    X"051218322001", -- 1254
    X"d2002081001a", -- 1255
    X"061218322001", -- 1256
    X"8ff5fb80f40b", -- 1257
    X"d114858ff6eb", -- 1258
    X"72200ad20004", -- 1259
    X"01120202230c", -- 1260
    X"d1043f8ff1db", -- 1261
    X"81f14a8ff1cb", -- 1262
    X"d114d58ff1bb", -- 1263
    X"02230cd2000a", -- 1264
    X"8ff1ab011202", -- 1265
    X"81f14abe0354", -- 1266
    X"d1047280f10b", -- 1267
    X"d1000a8ff1fb", -- 1268
    X"be00008ff1eb", -- 1269
    X"80130bd10471", -- 1270
    X"d10472c0a0f8", -- 1271
    X"81f14a80f10b", -- 1272
    X"d1000a8ff1fb", -- 1273
    X"be00008ff1eb", -- 1274
    X"83100ad10471", -- 1275
    X"80f10bd10472", -- 1276
    X"8ff1fb11f009", -- 1277
    X"d20004d11485", -- 1278
    X"02230c72200a", -- 1279
    X"8ff1eb011202", -- 1280
    X"8ff1dbd1043f", -- 1281
    X"d2000ad114e9", -- 1282
    X"01120202230c", -- 1283
    X"be01ce8ff1cb", -- 1284
    X"80f10b11f009", -- 1285
    X"8ff1fbd1043f", -- 1286
    X"80f01abe03e9", -- 1287
    X"82f03a81f02a", -- 1288
    X"84f05a83f04a", -- 1289
    X"86f07a85f06a", -- 1290
    X"1ff0158ef08a", -- 1291
    X"3ff01000e01a", -- 1292
    X"80f12b80f01b", -- 1293
    X"80f10a80fe3b", -- 1294
    X"10f00480f00b", -- 1295
    X"80f0ea8ff0fb", -- 1296
    X"be09b48ff0eb", -- 1297
    X"80f00b10f004", -- 1298
    X"8ff0fb80f0fa", -- 1299
    X"80f01abe0594", -- 1300
    X"8ef03a81f02a", -- 1301
    X"00e01a1ff010", -- 1302
    X"80f01b3ff00a", -- 1303
    X"80f23b80f12b", -- 1304
    X"80f45b80f34b", -- 1305
    X"83f07a82f08a", -- 1306
    X"c0015280f09a", -- 1307
    X"3100c580f0aa", -- 1308
    X"110002c010d6", -- 1309
    X"01140ad42aab", -- 1310
    X"80210b111013", -- 1311
    X"011102141000", -- 1312
    X"010106011402", -- 1313
    X"80310b11103a", -- 1314
    X"310070c0a638", -- 1315
    X"d1000080210b", -- 1316
    X"c0a63880310b", -- 1317
    X"81100a81f08a", -- 1318
    X"341014311005", -- 1319
    X"d10014c04026", -- 1320
    X"35408f141009", -- 1321
    X"d4008fc05030", -- 1322
    X"80f0aa314009", -- 1323
    X"d42aab150002", -- 1324
    X"35500105540a", -- 1325
    X"80240b045102", -- 1326
    X"054502045502", -- 1327
    X"044506340002", -- 1328
    X"80f01a80340b", -- 1329
    X"82f03a81f02a", -- 1330
    X"84f05a83f04a", -- 1331
    X"1ff00a85f06a", -- 1332
    X"3ff00600e01a", -- 1333
    X"80f12b80f01b", -- 1334
    X"80f34b80f23b", -- 1335
    X"80400ad405fc", -- 1336
    X"00020bd27c4d", -- 1337
    X"d23619800013", -- 1338
    X"000203d30000", -- 1339
    X"80f06b80400b", -- 1340
    X"81f02a80f01a", -- 1341
    X"83f04a82f03a", -- 1342
    X"1ff00684f05a", -- 1343
    X"3ff00f00e01a", -- 1344
    X"80f12b80f01b", -- 1345
    X"80f34b80f23b", -- 1346
    X"80f56b80f45b", -- 1347
    X"81f0ea10f009", -- 1348
    X"021318d30007", -- 1349
    X"022302832020", -- 1350
    X"81103280020b", -- 1351
    X"021318d30007", -- 1352
    X"022302832020", -- 1353
    X"80021b122001", -- 1354
    X"d30007811032", -- 1355
    X"832020021318", -- 1356
    X"122002022302", -- 1357
    X"81103280022b", -- 1358
    X"041318d30001", -- 1359
    X"d30007811012", -- 1360
    X"832020021318", -- 1361
    X"122003022302", -- 1362
    X"80023b022402", -- 1363
    X"c0aaeac0aad9", -- 1364
    X"82f0dac0028b", -- 1365
    X"80230bd30000", -- 1366
    X"c0ab69122001", -- 1367
    X"c0004bc0ac1a", -- 1368
    X"d5e000d21fff", -- 1369
    X"81f0fa84f0da", -- 1370
    X"021318d30001", -- 1371
    X"83000a811012", -- 1372
    X"054302100001", -- 1373
    X"802338d30000", -- 1374
    X"c0ac18d21fff", -- 1375
    X"80520bd2e000", -- 1376
    X"81f02a80f01a", -- 1377
    X"83f04a82f03a", -- 1378
    X"85f06a84f05a", -- 1379
    X"00e01a1ff00f", -- 1380
    X"80f01b3ff014", -- 1381
    X"80f23b80f12b", -- 1382
    X"80f45b80f34b", -- 1383
    X"80f67b80f56b", -- 1384
    X"80f89b80f78b", -- 1385
    X"80fabb80f9ab", -- 1386
    X"80fcdb80fbcb", -- 1387
    X"80fefb80fdeb", -- 1388
    X"d1000080f12a", -- 1389
    X"82f11a810128", -- 1390
    X"d1733380200a", -- 1391
    X"03010600010a", -- 1392
    X"d07333c03020", -- 1393
    X"82f10a80200b", -- 1394
    X"d17d6f80200a", -- 1395
    X"80200b00010a", -- 1396
    X"80f00bd005fd", -- 1397
    X"c0b248be0b35", -- 1398
    X"81004280f14a", -- 1399
    X"011302d3157c", -- 1400
    X"d2001081100a", -- 1401
    X"020218322001", -- 1402
    X"022302d31584", -- 1403
    X"73100282200a", -- 1404
    X"030302d01520", -- 1405
    X"74200283300a", -- 1406
    X"040402d01530", -- 1407
    X"03340284400a", -- 1408
    X"80530b85f11a", -- 1409
    X"80f50bd505fd", -- 1410
    X"8ff5fbd5065c", -- 1411
    X"83ffeabe05c4", -- 1412
    X"76100284ffda", -- 1413
    X"d01520166001", -- 1414
    X"86600a060602", -- 1415
    X"782002d70000", -- 1416
    X"d01530188001", -- 1417
    X"88800a080802", -- 1418
    X"066803d90000", -- 1419
    X"08830b886013", -- 1420
    X"155004054004", -- 1421
    X"85f10a08850e", -- 1422
    X"d505fd80590b", -- 1423
    X"8ff7fb80f50b", -- 1424
    X"be067f8ff6eb", -- 1425
    X"81f02a80f01a", -- 1426
    X"83f04a82f03a", -- 1427
    X"85f06a84f05a", -- 1428
    X"87f08a86f07a", -- 1429
    X"89f0aa88f09a", -- 1430
    X"8bf0ca8af0ba", -- 1431
    X"8df0ea8cf0da", -- 1432
    X"1ff0148ef0fa", -- 1433
    X"3ff00800e01a", -- 1434
    X"80f12b80f01b", -- 1435
    X"80f34b80f23b", -- 1436
    X"d0000080f45b", -- 1437
    X"c0b419d10000", -- 1438
    X"c0004bc0b47a", -- 1439
    X"82400a84f08a", -- 1440
    X"c02036144001", -- 1441
    X"c0b478d3ffff", -- 1442
    X"000203d30000", -- 1443
    X"d41000800023", -- 1444
    X"d1c800000406", -- 1445
    X"c01026010106", -- 1446
    X"c0b549d0c800", -- 1447
    X"c0003bc0b56a", -- 1448
    X"12200382f08a", -- 1449
    X"322001812ffa", -- 1450
    X"80200b80211b", -- 1451
    X"81f02a80f01a", -- 1452
    X"83f04a82f03a", -- 1453
    X"1ff00884f05a", -- 1454
    X"3ff00700e01a", -- 1455
    X"80f12b80f01b", -- 1456
    X"80f34b80f23b", -- 1457
    X"80f56b80f45b", -- 1458
    X"c0b6e980fe7b", -- 1459
    X"d0008fc0b6fa", -- 1460
    X"00001e10000b", -- 1461
    X"d10000d0033d", -- 1462
    X"10000180010b", -- 1463
    X"c0b76ac0b759", -- 1464
    X"d00431c000ab", -- 1465
    X"80010bd10000", -- 1466
    X"d0043b100001", -- 1467
    X"80010bd10ccd", -- 1468
    X"d1003cd0043c", -- 1469
    X"d1000080010b", -- 1470
    X"80010bd0043d", -- 1471
    X"80010bd0043e", -- 1472
    X"d2043fd10467", -- 1473
    X"d50004d4043f", -- 1474
    X"04450275500a", -- 1475
    X"d3000a80f10b", -- 1476
    X"8ff2fb8ff3eb", -- 1477
    X"12200abe0000", -- 1478
    X"d204728f24d9", -- 1479
    X"be00008ff2fb", -- 1480
    X"81f02a80f01a", -- 1481
    X"83f04a82f03a", -- 1482
    X"85f06a84f05a", -- 1483
    X"1ff0078ef07a", -- 1484
    X"d0069000e01a", -- 1485
    X"10000181000a", -- 1486
    X"d2068480f00b", -- 1487
    X"d2065b8ff2fb", -- 1488
    X"02120282200a", -- 1489
    X"be0a198ff2eb", -- 1490
    X"d20427100002", -- 1491
    X"d2068480f20b", -- 1492
    X"d206a18ff2fb", -- 1493
    X"be04488ff2eb", -- 1494
    X"80f20bd20684", -- 1495
    X"8ff2fbd20427", -- 1496
    X"8ff2ebd2000a", -- 1497
    X"d206a1be0000", -- 1498
    X"d806b7d30000", -- 1499
    X"12200a00001d", -- 1500
    X"133028122001", -- 1501
    X"d0033d00001d", -- 1502
    X"80f00b100050", -- 1503
    X"8ff0fbd0033d", -- 1504
    X"10000bd0008f", -- 1505
    X"be00008ff0eb", -- 1506
    X"84000a00001d", -- 1507
    X"c03212100001", -- 1508
    X"10000185000a", -- 1509
    X"c050f2051502", -- 1510
    X"8ff3fb80f40b", -- 1511
    X"8ff6ebd6068e", -- 1512
    X"8ff6dbd6068f", -- 1513
    X"d6068ebe0a2e", -- 1514
    X"d6068f85600a", -- 1515
    X"d6043c87600a", -- 1516
    X"c0c06880650b", -- 1517
    X"85600ad6043c", -- 1518
    X"80650bd6068e", -- 1519
    X"d70000d6068f", -- 1520
    X"15500180670b", -- 1521
    X"c0702037508f", -- 1522
    X"d6043cd5008f", -- 1523
    X"c0c06880650b", -- 1524
    X"80f40bc010f2", -- 1525
    X"d6068e8ff3fb", -- 1526
    X"d6068f8ff6eb", -- 1527
    X"be0a2e8ff6db", -- 1528
    X"85600ad6068e", -- 1529
    X"87600ad6068f", -- 1530
    X"80650bd6043c", -- 1531
    X"d6043cc0c068", -- 1532
    X"d6068e85600a", -- 1533
    X"d6068f80650b", -- 1534
    X"80670bd70000", -- 1535
    X"37508f155001", -- 1536
    X"d5008fc07020", -- 1537
    X"80650bd6043c", -- 1538
    X"85600ad6068e", -- 1539
    X"18800180850b", -- 1540
    X"066302d603d7", -- 1541
    X"d6068e80f60b", -- 1542
    X"8ff6fb86600a", -- 1543
    X"86600ad6068f", -- 1544
    X"be05528ff6eb", -- 1545
    X"8017b8d70000", -- 1546
    X"85f00abe0a6b", -- 1547
    X"055718d71fff", -- 1548
    X"be0a6b80050b", -- 1549
    X"d7000f86f00a", -- 1550
    X"80061b066718", -- 1551
    --X"80f60b86001a", -- 1552
    X"8ff5fb85000a", -- 1553
    X"8ff7ebd7065c", -- 1554
    X"80f60b86001a", -- 1552 // fix
    X"100002be0a81", -- 1555
    X"87600ad6043b", -- 1556
    X"d6068e877010", -- 1557
    X"35602886600a", -- 1558
    X"c0c359c050e6", -- 1559
    X"055004c0c3ba", -- 1560
    X"d5065c00501e", -- 1561
    X"89500a065602", -- 1562
    X"09970a155001", -- 1563
    X"09a9028a600a", -- 1564
    X"16600180690b", -- 1565
    X"10000184000a", -- 1566
    X"d6065c80f40b", -- 1567
    X"8ff1eb8ff6fb", -- 1568
    X"8ff6dbd6043e", -- 1569
    X"8ff6cbd6043d", -- 1570
    X"85ffdabe0aca", -- 1571
    X"85600ad6043e", -- 1572
    X"87600ad6043d", -- 1573
    X"80650bd6043b", -- 1574
    X"065906d932d9", -- 1575
    X"d6043bc06030", -- 1576
    X"d90ccd80690b", -- 1577
    X"c06036065906", -- 1578
    X"80690bd6043b", -- 1579
    X"c0c67ac0c5e9", -- 1580
    X"d603d7c0028b", -- 1581
    X"dc065c066302", -- 1582
    X"0a950b89600a", -- 1583
    X"89c00a00a023", -- 1584
    X"0a97131cc001", -- 1585
    X"09a0098aa011", -- 1586
    X"16600180690b", -- 1587
    X"80f20b000021", -- 1588
    X"066302d603d7", -- 1589
    X"d6060b8ff6fb", -- 1590
    X"8ff6eb066302", -- 1591
    X"8ff6dbd60028", -- 1592
    X"8ff6cbd60431", -- 1593
    X"8ff6bbd60000", -- 1594
    X"060020be0075", -- 1595
    X"8169b8d90000", -- 1596
    X"c0c84ac0c819", -- 1597
    X"16600bd6008f", -- 1598
    X"00601e166050", -- 1599
    X"89600ad6033d", -- 1600
    X"80690b899022", -- 1601
    X"80f20b166001", -- 1602
    X"066302d603d7", -- 1603
    X"d6060b8ff6fb", -- 1604
    X"8ff6eb066302", -- 1605
    X"8ff6dbd60028", -- 1606
    X"8ff6cbd60431", -- 1607
    X"8ff6bbd60001", -- 1608
    X"c0c9e8be0075", -- 1609
    X"066302d6060b", -- 1610
    X"36600a166028", -- 1611
    X"d6043180f60b", -- 1612
    X"d6000a8ff6fb", -- 1613
    X"be00008ff6eb", -- 1614
    X"3ff00700001d", -- 1615
    X"80f12b80f01b", -- 1616
    X"80f34b80f23b", -- 1617
    X"80001280f07a", -- 1618
    X"c0cab9d10001", -- 1619
    X"c0006bc0cada", -- 1620
    X"800012d20001", -- 1621
    X"011302030218", -- 1622
    X"01100280f06a", -- 1623
    X"80f15b011218", -- 1624
    X"81f02a80f01a", -- 1625
    X"83f04a82f03a", -- 1626
    X"00e01a1ff007", -- 1627
    X"80f01b3ff008", -- 1628
    X"80f23b80f12b", -- 1629
    X"80f45b80f34b", -- 1630
    X"80f08a80f56b", -- 1631
    X"81000ad40690", -- 1632
    X"d200ff831082", -- 1633
    X"80421b023218", -- 1634
    X"031218d200ff", -- 1635
    X"8510e281001a", -- 1636
    X"025218d20003", -- 1637
    X"023219833020", -- 1638
    X"d23fff80422b", -- 1639
    X"853062031218", -- 1640
    X"025218d200ff", -- 1641
    X"d2003f80423b", -- 1642
    X"853052031218", -- 1643
    X"025218d20001", -- 1644
    X"d2001f80424b", -- 1645
    X"81002a031218", -- 1646
    X"d200ff851082", -- 1647
    X"833080025218", -- 1648
    X"80425b023219", -- 1649
    X"031218d200ff", -- 1650
    X"d2000f853042", -- 1651
    X"80426b025218", -- 1652
    X"031218d2000f", -- 1653
    X"8510d281003a", -- 1654
    X"025218d20007", -- 1655
    X"023219833030", -- 1656
    X"d21fff80427b", -- 1657
    X"853082031218", -- 1658
    X"025218d2001f", -- 1659
    X"d200ff80428b", -- 1660
    X"81004a031218", -- 1661
    X"d2001f8510b2", -- 1662
    X"833050025218", -- 1663
    X"80429b023219", -- 1664
    X"031218d207ff", -- 1665
    X"d2000f853072", -- 1666
    X"8042ab025218", -- 1667
    X"031218d2007f", -- 1668
    X"81000a8043bb", -- 1669
    X"01121982001a", -- 1670
    X"01121982002a", -- 1671
    X"01121982003a", -- 1672
    X"01121982004a", -- 1673
    X"d2000083f07a", -- 1674
    X"d20001801229", -- 1675
    X"80f01a80320b", -- 1676
    X"82f03a81f02a", -- 1677
    X"84f05a83f04a", -- 1678
    X"1ff00885f06a", -- 1679
    X"d0069c00e01a", -- 1680
    X"d0069080f00b", -- 1681
    X"be0cb88ff0fb", -- 1682
    X"80f10b81003a", -- 1683
    X"8ff1fb81004a", -- 1684
    X"81ffeabe0c9f", -- 1685
    X"00001d80014b", -- 1686
    X"d006b7000024", -- 1687
    X"81001a81000a", -- 1688
    X"80f00bd0060b", -- 1689
    X"8ff0fbd006a1", -- 1690
    X"8ff0ebd006b7", -- 1691
    X"d0060bbe0893", -- 1692
    X"be06ee80f00b", -- 1693
    X"3ff00900001d", -- 1694
    X"80f12b80f01b", -- 1695
    X"80f09a80f23b", -- 1696
    X"00010b81f07a", -- 1697
    X"80f09a000023", -- 1698
    X"02010a81f06a", -- 1699
    X"80f08a902001", -- 1700
    X"02010a81f07a", -- 1701
    X"80f04b902001", -- 1702
    X"80f01a80f15b", -- 1703
    X"82f03a81f02a", -- 1704
    X"00e01a1ff009", -- 1705
    X"80f01b3ff00c", -- 1706
    X"80f23b80f12b", -- 1707
    X"80f45b80f34b", -- 1708
    X"d03fff80fe6b", -- 1709
    X"80f0ca80f00b", -- 1710
    X"be00cf8ff0fb", -- 1711
    X"80f0ba84ffea", -- 1712
    X"00041781f0ca", -- 1713
    X"d37fffd2ffff", -- 1714
    X"000008002007", -- 1715
    X"000008000417", -- 1716
    X"83f0aa82f09a", -- 1717
    X"80f30b022008", -- 1718
    X"8ff1eb8ff2fb", -- 1719
    X"be0d3d8ff0db", -- 1720
    X"80ffba81ffca", -- 1721
    X"80f07b800021", -- 1722
    X"80f01a80f18b", -- 1723
    X"82f03a81f02a", -- 1724
    X"84f05a83f04a", -- 1725
    X"1ff00c8ef06a", -- 1726
    X"df0bff00e01a", -- 1727
    X"d10000d00000", -- 1728
    X"d30000d20000", -- 1729
    X"d50000d40000", -- 1730
    X"d70000d60000", -- 1731
    X"d90000d80000", -- 1732
    X"db0000da0000", -- 1733
    X"dd0000dc0000", -- 1734
    X"d102b9de0000", -- 1735
    X"80120bd27530", -- 1736
    X"80121bd26590", -- 1737
    X"80122bd25208", -- 1738
    X"80123bd23a98", -- 1739
    X"80124bd21f40", -- 1740
    X"80125bd20000", -- 1741
    X"80126bd2e0c0", -- 1742
    X"80127bd2c568", -- 1743
    X"80128bd2adf8", -- 1744
    X"80129bd29a70", -- 1745
    X"d10000d00000", -- 1746
    X"c0daaac0da99", -- 1747
    X"80100bc00f0b", -- 1748
    X"d101cf111001", -- 1749
    X"c0db2ac0db19", -- 1750
    X"12208fd20050", -- 1751
    X"80100b00201e", -- 1752
    X"d100f0111001", -- 1753
    X"c0dbbac0dba9", -- 1754
    X"12208fd20050", -- 1755
    X"00201e12200b", -- 1756
    X"11100180100b", -- 1757
    X"d202d7d102d7", -- 1758
    X"80100b12200a", -- 1759
    X"8f12e9111001", -- 1760
    X"d202cdd102cd", -- 1761
    X"80100b12200a", -- 1762
    X"8f12e9111001", -- 1763
    X"d202e1d102e1", -- 1764
    X"80100b12200a", -- 1765
    X"8f12e9111001", -- 1766
    X"d002ebd10ccd", -- 1767
    X"d102b980010b", -- 1768
    X"d102c380f10b", -- 1769
    X"d1000a8ff1fb", -- 1770
    X"be00008ff1eb", -- 1771
    X"d20923d1032b", -- 1772
    X"d2124780120b", -- 1773
    X"d21b6a80121b", -- 1774
    X"d2248e80122b", -- 1775
    X"d22db280123b", -- 1776
    X"d236d580124b", -- 1777
    X"d23ff980125b", -- 1778
    X"d2491d80126b", -- 1779
    X"d2524080127b", -- 1780
    X"d25b6480128b", -- 1781
    X"d1032b80129b", -- 1782
    X"d40303d20303", -- 1783
    X"75500ad50004", -- 1784
    X"80f10b044502", -- 1785
    X"8ff3ebd3000a", -- 1786
    X"be00008ff2fb", -- 1787
    X"8f24d912200a", -- 1788
    X"d10000d04000", -- 1789
    X"80200bd20335", -- 1790
    X"80202b80211b", -- 1791
    X"80204b80213b", -- 1792
    X"80206b80215b", -- 1793
    X"d002ff80217b", -- 1794
    X"80010bd1c800", -- 1795
    X"80012b80011b", -- 1796
    X"be0e0d80013b", -- 1797
    X"3ff00200001d", -- 1798
    X"80f12b80f01b", -- 1799
    X"d00000d102f9", -- 1800
    X"80101b80100b", -- 1801
    X"80103b80102b", -- 1802
    X"80105b80104b", -- 1803
    X"81f02a80f01a", -- 1804
    X"00e01a1ff002", -- 1805
    X"80f01b3ff00f", -- 1806
    X"80f23b80f12b", -- 1807
    X"80f45b80f34b", -- 1808
    X"80f67b80f56b", -- 1809
    X"80f9ab80f89b", -- 1810
    X"80fbcb80fabb", -- 1811
    X"80fdeb80fcdb", -- 1812
    X"80600ad602f9", -- 1813
    X"82602a81601a", -- 1814
    X"84604a83603a", -- 1815
    X"89f0fa85605a", -- 1816
    X"c0e47ac0e359", -- 1817
    X"d81e7fc0050b", -- 1818
    X"0a281786900a", -- 1819
    X"0c4817d8f16b", -- 1820
    X"242000d8f12a", -- 1821
    X"00a0230aac03", -- 1822
    X"0a08139a676b", -- 1823
    X"1100009a176b", -- 1824
    X"8aa031106000", -- 1825
    X"02a00806a009", -- 1826
    X"19900180960b", -- 1827
    X"80600bd602f9", -- 1828
    X"80622b80611b", -- 1829
    X"80644b80633b", -- 1830
    X"80f01a80655b", -- 1831
    X"82f03a81f02a", -- 1832
    X"84f05a83f04a", -- 1833
    X"87f08a85f06a", -- 1834
    X"89f0aa88f09a", -- 1835
    X"8bf0ca8af0ba", -- 1836
    X"8df0ea8cf0da", -- 1837
    X"00e01a1ff00f", -- 1838
    X"80f01b3ff0ff", -- 1839
    X"80f23b80f12b", -- 1840
    X"80f45b80f34b", -- 1841
    X"80f67b80f56b", -- 1842
    X"80f89b80f78b", -- 1843
    X"80fabb80f9ab", -- 1844
    X"d00c0080fbcb", -- 1845
    X"82200a12f0ff", -- 1846
    X"c0e72917f00d", -- 1847
    X"c00f0bc0e78a", -- 1848
    X"84000a85200a", -- 1849
    X"122001100001", -- 1850
    X"80760b065415", -- 1851
    X"000021177001", -- 1852
    X"d10000d00001", -- 1853
    X"12f00d000023", -- 1854
    X"c0e89ac0e819", -- 1855
    X"85200ac003cb", -- 1856
    X"8b202a8a201a", -- 1857
    X"1220048c203a", -- 1858
    X"04aa13045513", -- 1859
    X"04cc1304bb13", -- 1860
    X"c00130000020", -- 1861
    X"c0e90912f00d", -- 1862
    X"c003cbc0e9ca", -- 1863
    X"8a201a84200a", -- 1864
    X"8c203a8b202a", -- 1865
    X"8aa022844022", -- 1866
    X"8cc0228bb022", -- 1867
    X"802a1b80240b", -- 1868
    X"802c3b802b2b", -- 1869
    X"c0e798122004", -- 1870
    X"d2000a004012", -- 1871
    X"d1079904400e", -- 1872
    X"044008122001", -- 1873
    X"d107a480140b", -- 1874
    X"80150bd400f0", -- 1875
    X"d60000d10001", -- 1876
    X"006023d70000", -- 1877
    X"34400113f00d", -- 1878
    X"c0ebc9063102", -- 1879
    X"d50001c0ec3a", -- 1880
    X"c05060054518", -- 1881
    X"85600a87300a", -- 1882
    X"166001133001", -- 1883
    X"854012087513", -- 1884
    X"00002400501e", -- 1885
    X"85600a87300a", -- 1886
    X"8b601a8a301a", -- 1887
    X"166002133002", -- 1888
    X"08ab13087513", -- 1889
    X"d70799000024", -- 1890
    X"07710208800e", -- 1891
    X"80780b088008", -- 1892
    X"077102d707a4", -- 1893
    X"80790b111001", -- 1894
    X"80f01a8d12b9", -- 1895
    X"82f03a81f02a", -- 1896
    X"84f05a83f04a", -- 1897
    X"86f07a85f06a", -- 1898
    X"88f09a87f08a", -- 1899
    X"8af0ba89f0aa", -- 1900
    X"1ff0ff8bf0ca", -- 1901
    X"3ff00a00e01a", -- 1902
    X"80f12b80f01b", -- 1903
    X"80f34b80f23b", -- 1904
    X"80f56b80f45b", -- 1905
    X"80f08a80fe7b", -- 1906
    X"c0f00ac0eef9", -- 1907
    X"80f09a00001e", -- 1908
    X"81f0aa100001", -- 1909
    X"d20cf0111001", -- 1910
    X"84000ad30cfa", -- 1911
    X"84100a80f40b", -- 1912
    X"84200a8ff4fb", -- 1913
    X"8ff4eb122001", -- 1914
    X"13300184300a", -- 1915
    X"be0d3d8ff4db", -- 1916
    X"85ffca84ffba", -- 1917
    X"80140b044008", -- 1918
    X"80050b111001", -- 1919
    X"80f01a100001", -- 1920
    X"82f03a81f02a", -- 1921
    X"84f05a83f04a", -- 1922
    X"8ef07a85f06a", -- 1923
    X"00e01a1ff00a", -- 1924
    X"80f01b3ff040", -- 1925
    X"80f23b80f12b", -- 1926
    X"80f45b80f34b", -- 1927
    X"80f67b80f56b", -- 1928
    X"80f89b80f78b", -- 1929
    X"80fabb80f9ab", -- 1930
    X"80fcdb80fbcb", -- 1931
    X"80fefb80fdeb", -- 1932
    X"82201a82f3fa", -- 1933
    X"d80000622001", -- 1934
    X"89901a89f40a", -- 1935
    X"042001022803", -- 1936
    X"86600a86f3fa", -- 1937
    X"87700a87f40a", -- 1938
    X"8ff6fb80f70b", -- 1939
    X"8ff4db8ff5eb", -- 1940
    X"80ffbabe0d54", -- 1941
    X"c0202181ffca", -- 1942
    X"080008000005", -- 1943
    X"80690b86f3da", -- 1944
    X"000008800043", -- 1945
    X"80601b16f01c", -- 1946
    X"80611b16f011", -- 1947
    X"8ff8fb80f90b", -- 1948
    X"8ff8db8ff9eb", -- 1949
    X"80ffbabe0d3d", -- 1950
    X"00000181ffca", -- 1951
    X"d77fffd6ffff", -- 1952
    X"000008006007", -- 1953
    X"86600a86f3fa", -- 1954
    X"87700a87f40a", -- 1955
    X"8ff6db8ff7eb", -- 1956
    X"8ff0fb80f10b", -- 1957
    X"80ffbabe0d3d", -- 1958
    X"0c001281ffca", -- 1959
    X"0a0008000c0e", -- 1960
    X"d00000d60002", -- 1961
    X"c0f5a9d10000", -- 1962
    X"376001c0f70a", -- 1963
    X"d7000100701e", -- 1964
    X"02270282f3fa", -- 1965
    X"83f40a82200a", -- 1966
    X"83300a033702", -- 1967
    X"8ff2fb80f30b", -- 1968
    X"02260212f01c", -- 1969
    X"82200a022706", -- 1970
    X"03360213f011", -- 1971
    X"83300a033706", -- 1972
    X"8ff2db8ff3eb", -- 1973
    X"84ffbabe0d3d", -- 1974
    X"00040385ffca", -- 1975
    X"800041177001", -- 1976
    X"82f3fa81fc0b", -- 1977
    X"82200a022602", -- 1978
    X"8df40a622001", -- 1979
    X"8dd00a0dd602", -- 1980
    X"022c03dc0000", -- 1981
    X"0002038cf10a", -- 1982
    X"80fb0b020001", -- 1983
    X"8ff3eb8ffafb", -- 1984
    X"be0d548ff2db", -- 1985
    X"85ffca84ffba", -- 1986
    X"044005c00021", -- 1987
    X"084008044c0e", -- 1988
    X"07760287f3da", -- 1989
    X"0290008f79fb", -- 1990
    X"022706d77fee", -- 1991
    X"c0f969c02130", -- 1992
    X"c000abc0f99a", -- 1993
    X"d102ec80f3ea", -- 1994
    X"11100182100a", -- 1995
    X"12200180200b", -- 1996
    X"80000a80f3da", -- 1997
    X"80100bd102f7", -- 1998
    X"80001a80f3da", -- 1999
    X"80101bd102f7", -- 2000
    X"c0fa89c10258", -- 2001
    X"376001c0fcaa", -- 2002
    X"d7000100701e", -- 2003
    X"8ff8fb80f90b", -- 2004
    X"00060210f011", -- 2005
    X"80000a000706", -- 2006
    X"10f01c8ff0eb", -- 2007
    X"000706000602", -- 2008
    X"8ff0db80000a", -- 2009
    X"80ffbabe0d3d", -- 2010
    X"81fc0b81ffca", -- 2011
    X"0cc7021cf01c", -- 2012
    X"6cc0018cc00a", -- 2013
    X"03370213f011", -- 2014
    X"d2000083300a", -- 2015
    X"8cf10a022c03", -- 2016
    X"000008000203", -- 2017
    X"02270212f032", -- 2018
    X"13f02780200b", -- 2019
    X"80310b033702", -- 2020
    X"844043177001", -- 2021
    X"12f032044008", -- 2022
    X"80240b022602", -- 2023
    X"03360213f027", -- 2024
    X"80f90b80350b", -- 2025
    X"8ff9eb8ff8fb", -- 2026
    X"be0d3d8ff8db", -- 2027
    X"81ffca80ffba", -- 2028
    X"d2ffff000001", -- 2029
    X"002007d37fff", -- 2030
    X"80fb0b000008", -- 2031
    X"8ff1eb8ffafb", -- 2032
    X"be0d3d8ff0db", -- 2033
    X"81ffca80ffba", -- 2034
    X"00070e070012", -- 2035
    X"0cc7020a0008", -- 2036
    X"c0ffcac0ff59", -- 2037
    X"12f03200601e", -- 2038
    X"13f027122001", -- 2039
    X"14f01c133001", -- 2040
    X"15f011144001", -- 2041
    X"87200a155001", -- 2042
    X"80470b122001", -- 2043
    X"87300a144001", -- 2044
    X"80570b133001", -- 2045
    X"166001155001", -- 2046
    X"177001d7000a", -- 2047
    X"c0f538806728", -- 2048
    X"d6100087f3ea", -- 2049
    X"c1010980760b", -- 2050
    X"c000abc101ca", -- 2051
    X"12200112f01c", -- 2052
    X"13300113f011", -- 2053
    X"14400184f3ea", -- 2054
    X"155001d502ec", -- 2055
    X"12200180200a", -- 2056
    X"8d300a600001", -- 2057
    X"dc0000133001", -- 2058
    X"800011000c03", -- 2059
    X"80400b000009", -- 2060
    X"80500b144001", -- 2061
    X"80f3da155001", -- 2062
    X"d102f780000a", -- 2063
    X"80f3da80100b", -- 2064
    X"d102f780001a", -- 2065
    X"80f01a80101b", -- 2066
    X"82f03a81f02a", -- 2067
    X"84f05a83f04a", -- 2068
    X"86f07a85f06a", -- 2069
    X"88f09a87f08a", -- 2070
    X"8af0ba89f0aa", -- 2071
    X"8cf0da8bf0ca", -- 2072
    X"8ef0fa8df0ea", -- 2073
    X"00e01a1ff040", -- 2074
    X"80f01b3ff00f", -- 2075
    X"80f23b80f12b", -- 2076
    X"80f45b80f34b", -- 2077
    X"80f67b80f56b", -- 2078
    X"80f89b80f78b", -- 2079
    X"80fabb80f9ab", -- 2080
    X"d1000080f0da", -- 2081
    X"d20000830109", -- 2082
    X"84f0fad30080", -- 2083
    X"000023604100", -- 2084
    X"84401a84f0ea", -- 2085
    X"004513d51000", -- 2086
    X"c10559040008", -- 2087
    X"d80005c1066a", -- 2088
    X"00801e388002", -- 2089
    X"89f0fad80002", -- 2090
    X"800011004917", -- 2091
    X"d98000000023", -- 2092
    X"a02001003913", -- 2093
    X"09980289f0ea", -- 2094
    X"da100089900a", -- 2095
    X"060008009a13", -- 2096
    X"135000124000", -- 2097
    X"157000146000", -- 2098
    X"89f0fa188001", -- 2099
    X"000023004917", -- 2100
    X"003913d98000", -- 2101
    X"89f0eaa02001", -- 2102
    X"89900a099802", -- 2103
    X"009a13da0800", -- 2104
    X"c10a28800071", -- 2105
    X"d30100d20000", -- 2106
    X"60420084f0fa", -- 2107
    X"84f0ea000023", -- 2108
    X"d5100084401a", -- 2109
    X"040008004513", -- 2110
    X"c1095ac10849", -- 2111
    X"388002d80005", -- 2112
    X"d8000200801e", -- 2113
    X"00491789f0fa", -- 2114
    X"000023800011", -- 2115
    X"003913d98000", -- 2116
    X"89f0eaa02001", -- 2117
    X"89900a099802", -- 2118
    X"009a13da1000", -- 2119
    X"124000060008", -- 2120
    X"146000135000", -- 2121
    X"188001157000", -- 2122
    X"00491789f0fa", -- 2123
    X"d98000000023", -- 2124
    X"a02001003913", -- 2125
    X"09980289f0ea", -- 2126
    X"da080089900a", -- 2127
    X"800061009a13", -- 2128
    X"80f01a80f1cb", -- 2129
    X"82f03a81f02a", -- 2130
    X"84f05a83f04a", -- 2131
    X"86f07a85f06a", -- 2132
    X"88f09a87f08a", -- 2133
    X"8af0ba89f0aa", -- 2134
    X"00e01a1ff00f", -- 2135
    X"80f01b3ff024", -- 2136
    X"80f23b80f12b", -- 2137
    X"80f45b80f34b", -- 2138
    X"80f67b80f56b", -- 2139
    X"80f89b80f78b", -- 2140
    X"80fabb80f9ab", -- 2141
    X"80fcdb80fbcb", -- 2142
    X"80fefb80fdeb", -- 2143
    X"dd0001dc0000", -- 2144
    X"81f10bd10800", -- 2145
    X"c10c9981f16b", -- 2146
    X"c0005bc10f9a", -- 2147
    X"000021d40000", -- 2148
    X"00040280f22a", -- 2149
    X"d1400080001a", -- 2150
    X"82f22a00010b", -- 2151
    X"8220aa022406", -- 2152
    X"000023d34000", -- 2153
    X"020020002313", -- 2154
    X"dc0001c02020", -- 2155
    X"12f010000021", -- 2156
    X"83200a022402", -- 2157
    X"80231b031306", -- 2158
    X"c02020020020", -- 2159
    X"000021dc0001", -- 2160
    X"00040280f22a", -- 2161
    X"d1400080001a", -- 2162
    X"82f22a00010b", -- 2163
    X"8220aa022406", -- 2164
    X"000023d34000", -- 2165
    X"020020002314", -- 2166
    X"dc0001c02020", -- 2167
    X"12f016000021", -- 2168
    X"83200a022402", -- 2169
    X"80231b031302", -- 2170
    X"c02020020020", -- 2171
    X"144001dc0001", -- 2172
    X"dd0000c0c2b0", -- 2173
    X"81f10bd10400", -- 2174
    X"c1103981f16b", -- 2175
    X"c0005bc1124a", -- 2176
    X"000021d40000", -- 2177
    X"00040280f22a", -- 2178
    X"d1200080001a", -- 2179
    X"82f22a00010b", -- 2180
    X"8220aa022406", -- 2181
    X"000023d32000", -- 2182
    X"12f010002313", -- 2183
    X"83200a022402", -- 2184
    X"80231b031306", -- 2185
    X"00040280f22a", -- 2186
    X"d1200080001a", -- 2187
    X"82f22a00010b", -- 2188
    X"8220aa022406", -- 2189
    X"000023d32000", -- 2190
    X"12f016002314", -- 2191
    X"83200a022402", -- 2192
    X"80231b031302", -- 2193
    X"d00000144001", -- 2194
    X"12f010d10000", -- 2195
    X"83300ad316b7", -- 2196
    X"8ff2fb80f30b", -- 2197
    X"be10368ffdeb", -- 2198
    X"d5000084ffda", -- 2199
    X"8407e8d7000a", -- 2200
    X"8457c8d70033", -- 2201
    X"163000155001", -- 2202
    X"d316b7174000", -- 2203
    X"83300a033502", -- 2204
    X"8ff2fb80f30b", -- 2205
    X"be10368ffdeb", -- 2206
    X"08470b84ffda", -- 2207
    X"c11449c083e3", -- 2208
    X"c0002bc1153a", -- 2209
    X"8b60128a3012", -- 2210
    X"80fc0b0cab02", -- 2211
    X"8ffdeb8ff2fb", -- 2212
    X"8affdabe1036", -- 2213
    X"c08043084a0b", -- 2214
    X"16c00017a000", -- 2215
    X"14a000c11538", -- 2216
    X"00002413c000", -- 2217
    X"077406066306", -- 2218
    X"807839d80000", -- 2219
    X"c116d8183000", -- 2220
    X"077000197000", -- 2221
    X"077c0d0c7011", -- 2222
    X"80f80bd83fff", -- 2223
    X"be00cf8ff7fb", -- 2224
    X"0a670b87ffea", -- 2225
    X"088c06d80014", -- 2226
    X"17a0000aa810", -- 2227
    X"077004c09026", -- 2228
    X"8aa0b30a470b", -- 2229
    X"87f23a083a06", -- 2230
    X"80780b077002", -- 2231
    X"100001138000", -- 2232
    X"801749d70000", -- 2233
    X"12f016d10001", -- 2234
    X"d10000c11798", -- 2235
    X"80f30b12f010", -- 2236
    X"8ffdeb8ff2fb", -- 2237
    X"84ffdabe1036", -- 2238
    X"37000ac11308", -- 2239
    X"c11869c070a6", -- 2240
    X"c000abc1189a", -- 2241
    X"81f23a80f24a", -- 2242
    X"10000182000a", -- 2243
    X"11100180120b", -- 2244
    X"81f02a80f01a", -- 2245
    X"83f04a82f03a", -- 2246
    X"85f06a84f05a", -- 2247
    X"87f08a86f07a", -- 2248
    X"89f0aa88f09a", -- 2249
    X"8bf0ca8af0ba", -- 2250
    X"8df0ea8cf0da", -- 2251
    X"1ff0248ef0fa", -- 2252
    X"3ff00b00e01a", -- 2253
    X"80f12b80f01b", -- 2254
    X"80f34b80f23b", -- 2255
    X"80f56b80f45b", -- 2256
    X"80f78b80f67b", -- 2257
    X"d0003f80f89b", -- 2258
    X"c11c6ac11b19", -- 2259
    X"d10d85c000ab", -- 2260
    X"82f0ba11103f", -- 2261
    X"32200112200a", -- 2262
    X"13300a83f0aa", -- 2263
    X"85200a333001", -- 2264
    X"04450684100a", -- 2265
    X"300001c04056", -- 2266
    X"c00020311001", -- 2267
    X"84100ac11b28", -- 2268
    X"d60e05045406", -- 2269
    X"86600a066002", -- 2270
    X"8660c306640b", -- 2271
    X"056402840090", -- 2272
    X"05540ad46488", -- 2273
    X"32200180350b", -- 2274
    X"80f01a333001", -- 2275
    X"82f03a81f02a", -- 2276
    X"84f05a83f04a", -- 2277
    X"86f07a85f06a", -- 2278
    X"88f09a87f08a", -- 2279
    X"00e01a1ff00b", -- 2280
    X"80f01b3ff016", -- 2281
    X"80f23b80f12b", -- 2282
    X"80f45b80f34b", -- 2283
    X"80f67b80f56b", -- 2284
    X"80f89b80f78b", -- 2285
    X"80f16a80f9ab", -- 2286
    X"d1040580001a", -- 2287
    X"011202d22000", -- 2288
    X"80f0bb000106", -- 2289
    X"c11f4ac11ee9", -- 2290
    X"300002d0000a", -- 2291
    X"d0000100001e", -- 2292
    X"14400114f00b", -- 2293
    X"d6200085f16a", -- 2294
    X"83500a82502a", -- 2295
    X"012306155001", -- 2296
    X"80410b011606", -- 2297
    X"d15c7d144001", -- 2298
    X"83500a011606", -- 2299
    X"011306155001", -- 2300
    X"c1202980410b", -- 2301
    X"c000abc120fa", -- 2302
    X"85f15a14f00b", -- 2303
    X"d70800d65000", -- 2304
    X"14400180400a", -- 2305
    X"80570bc00040", -- 2306
    X"c120f8155001", -- 2307
    X"82202102000b", -- 2308
    X"82202102360b", -- 2309
    X"80510b013702", -- 2310
    X"000024155001", -- 2311
    X"80504a85f15a", -- 2312
    X"02060bd64ccd", -- 2313
    X"80534b822011", -- 2314
    X"02060b80505a", -- 2315
    X"80535b822011", -- 2316
    X"c121f9d00000", -- 2317
    X"c000abc1224a", -- 2318
    X"81500a85f15a", -- 2319
    X"021006155001", -- 2320
    X"101000c02020", -- 2321
    X"000011000024", -- 2322
    X"c122dac122a9", -- 2323
    X"85f15ac000ab", -- 2324
    X"01100d81500a", -- 2325
    X"15500180510b", -- 2326
    X"81f02a80f01a", -- 2327
    X"83f04a82f03a", -- 2328
    X"85f06a84f05a", -- 2329
    X"87f08a86f07a", -- 2330
    X"89f0aa88f09a", -- 2331
    X"00e01a1ff016", -- 2332
    X"80f02b3ff017", -- 2333
    X"80f24b80f13b", -- 2334
    X"80f46b80f35b", -- 2335
    X"80f68b80f57b", -- 2336
    X"80f8ab80f79b", -- 2337
    X"80f00b80f17a", -- 2338
    X"8ff0fb10f00b", -- 2339
    X"be11d280fe1b", -- 2340
    X"80f00b80f17a", -- 2341
    X"8ff0fb10f00b", -- 2342
    X"8ff0eb80f16a", -- 2343
    X"8ff0db80f15a", -- 2344
    X"8ef01abe00fd", -- 2345
    X"81f03a80f02a", -- 2346
    X"83f05a82f04a", -- 2347
    X"85f07a84f06a", -- 2348
    X"87f09a86f08a", -- 2349
    X"1ff01788f0aa", -- 2350
    X"3ff01a00e01a", -- 2351
    X"80f12b80f01b", -- 2352
    X"80f1aa80fe3b", -- 2353
    X"10f00e80f00b", -- 2354
    X"be119b8ff0fb", -- 2355
    X"80f00b10f00e", -- 2356
    X"8ff0fb10f004", -- 2357
    X"8ff0ebd00690", -- 2358
    X"10f004be123a", -- 2359
    X"80f19a80f00b", -- 2360
    X"be05948ff0fb", -- 2361
    X"100002d00690", -- 2362
    X"80100b81f18a", -- 2363
    X"81f02a80f01a", -- 2364
    X"1ff01a8ef03a", -- 2365
    X"3ff0f300e01a", -- 2366
    X"80f02b80fe1b", -- 2367
    X"80f24b80f13b", -- 2368
    X"80f46b80f35b", -- 2369
    X"80f68b80f57b", -- 2370
    X"80f8ab80f79b", -- 2371
    X"80facb80f9bb", -- 2372
    X"d00000000021", -- 2373
    X"000023d10000", -- 2374
    X"82200a12f0f3", -- 2375
    X"d0008f32208f", -- 2376
    X"800012100050", -- 2377
    X"c12989100001", -- 2378
    X"00001ec129aa", -- 2379
    X"12200283200a", -- 2380
    X"020020003313", -- 2381
    X"c12a69c02100", -- 2382
    X"d3008fc12aaa", -- 2383
    X"00301e133050", -- 2384
    X"82200a12f0f3", -- 2385
    X"13f00e32208f", -- 2386
    X"12200184200a", -- 2387
    X"80340b844032", -- 2388
    X"c12cc8133001", -- 2389
    X"d70010d60000", -- 2390
    X"c06107060607", -- 2391
    X"c12bdac12b99", -- 2392
    X"133050d3008f", -- 2393
    X"12f0f300301e", -- 2394
    X"32208f82200a", -- 2395
    X"84200a13f00e", -- 2396
    X"844030122001", -- 2397
    X"13300180340b", -- 2398
    X"c12c89c12cc8", -- 2399
    X"d3008fc12cba", -- 2400
    X"00301e133050", -- 2401
    X"82200a12f0f3", -- 2402
    X"13f00e32208f", -- 2403
    X"12200184200a", -- 2404
    X"13300180340b", -- 2405
    X"d78000d60000", -- 2406
    X"da0028d00014", -- 2407
    X"13308f13f00e", -- 2408
    X"12208f12f00e", -- 2409
    X"d40000022006", -- 2410
    X"004023d50000", -- 2411
    X"c12dfac12db9", -- 2412
    X"84300ac0028b", -- 2413
    X"13300285200a", -- 2414
    X"044513122002", -- 2415
    X"c08041084607", -- 2416
    X"11f0f2264000", -- 2417
    X"10000180100b", -- 2418
    X"d400018e0aa9", -- 2419
    X"004023d50000", -- 2420
    X"81100a11f0f2", -- 2421
    X"12208f12f00e", -- 2422
    X"c12f29022106", -- 2423
    X"c0028bc12f4a", -- 2424
    X"04441384200a", -- 2425
    X"80f50b122002", -- 2426
    X"be06a48ff4fb", -- 2427
    X"84ffda85ffea", -- 2428
    X"044008066008", -- 2429
    X"8ff6fb80f70b", -- 2430
    X"8ff4db8ff5eb", -- 2431
    X"85ffcabe0d3d", -- 2432
    X"1bf0f184ffba", -- 2433
    X"d6000080b40b", -- 2434
    X"d00028d78000", -- 2435
    X"d40000da0050", -- 2436
    X"004023d50000", -- 2437
    X"12208f12f00e", -- 2438
    X"13308f13f00e", -- 2439
    X"c13149033006", -- 2440
    X"c0014bc131ba", -- 2441
    X"85300a84200a", -- 2442
    X"89302a88202a", -- 2443
    X"133004122004", -- 2444
    X"048913044513", -- 2445
    X"084607000024", -- 2446
    X"264000c08041", -- 2447
    X"80100b11f0f0", -- 2448
    X"8e0a69100001", -- 2449
    X"d40001266000", -- 2450
    X"004023d50000", -- 2451
    X"81100a11f0f0", -- 2452
    X"12208f12f00e", -- 2453
    X"c13309022106", -- 2454
    X"c0028bc1332a", -- 2455
    X"12200284200a", -- 2456
    X"80f50b044413", -- 2457
    X"be06a48ff4fb", -- 2458
    X"84ffda85ffea", -- 2459
    X"044008066008", -- 2460
    X"8ff6fb80f70b", -- 2461
    X"8ff4db8ff5eb", -- 2462
    X"85ffcabe0d3d", -- 2463
    X"1bf0ef84ffba", -- 2464
    X"d6000080b40b", -- 2465
    X"d00050d78000", -- 2466
    X"d40000da0090", -- 2467
    X"004023d50000", -- 2468
    X"12208f12f00e", -- 2469
    X"13308f13f00e", -- 2470
    X"c13529033006", -- 2471
    X"c0014bc1359a", -- 2472
    X"85300a84200a", -- 2473
    X"89302a88202a", -- 2474
    X"133004122004", -- 2475
    X"048913044513", -- 2476
    X"084607000024", -- 2477
    X"264000c08041", -- 2478
    X"80100b11f0ee", -- 2479
    X"8e0a69100002", -- 2480
    X"80000a10f0ee", -- 2481
    X"d50000d40000", -- 2482
    X"12f00e004023", -- 2483
    X"13f00e12208f", -- 2484
    X"03300613308f", -- 2485
    X"c13709333001", -- 2486
    X"c0028bc1374a", -- 2487
    X"85300a84200a", -- 2488
    X"122002044513", -- 2489
    X"084607133002", -- 2490
    X"264000c08051", -- 2491
    X"14000111f0ee", -- 2492
    X"d4000080140b", -- 2493
    X"004023d50000", -- 2494
    X"12208f12f00e", -- 2495
    X"13308f13f00e", -- 2496
    X"133001033006", -- 2497
    X"c138bac13879", -- 2498
    X"84200ac0028b", -- 2499
    X"04451385300a", -- 2500
    X"133002122002", -- 2501
    X"c08051084607", -- 2502
    X"11f0ee264000", -- 2503
    X"80140b340001", -- 2504
    X"d50000d40001", -- 2505
    X"11f0ee004023", -- 2506
    X"12f00e81100a", -- 2507
    X"02210612208f", -- 2508
    X"c139fac139d9", -- 2509
    X"84200ac0028b", -- 2510
    X"122002044413", -- 2511
    X"8ff4fb80f50b", -- 2512
    X"85ffeabe06a4", -- 2513
    X"06600884ffda", -- 2514
    X"80f70b044008", -- 2515
    X"8ff5eb8ff6fb", -- 2516
    X"be0d3d8ff4db", -- 2517
    X"84ffba85ffca", -- 2518
    X"80b40b1bf0eb", -- 2519
    X"80b00a1bf0f0", -- 2520
    X"1bf0ee800010", -- 2521
    X"02010681b00a", -- 2522
    X"333005032000", -- 2523
    X"1bf0efc03096", -- 2524
    X"1bf0eb83b00a", -- 2525
    X"84402284b00a", -- 2526
    X"1bf0ef033402", -- 2527
    X"1bf0f080b30b", -- 2528
    X"02200280b00a", -- 2529
    X"333007032000", -- 2530
    X"1bf0efc03096", -- 2531
    X"1bf0eb83b00a", -- 2532
    X"84402284b00a", -- 2533
    X"1bf0ef033402", -- 2534
    X"1bf0f280b30b", -- 2535
    X"80001080b00a", -- 2536
    X"81b00a1bf0f0", -- 2537
    X"032000020106", -- 2538
    X"c030a6333005", -- 2539
    X"83b00a1bf0f1", -- 2540
    X"84b00a1bf0ef", -- 2541
    X"044b0adb199a", -- 2542
    X"1bf0f1033402", -- 2543
    X"1bf0f280b30b", -- 2544
    X"02200280b00a", -- 2545
    X"333007032000", -- 2546
    X"1bf0f1c030a6", -- 2547
    X"1bf0ef83b00a", -- 2548
    X"db199a84b00a", -- 2549
    X"033402044b0a", -- 2550
    X"80b30b1bf0f1", -- 2551
    X"80b00a1bf0f1", -- 2552
    X"81b00a1bf0ef", -- 2553
    X"c02076020106", -- 2554
    X"80b10b1bf0f1", -- 2555
    X"82b00a1bf0f0", -- 2556
    X"80b20b1bf0f2", -- 2557
    X"81b00a1bf0eb", -- 2558
    X"80b00a1bf0f1", -- 2559
    X"c02056020106", -- 2560
    X"82b00a1bf0ee", -- 2561
    X"80b20b1bf0f2", -- 2562
    X"80f02a8ef01a", -- 2563
    X"82f04a81f03a", -- 2564
    X"84f06a83f05a", -- 2565
    X"86f08a85f07a", -- 2566
    X"88f0aa87f09a", -- 2567
    X"8af0ca89f0ba", -- 2568
    X"00e01a1ff0f3", -- 2569
    X"d106b1d0069b", -- 2570
    X"d40000d307c5", -- 2571
    X"00001d80340b", -- 2572
    X"10000110000a", -- 2573
    X"11100111100a", -- 2574
    X"82300ad307c5", -- 2575
    X"80320b122028", -- 2576
    X"d306c700001d", -- 2577
    X"80340bd41000", -- 2578
    X"d40028133001", -- 2579
    X"c142d9344001", -- 2580
    X"00401ec142ea", -- 2581
    X"80340bd40000", -- 2582
    X"80f10b133001", -- 2583
    X"8ff3fbd306c7", -- 2584
    X"d300288ff3eb", -- 2585
    X"d306c78ff3db", -- 2586
    X"8ff3cb133001", -- 2587
    X"8ff3bbd30000", -- 2588
    X"d306c7be0075", -- 2589
    X"d307ce80f30b", -- 2590
    X"d300288ff3fb", -- 2591
    X"be00008ff3eb", -- 2592
    X"d207c580f10b", -- 2593
    X"d3026982200a", -- 2594
    X"8ff3fb033202", -- 2595
    X"8ff3ebd306ef", -- 2596
    X"8ff3dbd30028", -- 2597
    X"8ff3cbd302cd", -- 2598
    X"8ff3bbd30000", -- 2599
    X"d306efbe0075", -- 2600
    X"d307ce80f30b", -- 2601
    X"8ff3fb133028", -- 2602
    X"8ff3ebd30028", -- 2603
    X"d207c5be0000", -- 2604
    X"d3026982200a", -- 2605
    X"80f30b033202", -- 2606
    X"8ff3fbd306ef", -- 2607
    X"8ff3ebd306c7", -- 2608
    X"83300ad307c3", -- 2609
    X"d307c48ff3db", -- 2610
    X"8ff3cb83300a", -- 2611
    X"82200ad207c5", -- 2612
    X"be15928ff2bb", -- 2613
    X"d2068e83ff9a", -- 2614
    X"84ffaa80230b", -- 2615
    X"80240bd2068f", -- 2616
    X"8ff4fb80f30b", -- 2617
    X"8ff3ebd307c3", -- 2618
    X"8ff3dbd307c4", -- 2619
    X"82200ad207c5", -- 2620
    X"be16918ff2cb", -- 2621
    X"d307c684ffba", -- 2622
    X"80240b82300a", -- 2623
    X"80320b122001", -- 2624
    X"d207c5d30269", -- 2625
    X"03320282200a", -- 2626
    X"c148aac14899", -- 2627
    X"82300ac0028b", -- 2628
    X"d20000133001", -- 2629
    X"83300ad307c5", -- 2630
    X"80f40b803299", -- 2631
    X"84fffabe16c3", -- 2632
    X"82300ad307c6", -- 2633
    X"12200180240b", -- 2634
    X"d3026980320b", -- 2635
    X"82200ad207c5", -- 2636
    X"c149e9033202", -- 2637
    X"c0028bc149fa", -- 2638
    X"13300182300a", -- 2639
    X"d3026980f10b", -- 2640
    X"82200ad207c5", -- 2641
    X"8ff3fb033202", -- 2642
    X"8ff3ebd3073f", -- 2643
    X"8ff3dbd30028", -- 2644
    X"8ff3cbd302e1", -- 2645
    X"8ff3bbd30000", -- 2646
    X"d306efbe0075", -- 2647
    X"d3073f80f30b", -- 2648
    X"d307c78ff3fb", -- 2649
    X"be16de8ff3eb", -- 2650
    X"d307cb84ffda", -- 2651
    X"d3068e80340b", -- 2652
    X"80f30b83300a", -- 2653
    X"83300ad3068f", -- 2654
    X"be17608ff3fb", -- 2655
    X"d307cd85ffea", -- 2656
    X"d2000180350b", -- 2657
    X"d53ccc805279", -- 2658
    X"c05040054506", -- 2659
    X"d307cbd43ccc", -- 2660
    X"d2073f80340b", -- 2661
    X"133050d307ce", -- 2662
    X"d306ef80342b", -- 2663
    X"c14d49d50717", -- 2664
    X"c0028bc14dca", -- 2665
    X"12200186200a", -- 2666
    X"13300187300a", -- 2667
    X"88801108640b", -- 2668
    X"80590b097906", -- 2669
    X"d30717155001", -- 2670
    X"d306c780f30b", -- 2671
    X"d3068e8ff3fb", -- 2672
    X"8ff3eb83300a", -- 2673
    X"83300ad302eb", -- 2674
    X"d3065c8ff3db", -- 2675
    X"d307678ff3cb", -- 2676
    X"be17a48ff3bb", -- 2677
    X"85ffaa84ff9a", -- 2678
    X"82300ad307c6", -- 2679
    X"12200180240b", -- 2680
    X"d307c680320b", -- 2681
    X"80250b82300a", -- 2682
    X"80320b122001", -- 2683
    X"84200ad207c7", -- 2684
    X"80340bd3078f", -- 2685
    X"04400484201a", -- 2686
    X"80340bd30794", -- 2687
    X"04400484202a", -- 2688
    X"80341bd3078f", -- 2689
    X"14400184203a", -- 2690
    X"d30794044004", -- 2691
    X"d306ef80341b", -- 2692
    X"d3073f80f30b", -- 2693
    X"d307678ff3fb", -- 2694
    X"d3078f8ff3eb", -- 2695
    X"d307948ff3db", -- 2696
    X"be1d878ff3cb", -- 2697
    X"80f30bd3065c", -- 2698
    X"8ff3fbd3078f", -- 2699
    X"8ff3ebd30794", -- 2700
    X"83300ad307cd", -- 2701
    X"be1ee18ff3bb", -- 2702
    X"d207cb83ffda", -- 2703
    X"83ffca80230b", -- 2704
    X"80230bd207cc", -- 2705
    X"d307c684ffaa", -- 2706
    X"80240b82300a", -- 2707
    X"80320b122001", -- 2708
    X"82200ad207cb", -- 2709
    X"d432d9d302eb", -- 2710
    X"c04030042406", -- 2711
    X"c15368d232d9", -- 2712
    X"042406d40ccd", -- 2713
    X"d20ccdc04026", -- 2714
    X"c1545980320b", -- 2715
    X"c0028bc154ea", -- 2716
    X"d307c5d20269", -- 2717
    X"02230283300a", -- 2718
    X"83300ad307cb", -- 2719
    X"84400ad407cc", -- 2720
    X"d50000d7065c", -- 2721
    X"88600a062502", -- 2722
    X"00802308830b", -- 2723
    X"17700188700a", -- 2724
    X"888011088413", -- 2725
    X"80680b088009", -- 2726
    X"d207cb166001", -- 2727
    X"80f20b82200a", -- 2728
    X"82200ad2068e", -- 2729
    X"be1e828ff2fb", -- 2730
    X"c1575ac15679", -- 2731
    X"d207cbc000ab", -- 2732
    X"d307cc82200a", -- 2733
    X"d4073f83300a", -- 2734
    X"34400a144028", -- 2735
    X"155028d50767", -- 2736
    X"d606ef35500a", -- 2737
    X"36600a166028", -- 2738
    X"87400adb02cd", -- 2739
    X"08720b144001", -- 2740
    X"1a9000888011", -- 2741
    X"15500187500a", -- 2742
    X"88802108730b", -- 2743
    X"87600a08a902", -- 2744
    X"087806166001", -- 2745
    X"1bb00180b80b", -- 2746
    X"d1000000001d", -- 2747
    X"80f10b111050", -- 2748
    X"8ff1fbd10000", -- 2749
    X"311050d100f0", -- 2750
    X"be00008ff1eb", -- 2751
    X"111050d100f0", -- 2752
    X"d100f080f10b", -- 2753
    X"d1008f8ff1fb", -- 2754
    X"be00008ff1eb", -- 2755
    X"111050d101cf", -- 2756
    X"d101cf80f10b", -- 2757
    X"d1008f8ff1fb", -- 2758
    X"8ff1eb11100b", -- 2759
    X"00001dbe0000", -- 2760
    X"80f01b3ff063", -- 2761
    X"80f23b80f12b", -- 2762
    X"80f45b80f34b", -- 2763
    X"80f67b80f56b", -- 2764
    X"80f89b80f78b", -- 2765
    X"80febb80f9ab", -- 2766
    X"80f00b80f61a", -- 2767
    X"8ff0fb80f62a", -- 2768
    X"8ff0eb10f00c", -- 2769
    X"d00000be161e", -- 2770
    X"82f60ad18000", -- 2771
    X"13300183f5fa", -- 2772
    X"80f40b14f00c", -- 2773
    X"04420684f63a", -- 2774
    X"be16778ff4fb", -- 2775
    X"84ffda85ffea", -- 2776
    X"c06041064007", -- 2777
    X"115000104000", -- 2778
    X"122001182000", -- 2779
    X"80f63a8f2329", -- 2780
    X"8ff8fb80f00b", -- 2781
    X"8ff0ebd00000", -- 2782
    X"10f00cbe0552", -- 2783
    X"80f63a80f00b", -- 2784
    X"be16778ff0fb", -- 2785
    X"84ffda85ffea", -- 2786
    X"85f0dbd00000", -- 2787
    X"d1000080f5ea", -- 2788
    X"318054800149", -- 2789
    X"c16108c01020", -- 2790
    X"11f03480f63a", -- 2791
    X"c15d6ac15d39", -- 2792
    X"82000ac0028b", -- 2793
    X"80120b100001", -- 2794
    X"80f63a111001", -- 2795
    X"8ff8fb80f00b", -- 2796
    X"8ff0ebd0ffff", -- 2797
    X"10f00cbe0552", -- 2798
    X"80f63a80f00b", -- 2799
    X"be16778ff0fb", -- 2800
    X"86ffda87ffea", -- 2801
    X"c000e1006407", -- 2802
    X"157000146000", -- 2803
    X"85f0dbd0ffff", -- 2804
    X"11f03480f63a", -- 2805
    X"c15f2ac15ef9", -- 2806
    X"82000ac0028b", -- 2807
    X"80120b100001", -- 2808
    X"80f63a111001", -- 2809
    X"8ff8fb80f00b", -- 2810
    X"8ff0ebd00001", -- 2811
    X"10f00cbe0552", -- 2812
    X"80f63a80f00b", -- 2813
    X"be16778ff0fb", -- 2814
    X"86ffda87ffea", -- 2815
    X"c00061006407", -- 2816
    X"157000146000", -- 2817
    X"85f0dbd00001", -- 2818
    X"10f034c16108", -- 2819
    X"c160c981f63a", -- 2820
    X"c0028bc160fa", -- 2821
    X"10000182000a", -- 2822
    X"11100180120b", -- 2823
    X"80f01a85f8cb", -- 2824
    X"82f03a81f02a", -- 2825
    X"84f05a83f04a", -- 2826
    X"86f07a85f06a", -- 2827
    X"88f09a87f08a", -- 2828
    X"8ef0ba89f0aa", -- 2829
    X"00e01a1ff063", -- 2830
    X"80f01b3ff05e", -- 2831
    X"80f23b80f12b", -- 2832
    X"80f45b80f34b", -- 2833
    X"80f67b80f56b", -- 2834
    X"80f89b80f78b", -- 2835
    X"80fabb80f9ab", -- 2836
    X"d10000d00000", -- 2837
    X"d50028d40000", -- 2838
    X"c1644918f00c", -- 2839
    X"82f5eac164ba", -- 2840
    X"03340283f5da", -- 2841
    X"d70000d60000", -- 2842
    X"d90028006023", -- 2843
    X"da0001099406", -- 2844
    X"c0a0600a9a18", -- 2845
    X"87300a86200a", -- 2846
    X"133001122001", -- 2847
    X"899012066713", -- 2848
    X"00901ec090b0", -- 2849
    X"87300a86200a", -- 2850
    X"8a301a89201a", -- 2851
    X"133002122002", -- 2852
    X"069a13066713", -- 2853
    X"80860b000024", -- 2854
    X"80870b188001", -- 2855
    X"066001188001", -- 2856
    X"c02031026007", -- 2857
    X"117000106000", -- 2858
    X"8d45a9144001", -- 2859
    X"332010020012", -- 2860
    X"d20010c03020", -- 2861
    X"023206d30012", -- 2862
    X"81f5ca10f00c", -- 2863
    X"c1669ac16639", -- 2864
    X"84000ac0028b", -- 2865
    X"85000a100001", -- 2866
    X"044210100001", -- 2867
    X"11100180140b", -- 2868
    X"81f02a80f01a", -- 2869
    X"83f04a82f03a", -- 2870
    X"85f06a84f05a", -- 2871
    X"87f08a86f07a", -- 2872
    X"89f0aa88f09a", -- 2873
    X"1ff05e8af0ba", -- 2874
    X"3ff00800e01a", -- 2875
    X"80f12b80f01b", -- 2876
    X"80f34b80f23b", -- 2877
    X"d10000d00000", -- 2878
    X"80f08a000023", -- 2879
    X"c1684981f07a", -- 2880
    X"c0028bc1688a", -- 2881
    X"83100a82000a", -- 2882
    X"111001100001", -- 2883
    X"80f25b022313", -- 2884
    X"80f01a80f36b", -- 2885
    X"82f03a81f02a", -- 2886
    X"1ff00883f04a", -- 2887
    X"3ff01100e01a", -- 2888
    X"80f12b80f01b", -- 2889
    X"80f34b80f23b", -- 2890
    X"80f0dad10000", -- 2891
    X"80f11a8001a8", -- 2892
    X"81100a81f0fa", -- 2893
    X"81f10a020106", -- 2894
    X"122002722003", -- 2895
    X"c16bc8022102", -- 2896
    X"31005580f11a", -- 2897
    X"120070c01030", -- 2898
    X"81f10ac16ab8", -- 2899
    X"32203a720003", -- 2900
    X"330005022102", -- 2901
    X"80130b81f0fa", -- 2902
    X"c01026313014", -- 2903
    X"81f0fad30014", -- 2904
    X"13300980130b", -- 2905
    X"c0105031308f", -- 2906
    X"303009d3008f", -- 2907
    X"80100b81f0fa", -- 2908
    X"80130b81f0ea", -- 2909
    X"80f01a80f2cb", -- 2910
    X"82f03a81f02a", -- 2911
    X"1ff01183f04a", -- 2912
    X"3ff00d00e01a", -- 2913
    X"80f12b80f01b", -- 2914
    X"80f34b80f23b", -- 2915
    X"80f0da80f45b", -- 2916
    X"d10001800012", -- 2917
    X"d30006d20000", -- 2918
    X"d40001800012", -- 2919
    X"011402040418", -- 2920
    X"8f23b9122001", -- 2921
    X"011218d20001", -- 2922
    X"80f01a80f1cb", -- 2923
    X"82f03a81f02a", -- 2924
    X"84f05a83f04a", -- 2925
    X"00e01a1ff00d", -- 2926
    X"80f01b3ff037", -- 2927
    X"80f23b80f12b", -- 2928
    X"80f45b80f34b", -- 2929
    X"80f67b80f56b", -- 2930
    X"80febb80f78b", -- 2931
    X"c16f1ac16ed9", -- 2932
    X"80f36ac0028b", -- 2933
    X"82000a11f00c", -- 2934
    X"822022100001", -- 2935
    X"11100180120b", -- 2936
    X"d40001000021", -- 2937
    X"004023d50000", -- 2938
    X"c16fcac16fa9", -- 2939
    X"80f36ac0028b", -- 2940
    X"10000182000a", -- 2941
    X"000020042213", -- 2942
    X"034012c00052", -- 2943
    X"02400904430e", -- 2944
    X"d40001c17118", -- 2945
    X"004023d50000", -- 2946
    X"c170cac170a9", -- 2947
    X"10f00cc0028b", -- 2948
    X"10000182000a", -- 2949
    X"034012042213", -- 2950
    X"02400904430e", -- 2951
    X"80f35a333004", -- 2952
    X"17300080020b", -- 2953
    X"03300433300f", -- 2954
    X"00002180031b", -- 2955
    X"d50000d40000", -- 2956
    X"c17209004023", -- 2957
    X"c0028bc1724a", -- 2958
    X"81f36a80f37a", -- 2959
    X"10000182000a", -- 2960
    X"11100183100a", -- 2961
    X"000020042313", -- 2962
    X"034012c00052", -- 2963
    X"02400904430e", -- 2964
    X"d40000c173c8", -- 2965
    X"004023d50000", -- 2966
    X"c1737ac17339", -- 2967
    X"80f37ac0028b", -- 2968
    X"82000a11f00c", -- 2969
    X"83100a100001", -- 2970
    X"042313111001", -- 2971
    X"04430e034012", -- 2972
    X"333002024009", -- 2973
    X"80022b80f35a", -- 2974
    X"33300f153000", -- 2975
    X"80033b033004", -- 2976
    X"d3fff1c02052", -- 2977
    X"d6000080033b", -- 2978
    X"822012c17548", -- 2979
    X"81f35a80f20b", -- 2980
    X"8ff1fb81100a", -- 2981
    X"82ffeabe00cf", -- 2982
    X"06230f035706", -- 2983
    X"036306d34ccd", -- 2984
    X"d64ccdc03020", -- 2985
    X"80f01a83f64b", -- 2986
    X"82f03a81f02a", -- 2987
    X"84f05a83f04a", -- 2988
    X"86f07a85f06a", -- 2989
    X"8ef0ba87f08a", -- 2990
    X"00e01a1ff037", -- 2991
    X"80f01b3ff00e", -- 2992
    X"80f23b80f12b", -- 2993
    X"80f45b80f34b", -- 2994
    X"80f67b80f56b", -- 2995
    X"80f89b80f78b", -- 2996
    X"80f0ea80f9ab", -- 2997
    X"c0103081f0da", -- 2998
    X"c17718120001", -- 2999
    X"d00028120000", -- 3000
    X"00200610000a", -- 3001
    X"d00000c00026", -- 3002
    X"033002d3161e", -- 3003
    X"d0000a81300a", -- 3004
    X"002002300002", -- 3005
    X"033002d3161e", -- 3006
    X"d4ffff82300a", -- 3007
    X"132000d5ffff", -- 3008
    X"133001032106", -- 3009
    X"c178c9c030e0", -- 3010
    X"00301ec1791a", -- 3011
    X"d00335d30000", -- 3012
    X"000202022202", -- 3013
    X"87001a86000a", -- 3014
    X"c08021086407", -- 3015
    X"300002246000", -- 3016
    X"d73a98d60000", -- 3017
    X"c08021084607", -- 3018
    X"80f3cbd30001", -- 3019
    X"81f02a80f01a", -- 3020
    X"83f04a82f03a", -- 3021
    X"85f06a84f05a", -- 3022
    X"87f08a86f07a", -- 3023
    X"89f0aa88f09a", -- 3024
    X"00e01a1ff00e", -- 3025
    X"80f01b3ff2a3", -- 3026
    X"80f23b80f12b", -- 3027
    X"80f45b80f34b", -- 3028
    X"80f67b80f56b", -- 3029
    X"80f89b80f78b", -- 3030
    X"80febb80f9ab", -- 3031
    X"00f002d002a0", -- 3032
    X"80001080000a", -- 3033
    X"01f102d102a1", -- 3034
    X"32102881100a", -- 3035
    X"d20028c02146", -- 3036
    X"c17c59022106", -- 3037
    X"00201ec17cba", -- 3038
    X"02f202d202a2", -- 3039
    X"02210282200a", -- 3040
    X"03f302d302a2", -- 3041
    X"84300a83300a", -- 3042
    X"04400a133001", -- 3043
    X"04450285200a", -- 3044
    X"12200180240b", -- 3045
    X"03f302d302a2", -- 3046
    X"80f30b83300a", -- 3047
    X"8ff3fb13f034", -- 3048
    X"d302a2be1819", -- 3049
    X"83300a03f302", -- 3050
    X"d302a380f30b", -- 3051
    X"83300a03f302", -- 3052
    X"13f00c8ff3fb", -- 3053
    X"be161e8ff3eb", -- 3054
    X"80f30b13f00c", -- 3055
    X"8ff3fb13f034", -- 3056
    X"03f302d302a2", -- 3057
    X"8ff3eb83300a", -- 3058
    X"03f302d3029f", -- 3059
    X"8ff3db83300a", -- 3060
    X"03f302d3029e", -- 3061
    X"8ff3cb83300a", -- 3062
    X"86ffbabe1a06", -- 3063
    X"03f302d3029d", -- 3064
    X"86ffaa80360b", -- 3065
    X"03f302d3029c", -- 3066
    X"32102880360b", -- 3067
    X"d20028c02146", -- 3068
    X"c18059022106", -- 3069
    X"00201ec180ba", -- 3070
    X"02f202d2029f", -- 3071
    X"02210282200a", -- 3072
    X"03f302d3029f", -- 3073
    X"84300a83300a", -- 3074
    X"04400a133001", -- 3075
    X"04450285200a", -- 3076
    X"12200180240b", -- 3077
    X"81f02a80f01a", -- 3078
    X"83f04a82f03a", -- 3079
    X"85f06a84f05a", -- 3080
    X"87f08a86f07a", -- 3081
    X"89f0aa88f09a", -- 3082
    X"1ff2a38ef0ba", -- 3083
    X"3ff04700e01a", -- 3084
    X"80f12b80f01b", -- 3085
    X"80f34b80f23b", -- 3086
    X"80f56b80f45b", -- 3087
    X"80f78b80f67b", -- 3088
    X"80f9ab80f89b", -- 3089
    X"80fbcb80fabb", -- 3090
    X"80fdeb80fcdb", -- 3091
    X"d0000080fefb", -- 3092
    X"000023d10000", -- 3093
    X"c1830982f47a", -- 3094
    X"c0028bc1832a", -- 3095
    X"12200183200a", -- 3096
    X"d27d00003313", -- 3097
    X"c020c0021206", -- 3098
    X"14f01082f47a", -- 3099
    X"c183fac183b9", -- 3100
    X"83200ac0028b", -- 3101
    X"833012122001", -- 3102
    X"14400180430b", -- 3103
    X"050012c184d8", -- 3104
    X"82f47a855012", -- 3105
    X"c1848914f010", -- 3106
    X"c0028bc184ca", -- 3107
    X"12200183200a", -- 3108
    X"80430b03350d", -- 3109
    X"10f038144001", -- 3110
    X"80020b82f46a", -- 3111
    X"80021b122008", -- 3112
    X"80022b122008", -- 3113
    X"80023b122008", -- 3114
    X"80024b122008", -- 3115
    X"80025b122008", -- 3116
    X"80026b122040", -- 3117
    X"80027b122040", -- 3118
    X"80028b122040", -- 3119
    X"80029b122040", -- 3120
    X"8002ab122040", -- 3121
    X"8002bb122040", -- 3122
    X"8002cb122040", -- 3123
    X"8002db122040", -- 3124
    X"80500a15f038", -- 3125
    X"300001100008", -- 3126
    X"11100881501a", -- 3127
    X"82502a311001", -- 3128
    X"322001122008", -- 3129
    X"13300883503a", -- 3130
    X"84504a333001", -- 3131
    X"344001144008", -- 3132
    X"d6000015f010", -- 3133
    X"006023d70000", -- 3134
    X"c1899ac18819", -- 3135
    X"88500ac0008b", -- 3136
    X"068813155001", -- 3137
    X"34400180470b", -- 3138
    X"15500188500a", -- 3139
    X"80370b068813", -- 3140
    X"88500a333001", -- 3141
    X"068813155001", -- 3142
    X"32200180270b", -- 3143
    X"15500188500a", -- 3144
    X"80170b068813", -- 3145
    X"88500a311001", -- 3146
    X"068813155001", -- 3147
    X"30000180070b", -- 3148
    X"344001d40040", -- 3149
    X"d80008354001", -- 3150
    X"19f010188001", -- 3151
    X"db00001a9001", -- 3152
    X"83c0ca1cf038", -- 3153
    X"82c09a033402", -- 3154
    X"81c05a022402", -- 3155
    X"80c08a011402", -- 3156
    X"d60000000502", -- 3157
    X"006023d70000", -- 3158
    X"1da0001c9000", -- 3159
    X"0eeb06de0008", -- 3160
    X"c0e2503ee001", -- 3161
    X"c18d7ac18b79", -- 3162
    X"86c00a00e01e", -- 3163
    X"87d00a1cc001", -- 3164
    X"0667131dd001", -- 3165
    X"1cc00186c00a", -- 3166
    X"1dd00187d00a", -- 3167
    X"80370b066713", -- 3168
    X"1cc00186c00a", -- 3169
    X"1dd00187d00a", -- 3170
    X"80270b066713", -- 3171
    X"1cc00186c00a", -- 3172
    X"1dd00187d00a", -- 3173
    X"80170b066713", -- 3174
    X"1cc00186c00a", -- 3175
    X"1dd00187d00a", -- 3176
    X"80070b066713", -- 3177
    X"022806033806", -- 3178
    X"000806011806", -- 3179
    X"1cc00186c00a", -- 3180
    X"1dd00187d00a", -- 3181
    X"86c00a066713", -- 3182
    X"87d00a1cc001", -- 3183
    X"0667131dd001", -- 3184
    X"86c00a80370b", -- 3185
    X"87d00a1cc001", -- 3186
    X"0667131dd001", -- 3187
    X"86c00a80270b", -- 3188
    X"87d00a1cc001", -- 3189
    X"0667131dd001", -- 3190
    X"34400880170b", -- 3191
    X"1aa005355001", -- 3192
    X"dc00081bb001", -- 3193
    X"19f0108abce9", -- 3194
    X"d800401a9002", -- 3195
    X"358001388001", -- 3196
    X"1cf038db0000", -- 3197
    X"04480284c0da", -- 3198
    X"03380283c0aa", -- 3199
    X"02280282c06a", -- 3200
    X"01150281c0ba", -- 3201
    X"00050280c07a", -- 3202
    X"d70000d60000", -- 3203
    X"1c9000006023", -- 3204
    X"de00081da000", -- 3205
    X"3ee0010eeb06", -- 3206
    X"c19129c0e2c0", -- 3207
    X"00e01ec1939a", -- 3208
    X"1cc00186c00a", -- 3209
    X"1dd00187d00a", -- 3210
    X"80470b066713", -- 3211
    X"1cc00186c00a", -- 3212
    X"1dd00187d00a", -- 3213
    X"80370b066713", -- 3214
    X"1cc00186c00a", -- 3215
    X"1dd00187d00a", -- 3216
    X"80270b066713", -- 3217
    X"1cc00186c00a", -- 3218
    X"1dd00187d00a", -- 3219
    X"80170b066713", -- 3220
    X"1cc00186c00a", -- 3221
    X"1dd00187d00a", -- 3222
    X"80070b066713", -- 3223
    X"344001344008", -- 3224
    X"333001333008", -- 3225
    X"322001322008", -- 3226
    X"311001311008", -- 3227
    X"300001300008", -- 3228
    X"1cc00186c00a", -- 3229
    X"1dd00187d00a", -- 3230
    X"80470b066713", -- 3231
    X"1cc00186c00a", -- 3232
    X"1dd00187d00a", -- 3233
    X"80370b066713", -- 3234
    X"1cc00186c00a", -- 3235
    X"1dd00187d00a", -- 3236
    X"80270b066713", -- 3237
    X"355001388008", -- 3238
    X"1bb0011aa005", -- 3239
    X"8abca9dc0008", -- 3240
    X"1a900319f010", -- 3241
    X"388001d80040", -- 3242
    X"db0000358001", -- 3243
    X"84c0ba1cf038", -- 3244
    X"83c07a044802", -- 3245
    X"82c0da033802", -- 3246
    X"81c0aa022502", -- 3247
    X"80c06a011502", -- 3248
    X"d60000000502", -- 3249
    X"006023d70000", -- 3250
    X"1da0001c9000", -- 3251
    X"0eeb06de0008", -- 3252
    X"c0e2c03ee001", -- 3253
    X"c1996ac196f9", -- 3254
    X"86c00a00e01e", -- 3255
    X"87d00a1cc001", -- 3256
    X"0667131dd001", -- 3257
    X"86c00a80470b", -- 3258
    X"87d00a1cc001", -- 3259
    X"0667131dd001", -- 3260
    X"86c00a80370b", -- 3261
    X"87d00a1cc001", -- 3262
    X"0667131dd001", -- 3263
    X"86c00a80270b", -- 3264
    X"87d00a1cc001", -- 3265
    X"0667131dd001", -- 3266
    X"86c00a80170b", -- 3267
    X"87d00a1cc001", -- 3268
    X"0667131dd001", -- 3269
    X"34400880070b", -- 3270
    X"333008344001", -- 3271
    X"322008333001", -- 3272
    X"311008322001", -- 3273
    X"300008311001", -- 3274
    X"86c00a300001", -- 3275
    X"87d00a1cc001", -- 3276
    X"0667131dd001", -- 3277
    X"86c00a80470b", -- 3278
    X"87d00a1cc001", -- 3279
    X"0667131dd001", -- 3280
    X"38800880370b", -- 3281
    X"1aa005355001", -- 3282
    X"dc00081bb001", -- 3283
    X"19f0108bbc09", -- 3284
    X"d800401a9004", -- 3285
    X"358001388001", -- 3286
    X"1cf038db0000", -- 3287
    X"03380283c08a", -- 3288
    X"02250282c0ca", -- 3289
    X"01150281c09a", -- 3290
    X"00050280c05a", -- 3291
    X"d70000d60000", -- 3292
    X"1c9000006023", -- 3293
    X"de00081da000", -- 3294
    X"3ee0010eeb06", -- 3295
    X"c19c49c0e290", -- 3296
    X"00e01ec19e8a", -- 3297
    X"1cc00186c00a", -- 3298
    X"1dd00187d00a", -- 3299
    X"80370b066713", -- 3300
    X"1cc00186c00a", -- 3301
    X"1dd00187d00a", -- 3302
    X"86c00a066713", -- 3303
    X"87d00a1cc001", -- 3304
    X"0667131dd001", -- 3305
    X"86c00a80270b", -- 3306
    X"87d00a1cc001", -- 3307
    X"0667131dd001", -- 3308
    X"86c00a80170b", -- 3309
    X"87d00a1cc001", -- 3310
    X"0667131dd001", -- 3311
    X"33300880070b", -- 3312
    X"322008333001", -- 3313
    X"311008322001", -- 3314
    X"300008311001", -- 3315
    X"86c00a300001", -- 3316
    X"87d00a1cc001", -- 3317
    X"0667131dd001", -- 3318
    X"38800880370b", -- 3319
    X"1aa005355001", -- 3320
    X"dc00081bb001", -- 3321
    X"80f01a8bbcb9", -- 3322
    X"82f03a81f02a", -- 3323
    X"84f05a83f04a", -- 3324
    X"86f07a85f06a", -- 3325
    X"88f09a87f08a", -- 3326
    X"8af0ba89f0aa", -- 3327
    X"8cf0da8bf0ca", -- 3328
    X"8ef0fa8df0ea", -- 3329
    X"00e01a1ff047", -- 3330
    X"80f01b3ff09a", -- 3331
    X"80f23b80f12b", -- 3332
    X"80f45b80f34b", -- 3333
    X"80f67b80f56b", -- 3334
    X"80f89b80f78b", -- 3335
    X"80fabb80f9ab", -- 3336
    X"80fcdb80fbcb", -- 3337
    X"80fefb80fdeb", -- 3338
    X"12f09910f02e", -- 3339
    X"80020b82200a", -- 3340
    X"80021b122008", -- 3341
    X"80022b122008", -- 3342
    X"80023b122008", -- 3343
    X"80024b122008", -- 3344
    X"80025b122008", -- 3345
    X"80026b122040", -- 3346
    X"80027b122040", -- 3347
    X"80028b122040", -- 3348
    X"80029b122040", -- 3349
    X"8002ab122040", -- 3350
    X"8002bb122040", -- 3351
    X"8002cb122040", -- 3352
    X"8002db122040", -- 3353
    X"80000a10f09a", -- 3354
    X"12f04411f06c", -- 3355
    X"d58000d47fff", -- 3356
    X"c1a4aac1a3d9", -- 3357
    X"83000ac0028b", -- 3358
    X"80140bc03064", -- 3359
    X"80250b111001", -- 3360
    X"c1a4a8122001", -- 3361
    X"11100180150b", -- 3362
    X"12200180240b", -- 3363
    X"80030b033004", -- 3364
    X"14f02e100001", -- 3365
    X"81406a80405a", -- 3366
    X"83408a82407a", -- 3367
    X"d80028d40000", -- 3368
    X"06540215f06c", -- 3369
    X"c0602686600a", -- 3370
    X"15500115f044", -- 3371
    X"86500a195028", -- 3372
    X"06670a87000a", -- 3373
    X"80060b87100a", -- 3374
    X"10000186501a", -- 3375
    X"87200a06670a", -- 3376
    X"86502a80160b", -- 3377
    X"06670a111001", -- 3378
    X"80260b87300a", -- 3379
    X"12200186503a", -- 3380
    X"06670a155005", -- 3381
    X"13300180360b", -- 3382
    X"1440058e59b9", -- 3383
    X"14f02e8e4829", -- 3384
    X"8140aa80409a", -- 3385
    X"d400018240ba", -- 3386
    X"06540215f06c", -- 3387
    X"c0602686600a", -- 3388
    X"15500215f044", -- 3389
    X"86500a195028", -- 3390
    X"06670a87000a", -- 3391
    X"80060b87100a", -- 3392
    X"10000186501a", -- 3393
    X"87200a06670a", -- 3394
    X"86502a80160b", -- 3395
    X"155005111001", -- 3396
    X"80260b06670a", -- 3397
    X"8f5909122001", -- 3398
    X"384028144005", -- 3399
    X"14f02ecf8e64", -- 3400
    X"8140da8040ca", -- 3401
    X"15f06cd40002", -- 3402
    X"86600a065402", -- 3403
    X"15f044c06026", -- 3404
    X"195028155003", -- 3405
    X"87000a86500a", -- 3406
    X"87100a06670a", -- 3407
    X"86501a80060b", -- 3408
    X"155005100001", -- 3409
    X"80160b06670a", -- 3410
    X"8f5959111001", -- 3411
    X"384028144005", -- 3412
    X"d0ffffcf8eb4", -- 3413
    X"d0000181f00b", -- 3414
    X"10f02e81f01b", -- 3415
    X"80000a100007", -- 3416
    X"10f02e81f02b", -- 3417
    X"80000a10000a", -- 3418
    X"10f02e81f03b", -- 3419
    X"80000a10000c", -- 3420
    X"10f02e81f04b", -- 3421
    X"80000a100003", -- 3422
    X"d0000381f05b", -- 3423
    X"d1ffff82f01b", -- 3424
    X"d1000181f1db", -- 3425
    X"d3ffff81f1eb", -- 3426
    X"d5ffffd40000", -- 3427
    X"87700a17f09a", -- 3428
    X"c1acf9177002", -- 3429
    X"c0008bc1ad8a", -- 3430
    X"88700ad20002", -- 3431
    X"c09060098506", -- 3432
    X"da0000093206", -- 3433
    X"158000809a38", -- 3434
    X"122005102000", -- 3435
    X"130000177005", -- 3436
    X"d5199a81f0fb", -- 3437
    X"12f02e05050a", -- 3438
    X"81200a122002", -- 3439
    X"16f09a011502", -- 3440
    X"06600286600a", -- 3441
    X"88100a86600a", -- 3442
    X"08890bd92000", -- 3443
    X"85503081f14a", -- 3444
    X"12f015011502", -- 3445
    X"15f09a82200a", -- 3446
    X"10f02185500a", -- 3447
    X"05500280000a", -- 3448
    X"c1b14ac1af59", -- 3449
    X"83500ac0008b", -- 3450
    X"008023036302", -- 3451
    X"11100187100a", -- 3452
    X"0a7b13db4000", -- 3453
    X"12200187200a", -- 3454
    X"0a7b13db2000", -- 3455
    X"0b330a0aa009", -- 3456
    X"87700a17f01e", -- 3457
    X"17f01d0c7b0b", -- 3458
    X"00c02387700a", -- 3459
    X"c0c0a10c7a14", -- 3460
    X"807b0b17f01d", -- 3461
    X"80730b17f01c", -- 3462
    X"807a0b17f01e", -- 3463
    X"81f7ab87f1fa", -- 3464
    X"10000581f0bb", -- 3465
    X"144001155005", -- 3466
    X"d7000283f1fa", -- 3467
    X"87f1aa8a47f9", -- 3468
    X"87f1ba81f7fb", -- 3469
    X"8df1ca82f70b", -- 3470
    X"800d0b10f095", -- 3471
    X"d7200086f1ea", -- 3472
    X"d0ffff06670b", -- 3473
    X"d0000181f0db", -- 3474
    X"15f02e81f0eb", -- 3475
    X"80f1fa85509a", -- 3476
    X"00040ad4199a", -- 3477
    X"85f13a000502", -- 3478
    X"01140a81f20a", -- 3479
    X"15f02e011502", -- 3480
    X"13f03c82501a", -- 3481
    X"c1b45ac1b379", -- 3482
    X"88000ac0008b", -- 3483
    X"d42000100008", -- 3484
    X"00802308840b", -- 3485
    X"11100888100a", -- 3486
    X"88200a088413", -- 3487
    X"d41000122001", -- 3488
    X"088009088413", -- 3489
    X"13300180380b", -- 3490
    X"85506a15f02e", -- 3491
    X"d4199a80f1fa", -- 3492
    X"00050200040a", -- 3493
    X"81f20a85f12a", -- 3494
    X"01150201140a", -- 3495
    X"82500a15f02e", -- 3496
    X"83505a15f02e", -- 3497
    X"1af09ad50000", -- 3498
    X"0aa5028aa00a", -- 3499
    X"1df0958aa00a", -- 3500
    X"0dad028dd00a", -- 3501
    X"88000a006023", -- 3502
    X"d41000100008", -- 3503
    X"88100a088413", -- 3504
    X"088413111008", -- 3505
    X"12200188200a", -- 3506
    X"088413d40800", -- 3507
    X"82f62b14f03c", -- 3508
    X"dc000182f73b", -- 3509
    X"c1b89ac1b6f9", -- 3510
    X"16f09ac0008b", -- 3511
    X"db10008a300a", -- 3512
    X"86600a008023", -- 3513
    X"0aab13133001", -- 3514
    X"8a400a066c02", -- 3515
    X"86600adb4000", -- 3516
    X"0aab13144001", -- 3517
    X"07a009066d02", -- 3518
    X"06660a8af1ea", -- 3519
    X"00a0230aa60b", -- 3520
    X"0aa7148af1da", -- 3521
    X"81f6dbc0a051", -- 3522
    X"81f5ab81f7eb", -- 3523
    X"1cc00581fcbb", -- 3524
    X"86f22a155005", -- 3525
    X"da002887f23a", -- 3526
    X"8af11a8c5a79", -- 3527
    X"0aab0b8bf1da", -- 3528
    X"8af10a00a023", -- 3529
    X"0aab148bf1ea", -- 3530
    X"8af1dac0a0d1", -- 3531
    X"8af1ea81fa0b", -- 3532
    X"8af1fa81fa1b", -- 3533
    X"8af20a81fa8b", -- 3534
    X"8af1aa81fa9b", -- 3535
    X"8af1ba81fa6b", -- 3536
    X"d0ffff81fa7b", -- 3537
    X"d0000181f0db", -- 3538
    X"d1ffff81f0eb", -- 3539
    X"d2ffffd00000", -- 3540
    X"c1bb9ac1bb09", -- 3541
    X"83f21ac0008b", -- 3542
    X"84400a14f09a", -- 3543
    X"86600a064302", -- 3544
    X"c05060056206", -- 3545
    X"d70000051306", -- 3546
    X"126000805738", -- 3547
    X"13300581f3fb", -- 3548
    X"d4199a81f1fa", -- 3549
    X"84f15a03140a", -- 3550
    X"15f09a044302", -- 3551
    X"05510285500a", -- 3552
    X"82f52b85500a", -- 3553
    X"d7200086400a", -- 3554
    X"84f12a06670b", -- 3555
    X"15f02e044302", -- 3556
    X"c1bd0985500a", -- 3557
    X"c0008bc1beda", -- 3558
    X"83300a13f09a", -- 3559
    X"88f22a82300a", -- 3560
    X"006023028202", -- 3561
    X"14400888400a", -- 3562
    X"088913d94000", -- 3563
    X"15500188500a", -- 3564
    X"088913d92000", -- 3565
    X"09220a088009", -- 3566
    X"0aa90b8af1ea", -- 3567
    X"8af1da00a023", -- 3568
    X"c0a0a10aa814", -- 3569
    X"81f2cb81f9db", -- 3570
    X"82f1fa81f8eb", -- 3571
    X"12f09a81f2ab", -- 3572
    X"02320682200a", -- 3573
    X"13300581f2bb", -- 3574
    X"d20002100001", -- 3575
    X"80f1aa8b0299", -- 3576
    X"80f1ba81f0fb", -- 3577
    X"d2199a82f00b", -- 3578
    X"84403004020a", -- 3579
    X"86f1ea85f1ca", -- 3580
    X"06670bd72000", -- 3581
    X"81f0dbd0ffff", -- 3582
    X"81f0ebd00001", -- 3583
    X"81f14a80f1fa", -- 3584
    X"00020ad2199a", -- 3585
    X"11f02e001002", -- 3586
    X"01140281106a", -- 3587
    X"82202a12f02e", -- 3588
    X"c1c0e913f03c", -- 3589
    X"c0008bc1c1da", -- 3590
    X"10000888000a", -- 3591
    X"08890bd92000", -- 3592
    X"88100a008023", -- 3593
    X"d92000111001", -- 3594
    X"88200a088913", -- 3595
    X"d91000122001", -- 3596
    X"088009088913", -- 3597
    X"13300180380b", -- 3598
    X"81f13a80f1fa", -- 3599
    X"00020ad2199a", -- 3600
    X"11f02e001002", -- 3601
    X"01140281105a", -- 3602
    X"82201a12f02e", -- 3603
    X"83309a13f02e", -- 3604
    X"84400a14f09a", -- 3605
    X"8c400a144001", -- 3606
    X"0060230c5c02", -- 3607
    X"10000888000a", -- 3608
    X"088913d91000", -- 3609
    X"11100188100a", -- 3610
    X"088913d91000", -- 3611
    X"12200188200a", -- 3612
    X"088913d90800", -- 3613
    X"82f73b82f62b", -- 3614
    X"c1c45916f03c", -- 3615
    X"c0008bc1c62a", -- 3616
    X"87700a17f09a", -- 3617
    X"8d700a177002", -- 3618
    X"db10008a300a", -- 3619
    X"0dcd02008023", -- 3620
    X"0aab13133001", -- 3621
    X"db40008a600a", -- 3622
    X"1660010ddd0a", -- 3623
    X"0ea0090aab13", -- 3624
    X"0aad0b8af1ea", -- 3625
    X"8af1da00a023", -- 3626
    X"c0a0b10aae14", -- 3627
    X"81feeb81fddb", -- 3628
    X"8aa00a1af09a", -- 3629
    X"81faab0a4a06", -- 3630
    X"8aa00a1af09a", -- 3631
    X"81fabb0a7a06", -- 3632
    X"86f22a177005", -- 3633
    X"14400587f23a", -- 3634
    X"8aa00a1af09a", -- 3635
    X"1aa0011aa028", -- 3636
    X"8af11a8c4a39", -- 3637
    X"0aab0b8bf1da", -- 3638
    X"8af10a00a023", -- 3639
    X"0aab148bf1ea", -- 3640
    X"8af1dac0a0d1", -- 3641
    X"8af1ea81fa0b", -- 3642
    X"8af1fa81fa1b", -- 3643
    X"8af20a81fa9b", -- 3644
    X"8af1aa81fa6b", -- 3645
    X"8af1ba81fa7b", -- 3646
    X"1bf02e81fa8b", -- 3647
    X"81fa2b8ab08a", -- 3648
    X"81fa3b8ab0ba", -- 3649
    X"81fa4b8ab0da", -- 3650
    X"81fa5b8ab04a", -- 3651
    X"10000180f21a", -- 3652
    X"31000582f01b", -- 3653
    X"14f06cce1354", -- 3654
    X"05450285f16a", -- 3655
    X"85f17a80500a", -- 3656
    X"81500a054502", -- 3657
    X"05450285f18a", -- 3658
    X"85f19a82500a", -- 3659
    X"83500a054502", -- 3660
    X"84400a14f097", -- 3661
    X"c1ca09d50000", -- 3662
    X"c0028bc1ca1a", -- 3663
    X"14400180450b", -- 3664
    X"84400a14f097", -- 3665
    X"86f16a850022", -- 3666
    X"80650b064602", -- 3667
    X"86f17a851022", -- 3668
    X"80650b064602", -- 3669
    X"86f18a852022", -- 3670
    X"80650b064602", -- 3671
    X"86f19a853022", -- 3672
    X"80650b064602", -- 3673
    X"84400a14f096", -- 3674
    X"c0507085f16a", -- 3675
    X"c1cbdac1cbc9", -- 3676
    X"d5000000501e", -- 3677
    X"14400180450b", -- 3678
    X"c1cca9c00110", -- 3679
    X"86f16ac1ccda", -- 3680
    X"077606d70028", -- 3681
    X"14f09800701e", -- 3682
    X"15f09684400a", -- 3683
    X"05560285500a", -- 3684
    X"14400187400a", -- 3685
    X"15500180570b", -- 3686
    X"c1cda9c1cdf8", -- 3687
    X"86f16ac1cdea", -- 3688
    X"077606d70028", -- 3689
    X"14f09800701e", -- 3690
    X"15f09684400a", -- 3691
    X"05560285500a", -- 3692
    X"14400187400a", -- 3693
    X"80570b077004", -- 3694
    X"c01130155001", -- 3695
    X"c1cf0ac1ceb9", -- 3696
    X"d7002886f17a", -- 3697
    X"00701e077606", -- 3698
    X"84400a14f098", -- 3699
    X"85500a15f096", -- 3700
    X"87400a055602", -- 3701
    X"86500a144001", -- 3702
    X"80570b076702", -- 3703
    X"c1d038155001", -- 3704
    X"c1d02ac1cfd9", -- 3705
    X"d7002886f17a", -- 3706
    X"00701e077606", -- 3707
    X"84400a14f098", -- 3708
    X"85500a15f096", -- 3709
    X"87400a055602", -- 3710
    X"86500a144001", -- 3711
    X"80570b076706", -- 3712
    X"c02130155001", -- 3713
    X"c1d14ac1d0f9", -- 3714
    X"d7002886f18a", -- 3715
    X"00701e077606", -- 3716
    X"84400a14f098", -- 3717
    X"85500a15f096", -- 3718
    X"87400a055602", -- 3719
    X"86500a144001", -- 3720
    X"80570b076702", -- 3721
    X"c1d278155001", -- 3722
    X"c1d26ac1d219", -- 3723
    X"d7002886f18a", -- 3724
    X"00701e077606", -- 3725
    X"84400a14f098", -- 3726
    X"85500a15f096", -- 3727
    X"87400a055602", -- 3728
    X"86500a144001", -- 3729
    X"80570b076706", -- 3730
    X"c03130155001", -- 3731
    X"c1d38ac1d339", -- 3732
    X"d7002886f19a", -- 3733
    X"00701e077606", -- 3734
    X"84400a14f098", -- 3735
    X"85500a15f096", -- 3736
    X"87400a055602", -- 3737
    X"86500a144001", -- 3738
    X"80570b076702", -- 3739
    X"c1d4b8155001", -- 3740
    X"c1d4aac1d459", -- 3741
    X"d7002886f19a", -- 3742
    X"00701e077606", -- 3743
    X"84400a14f098", -- 3744
    X"85500a15f096", -- 3745
    X"87400a055602", -- 3746
    X"86500a144001", -- 3747
    X"80570b076706", -- 3748
    X"d40000155001", -- 3749
    X"144001c00020", -- 3750
    X"144002c01020", -- 3751
    X"144004c02020", -- 3752
    X"144008c03020", -- 3753
    X"80540b15f095", -- 3754
    X"85f16ad7199a", -- 3755
    X"81f56b05570a", -- 3756
    X"05570a85f17a", -- 3757
    X"85f18a81f57b", -- 3758
    X"81f58b05570a", -- 3759
    X"04570a85f19a", -- 3760
    X"054502854020", -- 3761
    X"15500386f19a", -- 3762
    X"864010056506", -- 3763
    X"81f59b055602", -- 3764
    X"84f16a85f17a", -- 3765
    X"044502855030", -- 3766
    X"85506085f18a", -- 3767
    X"85f19a044502", -- 3768
    X"044502855090", -- 3769
    X"80540b15f094", -- 3770
    X"81f02a80f01a", -- 3771
    X"83f04a82f03a", -- 3772
    X"85f06a84f05a", -- 3773
    X"87f08a86f07a", -- 3774
    X"89f0aa88f09a", -- 3775
    X"8bf0ca8af0ba", -- 3776
    X"8df0ea8cf0da", -- 3777
    X"1ff09a8ef0fa", -- 3778
    X"3ff03800e01a", -- 3779
    X"80f12b80f01b", -- 3780
    X"80f34b80f23b", -- 3781
    X"c1d92980f45b", -- 3782
    X"c0028bc1d96a", -- 3783
    X"11f00c80f36a", -- 3784
    X"10000182000a", -- 3785
    X"80120b822032", -- 3786
    X"c1d9e9111001", -- 3787
    X"c0028bc1da0a", -- 3788
    X"d2000110f00c", -- 3789
    X"002023d30000", -- 3790
    X"10000181000a", -- 3791
    X"002012021113", -- 3792
    X"01200902200e", -- 3793
    X"84f35a120003", -- 3794
    X"84f34a80412b", -- 3795
    X"c1db1980422b", -- 3796
    X"c0028bc1db5a", -- 3797
    X"81f38a10f00c", -- 3798
    X"d30000d20001", -- 3799
    X"82000a002023", -- 3800
    X"83100a100001", -- 3801
    X"022313111001", -- 3802
    X"02200e002012", -- 3803
    X"120ffa012009", -- 3804
    X"01100484f35a", -- 3805
    X"84f34a80413b", -- 3806
    X"80423b322001", -- 3807
    X"c1dccac1dc89", -- 3808
    X"10f00cc0028b", -- 3809
    X"d2000181f37a", -- 3810
    X"002023d30000", -- 3811
    X"10000182000a", -- 3812
    X"11100183100a", -- 3813
    X"002012022313", -- 3814
    X"01200902200e", -- 3815
    X"84f35a120ffa", -- 3816
    X"84f34a80414b", -- 3817
    X"80424b322001", -- 3818
    X"81f02a80f01a", -- 3819
    X"83f04a82f03a", -- 3820
    X"1ff03884f05a", -- 3821
    X"3ff00400e01a", -- 3822
    X"80f12b80f01b", -- 3823
    X"80f34b80f23b", -- 3824
    X"c1de99000026", -- 3825
    X"c0050bc1deda", -- 3826
    X"d1fffed0ffff", -- 3827
    X"83000ad200a0", -- 3828
    X"83100acf3ff0", -- 3829
    X"12200180230b", -- 3830
    X"80f01a000025", -- 3831
    X"82f03a81f02a", -- 3832
    X"1ff00483f04a", -- 3833
    X"3ff01000001d", -- 3834
    X"80f12b80f01b", -- 3835
    X"80f34b80f23b", -- 3836
    X"80f56b80f45b", -- 3837
    X"80f78b80f67b", -- 3838
    X"80f9ab80f89b", -- 3839
    X"80fbcb80fabb", -- 3840
    X"80000ad01568", -- 3841
    X"81100a81f10a", -- 3842
    X"26000000010b", -- 3843
    X"d36ca8d2afc0", -- 3844
    X"0220038220f3", -- 3845
    X"81f0da103000", -- 3846
    X"84f10a00010b", -- 3847
    X"c0403484401a", -- 3848
    X"c1e158d50000", -- 3849
    X"824071d5ffff", -- 3850
    X"822021022007", -- 3851
    X"d5bd31143000", -- 3852
    X"d2488004450b", -- 3853
    X"8220a3d36730", -- 3854
    X"183000026207", -- 3855
    X"08890a89f0da", -- 3856
    X"80002ad01568", -- 3857
    X"d0156806800b", -- 3858
    X"81f10a80000a", -- 3859
    X"00010b81101a", -- 3860
    X"026007800033", -- 3861
    X"183000822021", -- 3862
    X"0a8b0bdbbd31", -- 3863
    X"08890a89f0da", -- 3864
    X"d80000c09220", -- 3865
    X"d2000880f8fb", -- 3866
    X"d01570322004", -- 3867
    X"80000a000802", -- 3868
    X"80003300090b", -- 3869
    X"c0002300a007", -- 3870
    X"188001c1e438", -- 3871
    X"03820680f8fb", -- 3872
    X"d60000cf3f54", -- 3873
    X"d2001080f6eb", -- 3874
    X"d01574322008", -- 3875
    X"80000a000602", -- 3876
    X"80005300090b", -- 3877
    X"c00023004007", -- 3878
    X"166001c1e748", -- 3879
    X"03620680f6eb", -- 3880
    X"c1e748cf3f54", -- 3881
    X"80f8fbd80000", -- 3882
    X"322004d20008", -- 3883
    X"108000d01570", -- 3884
    X"00090b80000a", -- 3885
    X"00a007800033", -- 3886
    X"c1e648c00025", -- 3887
    X"80f8fb188001", -- 3888
    X"cf3f52038206", -- 3889
    X"80f6ebd60000", -- 3890
    X"322008d20010", -- 3891
    X"106000d01574", -- 3892
    X"00090b80000a", -- 3893
    X"004007800053", -- 3894
    X"c1e748c00027", -- 3895
    X"80f6eb166001", -- 3896
    X"cf3f54036206", -- 3897
    X"81f02a80f01a", -- 3898
    X"83f04a82f03a", -- 3899
    X"85f06a84f05a", -- 3900
    X"87f08a86f07a", -- 3901
    X"89f0aa88f09a", -- 3902
    X"8bf0ca8af0ba", -- 3903
    X"00e01a1ff010", -- 3904
    X"80f01b3ff00b", -- 3905
    X"80f23b80f12b", -- 3906
    X"80f45b80f34b", -- 3907
    X"80f67b80f56b", -- 3908
    X"80f89b80f78b", -- 3909
    X"d1ffffd0ffff", -- 3910
    X"32202882f0aa", -- 3911
    X"c02186182000", -- 3912
    X"84200ad20335", -- 3913
    X"04400885201a", -- 3914
    X"04421782f0ba", -- 3915
    X"d64000844011", -- 3916
    X"044603d70000", -- 3917
    X"c02021024007", -- 3918
    X"044008204000", -- 3919
    X"04421782f0ba", -- 3920
    X"d64000844011", -- 3921
    X"044603d70000", -- 3922
    X"c02021024007", -- 3923
    X"d2161e204000", -- 3924
    X"82200a022802", -- 3925
    X"33300183f0aa", -- 3926
    X"033402d4161e", -- 3927
    X"04320683300a", -- 3928
    X"144001c04154", -- 3929
    X"c1ec6ac1eba9", -- 3930
    X"d4033500401e", -- 3931
    X"044202044202", -- 3932
    X"83401a82400a", -- 3933
    X"85f0ba022008", -- 3934
    X"822011022517", -- 3935
    X"d70000d64000", -- 3936
    X"062007022603", -- 3937
    X"202000c06021", -- 3938
    X"d40335144002", -- 3939
    X"83405a82404a", -- 3940
    X"80437b80426b", -- 3941
    X"83403a82402a", -- 3942
    X"80435b80424b", -- 3943
    X"83401a82400a", -- 3944
    X"80433b80422b", -- 3945
    X"80411b80400b", -- 3946
    X"81f02a80f01a", -- 3947
    X"83f04a82f03a", -- 3948
    X"85f06a84f05a", -- 3949
    X"87f08a86f07a", -- 3950
    X"1ff00b88f09a", -- 3951
    X"3ff03300e01a", -- 3952
    X"80f12b80f01b", -- 3953
    X"80f34b80f23b", -- 3954
    X"80f56b80f45b", -- 3955
    X"80f78b80f67b", -- 3956
    X"80f9ab80f89b", -- 3957
    X"80fbcb80fabb", -- 3958
    X"80fdeb80fcdb", -- 3959
    X"d002ff80fefb", -- 3960
    X"d0065c80f00b", -- 3961
    X"be05c48ff0fb", -- 3962
    X"81ffda80ffea", -- 3963
    X"82f32a82f1db", -- 3964
    X"85202a84200a", -- 3965
    X"86204a04450b", -- 3966
    X"83f31a06660b", -- 3967
    X"89302a88300a", -- 3968
    X"388001088902", -- 3969
    X"09990289304a", -- 3970
    X"0a8906199001", -- 3971
    X"0c4a10c0a050", -- 3972
    X"1b90000cc607", -- 3973
    X"0aa004c1f118", -- 3974
    X"0c4c070c6a10", -- 3975
    X"04c0121b8000", -- 3976
    X"06b40206c40e", -- 3977
    X"d44000366010", -- 3978
    X"8ff7fb80f40b", -- 3979
    X"87ffeabe00cf", -- 3980
    X"81f7ab077004", -- 3981
    X"06600436601d", -- 3982
    X"84202a81f6bb", -- 3983
    X"04450b85201a", -- 3984
    X"87204a86203a", -- 3985
    X"88302a06670b", -- 3986
    X"08890289301a", -- 3987
    X"8a304a89303a", -- 3988
    X"199001099a02", -- 3989
    X"c0a0700a8906", -- 3990
    X"044a101aa001", -- 3991
    X"0c4607866013", -- 3992
    X"c1f3a83b9001", -- 3993
    X"1aa0010aa004", -- 3994
    X"844013066a10", -- 3995
    X"3b80010c4607", -- 3996
    X"06c40e04c012", -- 3997
    X"36601006b402", -- 3998
    X"04650285f1ba", -- 3999
    X"85f1aa344018", -- 4000
    X"06641006750b", -- 4001
    X"84f2ea81f7cb", -- 4002
    X"804559d50001", -- 4003
    X"047506d501e1", -- 4004
    X"81f5cbc04020", -- 4005
    X"85203a84200a", -- 4006
    X"86201a04450b", -- 4007
    X"06670b87204a", -- 4008
    X"89303a88300a", -- 4009
    X"89301a088902", -- 4010
    X"099a028a304a", -- 4011
    X"0a8906199001", -- 4012
    X"1aa001c0a070", -- 4013
    X"866013044a10", -- 4014
    X"3b90010c4607", -- 4015
    X"0aa004c1f678", -- 4016
    X"066a101aa001", -- 4017
    X"0c4607844013", -- 4018
    X"04c0123b8001", -- 4019
    X"06b40206c40e", -- 4020
    X"85f1ba366010", -- 4021
    X"344011046502", -- 4022
    X"06750b85f1aa", -- 4023
    X"15f01c066410", -- 4024
    X"35100480571b", -- 4025
    X"02050fc05034", -- 4026
    X"140000c1f7d8", -- 4027
    X"331014d50000", -- 4028
    X"04430e033004", -- 4029
    X"14f01c125000", -- 4030
    X"8ff2db80f40b", -- 4031
    X"82fffabe1df5", -- 4032
    X"81f20b83ffea", -- 4033
    X"14f01e81f31b", -- 4034
    X"86500a85f31a", -- 4035
    X"80460b16600d", -- 4036
    X"16600e86501a", -- 4037
    X"87101080461b", -- 4038
    X"86502a377015", -- 4039
    X"80462b066702", -- 4040
    X"86503a371003", -- 4041
    X"80463b066702", -- 4042
    X"86504a371004", -- 4043
    X"80464b066702", -- 4044
    X"14400186400a", -- 4045
    X"c1fa4ac1f9f9", -- 4046
    X"85400ac0004b", -- 4047
    X"075606144001", -- 4048
    X"165000c07026", -- 4049
    X"c1fac9000024", -- 4050
    X"c0005bc1fb7a", -- 4051
    X"85f32a14f01e", -- 4052
    X"1cf0231bf028", -- 4053
    X"1440018a400a", -- 4054
    X"d8000007a606", -- 4055
    X"15500189500a", -- 4056
    X"088008088710", -- 4057
    X"1bb00180b90b", -- 4058
    X"1cc00180c80b", -- 4059
    X"d57fffd4ffff", -- 4060
    X"81f57b81f46b", -- 4061
    X"d9000188f2ea", -- 4062
    X"d800008489e9", -- 4063
    X"c2007ac1fc49", -- 4064
    X"d90000c0008b", -- 4065
    X"02280282f10a", -- 4066
    X"d61520722002", -- 4067
    X"83f11a022602", -- 4068
    X"733002033902", -- 4069
    X"033602d61530", -- 4070
    X"87300a86200a", -- 4071
    X"d73fff016702", -- 4072
    X"c07346071706", -- 4073
    X"d7000086201a", -- 4074
    X"db00008a301a", -- 4075
    X"866013066a03", -- 4076
    X"07110a06060a", -- 4077
    X"0b610a0a660a", -- 4078
    X"15f02314f028", -- 4079
    X"81f33b81f22b", -- 4080
    X"81f95b81f84b", -- 4081
    X"8d400a8c500a", -- 4082
    X"8c501a02c717", -- 4083
    X"08c1178d401a", -- 4084
    X"8c502a022803", -- 4085
    X"08ca178d402a", -- 4086
    X"8c503a022803", -- 4087
    X"08c6178d403a", -- 4088
    X"8c504a022803", -- 4089
    X"08cb178d404a", -- 4090
    X"82f12a0c2803", -- 4091
    X"88f14a83f13a", -- 4092
    X"84f16a89f15a", -- 4093
    X"04c40785f17a", -- 4094
    X"81fc6bc04097", -- 4095
    X"82f10a81fd7b", -- 4096
    X"81f48b042802", -- 4097
    X"05390283f11a", -- 4098
    X"19900181f59b", -- 4099
    X"d90004188001", -- 4100
    X"c205588b8969", -- 4101
    X"c20119d80000", -- 4102
    X"c0008bc2051a", -- 4103
    X"82f10ad90000", -- 4104
    X"722002022802", -- 4105
    X"022602d61520", -- 4106
    X"03390283f11a", -- 4107
    X"d71530733002", -- 4108
    X"86200a033702", -- 4109
    X"01670287300a", -- 4110
    X"d7000086201a", -- 4111
    X"db00008a301a", -- 4112
    X"866013066a03", -- 4113
    X"07110a06060a", -- 4114
    X"0b610a0a660a", -- 4115
    X"15f02314f028", -- 4116
    X"81f33b81f22b", -- 4117
    X"81f95b81f84b", -- 4118
    X"8d400a8c500a", -- 4119
    X"8c501a02c717", -- 4120
    X"08c1178d401a", -- 4121
    X"8c502a022803", -- 4122
    X"08ca178d402a", -- 4123
    X"8c503a022803", -- 4124
    X"08c6178d403a", -- 4125
    X"8c504a022803", -- 4126
    X"08cb178d404a", -- 4127
    X"82f12a0c2803", -- 4128
    X"88f14a83f13a", -- 4129
    X"84f16a89f15a", -- 4130
    X"04c40785f17a", -- 4131
    X"81fc6bc04097", -- 4132
    X"82f10a81fd7b", -- 4133
    X"81f48b042802", -- 4134
    X"05390283f11a", -- 4135
    X"19900181f59b", -- 4136
    X"d90004188001", -- 4137
    X"82f18a8b8999", -- 4138
    X"d41520722002", -- 4139
    X"83f19a022402", -- 4140
    X"d51530733002", -- 4141
    X"84200a033502", -- 4142
    X"06450285300a", -- 4143
    X"84201a83f60b", -- 4144
    X"86301ad50000", -- 4145
    X"084603d70000", -- 4146
    X"04600b868013", -- 4147
    X"06600486f2da", -- 4148
    X"04460e166004", -- 4149
    X"d002ff82f5fb", -- 4150
    X"8ff9fb80f00b", -- 4151
    X"be067f8ff8eb", -- 4152
    X"d0155081f18a", -- 4153
    X"81100a010102", -- 4154
    X"82f19a711010", -- 4155
    X"020202d01558", -- 4156
    X"00120282200a", -- 4157
    X"80f01a82f0db", -- 4158
    X"82f03a81f02a", -- 4159
    X"84f05a83f04a", -- 4160
    X"86f07a85f06a", -- 4161
    X"88f09a87f08a", -- 4162
    X"8af0ba89f0aa", -- 4163
    X"8cf0da8bf0ca", -- 4164
    X"8ef0fa8df0ea", -- 4165
    X"00e01a1ff033", -- 4166
    X"80f01b3ff008", -- 4167
    X"80f23b80f12b", -- 4168
    X"80f45b80f34b", -- 4169
    X"80f08a80f56b", -- 4170
    X"81000a84f07a", -- 4171
    X"021518d50080", -- 4172
    X"d500ffc02042", -- 4173
    X"c20a08011518", -- 4174
    X"011519d5ff00", -- 4175
    X"81001a821080", -- 4176
    X"d500ff831022", -- 4177
    X"022319033518", -- 4178
    X"d5000280420b", -- 4179
    X"c02042021518", -- 4180
    X"011518d50003", -- 4181
    X"d5fffcc20af8", -- 4182
    X"8210e0011519", -- 4183
    X"83106081002a", -- 4184
    X"033518d53fff", -- 4185
    X"81003a022319", -- 4186
    X"031518d50800", -- 4187
    X"d5001fc03042", -- 4188
    X"c20be8011518", -- 4189
    X"011519d5ffe0", -- 4190
    X"d507ff831050", -- 4191
    X"022319033518", -- 4192
    X"83108281004a", -- 4193
    X"033518d507ff", -- 4194
    X"80421b022319", -- 4195
    X"021518d50080", -- 4196
    X"d500ffc02042", -- 4197
    X"c20d08011518", -- 4198
    X"011519d5ff00", -- 4199
    X"81005a821080", -- 4200
    X"d500ff831040", -- 4201
    X"022319033518", -- 4202
    X"83103281006a", -- 4203
    X"033518d5000f", -- 4204
    X"80422b022319", -- 4205
    X"021518d50004", -- 4206
    X"d50007c02042", -- 4207
    X"c20e48011518", -- 4208
    X"011519d5fff8", -- 4209
    X"81007a8210d0", -- 4210
    X"d51fff831080", -- 4211
    X"022319033518", -- 4212
    X"83105281008a", -- 4213
    X"033518d500ff", -- 4214
    X"80423b022319", -- 4215
    X"021518d50010", -- 4216
    X"d5001fc02042", -- 4217
    X"c20f88011518", -- 4218
    X"011519d5ffe0", -- 4219
    X"81009a8210b0", -- 4220
    X"d507ff831070", -- 4221
    X"022319033518", -- 4222
    X"d5007f8100aa", -- 4223
    X"022319031518", -- 4224
    X"80f01a80424b", -- 4225
    X"82f03a81f02a", -- 4226
    X"84f05a83f04a", -- 4227
    X"1ff00885f06a", -- 4228
    X"d000a000e01a", -- 4229
    X"be0e1c80f00b", -- 4230
    X"80f00bd00000", -- 4231
    X"8ff0fbd007a4", -- 4232
    X"8ff0ebd00799", -- 4233
    X"d00799be0e5e", -- 4234
    X"d007a480f00b", -- 4235
    X"d0000a8ff0fb", -- 4236
    X"be0edd8ff0eb", -- 4237
    X"80f00bd007a4", -- 4238
    X"8ff0fbd00799", -- 4239
    X"8ff0ebd006b1", -- 4240
    X"8ff0dbd007af", -- 4241
    X"d002b9be0f0a", -- 4242
    X"d0068480f00b", -- 4243
    X"d006b18ff0fb", -- 4244
    X"be10b08ff0eb", -- 4245
    X"80f00bd00684", -- 4246
    X"8ff0fbd007b9", -- 4247
    X"8ff0ebd007c6", -- 4248
    X"d002c3be125f", -- 4249
    X"d007b980f00b", -- 4250
    X"d0069b8ff0fb", -- 4251
    X"be04488ff0eb", -- 4252
    X"80f00bd0069b", -- 4253
    X"8ff0fbd06000", -- 4254
    X"8ff0ebd0000a", -- 4255
    X"8ff0dbd006b1", -- 4256
    X"d0069bbe0015", -- 4257
    X"10000110000a", -- 4258
    X"d0600080f00b", -- 4259
    X"d0000a8ff0fb", -- 4260
    X"d006b18ff0eb", -- 4261
    X"10000110000a", -- 4262
    X"be00158ff0db", -- 4263
    X"80f00bd00684", -- 4264
    X"8ff0fbd002b9", -- 4265
    X"8ff0ebd0000a", -- 4266
    X"d007b9be0000", -- 4267
    X"d002c380f00b", -- 4268
    X"d0000a8ff0fb", -- 4269
    X"be00008ff0eb", -- 4270
    X"d0069b3ff00b", -- 4271
    X"d0007880f00b", -- 4272
    X"d002698ff0fb", -- 4273
    X"be003e8ff0eb", -- 4274
    X"10000ad0069b", -- 4275
    X"80f00b100001", -- 4276
    X"100028d00078", -- 4277
    X"d002698ff0fb", -- 4278
    X"8ff0eb100028", -- 4279
    X"d006b1be003e", -- 4280
    X"11f001100001", -- 4281
    X"80120bd21000", -- 4282
    X"c217b9111001", -- 4283
    X"c000abc2181a", -- 4284
    X"840ffad3599a", -- 4285
    X"82000a04430a", -- 4286
    X"022406100001", -- 4287
    X"11100180120b", -- 4288
    X"80f40b14f001", -- 4289
    X"8ff4fbd40269", -- 4290
    X"8ff4ebd4017f", -- 4291
    X"8ff4dbd40028", -- 4292
    X"8ff4cbd402d7", -- 4293
    X"8ff4bbd40001", -- 4294
    X"100001be0075", -- 4295
    X"11100111f001", -- 4296
    X"c219bac21959", -- 4297
    X"840ffac000ab", -- 4298
    X"82000a04430a", -- 4299
    X"022406100001", -- 4300
    X"11100180120b", -- 4301
    X"80f40b14f001", -- 4302
    X"144028d40269", -- 4303
    X"d4017f8ff4fb", -- 4304
    X"8ff4eb144028", -- 4305
    X"8ff4dbd40028", -- 4306
    X"8ff4cbd402d7", -- 4307
    X"8ff4bbd40001", -- 4308
    X"1ff00bbe0075", -- 4309
    X"80f00bd0017f", -- 4310
    X"81fffabe127d", -- 4311
    X"31100384fffa", -- 4312
    X"c02026321014", -- 4313
    X"121006d10014", -- 4314
    X"c0303033208f", -- 4315
    X"312006d2008f", -- 4316
    X"1307c3d00000", -- 4317
    X"1307c480310b", -- 4318
    X"d007ce80320b", -- 4319
    X"80021b80010b", -- 4320
    X"00001d80042b", -- 4321
    X"80f00bd00690", -- 4322
    X"8ff0fbd0069c", -- 4323
    X"00001dbe208e", -- 4324
    X"c21d09000026", -- 4325
    X"00301ec21d4a", -- 4326
    X"d1fffcd0fffd", -- 4327
    X"cf4ff284000a", -- 4328
    X"12200184200a", -- 4329
    X"00002580140b", -- 4330
    X"3ff00500e01a", -- 4331
    X"80f12b80f01b", -- 4332
    X"80f34b80f23b", -- 4333
    X"d2069c80f45b", -- 4334
    X"be21cad30005", -- 4335
    X"81f02a80f01a", -- 4336
    X"83f04a82f03a", -- 4337
    X"1ff00584f05a", -- 4338
    X"3ff00500001d", -- 4339
    X"80f12b80f01b", -- 4340
    X"80f34b80f23b", -- 4341
    X"d2060b80f45b", -- 4342
    X"be21cad30050", -- 4343
    X"81f02a80f01a", -- 4344
    X"83f04a82f03a", -- 4345
    X"1ff00584f05a", -- 4346
    X"3ff00400001d", -- 4347
    X"80f12b80f01b", -- 4348
    X"80f34b80f23b", -- 4349
    X"c22039000026", -- 4350
    X"c0005bc2207a", -- 4351
    X"d1fffed0ffff", -- 4352
    X"83000ad2069c", -- 4353
    X"83100acf3ff0", -- 4354
    X"12200180230b", -- 4355
    X"80f01a000025", -- 4356
    X"82f03a81f02a", -- 4357
    X"1ff00483f04a", -- 4358
    X"3ff00400001d", -- 4359
    X"80f12b80f01b", -- 4360
    X"80f34b80f23b", -- 4361
    X"c221b9000026", -- 4362
    X"c068fbc221fa", -- 4363
    X"d1fffed0ffff", -- 4364
    X"83000ad20000", -- 4365
    X"83100acf3ff0", -- 4366
    X"12200180230b", -- 4367
    X"80f01a000025", -- 4368
    X"82f03a81f02a", -- 4369
    X"1ff00483f04a", -- 4370
    X"3ff00500001d", -- 4371
    X"80f12b80f01b", -- 4372
    X"80f34b80f23b", -- 4373
    X"d2000080f45b", -- 4374
    X"be21cad3068f", -- 4375
    X"81f02a80f01a", -- 4376
    X"83f04a82f03a", -- 4377
    X"1ff00584f05a", -- 4378
    X"00000000001d", -- 4379
    X"000000000000", -- 4380
    X"000000000000", -- 4381
    X"000000000000", -- 4382
    X"000000000000", -- 4383
    X"000000000000", -- 4384
    X"000000000000", -- 4385
    X"000000000000", -- 4386
    X"000000000000", -- 4387
    X"000000000000", -- 4388
    X"000000000000", -- 4389
    X"000000000000", -- 4390
    X"000000000000", -- 4391
    X"000000000000", -- 4392
    X"000000000000", -- 4393
    X"000000000000", -- 4394
    X"000000000000", -- 4395
    X"000000000000", -- 4396
    X"000000000000", -- 4397
    X"000000000000", -- 4398
    X"000000000000", -- 4399
    X"000000000000", -- 4400
    X"000000000000", -- 4401
    X"000000000000", -- 4402
    X"000000000000", -- 4403
    X"000000000000", -- 4404
    X"000000000000", -- 4405
    X"000000000000", -- 4406
    X"000000000000", -- 4407
    X"000000000000", -- 4408
    X"000000000000", -- 4409
    X"000000000000", -- 4410
    X"000000000000", -- 4411
    X"000000000000", -- 4412
    X"000000000000", -- 4413
    X"000000000000", -- 4414
    X"000000000000", -- 4415
    X"000000000000", -- 4416
    X"000000000000", -- 4417
    X"000000000000", -- 4418
    X"000000000000", -- 4419
    X"000000000000", -- 4420
    X"000000000000", -- 4421
    X"000000000000", -- 4422
    X"000000000000", -- 4423
    X"000000000000", -- 4424
    X"000000000000", -- 4425
    X"000000000000", -- 4426
    X"000000000000", -- 4427
    X"000000000000", -- 4428
    X"000000000000", -- 4429
    X"000000000000", -- 4430
    X"000000000000", -- 4431
    X"000000000000", -- 4432
    X"000000000000", -- 4433
    X"000000000000", -- 4434
    X"000000000000", -- 4435
    X"000000000000", -- 4436
    X"000000000000", -- 4437
    X"000000000000", -- 4438
    X"000000000000", -- 4439
    X"000000000000", -- 4440
    X"000000000000", -- 4441
    X"000000000000", -- 4442
    X"000000000000", -- 4443
    X"000000000000", -- 4444
    X"000000000000", -- 4445
    X"000000000000", -- 4446
    X"000000000000", -- 4447
    X"000000000000", -- 4448
    X"000000000000", -- 4449
    X"000000000000", -- 4450
    X"000000000000", -- 4451
    X"000000000000", -- 4452
    X"000000000000", -- 4453
    X"000000000000", -- 4454
    X"000000000000", -- 4455
    X"000000000000", -- 4456
    X"000000000000", -- 4457
    X"000000000000", -- 4458
    X"000000000000", -- 4459
    X"000000000000", -- 4460
    X"000000000000", -- 4461
    X"000000000000", -- 4462
    X"000000000000", -- 4463
    X"000000000000", -- 4464
    X"000000000000", -- 4465
    X"000000000000", -- 4466
    X"000000000000", -- 4467
    X"000000000000", -- 4468
    X"000000000000", -- 4469
    X"000000000000", -- 4470
    X"000000000000", -- 4471
    X"000000000000", -- 4472
    X"000000000000", -- 4473
    X"000000000000", -- 4474
    X"000000000000", -- 4475
    X"000000000000", -- 4476
    X"000000000000", -- 4477
    X"000000000000", -- 4478
    X"000000000000", -- 4479
    X"000000000000", -- 4480
    X"000000000000", -- 4481
    X"000000000000", -- 4482
    X"000000000000", -- 4483
    X"000000000000", -- 4484
    X"000000000000", -- 4485
    X"000000000000", -- 4486
    X"000000000000", -- 4487
    X"000000000000", -- 4488
    X"000000000000", -- 4489
    X"000000000000", -- 4490
    X"000000000000", -- 4491
    X"000000000000", -- 4492
    X"000000000000", -- 4493
    X"000000000000", -- 4494
    X"000000000000", -- 4495
    X"000000000000", -- 4496
    X"000000000000", -- 4497
    X"000000000000", -- 4498
    X"000000000000", -- 4499
    X"000000000000", -- 4500
    X"000000000000", -- 4501
    X"000000000000", -- 4502
    X"000000000000", -- 4503
    X"000000000000", -- 4504
    X"000000000000", -- 4505
    X"000000000000", -- 4506
    X"000000000000", -- 4507
    X"000000000000", -- 4508
    X"000000000000", -- 4509
    X"000000000000", -- 4510
    X"000000000000", -- 4511
    X"000000000000", -- 4512
    X"000000000000", -- 4513
    X"000000000000", -- 4514
    X"000000000000", -- 4515
    X"000000000000", -- 4516
    X"000000000000", -- 4517
    X"000000000000", -- 4518
    X"000000000000", -- 4519
    X"000000000000", -- 4520
    X"000000000000", -- 4521
    X"000000000000", -- 4522
    X"000000000000", -- 4523
    X"000000000000", -- 4524
    X"000000000000", -- 4525
    X"000000000000", -- 4526
    X"000000000000", -- 4527
    X"000000000000", -- 4528
    X"000000000000", -- 4529
    X"000000000000", -- 4530
    X"000000000000", -- 4531
    X"000000000000", -- 4532
    X"000000000000", -- 4533
    X"000000000000", -- 4534
    X"000000000000", -- 4535
    X"000000000000", -- 4536
    X"000000000000", -- 4537
    X"000000000000", -- 4538
    X"000000000000", -- 4539
    X"000000000000", -- 4540
    X"000000000000", -- 4541
    X"000000000000", -- 4542
    X"000000000000", -- 4543
    X"000000000000", -- 4544
    X"000000000000", -- 4545
    X"000000000000", -- 4546
    X"000000000000", -- 4547
    X"000000000000", -- 4548
    X"000000000000", -- 4549
    X"000000000000", -- 4550
    X"000000000000", -- 4551
    X"000000000000", -- 4552
    X"000000000000", -- 4553
    X"000000000000", -- 4554
    X"000000000000", -- 4555
    X"000000000000", -- 4556
    X"000000000000", -- 4557
    X"000000000000", -- 4558
    X"000000000000", -- 4559
    X"000000000000", -- 4560
    X"000000000000", -- 4561
    X"000000000000", -- 4562
    X"000000000000", -- 4563
    X"000000000000", -- 4564
    X"000000000000", -- 4565
    X"000000000000", -- 4566
    X"000000000000", -- 4567
    X"000000000000", -- 4568
    X"000000000000", -- 4569
    X"000000000000", -- 4570
    X"000000000000", -- 4571
    X"000000000000", -- 4572
    X"000000000000", -- 4573
    X"000000000000", -- 4574
    X"000000000000", -- 4575
    X"000000000000", -- 4576
    X"000000000000", -- 4577
    X"000000000000", -- 4578
    X"000000000000", -- 4579
    X"000000000000", -- 4580
    X"000000000000", -- 4581
    X"000000000000", -- 4582
    X"000000000000", -- 4583
    X"000000000000", -- 4584
    X"000000000000", -- 4585
    X"000000000000", -- 4586
    X"000000000000", -- 4587
    X"000000000000", -- 4588
    X"000000000000", -- 4589
    X"000000000000", -- 4590
    X"000000000000", -- 4591
    X"000000000000", -- 4592
    X"000000000000", -- 4593
    X"000000000000", -- 4594
    X"000000000000", -- 4595
    X"000000000000", -- 4596
    X"000000000000", -- 4597
    X"000000000000", -- 4598
    X"000000000000", -- 4599
    X"000000000000", -- 4600
    X"000000000000", -- 4601
    X"000000000000", -- 4602
    X"000000000000", -- 4603
    X"000000000000", -- 4604
    X"000000000000", -- 4605
    X"000000000000", -- 4606
    X"000000000000"  -- 4607
  );

--END;

end G729A_ASIP_ROMI_PKG;

package body G729A_ASIP_ROMI_PKG is

end G729A_ASIP_ROMI_PKG;

