// `include "encoder.v"

module design49_10_200_top #(parameter WIDTH=32,CHANNEL=10) (clk, rst, in, out);

	localparam OUT_BUS=CHANNEL*WIDTH;
	input clk,rst;
	input [WIDTH-1:0] in;
	output [WIDTH-1:0] out;

	reg [WIDTH-1:0] d_in0;
	reg [WIDTH-1:0] d_in1;
	reg [WIDTH-1:0] d_in2;
	reg [WIDTH-1:0] d_in3;
	reg [WIDTH-1:0] d_in4;
	reg [WIDTH-1:0] d_in5;
	reg [WIDTH-1:0] d_in6;
	reg [WIDTH-1:0] d_in7;
	reg [WIDTH-1:0] d_in8;
	reg [WIDTH-1:0] d_in9;
	wire [WIDTH-1:0] d_out0;
	wire [WIDTH-1:0] d_out1;
	wire [WIDTH-1:0] d_out2;
	wire [WIDTH-1:0] d_out3;
	wire [WIDTH-1:0] d_out4;
	wire [WIDTH-1:0] d_out5;
	wire [WIDTH-1:0] d_out6;
	wire [WIDTH-1:0] d_out7;
	wire [WIDTH-1:0] d_out8;
	wire [WIDTH-1:0] d_out9;

	reg [OUT_BUS-1:0] tmp;

	always @ (posedge clk or posedge rst) begin
		if (rst)
			tmp <= 0;
		else
			tmp <= {tmp[OUT_BUS-(WIDTH-1):0],in};
	end

	always @ (posedge clk) begin
		d_in0 <= tmp[WIDTH-1:0];
		d_in1 <= tmp[(WIDTH*2)-1:WIDTH*1];
		d_in2 <= tmp[(WIDTH*3)-1:WIDTH*2];
		d_in3 <= tmp[(WIDTH*4)-1:WIDTH*3];
		d_in4 <= tmp[(WIDTH*5)-1:WIDTH*4];
		d_in5 <= tmp[(WIDTH*6)-1:WIDTH*5];
		d_in6 <= tmp[(WIDTH*7)-1:WIDTH*6];
		d_in7 <= tmp[(WIDTH*8)-1:WIDTH*7];
		d_in8 <= tmp[(WIDTH*9)-1:WIDTH*8];
		d_in9 <= tmp[(WIDTH*10)-1:WIDTH*9];
	end

	design49_10_200 #(.WIDTH(WIDTH)) design49_10_200_inst(.d_in0(d_in0),.d_in1(d_in1),.d_in2(d_in2),.d_in3(d_in3),.d_in4(d_in4),.d_in5(d_in5),.d_in6(d_in6),.d_in7(d_in7),.d_in8(d_in8),.d_in9(d_in9),.d_out0(d_out0),.d_out1(d_out1),.d_out2(d_out2),.d_out3(d_out3),.d_out4(d_out4),.d_out5(d_out5),.d_out6(d_out6),.d_out7(d_out7),.d_out8(d_out8),.d_out9(d_out9),.clk(clk),.rst(rst));

	assign out = d_out0^d_out1^d_out2^d_out3^d_out4^d_out5^d_out6^d_out7^d_out8^d_out9;

endmodule

module design49_10_200 #(parameter WIDTH=32) (d_in0, d_in1, d_in2, d_in3, d_in4, d_in5, d_in6, d_in7, d_in8, d_in9, d_out0, d_out1, d_out2, d_out3, d_out4, d_out5, d_out6, d_out7, d_out8, d_out9, clk, rst);
	input clk;
	input rst;
	input [WIDTH-1:0] d_in0; 
	input [WIDTH-1:0] d_in1; 
	input [WIDTH-1:0] d_in2; 
	input [WIDTH-1:0] d_in3; 
	input [WIDTH-1:0] d_in4; 
	input [WIDTH-1:0] d_in5; 
	input [WIDTH-1:0] d_in6; 
	input [WIDTH-1:0] d_in7; 
	input [WIDTH-1:0] d_in8; 
	input [WIDTH-1:0] d_in9; 
	output [WIDTH-1:0] d_out0; 
	output [WIDTH-1:0] d_out1; 
	output [WIDTH-1:0] d_out2; 
	output [WIDTH-1:0] d_out3; 
	output [WIDTH-1:0] d_out4; 
	output [WIDTH-1:0] d_out5; 
	output [WIDTH-1:0] d_out6; 
	output [WIDTH-1:0] d_out7; 
	output [WIDTH-1:0] d_out8; 
	output [WIDTH-1:0] d_out9; 

	wire [WIDTH-1:0] wire_d0_0;
	wire [WIDTH-1:0] wire_d0_1;
	wire [WIDTH-1:0] wire_d0_2;
	wire [WIDTH-1:0] wire_d0_3;
	wire [WIDTH-1:0] wire_d0_4;
	wire [WIDTH-1:0] wire_d0_5;
	wire [WIDTH-1:0] wire_d0_6;
	wire [WIDTH-1:0] wire_d0_7;
	wire [WIDTH-1:0] wire_d0_8;
	wire [WIDTH-1:0] wire_d0_9;
	wire [WIDTH-1:0] wire_d0_10;
	wire [WIDTH-1:0] wire_d0_11;
	wire [WIDTH-1:0] wire_d0_12;
	wire [WIDTH-1:0] wire_d0_13;
	wire [WIDTH-1:0] wire_d0_14;
	wire [WIDTH-1:0] wire_d0_15;
	wire [WIDTH-1:0] wire_d0_16;
	wire [WIDTH-1:0] wire_d0_17;
	wire [WIDTH-1:0] wire_d0_18;
	wire [WIDTH-1:0] wire_d0_19;
	wire [WIDTH-1:0] wire_d0_20;
	wire [WIDTH-1:0] wire_d0_21;
	wire [WIDTH-1:0] wire_d0_22;
	wire [WIDTH-1:0] wire_d0_23;
	wire [WIDTH-1:0] wire_d0_24;
	wire [WIDTH-1:0] wire_d0_25;
	wire [WIDTH-1:0] wire_d0_26;
	wire [WIDTH-1:0] wire_d0_27;
	wire [WIDTH-1:0] wire_d0_28;
	wire [WIDTH-1:0] wire_d0_29;
	wire [WIDTH-1:0] wire_d0_30;
	wire [WIDTH-1:0] wire_d0_31;
	wire [WIDTH-1:0] wire_d0_32;
	wire [WIDTH-1:0] wire_d0_33;
	wire [WIDTH-1:0] wire_d0_34;
	wire [WIDTH-1:0] wire_d0_35;
	wire [WIDTH-1:0] wire_d0_36;
	wire [WIDTH-1:0] wire_d0_37;
	wire [WIDTH-1:0] wire_d0_38;
	wire [WIDTH-1:0] wire_d0_39;
	wire [WIDTH-1:0] wire_d0_40;
	wire [WIDTH-1:0] wire_d0_41;
	wire [WIDTH-1:0] wire_d0_42;
	wire [WIDTH-1:0] wire_d0_43;
	wire [WIDTH-1:0] wire_d0_44;
	wire [WIDTH-1:0] wire_d0_45;
	wire [WIDTH-1:0] wire_d0_46;
	wire [WIDTH-1:0] wire_d0_47;
	wire [WIDTH-1:0] wire_d0_48;
	wire [WIDTH-1:0] wire_d0_49;
	wire [WIDTH-1:0] wire_d0_50;
	wire [WIDTH-1:0] wire_d0_51;
	wire [WIDTH-1:0] wire_d0_52;
	wire [WIDTH-1:0] wire_d0_53;
	wire [WIDTH-1:0] wire_d0_54;
	wire [WIDTH-1:0] wire_d0_55;
	wire [WIDTH-1:0] wire_d0_56;
	wire [WIDTH-1:0] wire_d0_57;
	wire [WIDTH-1:0] wire_d0_58;
	wire [WIDTH-1:0] wire_d0_59;
	wire [WIDTH-1:0] wire_d0_60;
	wire [WIDTH-1:0] wire_d0_61;
	wire [WIDTH-1:0] wire_d0_62;
	wire [WIDTH-1:0] wire_d0_63;
	wire [WIDTH-1:0] wire_d0_64;
	wire [WIDTH-1:0] wire_d0_65;
	wire [WIDTH-1:0] wire_d0_66;
	wire [WIDTH-1:0] wire_d0_67;
	wire [WIDTH-1:0] wire_d0_68;
	wire [WIDTH-1:0] wire_d0_69;
	wire [WIDTH-1:0] wire_d0_70;
	wire [WIDTH-1:0] wire_d0_71;
	wire [WIDTH-1:0] wire_d0_72;
	wire [WIDTH-1:0] wire_d0_73;
	wire [WIDTH-1:0] wire_d0_74;
	wire [WIDTH-1:0] wire_d0_75;
	wire [WIDTH-1:0] wire_d0_76;
	wire [WIDTH-1:0] wire_d0_77;
	wire [WIDTH-1:0] wire_d0_78;
	wire [WIDTH-1:0] wire_d0_79;
	wire [WIDTH-1:0] wire_d0_80;
	wire [WIDTH-1:0] wire_d0_81;
	wire [WIDTH-1:0] wire_d0_82;
	wire [WIDTH-1:0] wire_d0_83;
	wire [WIDTH-1:0] wire_d0_84;
	wire [WIDTH-1:0] wire_d0_85;
	wire [WIDTH-1:0] wire_d0_86;
	wire [WIDTH-1:0] wire_d0_87;
	wire [WIDTH-1:0] wire_d0_88;
	wire [WIDTH-1:0] wire_d0_89;
	wire [WIDTH-1:0] wire_d0_90;
	wire [WIDTH-1:0] wire_d0_91;
	wire [WIDTH-1:0] wire_d0_92;
	wire [WIDTH-1:0] wire_d0_93;
	wire [WIDTH-1:0] wire_d0_94;
	wire [WIDTH-1:0] wire_d0_95;
	wire [WIDTH-1:0] wire_d0_96;
	wire [WIDTH-1:0] wire_d0_97;
	wire [WIDTH-1:0] wire_d0_98;
	wire [WIDTH-1:0] wire_d0_99;
	wire [WIDTH-1:0] wire_d0_100;
	wire [WIDTH-1:0] wire_d0_101;
	wire [WIDTH-1:0] wire_d0_102;
	wire [WIDTH-1:0] wire_d0_103;
	wire [WIDTH-1:0] wire_d0_104;
	wire [WIDTH-1:0] wire_d0_105;
	wire [WIDTH-1:0] wire_d0_106;
	wire [WIDTH-1:0] wire_d0_107;
	wire [WIDTH-1:0] wire_d0_108;
	wire [WIDTH-1:0] wire_d0_109;
	wire [WIDTH-1:0] wire_d0_110;
	wire [WIDTH-1:0] wire_d0_111;
	wire [WIDTH-1:0] wire_d0_112;
	wire [WIDTH-1:0] wire_d0_113;
	wire [WIDTH-1:0] wire_d0_114;
	wire [WIDTH-1:0] wire_d0_115;
	wire [WIDTH-1:0] wire_d0_116;
	wire [WIDTH-1:0] wire_d0_117;
	wire [WIDTH-1:0] wire_d0_118;
	wire [WIDTH-1:0] wire_d0_119;
	wire [WIDTH-1:0] wire_d0_120;
	wire [WIDTH-1:0] wire_d0_121;
	wire [WIDTH-1:0] wire_d0_122;
	wire [WIDTH-1:0] wire_d0_123;
	wire [WIDTH-1:0] wire_d0_124;
	wire [WIDTH-1:0] wire_d0_125;
	wire [WIDTH-1:0] wire_d0_126;
	wire [WIDTH-1:0] wire_d0_127;
	wire [WIDTH-1:0] wire_d0_128;
	wire [WIDTH-1:0] wire_d0_129;
	wire [WIDTH-1:0] wire_d0_130;
	wire [WIDTH-1:0] wire_d0_131;
	wire [WIDTH-1:0] wire_d0_132;
	wire [WIDTH-1:0] wire_d0_133;
	wire [WIDTH-1:0] wire_d0_134;
	wire [WIDTH-1:0] wire_d0_135;
	wire [WIDTH-1:0] wire_d0_136;
	wire [WIDTH-1:0] wire_d0_137;
	wire [WIDTH-1:0] wire_d0_138;
	wire [WIDTH-1:0] wire_d0_139;
	wire [WIDTH-1:0] wire_d0_140;
	wire [WIDTH-1:0] wire_d0_141;
	wire [WIDTH-1:0] wire_d0_142;
	wire [WIDTH-1:0] wire_d0_143;
	wire [WIDTH-1:0] wire_d0_144;
	wire [WIDTH-1:0] wire_d0_145;
	wire [WIDTH-1:0] wire_d0_146;
	wire [WIDTH-1:0] wire_d0_147;
	wire [WIDTH-1:0] wire_d0_148;
	wire [WIDTH-1:0] wire_d0_149;
	wire [WIDTH-1:0] wire_d0_150;
	wire [WIDTH-1:0] wire_d0_151;
	wire [WIDTH-1:0] wire_d0_152;
	wire [WIDTH-1:0] wire_d0_153;
	wire [WIDTH-1:0] wire_d0_154;
	wire [WIDTH-1:0] wire_d0_155;
	wire [WIDTH-1:0] wire_d0_156;
	wire [WIDTH-1:0] wire_d0_157;
	wire [WIDTH-1:0] wire_d0_158;
	wire [WIDTH-1:0] wire_d0_159;
	wire [WIDTH-1:0] wire_d0_160;
	wire [WIDTH-1:0] wire_d0_161;
	wire [WIDTH-1:0] wire_d0_162;
	wire [WIDTH-1:0] wire_d0_163;
	wire [WIDTH-1:0] wire_d0_164;
	wire [WIDTH-1:0] wire_d0_165;
	wire [WIDTH-1:0] wire_d0_166;
	wire [WIDTH-1:0] wire_d0_167;
	wire [WIDTH-1:0] wire_d0_168;
	wire [WIDTH-1:0] wire_d0_169;
	wire [WIDTH-1:0] wire_d0_170;
	wire [WIDTH-1:0] wire_d0_171;
	wire [WIDTH-1:0] wire_d0_172;
	wire [WIDTH-1:0] wire_d0_173;
	wire [WIDTH-1:0] wire_d0_174;
	wire [WIDTH-1:0] wire_d0_175;
	wire [WIDTH-1:0] wire_d0_176;
	wire [WIDTH-1:0] wire_d0_177;
	wire [WIDTH-1:0] wire_d0_178;
	wire [WIDTH-1:0] wire_d0_179;
	wire [WIDTH-1:0] wire_d0_180;
	wire [WIDTH-1:0] wire_d0_181;
	wire [WIDTH-1:0] wire_d0_182;
	wire [WIDTH-1:0] wire_d0_183;
	wire [WIDTH-1:0] wire_d0_184;
	wire [WIDTH-1:0] wire_d0_185;
	wire [WIDTH-1:0] wire_d0_186;
	wire [WIDTH-1:0] wire_d0_187;
	wire [WIDTH-1:0] wire_d0_188;
	wire [WIDTH-1:0] wire_d0_189;
	wire [WIDTH-1:0] wire_d0_190;
	wire [WIDTH-1:0] wire_d0_191;
	wire [WIDTH-1:0] wire_d0_192;
	wire [WIDTH-1:0] wire_d0_193;
	wire [WIDTH-1:0] wire_d0_194;
	wire [WIDTH-1:0] wire_d0_195;
	wire [WIDTH-1:0] wire_d0_196;
	wire [WIDTH-1:0] wire_d0_197;
	wire [WIDTH-1:0] wire_d0_198;
	wire [WIDTH-1:0] wire_d1_0;
	wire [WIDTH-1:0] wire_d1_1;
	wire [WIDTH-1:0] wire_d1_2;
	wire [WIDTH-1:0] wire_d1_3;
	wire [WIDTH-1:0] wire_d1_4;
	wire [WIDTH-1:0] wire_d1_5;
	wire [WIDTH-1:0] wire_d1_6;
	wire [WIDTH-1:0] wire_d1_7;
	wire [WIDTH-1:0] wire_d1_8;
	wire [WIDTH-1:0] wire_d1_9;
	wire [WIDTH-1:0] wire_d1_10;
	wire [WIDTH-1:0] wire_d1_11;
	wire [WIDTH-1:0] wire_d1_12;
	wire [WIDTH-1:0] wire_d1_13;
	wire [WIDTH-1:0] wire_d1_14;
	wire [WIDTH-1:0] wire_d1_15;
	wire [WIDTH-1:0] wire_d1_16;
	wire [WIDTH-1:0] wire_d1_17;
	wire [WIDTH-1:0] wire_d1_18;
	wire [WIDTH-1:0] wire_d1_19;
	wire [WIDTH-1:0] wire_d1_20;
	wire [WIDTH-1:0] wire_d1_21;
	wire [WIDTH-1:0] wire_d1_22;
	wire [WIDTH-1:0] wire_d1_23;
	wire [WIDTH-1:0] wire_d1_24;
	wire [WIDTH-1:0] wire_d1_25;
	wire [WIDTH-1:0] wire_d1_26;
	wire [WIDTH-1:0] wire_d1_27;
	wire [WIDTH-1:0] wire_d1_28;
	wire [WIDTH-1:0] wire_d1_29;
	wire [WIDTH-1:0] wire_d1_30;
	wire [WIDTH-1:0] wire_d1_31;
	wire [WIDTH-1:0] wire_d1_32;
	wire [WIDTH-1:0] wire_d1_33;
	wire [WIDTH-1:0] wire_d1_34;
	wire [WIDTH-1:0] wire_d1_35;
	wire [WIDTH-1:0] wire_d1_36;
	wire [WIDTH-1:0] wire_d1_37;
	wire [WIDTH-1:0] wire_d1_38;
	wire [WIDTH-1:0] wire_d1_39;
	wire [WIDTH-1:0] wire_d1_40;
	wire [WIDTH-1:0] wire_d1_41;
	wire [WIDTH-1:0] wire_d1_42;
	wire [WIDTH-1:0] wire_d1_43;
	wire [WIDTH-1:0] wire_d1_44;
	wire [WIDTH-1:0] wire_d1_45;
	wire [WIDTH-1:0] wire_d1_46;
	wire [WIDTH-1:0] wire_d1_47;
	wire [WIDTH-1:0] wire_d1_48;
	wire [WIDTH-1:0] wire_d1_49;
	wire [WIDTH-1:0] wire_d1_50;
	wire [WIDTH-1:0] wire_d1_51;
	wire [WIDTH-1:0] wire_d1_52;
	wire [WIDTH-1:0] wire_d1_53;
	wire [WIDTH-1:0] wire_d1_54;
	wire [WIDTH-1:0] wire_d1_55;
	wire [WIDTH-1:0] wire_d1_56;
	wire [WIDTH-1:0] wire_d1_57;
	wire [WIDTH-1:0] wire_d1_58;
	wire [WIDTH-1:0] wire_d1_59;
	wire [WIDTH-1:0] wire_d1_60;
	wire [WIDTH-1:0] wire_d1_61;
	wire [WIDTH-1:0] wire_d1_62;
	wire [WIDTH-1:0] wire_d1_63;
	wire [WIDTH-1:0] wire_d1_64;
	wire [WIDTH-1:0] wire_d1_65;
	wire [WIDTH-1:0] wire_d1_66;
	wire [WIDTH-1:0] wire_d1_67;
	wire [WIDTH-1:0] wire_d1_68;
	wire [WIDTH-1:0] wire_d1_69;
	wire [WIDTH-1:0] wire_d1_70;
	wire [WIDTH-1:0] wire_d1_71;
	wire [WIDTH-1:0] wire_d1_72;
	wire [WIDTH-1:0] wire_d1_73;
	wire [WIDTH-1:0] wire_d1_74;
	wire [WIDTH-1:0] wire_d1_75;
	wire [WIDTH-1:0] wire_d1_76;
	wire [WIDTH-1:0] wire_d1_77;
	wire [WIDTH-1:0] wire_d1_78;
	wire [WIDTH-1:0] wire_d1_79;
	wire [WIDTH-1:0] wire_d1_80;
	wire [WIDTH-1:0] wire_d1_81;
	wire [WIDTH-1:0] wire_d1_82;
	wire [WIDTH-1:0] wire_d1_83;
	wire [WIDTH-1:0] wire_d1_84;
	wire [WIDTH-1:0] wire_d1_85;
	wire [WIDTH-1:0] wire_d1_86;
	wire [WIDTH-1:0] wire_d1_87;
	wire [WIDTH-1:0] wire_d1_88;
	wire [WIDTH-1:0] wire_d1_89;
	wire [WIDTH-1:0] wire_d1_90;
	wire [WIDTH-1:0] wire_d1_91;
	wire [WIDTH-1:0] wire_d1_92;
	wire [WIDTH-1:0] wire_d1_93;
	wire [WIDTH-1:0] wire_d1_94;
	wire [WIDTH-1:0] wire_d1_95;
	wire [WIDTH-1:0] wire_d1_96;
	wire [WIDTH-1:0] wire_d1_97;
	wire [WIDTH-1:0] wire_d1_98;
	wire [WIDTH-1:0] wire_d1_99;
	wire [WIDTH-1:0] wire_d1_100;
	wire [WIDTH-1:0] wire_d1_101;
	wire [WIDTH-1:0] wire_d1_102;
	wire [WIDTH-1:0] wire_d1_103;
	wire [WIDTH-1:0] wire_d1_104;
	wire [WIDTH-1:0] wire_d1_105;
	wire [WIDTH-1:0] wire_d1_106;
	wire [WIDTH-1:0] wire_d1_107;
	wire [WIDTH-1:0] wire_d1_108;
	wire [WIDTH-1:0] wire_d1_109;
	wire [WIDTH-1:0] wire_d1_110;
	wire [WIDTH-1:0] wire_d1_111;
	wire [WIDTH-1:0] wire_d1_112;
	wire [WIDTH-1:0] wire_d1_113;
	wire [WIDTH-1:0] wire_d1_114;
	wire [WIDTH-1:0] wire_d1_115;
	wire [WIDTH-1:0] wire_d1_116;
	wire [WIDTH-1:0] wire_d1_117;
	wire [WIDTH-1:0] wire_d1_118;
	wire [WIDTH-1:0] wire_d1_119;
	wire [WIDTH-1:0] wire_d1_120;
	wire [WIDTH-1:0] wire_d1_121;
	wire [WIDTH-1:0] wire_d1_122;
	wire [WIDTH-1:0] wire_d1_123;
	wire [WIDTH-1:0] wire_d1_124;
	wire [WIDTH-1:0] wire_d1_125;
	wire [WIDTH-1:0] wire_d1_126;
	wire [WIDTH-1:0] wire_d1_127;
	wire [WIDTH-1:0] wire_d1_128;
	wire [WIDTH-1:0] wire_d1_129;
	wire [WIDTH-1:0] wire_d1_130;
	wire [WIDTH-1:0] wire_d1_131;
	wire [WIDTH-1:0] wire_d1_132;
	wire [WIDTH-1:0] wire_d1_133;
	wire [WIDTH-1:0] wire_d1_134;
	wire [WIDTH-1:0] wire_d1_135;
	wire [WIDTH-1:0] wire_d1_136;
	wire [WIDTH-1:0] wire_d1_137;
	wire [WIDTH-1:0] wire_d1_138;
	wire [WIDTH-1:0] wire_d1_139;
	wire [WIDTH-1:0] wire_d1_140;
	wire [WIDTH-1:0] wire_d1_141;
	wire [WIDTH-1:0] wire_d1_142;
	wire [WIDTH-1:0] wire_d1_143;
	wire [WIDTH-1:0] wire_d1_144;
	wire [WIDTH-1:0] wire_d1_145;
	wire [WIDTH-1:0] wire_d1_146;
	wire [WIDTH-1:0] wire_d1_147;
	wire [WIDTH-1:0] wire_d1_148;
	wire [WIDTH-1:0] wire_d1_149;
	wire [WIDTH-1:0] wire_d1_150;
	wire [WIDTH-1:0] wire_d1_151;
	wire [WIDTH-1:0] wire_d1_152;
	wire [WIDTH-1:0] wire_d1_153;
	wire [WIDTH-1:0] wire_d1_154;
	wire [WIDTH-1:0] wire_d1_155;
	wire [WIDTH-1:0] wire_d1_156;
	wire [WIDTH-1:0] wire_d1_157;
	wire [WIDTH-1:0] wire_d1_158;
	wire [WIDTH-1:0] wire_d1_159;
	wire [WIDTH-1:0] wire_d1_160;
	wire [WIDTH-1:0] wire_d1_161;
	wire [WIDTH-1:0] wire_d1_162;
	wire [WIDTH-1:0] wire_d1_163;
	wire [WIDTH-1:0] wire_d1_164;
	wire [WIDTH-1:0] wire_d1_165;
	wire [WIDTH-1:0] wire_d1_166;
	wire [WIDTH-1:0] wire_d1_167;
	wire [WIDTH-1:0] wire_d1_168;
	wire [WIDTH-1:0] wire_d1_169;
	wire [WIDTH-1:0] wire_d1_170;
	wire [WIDTH-1:0] wire_d1_171;
	wire [WIDTH-1:0] wire_d1_172;
	wire [WIDTH-1:0] wire_d1_173;
	wire [WIDTH-1:0] wire_d1_174;
	wire [WIDTH-1:0] wire_d1_175;
	wire [WIDTH-1:0] wire_d1_176;
	wire [WIDTH-1:0] wire_d1_177;
	wire [WIDTH-1:0] wire_d1_178;
	wire [WIDTH-1:0] wire_d1_179;
	wire [WIDTH-1:0] wire_d1_180;
	wire [WIDTH-1:0] wire_d1_181;
	wire [WIDTH-1:0] wire_d1_182;
	wire [WIDTH-1:0] wire_d1_183;
	wire [WIDTH-1:0] wire_d1_184;
	wire [WIDTH-1:0] wire_d1_185;
	wire [WIDTH-1:0] wire_d1_186;
	wire [WIDTH-1:0] wire_d1_187;
	wire [WIDTH-1:0] wire_d1_188;
	wire [WIDTH-1:0] wire_d1_189;
	wire [WIDTH-1:0] wire_d1_190;
	wire [WIDTH-1:0] wire_d1_191;
	wire [WIDTH-1:0] wire_d1_192;
	wire [WIDTH-1:0] wire_d1_193;
	wire [WIDTH-1:0] wire_d1_194;
	wire [WIDTH-1:0] wire_d1_195;
	wire [WIDTH-1:0] wire_d1_196;
	wire [WIDTH-1:0] wire_d1_197;
	wire [WIDTH-1:0] wire_d1_198;
	wire [WIDTH-1:0] wire_d2_0;
	wire [WIDTH-1:0] wire_d2_1;
	wire [WIDTH-1:0] wire_d2_2;
	wire [WIDTH-1:0] wire_d2_3;
	wire [WIDTH-1:0] wire_d2_4;
	wire [WIDTH-1:0] wire_d2_5;
	wire [WIDTH-1:0] wire_d2_6;
	wire [WIDTH-1:0] wire_d2_7;
	wire [WIDTH-1:0] wire_d2_8;
	wire [WIDTH-1:0] wire_d2_9;
	wire [WIDTH-1:0] wire_d2_10;
	wire [WIDTH-1:0] wire_d2_11;
	wire [WIDTH-1:0] wire_d2_12;
	wire [WIDTH-1:0] wire_d2_13;
	wire [WIDTH-1:0] wire_d2_14;
	wire [WIDTH-1:0] wire_d2_15;
	wire [WIDTH-1:0] wire_d2_16;
	wire [WIDTH-1:0] wire_d2_17;
	wire [WIDTH-1:0] wire_d2_18;
	wire [WIDTH-1:0] wire_d2_19;
	wire [WIDTH-1:0] wire_d2_20;
	wire [WIDTH-1:0] wire_d2_21;
	wire [WIDTH-1:0] wire_d2_22;
	wire [WIDTH-1:0] wire_d2_23;
	wire [WIDTH-1:0] wire_d2_24;
	wire [WIDTH-1:0] wire_d2_25;
	wire [WIDTH-1:0] wire_d2_26;
	wire [WIDTH-1:0] wire_d2_27;
	wire [WIDTH-1:0] wire_d2_28;
	wire [WIDTH-1:0] wire_d2_29;
	wire [WIDTH-1:0] wire_d2_30;
	wire [WIDTH-1:0] wire_d2_31;
	wire [WIDTH-1:0] wire_d2_32;
	wire [WIDTH-1:0] wire_d2_33;
	wire [WIDTH-1:0] wire_d2_34;
	wire [WIDTH-1:0] wire_d2_35;
	wire [WIDTH-1:0] wire_d2_36;
	wire [WIDTH-1:0] wire_d2_37;
	wire [WIDTH-1:0] wire_d2_38;
	wire [WIDTH-1:0] wire_d2_39;
	wire [WIDTH-1:0] wire_d2_40;
	wire [WIDTH-1:0] wire_d2_41;
	wire [WIDTH-1:0] wire_d2_42;
	wire [WIDTH-1:0] wire_d2_43;
	wire [WIDTH-1:0] wire_d2_44;
	wire [WIDTH-1:0] wire_d2_45;
	wire [WIDTH-1:0] wire_d2_46;
	wire [WIDTH-1:0] wire_d2_47;
	wire [WIDTH-1:0] wire_d2_48;
	wire [WIDTH-1:0] wire_d2_49;
	wire [WIDTH-1:0] wire_d2_50;
	wire [WIDTH-1:0] wire_d2_51;
	wire [WIDTH-1:0] wire_d2_52;
	wire [WIDTH-1:0] wire_d2_53;
	wire [WIDTH-1:0] wire_d2_54;
	wire [WIDTH-1:0] wire_d2_55;
	wire [WIDTH-1:0] wire_d2_56;
	wire [WIDTH-1:0] wire_d2_57;
	wire [WIDTH-1:0] wire_d2_58;
	wire [WIDTH-1:0] wire_d2_59;
	wire [WIDTH-1:0] wire_d2_60;
	wire [WIDTH-1:0] wire_d2_61;
	wire [WIDTH-1:0] wire_d2_62;
	wire [WIDTH-1:0] wire_d2_63;
	wire [WIDTH-1:0] wire_d2_64;
	wire [WIDTH-1:0] wire_d2_65;
	wire [WIDTH-1:0] wire_d2_66;
	wire [WIDTH-1:0] wire_d2_67;
	wire [WIDTH-1:0] wire_d2_68;
	wire [WIDTH-1:0] wire_d2_69;
	wire [WIDTH-1:0] wire_d2_70;
	wire [WIDTH-1:0] wire_d2_71;
	wire [WIDTH-1:0] wire_d2_72;
	wire [WIDTH-1:0] wire_d2_73;
	wire [WIDTH-1:0] wire_d2_74;
	wire [WIDTH-1:0] wire_d2_75;
	wire [WIDTH-1:0] wire_d2_76;
	wire [WIDTH-1:0] wire_d2_77;
	wire [WIDTH-1:0] wire_d2_78;
	wire [WIDTH-1:0] wire_d2_79;
	wire [WIDTH-1:0] wire_d2_80;
	wire [WIDTH-1:0] wire_d2_81;
	wire [WIDTH-1:0] wire_d2_82;
	wire [WIDTH-1:0] wire_d2_83;
	wire [WIDTH-1:0] wire_d2_84;
	wire [WIDTH-1:0] wire_d2_85;
	wire [WIDTH-1:0] wire_d2_86;
	wire [WIDTH-1:0] wire_d2_87;
	wire [WIDTH-1:0] wire_d2_88;
	wire [WIDTH-1:0] wire_d2_89;
	wire [WIDTH-1:0] wire_d2_90;
	wire [WIDTH-1:0] wire_d2_91;
	wire [WIDTH-1:0] wire_d2_92;
	wire [WIDTH-1:0] wire_d2_93;
	wire [WIDTH-1:0] wire_d2_94;
	wire [WIDTH-1:0] wire_d2_95;
	wire [WIDTH-1:0] wire_d2_96;
	wire [WIDTH-1:0] wire_d2_97;
	wire [WIDTH-1:0] wire_d2_98;
	wire [WIDTH-1:0] wire_d2_99;
	wire [WIDTH-1:0] wire_d2_100;
	wire [WIDTH-1:0] wire_d2_101;
	wire [WIDTH-1:0] wire_d2_102;
	wire [WIDTH-1:0] wire_d2_103;
	wire [WIDTH-1:0] wire_d2_104;
	wire [WIDTH-1:0] wire_d2_105;
	wire [WIDTH-1:0] wire_d2_106;
	wire [WIDTH-1:0] wire_d2_107;
	wire [WIDTH-1:0] wire_d2_108;
	wire [WIDTH-1:0] wire_d2_109;
	wire [WIDTH-1:0] wire_d2_110;
	wire [WIDTH-1:0] wire_d2_111;
	wire [WIDTH-1:0] wire_d2_112;
	wire [WIDTH-1:0] wire_d2_113;
	wire [WIDTH-1:0] wire_d2_114;
	wire [WIDTH-1:0] wire_d2_115;
	wire [WIDTH-1:0] wire_d2_116;
	wire [WIDTH-1:0] wire_d2_117;
	wire [WIDTH-1:0] wire_d2_118;
	wire [WIDTH-1:0] wire_d2_119;
	wire [WIDTH-1:0] wire_d2_120;
	wire [WIDTH-1:0] wire_d2_121;
	wire [WIDTH-1:0] wire_d2_122;
	wire [WIDTH-1:0] wire_d2_123;
	wire [WIDTH-1:0] wire_d2_124;
	wire [WIDTH-1:0] wire_d2_125;
	wire [WIDTH-1:0] wire_d2_126;
	wire [WIDTH-1:0] wire_d2_127;
	wire [WIDTH-1:0] wire_d2_128;
	wire [WIDTH-1:0] wire_d2_129;
	wire [WIDTH-1:0] wire_d2_130;
	wire [WIDTH-1:0] wire_d2_131;
	wire [WIDTH-1:0] wire_d2_132;
	wire [WIDTH-1:0] wire_d2_133;
	wire [WIDTH-1:0] wire_d2_134;
	wire [WIDTH-1:0] wire_d2_135;
	wire [WIDTH-1:0] wire_d2_136;
	wire [WIDTH-1:0] wire_d2_137;
	wire [WIDTH-1:0] wire_d2_138;
	wire [WIDTH-1:0] wire_d2_139;
	wire [WIDTH-1:0] wire_d2_140;
	wire [WIDTH-1:0] wire_d2_141;
	wire [WIDTH-1:0] wire_d2_142;
	wire [WIDTH-1:0] wire_d2_143;
	wire [WIDTH-1:0] wire_d2_144;
	wire [WIDTH-1:0] wire_d2_145;
	wire [WIDTH-1:0] wire_d2_146;
	wire [WIDTH-1:0] wire_d2_147;
	wire [WIDTH-1:0] wire_d2_148;
	wire [WIDTH-1:0] wire_d2_149;
	wire [WIDTH-1:0] wire_d2_150;
	wire [WIDTH-1:0] wire_d2_151;
	wire [WIDTH-1:0] wire_d2_152;
	wire [WIDTH-1:0] wire_d2_153;
	wire [WIDTH-1:0] wire_d2_154;
	wire [WIDTH-1:0] wire_d2_155;
	wire [WIDTH-1:0] wire_d2_156;
	wire [WIDTH-1:0] wire_d2_157;
	wire [WIDTH-1:0] wire_d2_158;
	wire [WIDTH-1:0] wire_d2_159;
	wire [WIDTH-1:0] wire_d2_160;
	wire [WIDTH-1:0] wire_d2_161;
	wire [WIDTH-1:0] wire_d2_162;
	wire [WIDTH-1:0] wire_d2_163;
	wire [WIDTH-1:0] wire_d2_164;
	wire [WIDTH-1:0] wire_d2_165;
	wire [WIDTH-1:0] wire_d2_166;
	wire [WIDTH-1:0] wire_d2_167;
	wire [WIDTH-1:0] wire_d2_168;
	wire [WIDTH-1:0] wire_d2_169;
	wire [WIDTH-1:0] wire_d2_170;
	wire [WIDTH-1:0] wire_d2_171;
	wire [WIDTH-1:0] wire_d2_172;
	wire [WIDTH-1:0] wire_d2_173;
	wire [WIDTH-1:0] wire_d2_174;
	wire [WIDTH-1:0] wire_d2_175;
	wire [WIDTH-1:0] wire_d2_176;
	wire [WIDTH-1:0] wire_d2_177;
	wire [WIDTH-1:0] wire_d2_178;
	wire [WIDTH-1:0] wire_d2_179;
	wire [WIDTH-1:0] wire_d2_180;
	wire [WIDTH-1:0] wire_d2_181;
	wire [WIDTH-1:0] wire_d2_182;
	wire [WIDTH-1:0] wire_d2_183;
	wire [WIDTH-1:0] wire_d2_184;
	wire [WIDTH-1:0] wire_d2_185;
	wire [WIDTH-1:0] wire_d2_186;
	wire [WIDTH-1:0] wire_d2_187;
	wire [WIDTH-1:0] wire_d2_188;
	wire [WIDTH-1:0] wire_d2_189;
	wire [WIDTH-1:0] wire_d2_190;
	wire [WIDTH-1:0] wire_d2_191;
	wire [WIDTH-1:0] wire_d2_192;
	wire [WIDTH-1:0] wire_d2_193;
	wire [WIDTH-1:0] wire_d2_194;
	wire [WIDTH-1:0] wire_d2_195;
	wire [WIDTH-1:0] wire_d2_196;
	wire [WIDTH-1:0] wire_d2_197;
	wire [WIDTH-1:0] wire_d2_198;
	wire [WIDTH-1:0] wire_d3_0;
	wire [WIDTH-1:0] wire_d3_1;
	wire [WIDTH-1:0] wire_d3_2;
	wire [WIDTH-1:0] wire_d3_3;
	wire [WIDTH-1:0] wire_d3_4;
	wire [WIDTH-1:0] wire_d3_5;
	wire [WIDTH-1:0] wire_d3_6;
	wire [WIDTH-1:0] wire_d3_7;
	wire [WIDTH-1:0] wire_d3_8;
	wire [WIDTH-1:0] wire_d3_9;
	wire [WIDTH-1:0] wire_d3_10;
	wire [WIDTH-1:0] wire_d3_11;
	wire [WIDTH-1:0] wire_d3_12;
	wire [WIDTH-1:0] wire_d3_13;
	wire [WIDTH-1:0] wire_d3_14;
	wire [WIDTH-1:0] wire_d3_15;
	wire [WIDTH-1:0] wire_d3_16;
	wire [WIDTH-1:0] wire_d3_17;
	wire [WIDTH-1:0] wire_d3_18;
	wire [WIDTH-1:0] wire_d3_19;
	wire [WIDTH-1:0] wire_d3_20;
	wire [WIDTH-1:0] wire_d3_21;
	wire [WIDTH-1:0] wire_d3_22;
	wire [WIDTH-1:0] wire_d3_23;
	wire [WIDTH-1:0] wire_d3_24;
	wire [WIDTH-1:0] wire_d3_25;
	wire [WIDTH-1:0] wire_d3_26;
	wire [WIDTH-1:0] wire_d3_27;
	wire [WIDTH-1:0] wire_d3_28;
	wire [WIDTH-1:0] wire_d3_29;
	wire [WIDTH-1:0] wire_d3_30;
	wire [WIDTH-1:0] wire_d3_31;
	wire [WIDTH-1:0] wire_d3_32;
	wire [WIDTH-1:0] wire_d3_33;
	wire [WIDTH-1:0] wire_d3_34;
	wire [WIDTH-1:0] wire_d3_35;
	wire [WIDTH-1:0] wire_d3_36;
	wire [WIDTH-1:0] wire_d3_37;
	wire [WIDTH-1:0] wire_d3_38;
	wire [WIDTH-1:0] wire_d3_39;
	wire [WIDTH-1:0] wire_d3_40;
	wire [WIDTH-1:0] wire_d3_41;
	wire [WIDTH-1:0] wire_d3_42;
	wire [WIDTH-1:0] wire_d3_43;
	wire [WIDTH-1:0] wire_d3_44;
	wire [WIDTH-1:0] wire_d3_45;
	wire [WIDTH-1:0] wire_d3_46;
	wire [WIDTH-1:0] wire_d3_47;
	wire [WIDTH-1:0] wire_d3_48;
	wire [WIDTH-1:0] wire_d3_49;
	wire [WIDTH-1:0] wire_d3_50;
	wire [WIDTH-1:0] wire_d3_51;
	wire [WIDTH-1:0] wire_d3_52;
	wire [WIDTH-1:0] wire_d3_53;
	wire [WIDTH-1:0] wire_d3_54;
	wire [WIDTH-1:0] wire_d3_55;
	wire [WIDTH-1:0] wire_d3_56;
	wire [WIDTH-1:0] wire_d3_57;
	wire [WIDTH-1:0] wire_d3_58;
	wire [WIDTH-1:0] wire_d3_59;
	wire [WIDTH-1:0] wire_d3_60;
	wire [WIDTH-1:0] wire_d3_61;
	wire [WIDTH-1:0] wire_d3_62;
	wire [WIDTH-1:0] wire_d3_63;
	wire [WIDTH-1:0] wire_d3_64;
	wire [WIDTH-1:0] wire_d3_65;
	wire [WIDTH-1:0] wire_d3_66;
	wire [WIDTH-1:0] wire_d3_67;
	wire [WIDTH-1:0] wire_d3_68;
	wire [WIDTH-1:0] wire_d3_69;
	wire [WIDTH-1:0] wire_d3_70;
	wire [WIDTH-1:0] wire_d3_71;
	wire [WIDTH-1:0] wire_d3_72;
	wire [WIDTH-1:0] wire_d3_73;
	wire [WIDTH-1:0] wire_d3_74;
	wire [WIDTH-1:0] wire_d3_75;
	wire [WIDTH-1:0] wire_d3_76;
	wire [WIDTH-1:0] wire_d3_77;
	wire [WIDTH-1:0] wire_d3_78;
	wire [WIDTH-1:0] wire_d3_79;
	wire [WIDTH-1:0] wire_d3_80;
	wire [WIDTH-1:0] wire_d3_81;
	wire [WIDTH-1:0] wire_d3_82;
	wire [WIDTH-1:0] wire_d3_83;
	wire [WIDTH-1:0] wire_d3_84;
	wire [WIDTH-1:0] wire_d3_85;
	wire [WIDTH-1:0] wire_d3_86;
	wire [WIDTH-1:0] wire_d3_87;
	wire [WIDTH-1:0] wire_d3_88;
	wire [WIDTH-1:0] wire_d3_89;
	wire [WIDTH-1:0] wire_d3_90;
	wire [WIDTH-1:0] wire_d3_91;
	wire [WIDTH-1:0] wire_d3_92;
	wire [WIDTH-1:0] wire_d3_93;
	wire [WIDTH-1:0] wire_d3_94;
	wire [WIDTH-1:0] wire_d3_95;
	wire [WIDTH-1:0] wire_d3_96;
	wire [WIDTH-1:0] wire_d3_97;
	wire [WIDTH-1:0] wire_d3_98;
	wire [WIDTH-1:0] wire_d3_99;
	wire [WIDTH-1:0] wire_d3_100;
	wire [WIDTH-1:0] wire_d3_101;
	wire [WIDTH-1:0] wire_d3_102;
	wire [WIDTH-1:0] wire_d3_103;
	wire [WIDTH-1:0] wire_d3_104;
	wire [WIDTH-1:0] wire_d3_105;
	wire [WIDTH-1:0] wire_d3_106;
	wire [WIDTH-1:0] wire_d3_107;
	wire [WIDTH-1:0] wire_d3_108;
	wire [WIDTH-1:0] wire_d3_109;
	wire [WIDTH-1:0] wire_d3_110;
	wire [WIDTH-1:0] wire_d3_111;
	wire [WIDTH-1:0] wire_d3_112;
	wire [WIDTH-1:0] wire_d3_113;
	wire [WIDTH-1:0] wire_d3_114;
	wire [WIDTH-1:0] wire_d3_115;
	wire [WIDTH-1:0] wire_d3_116;
	wire [WIDTH-1:0] wire_d3_117;
	wire [WIDTH-1:0] wire_d3_118;
	wire [WIDTH-1:0] wire_d3_119;
	wire [WIDTH-1:0] wire_d3_120;
	wire [WIDTH-1:0] wire_d3_121;
	wire [WIDTH-1:0] wire_d3_122;
	wire [WIDTH-1:0] wire_d3_123;
	wire [WIDTH-1:0] wire_d3_124;
	wire [WIDTH-1:0] wire_d3_125;
	wire [WIDTH-1:0] wire_d3_126;
	wire [WIDTH-1:0] wire_d3_127;
	wire [WIDTH-1:0] wire_d3_128;
	wire [WIDTH-1:0] wire_d3_129;
	wire [WIDTH-1:0] wire_d3_130;
	wire [WIDTH-1:0] wire_d3_131;
	wire [WIDTH-1:0] wire_d3_132;
	wire [WIDTH-1:0] wire_d3_133;
	wire [WIDTH-1:0] wire_d3_134;
	wire [WIDTH-1:0] wire_d3_135;
	wire [WIDTH-1:0] wire_d3_136;
	wire [WIDTH-1:0] wire_d3_137;
	wire [WIDTH-1:0] wire_d3_138;
	wire [WIDTH-1:0] wire_d3_139;
	wire [WIDTH-1:0] wire_d3_140;
	wire [WIDTH-1:0] wire_d3_141;
	wire [WIDTH-1:0] wire_d3_142;
	wire [WIDTH-1:0] wire_d3_143;
	wire [WIDTH-1:0] wire_d3_144;
	wire [WIDTH-1:0] wire_d3_145;
	wire [WIDTH-1:0] wire_d3_146;
	wire [WIDTH-1:0] wire_d3_147;
	wire [WIDTH-1:0] wire_d3_148;
	wire [WIDTH-1:0] wire_d3_149;
	wire [WIDTH-1:0] wire_d3_150;
	wire [WIDTH-1:0] wire_d3_151;
	wire [WIDTH-1:0] wire_d3_152;
	wire [WIDTH-1:0] wire_d3_153;
	wire [WIDTH-1:0] wire_d3_154;
	wire [WIDTH-1:0] wire_d3_155;
	wire [WIDTH-1:0] wire_d3_156;
	wire [WIDTH-1:0] wire_d3_157;
	wire [WIDTH-1:0] wire_d3_158;
	wire [WIDTH-1:0] wire_d3_159;
	wire [WIDTH-1:0] wire_d3_160;
	wire [WIDTH-1:0] wire_d3_161;
	wire [WIDTH-1:0] wire_d3_162;
	wire [WIDTH-1:0] wire_d3_163;
	wire [WIDTH-1:0] wire_d3_164;
	wire [WIDTH-1:0] wire_d3_165;
	wire [WIDTH-1:0] wire_d3_166;
	wire [WIDTH-1:0] wire_d3_167;
	wire [WIDTH-1:0] wire_d3_168;
	wire [WIDTH-1:0] wire_d3_169;
	wire [WIDTH-1:0] wire_d3_170;
	wire [WIDTH-1:0] wire_d3_171;
	wire [WIDTH-1:0] wire_d3_172;
	wire [WIDTH-1:0] wire_d3_173;
	wire [WIDTH-1:0] wire_d3_174;
	wire [WIDTH-1:0] wire_d3_175;
	wire [WIDTH-1:0] wire_d3_176;
	wire [WIDTH-1:0] wire_d3_177;
	wire [WIDTH-1:0] wire_d3_178;
	wire [WIDTH-1:0] wire_d3_179;
	wire [WIDTH-1:0] wire_d3_180;
	wire [WIDTH-1:0] wire_d3_181;
	wire [WIDTH-1:0] wire_d3_182;
	wire [WIDTH-1:0] wire_d3_183;
	wire [WIDTH-1:0] wire_d3_184;
	wire [WIDTH-1:0] wire_d3_185;
	wire [WIDTH-1:0] wire_d3_186;
	wire [WIDTH-1:0] wire_d3_187;
	wire [WIDTH-1:0] wire_d3_188;
	wire [WIDTH-1:0] wire_d3_189;
	wire [WIDTH-1:0] wire_d3_190;
	wire [WIDTH-1:0] wire_d3_191;
	wire [WIDTH-1:0] wire_d3_192;
	wire [WIDTH-1:0] wire_d3_193;
	wire [WIDTH-1:0] wire_d3_194;
	wire [WIDTH-1:0] wire_d3_195;
	wire [WIDTH-1:0] wire_d3_196;
	wire [WIDTH-1:0] wire_d3_197;
	wire [WIDTH-1:0] wire_d3_198;
	wire [WIDTH-1:0] wire_d4_0;
	wire [WIDTH-1:0] wire_d4_1;
	wire [WIDTH-1:0] wire_d4_2;
	wire [WIDTH-1:0] wire_d4_3;
	wire [WIDTH-1:0] wire_d4_4;
	wire [WIDTH-1:0] wire_d4_5;
	wire [WIDTH-1:0] wire_d4_6;
	wire [WIDTH-1:0] wire_d4_7;
	wire [WIDTH-1:0] wire_d4_8;
	wire [WIDTH-1:0] wire_d4_9;
	wire [WIDTH-1:0] wire_d4_10;
	wire [WIDTH-1:0] wire_d4_11;
	wire [WIDTH-1:0] wire_d4_12;
	wire [WIDTH-1:0] wire_d4_13;
	wire [WIDTH-1:0] wire_d4_14;
	wire [WIDTH-1:0] wire_d4_15;
	wire [WIDTH-1:0] wire_d4_16;
	wire [WIDTH-1:0] wire_d4_17;
	wire [WIDTH-1:0] wire_d4_18;
	wire [WIDTH-1:0] wire_d4_19;
	wire [WIDTH-1:0] wire_d4_20;
	wire [WIDTH-1:0] wire_d4_21;
	wire [WIDTH-1:0] wire_d4_22;
	wire [WIDTH-1:0] wire_d4_23;
	wire [WIDTH-1:0] wire_d4_24;
	wire [WIDTH-1:0] wire_d4_25;
	wire [WIDTH-1:0] wire_d4_26;
	wire [WIDTH-1:0] wire_d4_27;
	wire [WIDTH-1:0] wire_d4_28;
	wire [WIDTH-1:0] wire_d4_29;
	wire [WIDTH-1:0] wire_d4_30;
	wire [WIDTH-1:0] wire_d4_31;
	wire [WIDTH-1:0] wire_d4_32;
	wire [WIDTH-1:0] wire_d4_33;
	wire [WIDTH-1:0] wire_d4_34;
	wire [WIDTH-1:0] wire_d4_35;
	wire [WIDTH-1:0] wire_d4_36;
	wire [WIDTH-1:0] wire_d4_37;
	wire [WIDTH-1:0] wire_d4_38;
	wire [WIDTH-1:0] wire_d4_39;
	wire [WIDTH-1:0] wire_d4_40;
	wire [WIDTH-1:0] wire_d4_41;
	wire [WIDTH-1:0] wire_d4_42;
	wire [WIDTH-1:0] wire_d4_43;
	wire [WIDTH-1:0] wire_d4_44;
	wire [WIDTH-1:0] wire_d4_45;
	wire [WIDTH-1:0] wire_d4_46;
	wire [WIDTH-1:0] wire_d4_47;
	wire [WIDTH-1:0] wire_d4_48;
	wire [WIDTH-1:0] wire_d4_49;
	wire [WIDTH-1:0] wire_d4_50;
	wire [WIDTH-1:0] wire_d4_51;
	wire [WIDTH-1:0] wire_d4_52;
	wire [WIDTH-1:0] wire_d4_53;
	wire [WIDTH-1:0] wire_d4_54;
	wire [WIDTH-1:0] wire_d4_55;
	wire [WIDTH-1:0] wire_d4_56;
	wire [WIDTH-1:0] wire_d4_57;
	wire [WIDTH-1:0] wire_d4_58;
	wire [WIDTH-1:0] wire_d4_59;
	wire [WIDTH-1:0] wire_d4_60;
	wire [WIDTH-1:0] wire_d4_61;
	wire [WIDTH-1:0] wire_d4_62;
	wire [WIDTH-1:0] wire_d4_63;
	wire [WIDTH-1:0] wire_d4_64;
	wire [WIDTH-1:0] wire_d4_65;
	wire [WIDTH-1:0] wire_d4_66;
	wire [WIDTH-1:0] wire_d4_67;
	wire [WIDTH-1:0] wire_d4_68;
	wire [WIDTH-1:0] wire_d4_69;
	wire [WIDTH-1:0] wire_d4_70;
	wire [WIDTH-1:0] wire_d4_71;
	wire [WIDTH-1:0] wire_d4_72;
	wire [WIDTH-1:0] wire_d4_73;
	wire [WIDTH-1:0] wire_d4_74;
	wire [WIDTH-1:0] wire_d4_75;
	wire [WIDTH-1:0] wire_d4_76;
	wire [WIDTH-1:0] wire_d4_77;
	wire [WIDTH-1:0] wire_d4_78;
	wire [WIDTH-1:0] wire_d4_79;
	wire [WIDTH-1:0] wire_d4_80;
	wire [WIDTH-1:0] wire_d4_81;
	wire [WIDTH-1:0] wire_d4_82;
	wire [WIDTH-1:0] wire_d4_83;
	wire [WIDTH-1:0] wire_d4_84;
	wire [WIDTH-1:0] wire_d4_85;
	wire [WIDTH-1:0] wire_d4_86;
	wire [WIDTH-1:0] wire_d4_87;
	wire [WIDTH-1:0] wire_d4_88;
	wire [WIDTH-1:0] wire_d4_89;
	wire [WIDTH-1:0] wire_d4_90;
	wire [WIDTH-1:0] wire_d4_91;
	wire [WIDTH-1:0] wire_d4_92;
	wire [WIDTH-1:0] wire_d4_93;
	wire [WIDTH-1:0] wire_d4_94;
	wire [WIDTH-1:0] wire_d4_95;
	wire [WIDTH-1:0] wire_d4_96;
	wire [WIDTH-1:0] wire_d4_97;
	wire [WIDTH-1:0] wire_d4_98;
	wire [WIDTH-1:0] wire_d4_99;
	wire [WIDTH-1:0] wire_d4_100;
	wire [WIDTH-1:0] wire_d4_101;
	wire [WIDTH-1:0] wire_d4_102;
	wire [WIDTH-1:0] wire_d4_103;
	wire [WIDTH-1:0] wire_d4_104;
	wire [WIDTH-1:0] wire_d4_105;
	wire [WIDTH-1:0] wire_d4_106;
	wire [WIDTH-1:0] wire_d4_107;
	wire [WIDTH-1:0] wire_d4_108;
	wire [WIDTH-1:0] wire_d4_109;
	wire [WIDTH-1:0] wire_d4_110;
	wire [WIDTH-1:0] wire_d4_111;
	wire [WIDTH-1:0] wire_d4_112;
	wire [WIDTH-1:0] wire_d4_113;
	wire [WIDTH-1:0] wire_d4_114;
	wire [WIDTH-1:0] wire_d4_115;
	wire [WIDTH-1:0] wire_d4_116;
	wire [WIDTH-1:0] wire_d4_117;
	wire [WIDTH-1:0] wire_d4_118;
	wire [WIDTH-1:0] wire_d4_119;
	wire [WIDTH-1:0] wire_d4_120;
	wire [WIDTH-1:0] wire_d4_121;
	wire [WIDTH-1:0] wire_d4_122;
	wire [WIDTH-1:0] wire_d4_123;
	wire [WIDTH-1:0] wire_d4_124;
	wire [WIDTH-1:0] wire_d4_125;
	wire [WIDTH-1:0] wire_d4_126;
	wire [WIDTH-1:0] wire_d4_127;
	wire [WIDTH-1:0] wire_d4_128;
	wire [WIDTH-1:0] wire_d4_129;
	wire [WIDTH-1:0] wire_d4_130;
	wire [WIDTH-1:0] wire_d4_131;
	wire [WIDTH-1:0] wire_d4_132;
	wire [WIDTH-1:0] wire_d4_133;
	wire [WIDTH-1:0] wire_d4_134;
	wire [WIDTH-1:0] wire_d4_135;
	wire [WIDTH-1:0] wire_d4_136;
	wire [WIDTH-1:0] wire_d4_137;
	wire [WIDTH-1:0] wire_d4_138;
	wire [WIDTH-1:0] wire_d4_139;
	wire [WIDTH-1:0] wire_d4_140;
	wire [WIDTH-1:0] wire_d4_141;
	wire [WIDTH-1:0] wire_d4_142;
	wire [WIDTH-1:0] wire_d4_143;
	wire [WIDTH-1:0] wire_d4_144;
	wire [WIDTH-1:0] wire_d4_145;
	wire [WIDTH-1:0] wire_d4_146;
	wire [WIDTH-1:0] wire_d4_147;
	wire [WIDTH-1:0] wire_d4_148;
	wire [WIDTH-1:0] wire_d4_149;
	wire [WIDTH-1:0] wire_d4_150;
	wire [WIDTH-1:0] wire_d4_151;
	wire [WIDTH-1:0] wire_d4_152;
	wire [WIDTH-1:0] wire_d4_153;
	wire [WIDTH-1:0] wire_d4_154;
	wire [WIDTH-1:0] wire_d4_155;
	wire [WIDTH-1:0] wire_d4_156;
	wire [WIDTH-1:0] wire_d4_157;
	wire [WIDTH-1:0] wire_d4_158;
	wire [WIDTH-1:0] wire_d4_159;
	wire [WIDTH-1:0] wire_d4_160;
	wire [WIDTH-1:0] wire_d4_161;
	wire [WIDTH-1:0] wire_d4_162;
	wire [WIDTH-1:0] wire_d4_163;
	wire [WIDTH-1:0] wire_d4_164;
	wire [WIDTH-1:0] wire_d4_165;
	wire [WIDTH-1:0] wire_d4_166;
	wire [WIDTH-1:0] wire_d4_167;
	wire [WIDTH-1:0] wire_d4_168;
	wire [WIDTH-1:0] wire_d4_169;
	wire [WIDTH-1:0] wire_d4_170;
	wire [WIDTH-1:0] wire_d4_171;
	wire [WIDTH-1:0] wire_d4_172;
	wire [WIDTH-1:0] wire_d4_173;
	wire [WIDTH-1:0] wire_d4_174;
	wire [WIDTH-1:0] wire_d4_175;
	wire [WIDTH-1:0] wire_d4_176;
	wire [WIDTH-1:0] wire_d4_177;
	wire [WIDTH-1:0] wire_d4_178;
	wire [WIDTH-1:0] wire_d4_179;
	wire [WIDTH-1:0] wire_d4_180;
	wire [WIDTH-1:0] wire_d4_181;
	wire [WIDTH-1:0] wire_d4_182;
	wire [WIDTH-1:0] wire_d4_183;
	wire [WIDTH-1:0] wire_d4_184;
	wire [WIDTH-1:0] wire_d4_185;
	wire [WIDTH-1:0] wire_d4_186;
	wire [WIDTH-1:0] wire_d4_187;
	wire [WIDTH-1:0] wire_d4_188;
	wire [WIDTH-1:0] wire_d4_189;
	wire [WIDTH-1:0] wire_d4_190;
	wire [WIDTH-1:0] wire_d4_191;
	wire [WIDTH-1:0] wire_d4_192;
	wire [WIDTH-1:0] wire_d4_193;
	wire [WIDTH-1:0] wire_d4_194;
	wire [WIDTH-1:0] wire_d4_195;
	wire [WIDTH-1:0] wire_d4_196;
	wire [WIDTH-1:0] wire_d4_197;
	wire [WIDTH-1:0] wire_d4_198;
	wire [WIDTH-1:0] wire_d5_0;
	wire [WIDTH-1:0] wire_d5_1;
	wire [WIDTH-1:0] wire_d5_2;
	wire [WIDTH-1:0] wire_d5_3;
	wire [WIDTH-1:0] wire_d5_4;
	wire [WIDTH-1:0] wire_d5_5;
	wire [WIDTH-1:0] wire_d5_6;
	wire [WIDTH-1:0] wire_d5_7;
	wire [WIDTH-1:0] wire_d5_8;
	wire [WIDTH-1:0] wire_d5_9;
	wire [WIDTH-1:0] wire_d5_10;
	wire [WIDTH-1:0] wire_d5_11;
	wire [WIDTH-1:0] wire_d5_12;
	wire [WIDTH-1:0] wire_d5_13;
	wire [WIDTH-1:0] wire_d5_14;
	wire [WIDTH-1:0] wire_d5_15;
	wire [WIDTH-1:0] wire_d5_16;
	wire [WIDTH-1:0] wire_d5_17;
	wire [WIDTH-1:0] wire_d5_18;
	wire [WIDTH-1:0] wire_d5_19;
	wire [WIDTH-1:0] wire_d5_20;
	wire [WIDTH-1:0] wire_d5_21;
	wire [WIDTH-1:0] wire_d5_22;
	wire [WIDTH-1:0] wire_d5_23;
	wire [WIDTH-1:0] wire_d5_24;
	wire [WIDTH-1:0] wire_d5_25;
	wire [WIDTH-1:0] wire_d5_26;
	wire [WIDTH-1:0] wire_d5_27;
	wire [WIDTH-1:0] wire_d5_28;
	wire [WIDTH-1:0] wire_d5_29;
	wire [WIDTH-1:0] wire_d5_30;
	wire [WIDTH-1:0] wire_d5_31;
	wire [WIDTH-1:0] wire_d5_32;
	wire [WIDTH-1:0] wire_d5_33;
	wire [WIDTH-1:0] wire_d5_34;
	wire [WIDTH-1:0] wire_d5_35;
	wire [WIDTH-1:0] wire_d5_36;
	wire [WIDTH-1:0] wire_d5_37;
	wire [WIDTH-1:0] wire_d5_38;
	wire [WIDTH-1:0] wire_d5_39;
	wire [WIDTH-1:0] wire_d5_40;
	wire [WIDTH-1:0] wire_d5_41;
	wire [WIDTH-1:0] wire_d5_42;
	wire [WIDTH-1:0] wire_d5_43;
	wire [WIDTH-1:0] wire_d5_44;
	wire [WIDTH-1:0] wire_d5_45;
	wire [WIDTH-1:0] wire_d5_46;
	wire [WIDTH-1:0] wire_d5_47;
	wire [WIDTH-1:0] wire_d5_48;
	wire [WIDTH-1:0] wire_d5_49;
	wire [WIDTH-1:0] wire_d5_50;
	wire [WIDTH-1:0] wire_d5_51;
	wire [WIDTH-1:0] wire_d5_52;
	wire [WIDTH-1:0] wire_d5_53;
	wire [WIDTH-1:0] wire_d5_54;
	wire [WIDTH-1:0] wire_d5_55;
	wire [WIDTH-1:0] wire_d5_56;
	wire [WIDTH-1:0] wire_d5_57;
	wire [WIDTH-1:0] wire_d5_58;
	wire [WIDTH-1:0] wire_d5_59;
	wire [WIDTH-1:0] wire_d5_60;
	wire [WIDTH-1:0] wire_d5_61;
	wire [WIDTH-1:0] wire_d5_62;
	wire [WIDTH-1:0] wire_d5_63;
	wire [WIDTH-1:0] wire_d5_64;
	wire [WIDTH-1:0] wire_d5_65;
	wire [WIDTH-1:0] wire_d5_66;
	wire [WIDTH-1:0] wire_d5_67;
	wire [WIDTH-1:0] wire_d5_68;
	wire [WIDTH-1:0] wire_d5_69;
	wire [WIDTH-1:0] wire_d5_70;
	wire [WIDTH-1:0] wire_d5_71;
	wire [WIDTH-1:0] wire_d5_72;
	wire [WIDTH-1:0] wire_d5_73;
	wire [WIDTH-1:0] wire_d5_74;
	wire [WIDTH-1:0] wire_d5_75;
	wire [WIDTH-1:0] wire_d5_76;
	wire [WIDTH-1:0] wire_d5_77;
	wire [WIDTH-1:0] wire_d5_78;
	wire [WIDTH-1:0] wire_d5_79;
	wire [WIDTH-1:0] wire_d5_80;
	wire [WIDTH-1:0] wire_d5_81;
	wire [WIDTH-1:0] wire_d5_82;
	wire [WIDTH-1:0] wire_d5_83;
	wire [WIDTH-1:0] wire_d5_84;
	wire [WIDTH-1:0] wire_d5_85;
	wire [WIDTH-1:0] wire_d5_86;
	wire [WIDTH-1:0] wire_d5_87;
	wire [WIDTH-1:0] wire_d5_88;
	wire [WIDTH-1:0] wire_d5_89;
	wire [WIDTH-1:0] wire_d5_90;
	wire [WIDTH-1:0] wire_d5_91;
	wire [WIDTH-1:0] wire_d5_92;
	wire [WIDTH-1:0] wire_d5_93;
	wire [WIDTH-1:0] wire_d5_94;
	wire [WIDTH-1:0] wire_d5_95;
	wire [WIDTH-1:0] wire_d5_96;
	wire [WIDTH-1:0] wire_d5_97;
	wire [WIDTH-1:0] wire_d5_98;
	wire [WIDTH-1:0] wire_d5_99;
	wire [WIDTH-1:0] wire_d5_100;
	wire [WIDTH-1:0] wire_d5_101;
	wire [WIDTH-1:0] wire_d5_102;
	wire [WIDTH-1:0] wire_d5_103;
	wire [WIDTH-1:0] wire_d5_104;
	wire [WIDTH-1:0] wire_d5_105;
	wire [WIDTH-1:0] wire_d5_106;
	wire [WIDTH-1:0] wire_d5_107;
	wire [WIDTH-1:0] wire_d5_108;
	wire [WIDTH-1:0] wire_d5_109;
	wire [WIDTH-1:0] wire_d5_110;
	wire [WIDTH-1:0] wire_d5_111;
	wire [WIDTH-1:0] wire_d5_112;
	wire [WIDTH-1:0] wire_d5_113;
	wire [WIDTH-1:0] wire_d5_114;
	wire [WIDTH-1:0] wire_d5_115;
	wire [WIDTH-1:0] wire_d5_116;
	wire [WIDTH-1:0] wire_d5_117;
	wire [WIDTH-1:0] wire_d5_118;
	wire [WIDTH-1:0] wire_d5_119;
	wire [WIDTH-1:0] wire_d5_120;
	wire [WIDTH-1:0] wire_d5_121;
	wire [WIDTH-1:0] wire_d5_122;
	wire [WIDTH-1:0] wire_d5_123;
	wire [WIDTH-1:0] wire_d5_124;
	wire [WIDTH-1:0] wire_d5_125;
	wire [WIDTH-1:0] wire_d5_126;
	wire [WIDTH-1:0] wire_d5_127;
	wire [WIDTH-1:0] wire_d5_128;
	wire [WIDTH-1:0] wire_d5_129;
	wire [WIDTH-1:0] wire_d5_130;
	wire [WIDTH-1:0] wire_d5_131;
	wire [WIDTH-1:0] wire_d5_132;
	wire [WIDTH-1:0] wire_d5_133;
	wire [WIDTH-1:0] wire_d5_134;
	wire [WIDTH-1:0] wire_d5_135;
	wire [WIDTH-1:0] wire_d5_136;
	wire [WIDTH-1:0] wire_d5_137;
	wire [WIDTH-1:0] wire_d5_138;
	wire [WIDTH-1:0] wire_d5_139;
	wire [WIDTH-1:0] wire_d5_140;
	wire [WIDTH-1:0] wire_d5_141;
	wire [WIDTH-1:0] wire_d5_142;
	wire [WIDTH-1:0] wire_d5_143;
	wire [WIDTH-1:0] wire_d5_144;
	wire [WIDTH-1:0] wire_d5_145;
	wire [WIDTH-1:0] wire_d5_146;
	wire [WIDTH-1:0] wire_d5_147;
	wire [WIDTH-1:0] wire_d5_148;
	wire [WIDTH-1:0] wire_d5_149;
	wire [WIDTH-1:0] wire_d5_150;
	wire [WIDTH-1:0] wire_d5_151;
	wire [WIDTH-1:0] wire_d5_152;
	wire [WIDTH-1:0] wire_d5_153;
	wire [WIDTH-1:0] wire_d5_154;
	wire [WIDTH-1:0] wire_d5_155;
	wire [WIDTH-1:0] wire_d5_156;
	wire [WIDTH-1:0] wire_d5_157;
	wire [WIDTH-1:0] wire_d5_158;
	wire [WIDTH-1:0] wire_d5_159;
	wire [WIDTH-1:0] wire_d5_160;
	wire [WIDTH-1:0] wire_d5_161;
	wire [WIDTH-1:0] wire_d5_162;
	wire [WIDTH-1:0] wire_d5_163;
	wire [WIDTH-1:0] wire_d5_164;
	wire [WIDTH-1:0] wire_d5_165;
	wire [WIDTH-1:0] wire_d5_166;
	wire [WIDTH-1:0] wire_d5_167;
	wire [WIDTH-1:0] wire_d5_168;
	wire [WIDTH-1:0] wire_d5_169;
	wire [WIDTH-1:0] wire_d5_170;
	wire [WIDTH-1:0] wire_d5_171;
	wire [WIDTH-1:0] wire_d5_172;
	wire [WIDTH-1:0] wire_d5_173;
	wire [WIDTH-1:0] wire_d5_174;
	wire [WIDTH-1:0] wire_d5_175;
	wire [WIDTH-1:0] wire_d5_176;
	wire [WIDTH-1:0] wire_d5_177;
	wire [WIDTH-1:0] wire_d5_178;
	wire [WIDTH-1:0] wire_d5_179;
	wire [WIDTH-1:0] wire_d5_180;
	wire [WIDTH-1:0] wire_d5_181;
	wire [WIDTH-1:0] wire_d5_182;
	wire [WIDTH-1:0] wire_d5_183;
	wire [WIDTH-1:0] wire_d5_184;
	wire [WIDTH-1:0] wire_d5_185;
	wire [WIDTH-1:0] wire_d5_186;
	wire [WIDTH-1:0] wire_d5_187;
	wire [WIDTH-1:0] wire_d5_188;
	wire [WIDTH-1:0] wire_d5_189;
	wire [WIDTH-1:0] wire_d5_190;
	wire [WIDTH-1:0] wire_d5_191;
	wire [WIDTH-1:0] wire_d5_192;
	wire [WIDTH-1:0] wire_d5_193;
	wire [WIDTH-1:0] wire_d5_194;
	wire [WIDTH-1:0] wire_d5_195;
	wire [WIDTH-1:0] wire_d5_196;
	wire [WIDTH-1:0] wire_d5_197;
	wire [WIDTH-1:0] wire_d5_198;
	wire [WIDTH-1:0] wire_d6_0;
	wire [WIDTH-1:0] wire_d6_1;
	wire [WIDTH-1:0] wire_d6_2;
	wire [WIDTH-1:0] wire_d6_3;
	wire [WIDTH-1:0] wire_d6_4;
	wire [WIDTH-1:0] wire_d6_5;
	wire [WIDTH-1:0] wire_d6_6;
	wire [WIDTH-1:0] wire_d6_7;
	wire [WIDTH-1:0] wire_d6_8;
	wire [WIDTH-1:0] wire_d6_9;
	wire [WIDTH-1:0] wire_d6_10;
	wire [WIDTH-1:0] wire_d6_11;
	wire [WIDTH-1:0] wire_d6_12;
	wire [WIDTH-1:0] wire_d6_13;
	wire [WIDTH-1:0] wire_d6_14;
	wire [WIDTH-1:0] wire_d6_15;
	wire [WIDTH-1:0] wire_d6_16;
	wire [WIDTH-1:0] wire_d6_17;
	wire [WIDTH-1:0] wire_d6_18;
	wire [WIDTH-1:0] wire_d6_19;
	wire [WIDTH-1:0] wire_d6_20;
	wire [WIDTH-1:0] wire_d6_21;
	wire [WIDTH-1:0] wire_d6_22;
	wire [WIDTH-1:0] wire_d6_23;
	wire [WIDTH-1:0] wire_d6_24;
	wire [WIDTH-1:0] wire_d6_25;
	wire [WIDTH-1:0] wire_d6_26;
	wire [WIDTH-1:0] wire_d6_27;
	wire [WIDTH-1:0] wire_d6_28;
	wire [WIDTH-1:0] wire_d6_29;
	wire [WIDTH-1:0] wire_d6_30;
	wire [WIDTH-1:0] wire_d6_31;
	wire [WIDTH-1:0] wire_d6_32;
	wire [WIDTH-1:0] wire_d6_33;
	wire [WIDTH-1:0] wire_d6_34;
	wire [WIDTH-1:0] wire_d6_35;
	wire [WIDTH-1:0] wire_d6_36;
	wire [WIDTH-1:0] wire_d6_37;
	wire [WIDTH-1:0] wire_d6_38;
	wire [WIDTH-1:0] wire_d6_39;
	wire [WIDTH-1:0] wire_d6_40;
	wire [WIDTH-1:0] wire_d6_41;
	wire [WIDTH-1:0] wire_d6_42;
	wire [WIDTH-1:0] wire_d6_43;
	wire [WIDTH-1:0] wire_d6_44;
	wire [WIDTH-1:0] wire_d6_45;
	wire [WIDTH-1:0] wire_d6_46;
	wire [WIDTH-1:0] wire_d6_47;
	wire [WIDTH-1:0] wire_d6_48;
	wire [WIDTH-1:0] wire_d6_49;
	wire [WIDTH-1:0] wire_d6_50;
	wire [WIDTH-1:0] wire_d6_51;
	wire [WIDTH-1:0] wire_d6_52;
	wire [WIDTH-1:0] wire_d6_53;
	wire [WIDTH-1:0] wire_d6_54;
	wire [WIDTH-1:0] wire_d6_55;
	wire [WIDTH-1:0] wire_d6_56;
	wire [WIDTH-1:0] wire_d6_57;
	wire [WIDTH-1:0] wire_d6_58;
	wire [WIDTH-1:0] wire_d6_59;
	wire [WIDTH-1:0] wire_d6_60;
	wire [WIDTH-1:0] wire_d6_61;
	wire [WIDTH-1:0] wire_d6_62;
	wire [WIDTH-1:0] wire_d6_63;
	wire [WIDTH-1:0] wire_d6_64;
	wire [WIDTH-1:0] wire_d6_65;
	wire [WIDTH-1:0] wire_d6_66;
	wire [WIDTH-1:0] wire_d6_67;
	wire [WIDTH-1:0] wire_d6_68;
	wire [WIDTH-1:0] wire_d6_69;
	wire [WIDTH-1:0] wire_d6_70;
	wire [WIDTH-1:0] wire_d6_71;
	wire [WIDTH-1:0] wire_d6_72;
	wire [WIDTH-1:0] wire_d6_73;
	wire [WIDTH-1:0] wire_d6_74;
	wire [WIDTH-1:0] wire_d6_75;
	wire [WIDTH-1:0] wire_d6_76;
	wire [WIDTH-1:0] wire_d6_77;
	wire [WIDTH-1:0] wire_d6_78;
	wire [WIDTH-1:0] wire_d6_79;
	wire [WIDTH-1:0] wire_d6_80;
	wire [WIDTH-1:0] wire_d6_81;
	wire [WIDTH-1:0] wire_d6_82;
	wire [WIDTH-1:0] wire_d6_83;
	wire [WIDTH-1:0] wire_d6_84;
	wire [WIDTH-1:0] wire_d6_85;
	wire [WIDTH-1:0] wire_d6_86;
	wire [WIDTH-1:0] wire_d6_87;
	wire [WIDTH-1:0] wire_d6_88;
	wire [WIDTH-1:0] wire_d6_89;
	wire [WIDTH-1:0] wire_d6_90;
	wire [WIDTH-1:0] wire_d6_91;
	wire [WIDTH-1:0] wire_d6_92;
	wire [WIDTH-1:0] wire_d6_93;
	wire [WIDTH-1:0] wire_d6_94;
	wire [WIDTH-1:0] wire_d6_95;
	wire [WIDTH-1:0] wire_d6_96;
	wire [WIDTH-1:0] wire_d6_97;
	wire [WIDTH-1:0] wire_d6_98;
	wire [WIDTH-1:0] wire_d6_99;
	wire [WIDTH-1:0] wire_d6_100;
	wire [WIDTH-1:0] wire_d6_101;
	wire [WIDTH-1:0] wire_d6_102;
	wire [WIDTH-1:0] wire_d6_103;
	wire [WIDTH-1:0] wire_d6_104;
	wire [WIDTH-1:0] wire_d6_105;
	wire [WIDTH-1:0] wire_d6_106;
	wire [WIDTH-1:0] wire_d6_107;
	wire [WIDTH-1:0] wire_d6_108;
	wire [WIDTH-1:0] wire_d6_109;
	wire [WIDTH-1:0] wire_d6_110;
	wire [WIDTH-1:0] wire_d6_111;
	wire [WIDTH-1:0] wire_d6_112;
	wire [WIDTH-1:0] wire_d6_113;
	wire [WIDTH-1:0] wire_d6_114;
	wire [WIDTH-1:0] wire_d6_115;
	wire [WIDTH-1:0] wire_d6_116;
	wire [WIDTH-1:0] wire_d6_117;
	wire [WIDTH-1:0] wire_d6_118;
	wire [WIDTH-1:0] wire_d6_119;
	wire [WIDTH-1:0] wire_d6_120;
	wire [WIDTH-1:0] wire_d6_121;
	wire [WIDTH-1:0] wire_d6_122;
	wire [WIDTH-1:0] wire_d6_123;
	wire [WIDTH-1:0] wire_d6_124;
	wire [WIDTH-1:0] wire_d6_125;
	wire [WIDTH-1:0] wire_d6_126;
	wire [WIDTH-1:0] wire_d6_127;
	wire [WIDTH-1:0] wire_d6_128;
	wire [WIDTH-1:0] wire_d6_129;
	wire [WIDTH-1:0] wire_d6_130;
	wire [WIDTH-1:0] wire_d6_131;
	wire [WIDTH-1:0] wire_d6_132;
	wire [WIDTH-1:0] wire_d6_133;
	wire [WIDTH-1:0] wire_d6_134;
	wire [WIDTH-1:0] wire_d6_135;
	wire [WIDTH-1:0] wire_d6_136;
	wire [WIDTH-1:0] wire_d6_137;
	wire [WIDTH-1:0] wire_d6_138;
	wire [WIDTH-1:0] wire_d6_139;
	wire [WIDTH-1:0] wire_d6_140;
	wire [WIDTH-1:0] wire_d6_141;
	wire [WIDTH-1:0] wire_d6_142;
	wire [WIDTH-1:0] wire_d6_143;
	wire [WIDTH-1:0] wire_d6_144;
	wire [WIDTH-1:0] wire_d6_145;
	wire [WIDTH-1:0] wire_d6_146;
	wire [WIDTH-1:0] wire_d6_147;
	wire [WIDTH-1:0] wire_d6_148;
	wire [WIDTH-1:0] wire_d6_149;
	wire [WIDTH-1:0] wire_d6_150;
	wire [WIDTH-1:0] wire_d6_151;
	wire [WIDTH-1:0] wire_d6_152;
	wire [WIDTH-1:0] wire_d6_153;
	wire [WIDTH-1:0] wire_d6_154;
	wire [WIDTH-1:0] wire_d6_155;
	wire [WIDTH-1:0] wire_d6_156;
	wire [WIDTH-1:0] wire_d6_157;
	wire [WIDTH-1:0] wire_d6_158;
	wire [WIDTH-1:0] wire_d6_159;
	wire [WIDTH-1:0] wire_d6_160;
	wire [WIDTH-1:0] wire_d6_161;
	wire [WIDTH-1:0] wire_d6_162;
	wire [WIDTH-1:0] wire_d6_163;
	wire [WIDTH-1:0] wire_d6_164;
	wire [WIDTH-1:0] wire_d6_165;
	wire [WIDTH-1:0] wire_d6_166;
	wire [WIDTH-1:0] wire_d6_167;
	wire [WIDTH-1:0] wire_d6_168;
	wire [WIDTH-1:0] wire_d6_169;
	wire [WIDTH-1:0] wire_d6_170;
	wire [WIDTH-1:0] wire_d6_171;
	wire [WIDTH-1:0] wire_d6_172;
	wire [WIDTH-1:0] wire_d6_173;
	wire [WIDTH-1:0] wire_d6_174;
	wire [WIDTH-1:0] wire_d6_175;
	wire [WIDTH-1:0] wire_d6_176;
	wire [WIDTH-1:0] wire_d6_177;
	wire [WIDTH-1:0] wire_d6_178;
	wire [WIDTH-1:0] wire_d6_179;
	wire [WIDTH-1:0] wire_d6_180;
	wire [WIDTH-1:0] wire_d6_181;
	wire [WIDTH-1:0] wire_d6_182;
	wire [WIDTH-1:0] wire_d6_183;
	wire [WIDTH-1:0] wire_d6_184;
	wire [WIDTH-1:0] wire_d6_185;
	wire [WIDTH-1:0] wire_d6_186;
	wire [WIDTH-1:0] wire_d6_187;
	wire [WIDTH-1:0] wire_d6_188;
	wire [WIDTH-1:0] wire_d6_189;
	wire [WIDTH-1:0] wire_d6_190;
	wire [WIDTH-1:0] wire_d6_191;
	wire [WIDTH-1:0] wire_d6_192;
	wire [WIDTH-1:0] wire_d6_193;
	wire [WIDTH-1:0] wire_d6_194;
	wire [WIDTH-1:0] wire_d6_195;
	wire [WIDTH-1:0] wire_d6_196;
	wire [WIDTH-1:0] wire_d6_197;
	wire [WIDTH-1:0] wire_d6_198;
	wire [WIDTH-1:0] wire_d7_0;
	wire [WIDTH-1:0] wire_d7_1;
	wire [WIDTH-1:0] wire_d7_2;
	wire [WIDTH-1:0] wire_d7_3;
	wire [WIDTH-1:0] wire_d7_4;
	wire [WIDTH-1:0] wire_d7_5;
	wire [WIDTH-1:0] wire_d7_6;
	wire [WIDTH-1:0] wire_d7_7;
	wire [WIDTH-1:0] wire_d7_8;
	wire [WIDTH-1:0] wire_d7_9;
	wire [WIDTH-1:0] wire_d7_10;
	wire [WIDTH-1:0] wire_d7_11;
	wire [WIDTH-1:0] wire_d7_12;
	wire [WIDTH-1:0] wire_d7_13;
	wire [WIDTH-1:0] wire_d7_14;
	wire [WIDTH-1:0] wire_d7_15;
	wire [WIDTH-1:0] wire_d7_16;
	wire [WIDTH-1:0] wire_d7_17;
	wire [WIDTH-1:0] wire_d7_18;
	wire [WIDTH-1:0] wire_d7_19;
	wire [WIDTH-1:0] wire_d7_20;
	wire [WIDTH-1:0] wire_d7_21;
	wire [WIDTH-1:0] wire_d7_22;
	wire [WIDTH-1:0] wire_d7_23;
	wire [WIDTH-1:0] wire_d7_24;
	wire [WIDTH-1:0] wire_d7_25;
	wire [WIDTH-1:0] wire_d7_26;
	wire [WIDTH-1:0] wire_d7_27;
	wire [WIDTH-1:0] wire_d7_28;
	wire [WIDTH-1:0] wire_d7_29;
	wire [WIDTH-1:0] wire_d7_30;
	wire [WIDTH-1:0] wire_d7_31;
	wire [WIDTH-1:0] wire_d7_32;
	wire [WIDTH-1:0] wire_d7_33;
	wire [WIDTH-1:0] wire_d7_34;
	wire [WIDTH-1:0] wire_d7_35;
	wire [WIDTH-1:0] wire_d7_36;
	wire [WIDTH-1:0] wire_d7_37;
	wire [WIDTH-1:0] wire_d7_38;
	wire [WIDTH-1:0] wire_d7_39;
	wire [WIDTH-1:0] wire_d7_40;
	wire [WIDTH-1:0] wire_d7_41;
	wire [WIDTH-1:0] wire_d7_42;
	wire [WIDTH-1:0] wire_d7_43;
	wire [WIDTH-1:0] wire_d7_44;
	wire [WIDTH-1:0] wire_d7_45;
	wire [WIDTH-1:0] wire_d7_46;
	wire [WIDTH-1:0] wire_d7_47;
	wire [WIDTH-1:0] wire_d7_48;
	wire [WIDTH-1:0] wire_d7_49;
	wire [WIDTH-1:0] wire_d7_50;
	wire [WIDTH-1:0] wire_d7_51;
	wire [WIDTH-1:0] wire_d7_52;
	wire [WIDTH-1:0] wire_d7_53;
	wire [WIDTH-1:0] wire_d7_54;
	wire [WIDTH-1:0] wire_d7_55;
	wire [WIDTH-1:0] wire_d7_56;
	wire [WIDTH-1:0] wire_d7_57;
	wire [WIDTH-1:0] wire_d7_58;
	wire [WIDTH-1:0] wire_d7_59;
	wire [WIDTH-1:0] wire_d7_60;
	wire [WIDTH-1:0] wire_d7_61;
	wire [WIDTH-1:0] wire_d7_62;
	wire [WIDTH-1:0] wire_d7_63;
	wire [WIDTH-1:0] wire_d7_64;
	wire [WIDTH-1:0] wire_d7_65;
	wire [WIDTH-1:0] wire_d7_66;
	wire [WIDTH-1:0] wire_d7_67;
	wire [WIDTH-1:0] wire_d7_68;
	wire [WIDTH-1:0] wire_d7_69;
	wire [WIDTH-1:0] wire_d7_70;
	wire [WIDTH-1:0] wire_d7_71;
	wire [WIDTH-1:0] wire_d7_72;
	wire [WIDTH-1:0] wire_d7_73;
	wire [WIDTH-1:0] wire_d7_74;
	wire [WIDTH-1:0] wire_d7_75;
	wire [WIDTH-1:0] wire_d7_76;
	wire [WIDTH-1:0] wire_d7_77;
	wire [WIDTH-1:0] wire_d7_78;
	wire [WIDTH-1:0] wire_d7_79;
	wire [WIDTH-1:0] wire_d7_80;
	wire [WIDTH-1:0] wire_d7_81;
	wire [WIDTH-1:0] wire_d7_82;
	wire [WIDTH-1:0] wire_d7_83;
	wire [WIDTH-1:0] wire_d7_84;
	wire [WIDTH-1:0] wire_d7_85;
	wire [WIDTH-1:0] wire_d7_86;
	wire [WIDTH-1:0] wire_d7_87;
	wire [WIDTH-1:0] wire_d7_88;
	wire [WIDTH-1:0] wire_d7_89;
	wire [WIDTH-1:0] wire_d7_90;
	wire [WIDTH-1:0] wire_d7_91;
	wire [WIDTH-1:0] wire_d7_92;
	wire [WIDTH-1:0] wire_d7_93;
	wire [WIDTH-1:0] wire_d7_94;
	wire [WIDTH-1:0] wire_d7_95;
	wire [WIDTH-1:0] wire_d7_96;
	wire [WIDTH-1:0] wire_d7_97;
	wire [WIDTH-1:0] wire_d7_98;
	wire [WIDTH-1:0] wire_d7_99;
	wire [WIDTH-1:0] wire_d7_100;
	wire [WIDTH-1:0] wire_d7_101;
	wire [WIDTH-1:0] wire_d7_102;
	wire [WIDTH-1:0] wire_d7_103;
	wire [WIDTH-1:0] wire_d7_104;
	wire [WIDTH-1:0] wire_d7_105;
	wire [WIDTH-1:0] wire_d7_106;
	wire [WIDTH-1:0] wire_d7_107;
	wire [WIDTH-1:0] wire_d7_108;
	wire [WIDTH-1:0] wire_d7_109;
	wire [WIDTH-1:0] wire_d7_110;
	wire [WIDTH-1:0] wire_d7_111;
	wire [WIDTH-1:0] wire_d7_112;
	wire [WIDTH-1:0] wire_d7_113;
	wire [WIDTH-1:0] wire_d7_114;
	wire [WIDTH-1:0] wire_d7_115;
	wire [WIDTH-1:0] wire_d7_116;
	wire [WIDTH-1:0] wire_d7_117;
	wire [WIDTH-1:0] wire_d7_118;
	wire [WIDTH-1:0] wire_d7_119;
	wire [WIDTH-1:0] wire_d7_120;
	wire [WIDTH-1:0] wire_d7_121;
	wire [WIDTH-1:0] wire_d7_122;
	wire [WIDTH-1:0] wire_d7_123;
	wire [WIDTH-1:0] wire_d7_124;
	wire [WIDTH-1:0] wire_d7_125;
	wire [WIDTH-1:0] wire_d7_126;
	wire [WIDTH-1:0] wire_d7_127;
	wire [WIDTH-1:0] wire_d7_128;
	wire [WIDTH-1:0] wire_d7_129;
	wire [WIDTH-1:0] wire_d7_130;
	wire [WIDTH-1:0] wire_d7_131;
	wire [WIDTH-1:0] wire_d7_132;
	wire [WIDTH-1:0] wire_d7_133;
	wire [WIDTH-1:0] wire_d7_134;
	wire [WIDTH-1:0] wire_d7_135;
	wire [WIDTH-1:0] wire_d7_136;
	wire [WIDTH-1:0] wire_d7_137;
	wire [WIDTH-1:0] wire_d7_138;
	wire [WIDTH-1:0] wire_d7_139;
	wire [WIDTH-1:0] wire_d7_140;
	wire [WIDTH-1:0] wire_d7_141;
	wire [WIDTH-1:0] wire_d7_142;
	wire [WIDTH-1:0] wire_d7_143;
	wire [WIDTH-1:0] wire_d7_144;
	wire [WIDTH-1:0] wire_d7_145;
	wire [WIDTH-1:0] wire_d7_146;
	wire [WIDTH-1:0] wire_d7_147;
	wire [WIDTH-1:0] wire_d7_148;
	wire [WIDTH-1:0] wire_d7_149;
	wire [WIDTH-1:0] wire_d7_150;
	wire [WIDTH-1:0] wire_d7_151;
	wire [WIDTH-1:0] wire_d7_152;
	wire [WIDTH-1:0] wire_d7_153;
	wire [WIDTH-1:0] wire_d7_154;
	wire [WIDTH-1:0] wire_d7_155;
	wire [WIDTH-1:0] wire_d7_156;
	wire [WIDTH-1:0] wire_d7_157;
	wire [WIDTH-1:0] wire_d7_158;
	wire [WIDTH-1:0] wire_d7_159;
	wire [WIDTH-1:0] wire_d7_160;
	wire [WIDTH-1:0] wire_d7_161;
	wire [WIDTH-1:0] wire_d7_162;
	wire [WIDTH-1:0] wire_d7_163;
	wire [WIDTH-1:0] wire_d7_164;
	wire [WIDTH-1:0] wire_d7_165;
	wire [WIDTH-1:0] wire_d7_166;
	wire [WIDTH-1:0] wire_d7_167;
	wire [WIDTH-1:0] wire_d7_168;
	wire [WIDTH-1:0] wire_d7_169;
	wire [WIDTH-1:0] wire_d7_170;
	wire [WIDTH-1:0] wire_d7_171;
	wire [WIDTH-1:0] wire_d7_172;
	wire [WIDTH-1:0] wire_d7_173;
	wire [WIDTH-1:0] wire_d7_174;
	wire [WIDTH-1:0] wire_d7_175;
	wire [WIDTH-1:0] wire_d7_176;
	wire [WIDTH-1:0] wire_d7_177;
	wire [WIDTH-1:0] wire_d7_178;
	wire [WIDTH-1:0] wire_d7_179;
	wire [WIDTH-1:0] wire_d7_180;
	wire [WIDTH-1:0] wire_d7_181;
	wire [WIDTH-1:0] wire_d7_182;
	wire [WIDTH-1:0] wire_d7_183;
	wire [WIDTH-1:0] wire_d7_184;
	wire [WIDTH-1:0] wire_d7_185;
	wire [WIDTH-1:0] wire_d7_186;
	wire [WIDTH-1:0] wire_d7_187;
	wire [WIDTH-1:0] wire_d7_188;
	wire [WIDTH-1:0] wire_d7_189;
	wire [WIDTH-1:0] wire_d7_190;
	wire [WIDTH-1:0] wire_d7_191;
	wire [WIDTH-1:0] wire_d7_192;
	wire [WIDTH-1:0] wire_d7_193;
	wire [WIDTH-1:0] wire_d7_194;
	wire [WIDTH-1:0] wire_d7_195;
	wire [WIDTH-1:0] wire_d7_196;
	wire [WIDTH-1:0] wire_d7_197;
	wire [WIDTH-1:0] wire_d7_198;
	wire [WIDTH-1:0] wire_d8_0;
	wire [WIDTH-1:0] wire_d8_1;
	wire [WIDTH-1:0] wire_d8_2;
	wire [WIDTH-1:0] wire_d8_3;
	wire [WIDTH-1:0] wire_d8_4;
	wire [WIDTH-1:0] wire_d8_5;
	wire [WIDTH-1:0] wire_d8_6;
	wire [WIDTH-1:0] wire_d8_7;
	wire [WIDTH-1:0] wire_d8_8;
	wire [WIDTH-1:0] wire_d8_9;
	wire [WIDTH-1:0] wire_d8_10;
	wire [WIDTH-1:0] wire_d8_11;
	wire [WIDTH-1:0] wire_d8_12;
	wire [WIDTH-1:0] wire_d8_13;
	wire [WIDTH-1:0] wire_d8_14;
	wire [WIDTH-1:0] wire_d8_15;
	wire [WIDTH-1:0] wire_d8_16;
	wire [WIDTH-1:0] wire_d8_17;
	wire [WIDTH-1:0] wire_d8_18;
	wire [WIDTH-1:0] wire_d8_19;
	wire [WIDTH-1:0] wire_d8_20;
	wire [WIDTH-1:0] wire_d8_21;
	wire [WIDTH-1:0] wire_d8_22;
	wire [WIDTH-1:0] wire_d8_23;
	wire [WIDTH-1:0] wire_d8_24;
	wire [WIDTH-1:0] wire_d8_25;
	wire [WIDTH-1:0] wire_d8_26;
	wire [WIDTH-1:0] wire_d8_27;
	wire [WIDTH-1:0] wire_d8_28;
	wire [WIDTH-1:0] wire_d8_29;
	wire [WIDTH-1:0] wire_d8_30;
	wire [WIDTH-1:0] wire_d8_31;
	wire [WIDTH-1:0] wire_d8_32;
	wire [WIDTH-1:0] wire_d8_33;
	wire [WIDTH-1:0] wire_d8_34;
	wire [WIDTH-1:0] wire_d8_35;
	wire [WIDTH-1:0] wire_d8_36;
	wire [WIDTH-1:0] wire_d8_37;
	wire [WIDTH-1:0] wire_d8_38;
	wire [WIDTH-1:0] wire_d8_39;
	wire [WIDTH-1:0] wire_d8_40;
	wire [WIDTH-1:0] wire_d8_41;
	wire [WIDTH-1:0] wire_d8_42;
	wire [WIDTH-1:0] wire_d8_43;
	wire [WIDTH-1:0] wire_d8_44;
	wire [WIDTH-1:0] wire_d8_45;
	wire [WIDTH-1:0] wire_d8_46;
	wire [WIDTH-1:0] wire_d8_47;
	wire [WIDTH-1:0] wire_d8_48;
	wire [WIDTH-1:0] wire_d8_49;
	wire [WIDTH-1:0] wire_d8_50;
	wire [WIDTH-1:0] wire_d8_51;
	wire [WIDTH-1:0] wire_d8_52;
	wire [WIDTH-1:0] wire_d8_53;
	wire [WIDTH-1:0] wire_d8_54;
	wire [WIDTH-1:0] wire_d8_55;
	wire [WIDTH-1:0] wire_d8_56;
	wire [WIDTH-1:0] wire_d8_57;
	wire [WIDTH-1:0] wire_d8_58;
	wire [WIDTH-1:0] wire_d8_59;
	wire [WIDTH-1:0] wire_d8_60;
	wire [WIDTH-1:0] wire_d8_61;
	wire [WIDTH-1:0] wire_d8_62;
	wire [WIDTH-1:0] wire_d8_63;
	wire [WIDTH-1:0] wire_d8_64;
	wire [WIDTH-1:0] wire_d8_65;
	wire [WIDTH-1:0] wire_d8_66;
	wire [WIDTH-1:0] wire_d8_67;
	wire [WIDTH-1:0] wire_d8_68;
	wire [WIDTH-1:0] wire_d8_69;
	wire [WIDTH-1:0] wire_d8_70;
	wire [WIDTH-1:0] wire_d8_71;
	wire [WIDTH-1:0] wire_d8_72;
	wire [WIDTH-1:0] wire_d8_73;
	wire [WIDTH-1:0] wire_d8_74;
	wire [WIDTH-1:0] wire_d8_75;
	wire [WIDTH-1:0] wire_d8_76;
	wire [WIDTH-1:0] wire_d8_77;
	wire [WIDTH-1:0] wire_d8_78;
	wire [WIDTH-1:0] wire_d8_79;
	wire [WIDTH-1:0] wire_d8_80;
	wire [WIDTH-1:0] wire_d8_81;
	wire [WIDTH-1:0] wire_d8_82;
	wire [WIDTH-1:0] wire_d8_83;
	wire [WIDTH-1:0] wire_d8_84;
	wire [WIDTH-1:0] wire_d8_85;
	wire [WIDTH-1:0] wire_d8_86;
	wire [WIDTH-1:0] wire_d8_87;
	wire [WIDTH-1:0] wire_d8_88;
	wire [WIDTH-1:0] wire_d8_89;
	wire [WIDTH-1:0] wire_d8_90;
	wire [WIDTH-1:0] wire_d8_91;
	wire [WIDTH-1:0] wire_d8_92;
	wire [WIDTH-1:0] wire_d8_93;
	wire [WIDTH-1:0] wire_d8_94;
	wire [WIDTH-1:0] wire_d8_95;
	wire [WIDTH-1:0] wire_d8_96;
	wire [WIDTH-1:0] wire_d8_97;
	wire [WIDTH-1:0] wire_d8_98;
	wire [WIDTH-1:0] wire_d8_99;
	wire [WIDTH-1:0] wire_d8_100;
	wire [WIDTH-1:0] wire_d8_101;
	wire [WIDTH-1:0] wire_d8_102;
	wire [WIDTH-1:0] wire_d8_103;
	wire [WIDTH-1:0] wire_d8_104;
	wire [WIDTH-1:0] wire_d8_105;
	wire [WIDTH-1:0] wire_d8_106;
	wire [WIDTH-1:0] wire_d8_107;
	wire [WIDTH-1:0] wire_d8_108;
	wire [WIDTH-1:0] wire_d8_109;
	wire [WIDTH-1:0] wire_d8_110;
	wire [WIDTH-1:0] wire_d8_111;
	wire [WIDTH-1:0] wire_d8_112;
	wire [WIDTH-1:0] wire_d8_113;
	wire [WIDTH-1:0] wire_d8_114;
	wire [WIDTH-1:0] wire_d8_115;
	wire [WIDTH-1:0] wire_d8_116;
	wire [WIDTH-1:0] wire_d8_117;
	wire [WIDTH-1:0] wire_d8_118;
	wire [WIDTH-1:0] wire_d8_119;
	wire [WIDTH-1:0] wire_d8_120;
	wire [WIDTH-1:0] wire_d8_121;
	wire [WIDTH-1:0] wire_d8_122;
	wire [WIDTH-1:0] wire_d8_123;
	wire [WIDTH-1:0] wire_d8_124;
	wire [WIDTH-1:0] wire_d8_125;
	wire [WIDTH-1:0] wire_d8_126;
	wire [WIDTH-1:0] wire_d8_127;
	wire [WIDTH-1:0] wire_d8_128;
	wire [WIDTH-1:0] wire_d8_129;
	wire [WIDTH-1:0] wire_d8_130;
	wire [WIDTH-1:0] wire_d8_131;
	wire [WIDTH-1:0] wire_d8_132;
	wire [WIDTH-1:0] wire_d8_133;
	wire [WIDTH-1:0] wire_d8_134;
	wire [WIDTH-1:0] wire_d8_135;
	wire [WIDTH-1:0] wire_d8_136;
	wire [WIDTH-1:0] wire_d8_137;
	wire [WIDTH-1:0] wire_d8_138;
	wire [WIDTH-1:0] wire_d8_139;
	wire [WIDTH-1:0] wire_d8_140;
	wire [WIDTH-1:0] wire_d8_141;
	wire [WIDTH-1:0] wire_d8_142;
	wire [WIDTH-1:0] wire_d8_143;
	wire [WIDTH-1:0] wire_d8_144;
	wire [WIDTH-1:0] wire_d8_145;
	wire [WIDTH-1:0] wire_d8_146;
	wire [WIDTH-1:0] wire_d8_147;
	wire [WIDTH-1:0] wire_d8_148;
	wire [WIDTH-1:0] wire_d8_149;
	wire [WIDTH-1:0] wire_d8_150;
	wire [WIDTH-1:0] wire_d8_151;
	wire [WIDTH-1:0] wire_d8_152;
	wire [WIDTH-1:0] wire_d8_153;
	wire [WIDTH-1:0] wire_d8_154;
	wire [WIDTH-1:0] wire_d8_155;
	wire [WIDTH-1:0] wire_d8_156;
	wire [WIDTH-1:0] wire_d8_157;
	wire [WIDTH-1:0] wire_d8_158;
	wire [WIDTH-1:0] wire_d8_159;
	wire [WIDTH-1:0] wire_d8_160;
	wire [WIDTH-1:0] wire_d8_161;
	wire [WIDTH-1:0] wire_d8_162;
	wire [WIDTH-1:0] wire_d8_163;
	wire [WIDTH-1:0] wire_d8_164;
	wire [WIDTH-1:0] wire_d8_165;
	wire [WIDTH-1:0] wire_d8_166;
	wire [WIDTH-1:0] wire_d8_167;
	wire [WIDTH-1:0] wire_d8_168;
	wire [WIDTH-1:0] wire_d8_169;
	wire [WIDTH-1:0] wire_d8_170;
	wire [WIDTH-1:0] wire_d8_171;
	wire [WIDTH-1:0] wire_d8_172;
	wire [WIDTH-1:0] wire_d8_173;
	wire [WIDTH-1:0] wire_d8_174;
	wire [WIDTH-1:0] wire_d8_175;
	wire [WIDTH-1:0] wire_d8_176;
	wire [WIDTH-1:0] wire_d8_177;
	wire [WIDTH-1:0] wire_d8_178;
	wire [WIDTH-1:0] wire_d8_179;
	wire [WIDTH-1:0] wire_d8_180;
	wire [WIDTH-1:0] wire_d8_181;
	wire [WIDTH-1:0] wire_d8_182;
	wire [WIDTH-1:0] wire_d8_183;
	wire [WIDTH-1:0] wire_d8_184;
	wire [WIDTH-1:0] wire_d8_185;
	wire [WIDTH-1:0] wire_d8_186;
	wire [WIDTH-1:0] wire_d8_187;
	wire [WIDTH-1:0] wire_d8_188;
	wire [WIDTH-1:0] wire_d8_189;
	wire [WIDTH-1:0] wire_d8_190;
	wire [WIDTH-1:0] wire_d8_191;
	wire [WIDTH-1:0] wire_d8_192;
	wire [WIDTH-1:0] wire_d8_193;
	wire [WIDTH-1:0] wire_d8_194;
	wire [WIDTH-1:0] wire_d8_195;
	wire [WIDTH-1:0] wire_d8_196;
	wire [WIDTH-1:0] wire_d8_197;
	wire [WIDTH-1:0] wire_d8_198;
	wire [WIDTH-1:0] wire_d9_0;
	wire [WIDTH-1:0] wire_d9_1;
	wire [WIDTH-1:0] wire_d9_2;
	wire [WIDTH-1:0] wire_d9_3;
	wire [WIDTH-1:0] wire_d9_4;
	wire [WIDTH-1:0] wire_d9_5;
	wire [WIDTH-1:0] wire_d9_6;
	wire [WIDTH-1:0] wire_d9_7;
	wire [WIDTH-1:0] wire_d9_8;
	wire [WIDTH-1:0] wire_d9_9;
	wire [WIDTH-1:0] wire_d9_10;
	wire [WIDTH-1:0] wire_d9_11;
	wire [WIDTH-1:0] wire_d9_12;
	wire [WIDTH-1:0] wire_d9_13;
	wire [WIDTH-1:0] wire_d9_14;
	wire [WIDTH-1:0] wire_d9_15;
	wire [WIDTH-1:0] wire_d9_16;
	wire [WIDTH-1:0] wire_d9_17;
	wire [WIDTH-1:0] wire_d9_18;
	wire [WIDTH-1:0] wire_d9_19;
	wire [WIDTH-1:0] wire_d9_20;
	wire [WIDTH-1:0] wire_d9_21;
	wire [WIDTH-1:0] wire_d9_22;
	wire [WIDTH-1:0] wire_d9_23;
	wire [WIDTH-1:0] wire_d9_24;
	wire [WIDTH-1:0] wire_d9_25;
	wire [WIDTH-1:0] wire_d9_26;
	wire [WIDTH-1:0] wire_d9_27;
	wire [WIDTH-1:0] wire_d9_28;
	wire [WIDTH-1:0] wire_d9_29;
	wire [WIDTH-1:0] wire_d9_30;
	wire [WIDTH-1:0] wire_d9_31;
	wire [WIDTH-1:0] wire_d9_32;
	wire [WIDTH-1:0] wire_d9_33;
	wire [WIDTH-1:0] wire_d9_34;
	wire [WIDTH-1:0] wire_d9_35;
	wire [WIDTH-1:0] wire_d9_36;
	wire [WIDTH-1:0] wire_d9_37;
	wire [WIDTH-1:0] wire_d9_38;
	wire [WIDTH-1:0] wire_d9_39;
	wire [WIDTH-1:0] wire_d9_40;
	wire [WIDTH-1:0] wire_d9_41;
	wire [WIDTH-1:0] wire_d9_42;
	wire [WIDTH-1:0] wire_d9_43;
	wire [WIDTH-1:0] wire_d9_44;
	wire [WIDTH-1:0] wire_d9_45;
	wire [WIDTH-1:0] wire_d9_46;
	wire [WIDTH-1:0] wire_d9_47;
	wire [WIDTH-1:0] wire_d9_48;
	wire [WIDTH-1:0] wire_d9_49;
	wire [WIDTH-1:0] wire_d9_50;
	wire [WIDTH-1:0] wire_d9_51;
	wire [WIDTH-1:0] wire_d9_52;
	wire [WIDTH-1:0] wire_d9_53;
	wire [WIDTH-1:0] wire_d9_54;
	wire [WIDTH-1:0] wire_d9_55;
	wire [WIDTH-1:0] wire_d9_56;
	wire [WIDTH-1:0] wire_d9_57;
	wire [WIDTH-1:0] wire_d9_58;
	wire [WIDTH-1:0] wire_d9_59;
	wire [WIDTH-1:0] wire_d9_60;
	wire [WIDTH-1:0] wire_d9_61;
	wire [WIDTH-1:0] wire_d9_62;
	wire [WIDTH-1:0] wire_d9_63;
	wire [WIDTH-1:0] wire_d9_64;
	wire [WIDTH-1:0] wire_d9_65;
	wire [WIDTH-1:0] wire_d9_66;
	wire [WIDTH-1:0] wire_d9_67;
	wire [WIDTH-1:0] wire_d9_68;
	wire [WIDTH-1:0] wire_d9_69;
	wire [WIDTH-1:0] wire_d9_70;
	wire [WIDTH-1:0] wire_d9_71;
	wire [WIDTH-1:0] wire_d9_72;
	wire [WIDTH-1:0] wire_d9_73;
	wire [WIDTH-1:0] wire_d9_74;
	wire [WIDTH-1:0] wire_d9_75;
	wire [WIDTH-1:0] wire_d9_76;
	wire [WIDTH-1:0] wire_d9_77;
	wire [WIDTH-1:0] wire_d9_78;
	wire [WIDTH-1:0] wire_d9_79;
	wire [WIDTH-1:0] wire_d9_80;
	wire [WIDTH-1:0] wire_d9_81;
	wire [WIDTH-1:0] wire_d9_82;
	wire [WIDTH-1:0] wire_d9_83;
	wire [WIDTH-1:0] wire_d9_84;
	wire [WIDTH-1:0] wire_d9_85;
	wire [WIDTH-1:0] wire_d9_86;
	wire [WIDTH-1:0] wire_d9_87;
	wire [WIDTH-1:0] wire_d9_88;
	wire [WIDTH-1:0] wire_d9_89;
	wire [WIDTH-1:0] wire_d9_90;
	wire [WIDTH-1:0] wire_d9_91;
	wire [WIDTH-1:0] wire_d9_92;
	wire [WIDTH-1:0] wire_d9_93;
	wire [WIDTH-1:0] wire_d9_94;
	wire [WIDTH-1:0] wire_d9_95;
	wire [WIDTH-1:0] wire_d9_96;
	wire [WIDTH-1:0] wire_d9_97;
	wire [WIDTH-1:0] wire_d9_98;
	wire [WIDTH-1:0] wire_d9_99;
	wire [WIDTH-1:0] wire_d9_100;
	wire [WIDTH-1:0] wire_d9_101;
	wire [WIDTH-1:0] wire_d9_102;
	wire [WIDTH-1:0] wire_d9_103;
	wire [WIDTH-1:0] wire_d9_104;
	wire [WIDTH-1:0] wire_d9_105;
	wire [WIDTH-1:0] wire_d9_106;
	wire [WIDTH-1:0] wire_d9_107;
	wire [WIDTH-1:0] wire_d9_108;
	wire [WIDTH-1:0] wire_d9_109;
	wire [WIDTH-1:0] wire_d9_110;
	wire [WIDTH-1:0] wire_d9_111;
	wire [WIDTH-1:0] wire_d9_112;
	wire [WIDTH-1:0] wire_d9_113;
	wire [WIDTH-1:0] wire_d9_114;
	wire [WIDTH-1:0] wire_d9_115;
	wire [WIDTH-1:0] wire_d9_116;
	wire [WIDTH-1:0] wire_d9_117;
	wire [WIDTH-1:0] wire_d9_118;
	wire [WIDTH-1:0] wire_d9_119;
	wire [WIDTH-1:0] wire_d9_120;
	wire [WIDTH-1:0] wire_d9_121;
	wire [WIDTH-1:0] wire_d9_122;
	wire [WIDTH-1:0] wire_d9_123;
	wire [WIDTH-1:0] wire_d9_124;
	wire [WIDTH-1:0] wire_d9_125;
	wire [WIDTH-1:0] wire_d9_126;
	wire [WIDTH-1:0] wire_d9_127;
	wire [WIDTH-1:0] wire_d9_128;
	wire [WIDTH-1:0] wire_d9_129;
	wire [WIDTH-1:0] wire_d9_130;
	wire [WIDTH-1:0] wire_d9_131;
	wire [WIDTH-1:0] wire_d9_132;
	wire [WIDTH-1:0] wire_d9_133;
	wire [WIDTH-1:0] wire_d9_134;
	wire [WIDTH-1:0] wire_d9_135;
	wire [WIDTH-1:0] wire_d9_136;
	wire [WIDTH-1:0] wire_d9_137;
	wire [WIDTH-1:0] wire_d9_138;
	wire [WIDTH-1:0] wire_d9_139;
	wire [WIDTH-1:0] wire_d9_140;
	wire [WIDTH-1:0] wire_d9_141;
	wire [WIDTH-1:0] wire_d9_142;
	wire [WIDTH-1:0] wire_d9_143;
	wire [WIDTH-1:0] wire_d9_144;
	wire [WIDTH-1:0] wire_d9_145;
	wire [WIDTH-1:0] wire_d9_146;
	wire [WIDTH-1:0] wire_d9_147;
	wire [WIDTH-1:0] wire_d9_148;
	wire [WIDTH-1:0] wire_d9_149;
	wire [WIDTH-1:0] wire_d9_150;
	wire [WIDTH-1:0] wire_d9_151;
	wire [WIDTH-1:0] wire_d9_152;
	wire [WIDTH-1:0] wire_d9_153;
	wire [WIDTH-1:0] wire_d9_154;
	wire [WIDTH-1:0] wire_d9_155;
	wire [WIDTH-1:0] wire_d9_156;
	wire [WIDTH-1:0] wire_d9_157;
	wire [WIDTH-1:0] wire_d9_158;
	wire [WIDTH-1:0] wire_d9_159;
	wire [WIDTH-1:0] wire_d9_160;
	wire [WIDTH-1:0] wire_d9_161;
	wire [WIDTH-1:0] wire_d9_162;
	wire [WIDTH-1:0] wire_d9_163;
	wire [WIDTH-1:0] wire_d9_164;
	wire [WIDTH-1:0] wire_d9_165;
	wire [WIDTH-1:0] wire_d9_166;
	wire [WIDTH-1:0] wire_d9_167;
	wire [WIDTH-1:0] wire_d9_168;
	wire [WIDTH-1:0] wire_d9_169;
	wire [WIDTH-1:0] wire_d9_170;
	wire [WIDTH-1:0] wire_d9_171;
	wire [WIDTH-1:0] wire_d9_172;
	wire [WIDTH-1:0] wire_d9_173;
	wire [WIDTH-1:0] wire_d9_174;
	wire [WIDTH-1:0] wire_d9_175;
	wire [WIDTH-1:0] wire_d9_176;
	wire [WIDTH-1:0] wire_d9_177;
	wire [WIDTH-1:0] wire_d9_178;
	wire [WIDTH-1:0] wire_d9_179;
	wire [WIDTH-1:0] wire_d9_180;
	wire [WIDTH-1:0] wire_d9_181;
	wire [WIDTH-1:0] wire_d9_182;
	wire [WIDTH-1:0] wire_d9_183;
	wire [WIDTH-1:0] wire_d9_184;
	wire [WIDTH-1:0] wire_d9_185;
	wire [WIDTH-1:0] wire_d9_186;
	wire [WIDTH-1:0] wire_d9_187;
	wire [WIDTH-1:0] wire_d9_188;
	wire [WIDTH-1:0] wire_d9_189;
	wire [WIDTH-1:0] wire_d9_190;
	wire [WIDTH-1:0] wire_d9_191;
	wire [WIDTH-1:0] wire_d9_192;
	wire [WIDTH-1:0] wire_d9_193;
	wire [WIDTH-1:0] wire_d9_194;
	wire [WIDTH-1:0] wire_d9_195;
	wire [WIDTH-1:0] wire_d9_196;
	wire [WIDTH-1:0] wire_d9_197;
	wire [WIDTH-1:0] wire_d9_198;

	encoder #(.WIDTH(WIDTH)) encoder_instance100(.data_in(d_in0),.data_out(wire_d0_0),.clk(clk),.rst(rst));            //channel 1
	encoder #(.WIDTH(WIDTH)) encoder_instance101(.data_in(wire_d0_0),.data_out(wire_d0_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance102(.data_in(wire_d0_1),.data_out(wire_d0_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance103(.data_in(wire_d0_2),.data_out(wire_d0_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance104(.data_in(wire_d0_3),.data_out(wire_d0_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance105(.data_in(wire_d0_4),.data_out(wire_d0_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance106(.data_in(wire_d0_5),.data_out(wire_d0_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance107(.data_in(wire_d0_6),.data_out(wire_d0_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance108(.data_in(wire_d0_7),.data_out(wire_d0_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance109(.data_in(wire_d0_8),.data_out(wire_d0_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1010(.data_in(wire_d0_9),.data_out(wire_d0_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1011(.data_in(wire_d0_10),.data_out(wire_d0_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1012(.data_in(wire_d0_11),.data_out(wire_d0_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1013(.data_in(wire_d0_12),.data_out(wire_d0_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1014(.data_in(wire_d0_13),.data_out(wire_d0_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1015(.data_in(wire_d0_14),.data_out(wire_d0_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1016(.data_in(wire_d0_15),.data_out(wire_d0_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1017(.data_in(wire_d0_16),.data_out(wire_d0_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1018(.data_in(wire_d0_17),.data_out(wire_d0_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1019(.data_in(wire_d0_18),.data_out(wire_d0_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1020(.data_in(wire_d0_19),.data_out(wire_d0_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1021(.data_in(wire_d0_20),.data_out(wire_d0_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1022(.data_in(wire_d0_21),.data_out(wire_d0_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1023(.data_in(wire_d0_22),.data_out(wire_d0_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1024(.data_in(wire_d0_23),.data_out(wire_d0_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1025(.data_in(wire_d0_24),.data_out(wire_d0_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1026(.data_in(wire_d0_25),.data_out(wire_d0_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1027(.data_in(wire_d0_26),.data_out(wire_d0_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1028(.data_in(wire_d0_27),.data_out(wire_d0_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1029(.data_in(wire_d0_28),.data_out(wire_d0_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1030(.data_in(wire_d0_29),.data_out(wire_d0_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1031(.data_in(wire_d0_30),.data_out(wire_d0_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1032(.data_in(wire_d0_31),.data_out(wire_d0_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1033(.data_in(wire_d0_32),.data_out(wire_d0_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1034(.data_in(wire_d0_33),.data_out(wire_d0_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1035(.data_in(wire_d0_34),.data_out(wire_d0_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1036(.data_in(wire_d0_35),.data_out(wire_d0_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1037(.data_in(wire_d0_36),.data_out(wire_d0_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1038(.data_in(wire_d0_37),.data_out(wire_d0_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1039(.data_in(wire_d0_38),.data_out(wire_d0_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1040(.data_in(wire_d0_39),.data_out(wire_d0_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1041(.data_in(wire_d0_40),.data_out(wire_d0_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1042(.data_in(wire_d0_41),.data_out(wire_d0_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1043(.data_in(wire_d0_42),.data_out(wire_d0_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1044(.data_in(wire_d0_43),.data_out(wire_d0_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1045(.data_in(wire_d0_44),.data_out(wire_d0_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1046(.data_in(wire_d0_45),.data_out(wire_d0_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1047(.data_in(wire_d0_46),.data_out(wire_d0_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1048(.data_in(wire_d0_47),.data_out(wire_d0_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1049(.data_in(wire_d0_48),.data_out(wire_d0_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1050(.data_in(wire_d0_49),.data_out(wire_d0_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1051(.data_in(wire_d0_50),.data_out(wire_d0_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1052(.data_in(wire_d0_51),.data_out(wire_d0_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1053(.data_in(wire_d0_52),.data_out(wire_d0_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1054(.data_in(wire_d0_53),.data_out(wire_d0_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1055(.data_in(wire_d0_54),.data_out(wire_d0_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1056(.data_in(wire_d0_55),.data_out(wire_d0_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1057(.data_in(wire_d0_56),.data_out(wire_d0_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1058(.data_in(wire_d0_57),.data_out(wire_d0_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1059(.data_in(wire_d0_58),.data_out(wire_d0_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1060(.data_in(wire_d0_59),.data_out(wire_d0_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1061(.data_in(wire_d0_60),.data_out(wire_d0_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1062(.data_in(wire_d0_61),.data_out(wire_d0_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1063(.data_in(wire_d0_62),.data_out(wire_d0_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1064(.data_in(wire_d0_63),.data_out(wire_d0_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1065(.data_in(wire_d0_64),.data_out(wire_d0_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1066(.data_in(wire_d0_65),.data_out(wire_d0_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1067(.data_in(wire_d0_66),.data_out(wire_d0_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1068(.data_in(wire_d0_67),.data_out(wire_d0_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1069(.data_in(wire_d0_68),.data_out(wire_d0_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1070(.data_in(wire_d0_69),.data_out(wire_d0_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1071(.data_in(wire_d0_70),.data_out(wire_d0_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1072(.data_in(wire_d0_71),.data_out(wire_d0_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1073(.data_in(wire_d0_72),.data_out(wire_d0_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1074(.data_in(wire_d0_73),.data_out(wire_d0_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1075(.data_in(wire_d0_74),.data_out(wire_d0_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1076(.data_in(wire_d0_75),.data_out(wire_d0_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1077(.data_in(wire_d0_76),.data_out(wire_d0_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1078(.data_in(wire_d0_77),.data_out(wire_d0_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1079(.data_in(wire_d0_78),.data_out(wire_d0_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1080(.data_in(wire_d0_79),.data_out(wire_d0_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1081(.data_in(wire_d0_80),.data_out(wire_d0_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1082(.data_in(wire_d0_81),.data_out(wire_d0_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1083(.data_in(wire_d0_82),.data_out(wire_d0_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1084(.data_in(wire_d0_83),.data_out(wire_d0_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1085(.data_in(wire_d0_84),.data_out(wire_d0_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1086(.data_in(wire_d0_85),.data_out(wire_d0_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1087(.data_in(wire_d0_86),.data_out(wire_d0_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1088(.data_in(wire_d0_87),.data_out(wire_d0_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1089(.data_in(wire_d0_88),.data_out(wire_d0_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1090(.data_in(wire_d0_89),.data_out(wire_d0_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1091(.data_in(wire_d0_90),.data_out(wire_d0_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1092(.data_in(wire_d0_91),.data_out(wire_d0_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1093(.data_in(wire_d0_92),.data_out(wire_d0_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1094(.data_in(wire_d0_93),.data_out(wire_d0_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1095(.data_in(wire_d0_94),.data_out(wire_d0_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1096(.data_in(wire_d0_95),.data_out(wire_d0_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1097(.data_in(wire_d0_96),.data_out(wire_d0_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1098(.data_in(wire_d0_97),.data_out(wire_d0_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1099(.data_in(wire_d0_98),.data_out(wire_d0_99),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10100(.data_in(wire_d0_99),.data_out(wire_d0_100),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10101(.data_in(wire_d0_100),.data_out(wire_d0_101),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10102(.data_in(wire_d0_101),.data_out(wire_d0_102),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10103(.data_in(wire_d0_102),.data_out(wire_d0_103),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10104(.data_in(wire_d0_103),.data_out(wire_d0_104),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10105(.data_in(wire_d0_104),.data_out(wire_d0_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10106(.data_in(wire_d0_105),.data_out(wire_d0_106),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10107(.data_in(wire_d0_106),.data_out(wire_d0_107),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10108(.data_in(wire_d0_107),.data_out(wire_d0_108),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10109(.data_in(wire_d0_108),.data_out(wire_d0_109),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10110(.data_in(wire_d0_109),.data_out(wire_d0_110),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10111(.data_in(wire_d0_110),.data_out(wire_d0_111),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10112(.data_in(wire_d0_111),.data_out(wire_d0_112),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10113(.data_in(wire_d0_112),.data_out(wire_d0_113),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10114(.data_in(wire_d0_113),.data_out(wire_d0_114),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10115(.data_in(wire_d0_114),.data_out(wire_d0_115),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10116(.data_in(wire_d0_115),.data_out(wire_d0_116),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10117(.data_in(wire_d0_116),.data_out(wire_d0_117),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10118(.data_in(wire_d0_117),.data_out(wire_d0_118),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10119(.data_in(wire_d0_118),.data_out(wire_d0_119),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10120(.data_in(wire_d0_119),.data_out(wire_d0_120),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10121(.data_in(wire_d0_120),.data_out(wire_d0_121),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10122(.data_in(wire_d0_121),.data_out(wire_d0_122),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10123(.data_in(wire_d0_122),.data_out(wire_d0_123),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10124(.data_in(wire_d0_123),.data_out(wire_d0_124),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10125(.data_in(wire_d0_124),.data_out(wire_d0_125),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10126(.data_in(wire_d0_125),.data_out(wire_d0_126),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10127(.data_in(wire_d0_126),.data_out(wire_d0_127),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10128(.data_in(wire_d0_127),.data_out(wire_d0_128),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10129(.data_in(wire_d0_128),.data_out(wire_d0_129),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10130(.data_in(wire_d0_129),.data_out(wire_d0_130),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10131(.data_in(wire_d0_130),.data_out(wire_d0_131),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10132(.data_in(wire_d0_131),.data_out(wire_d0_132),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10133(.data_in(wire_d0_132),.data_out(wire_d0_133),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10134(.data_in(wire_d0_133),.data_out(wire_d0_134),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10135(.data_in(wire_d0_134),.data_out(wire_d0_135),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10136(.data_in(wire_d0_135),.data_out(wire_d0_136),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10137(.data_in(wire_d0_136),.data_out(wire_d0_137),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10138(.data_in(wire_d0_137),.data_out(wire_d0_138),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10139(.data_in(wire_d0_138),.data_out(wire_d0_139),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10140(.data_in(wire_d0_139),.data_out(wire_d0_140),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10141(.data_in(wire_d0_140),.data_out(wire_d0_141),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10142(.data_in(wire_d0_141),.data_out(wire_d0_142),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10143(.data_in(wire_d0_142),.data_out(wire_d0_143),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10144(.data_in(wire_d0_143),.data_out(wire_d0_144),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10145(.data_in(wire_d0_144),.data_out(wire_d0_145),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10146(.data_in(wire_d0_145),.data_out(wire_d0_146),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10147(.data_in(wire_d0_146),.data_out(wire_d0_147),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10148(.data_in(wire_d0_147),.data_out(wire_d0_148),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10149(.data_in(wire_d0_148),.data_out(wire_d0_149),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10150(.data_in(wire_d0_149),.data_out(wire_d0_150),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10151(.data_in(wire_d0_150),.data_out(wire_d0_151),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10152(.data_in(wire_d0_151),.data_out(wire_d0_152),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10153(.data_in(wire_d0_152),.data_out(wire_d0_153),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10154(.data_in(wire_d0_153),.data_out(wire_d0_154),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10155(.data_in(wire_d0_154),.data_out(wire_d0_155),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10156(.data_in(wire_d0_155),.data_out(wire_d0_156),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10157(.data_in(wire_d0_156),.data_out(wire_d0_157),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10158(.data_in(wire_d0_157),.data_out(wire_d0_158),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10159(.data_in(wire_d0_158),.data_out(wire_d0_159),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10160(.data_in(wire_d0_159),.data_out(wire_d0_160),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10161(.data_in(wire_d0_160),.data_out(wire_d0_161),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10162(.data_in(wire_d0_161),.data_out(wire_d0_162),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10163(.data_in(wire_d0_162),.data_out(wire_d0_163),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10164(.data_in(wire_d0_163),.data_out(wire_d0_164),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10165(.data_in(wire_d0_164),.data_out(wire_d0_165),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10166(.data_in(wire_d0_165),.data_out(wire_d0_166),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10167(.data_in(wire_d0_166),.data_out(wire_d0_167),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10168(.data_in(wire_d0_167),.data_out(wire_d0_168),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10169(.data_in(wire_d0_168),.data_out(wire_d0_169),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10170(.data_in(wire_d0_169),.data_out(wire_d0_170),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10171(.data_in(wire_d0_170),.data_out(wire_d0_171),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10172(.data_in(wire_d0_171),.data_out(wire_d0_172),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10173(.data_in(wire_d0_172),.data_out(wire_d0_173),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10174(.data_in(wire_d0_173),.data_out(wire_d0_174),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10175(.data_in(wire_d0_174),.data_out(wire_d0_175),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10176(.data_in(wire_d0_175),.data_out(wire_d0_176),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10177(.data_in(wire_d0_176),.data_out(wire_d0_177),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10178(.data_in(wire_d0_177),.data_out(wire_d0_178),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10179(.data_in(wire_d0_178),.data_out(wire_d0_179),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10180(.data_in(wire_d0_179),.data_out(wire_d0_180),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10181(.data_in(wire_d0_180),.data_out(wire_d0_181),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10182(.data_in(wire_d0_181),.data_out(wire_d0_182),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10183(.data_in(wire_d0_182),.data_out(wire_d0_183),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10184(.data_in(wire_d0_183),.data_out(wire_d0_184),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10185(.data_in(wire_d0_184),.data_out(wire_d0_185),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10186(.data_in(wire_d0_185),.data_out(wire_d0_186),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10187(.data_in(wire_d0_186),.data_out(wire_d0_187),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10188(.data_in(wire_d0_187),.data_out(wire_d0_188),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10189(.data_in(wire_d0_188),.data_out(wire_d0_189),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10190(.data_in(wire_d0_189),.data_out(wire_d0_190),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10191(.data_in(wire_d0_190),.data_out(wire_d0_191),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10192(.data_in(wire_d0_191),.data_out(wire_d0_192),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10193(.data_in(wire_d0_192),.data_out(wire_d0_193),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10194(.data_in(wire_d0_193),.data_out(wire_d0_194),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10195(.data_in(wire_d0_194),.data_out(wire_d0_195),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10196(.data_in(wire_d0_195),.data_out(wire_d0_196),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10197(.data_in(wire_d0_196),.data_out(wire_d0_197),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10198(.data_in(wire_d0_197),.data_out(wire_d0_198),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10199(.data_in(wire_d0_198),.data_out(d_out0),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance210(.data_in(d_in1),.data_out(wire_d1_0),.clk(clk),.rst(rst));            //channel 2
	encoder #(.WIDTH(WIDTH)) encoder_instance211(.data_in(wire_d1_0),.data_out(wire_d1_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212(.data_in(wire_d1_1),.data_out(wire_d1_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance213(.data_in(wire_d1_2),.data_out(wire_d1_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance214(.data_in(wire_d1_3),.data_out(wire_d1_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance215(.data_in(wire_d1_4),.data_out(wire_d1_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance216(.data_in(wire_d1_5),.data_out(wire_d1_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance217(.data_in(wire_d1_6),.data_out(wire_d1_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance218(.data_in(wire_d1_7),.data_out(wire_d1_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance219(.data_in(wire_d1_8),.data_out(wire_d1_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2110(.data_in(wire_d1_9),.data_out(wire_d1_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2111(.data_in(wire_d1_10),.data_out(wire_d1_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2112(.data_in(wire_d1_11),.data_out(wire_d1_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2113(.data_in(wire_d1_12),.data_out(wire_d1_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2114(.data_in(wire_d1_13),.data_out(wire_d1_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2115(.data_in(wire_d1_14),.data_out(wire_d1_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2116(.data_in(wire_d1_15),.data_out(wire_d1_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2117(.data_in(wire_d1_16),.data_out(wire_d1_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2118(.data_in(wire_d1_17),.data_out(wire_d1_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2119(.data_in(wire_d1_18),.data_out(wire_d1_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2120(.data_in(wire_d1_19),.data_out(wire_d1_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2121(.data_in(wire_d1_20),.data_out(wire_d1_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2122(.data_in(wire_d1_21),.data_out(wire_d1_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2123(.data_in(wire_d1_22),.data_out(wire_d1_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2124(.data_in(wire_d1_23),.data_out(wire_d1_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2125(.data_in(wire_d1_24),.data_out(wire_d1_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2126(.data_in(wire_d1_25),.data_out(wire_d1_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2127(.data_in(wire_d1_26),.data_out(wire_d1_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2128(.data_in(wire_d1_27),.data_out(wire_d1_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2129(.data_in(wire_d1_28),.data_out(wire_d1_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2130(.data_in(wire_d1_29),.data_out(wire_d1_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2131(.data_in(wire_d1_30),.data_out(wire_d1_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2132(.data_in(wire_d1_31),.data_out(wire_d1_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2133(.data_in(wire_d1_32),.data_out(wire_d1_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2134(.data_in(wire_d1_33),.data_out(wire_d1_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2135(.data_in(wire_d1_34),.data_out(wire_d1_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2136(.data_in(wire_d1_35),.data_out(wire_d1_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2137(.data_in(wire_d1_36),.data_out(wire_d1_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2138(.data_in(wire_d1_37),.data_out(wire_d1_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2139(.data_in(wire_d1_38),.data_out(wire_d1_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2140(.data_in(wire_d1_39),.data_out(wire_d1_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2141(.data_in(wire_d1_40),.data_out(wire_d1_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2142(.data_in(wire_d1_41),.data_out(wire_d1_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2143(.data_in(wire_d1_42),.data_out(wire_d1_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2144(.data_in(wire_d1_43),.data_out(wire_d1_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2145(.data_in(wire_d1_44),.data_out(wire_d1_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2146(.data_in(wire_d1_45),.data_out(wire_d1_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2147(.data_in(wire_d1_46),.data_out(wire_d1_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2148(.data_in(wire_d1_47),.data_out(wire_d1_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2149(.data_in(wire_d1_48),.data_out(wire_d1_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2150(.data_in(wire_d1_49),.data_out(wire_d1_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2151(.data_in(wire_d1_50),.data_out(wire_d1_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2152(.data_in(wire_d1_51),.data_out(wire_d1_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2153(.data_in(wire_d1_52),.data_out(wire_d1_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2154(.data_in(wire_d1_53),.data_out(wire_d1_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2155(.data_in(wire_d1_54),.data_out(wire_d1_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2156(.data_in(wire_d1_55),.data_out(wire_d1_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2157(.data_in(wire_d1_56),.data_out(wire_d1_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2158(.data_in(wire_d1_57),.data_out(wire_d1_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2159(.data_in(wire_d1_58),.data_out(wire_d1_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2160(.data_in(wire_d1_59),.data_out(wire_d1_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2161(.data_in(wire_d1_60),.data_out(wire_d1_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2162(.data_in(wire_d1_61),.data_out(wire_d1_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2163(.data_in(wire_d1_62),.data_out(wire_d1_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2164(.data_in(wire_d1_63),.data_out(wire_d1_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2165(.data_in(wire_d1_64),.data_out(wire_d1_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2166(.data_in(wire_d1_65),.data_out(wire_d1_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2167(.data_in(wire_d1_66),.data_out(wire_d1_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2168(.data_in(wire_d1_67),.data_out(wire_d1_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2169(.data_in(wire_d1_68),.data_out(wire_d1_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2170(.data_in(wire_d1_69),.data_out(wire_d1_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2171(.data_in(wire_d1_70),.data_out(wire_d1_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2172(.data_in(wire_d1_71),.data_out(wire_d1_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2173(.data_in(wire_d1_72),.data_out(wire_d1_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2174(.data_in(wire_d1_73),.data_out(wire_d1_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2175(.data_in(wire_d1_74),.data_out(wire_d1_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2176(.data_in(wire_d1_75),.data_out(wire_d1_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2177(.data_in(wire_d1_76),.data_out(wire_d1_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2178(.data_in(wire_d1_77),.data_out(wire_d1_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2179(.data_in(wire_d1_78),.data_out(wire_d1_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2180(.data_in(wire_d1_79),.data_out(wire_d1_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2181(.data_in(wire_d1_80),.data_out(wire_d1_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2182(.data_in(wire_d1_81),.data_out(wire_d1_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2183(.data_in(wire_d1_82),.data_out(wire_d1_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2184(.data_in(wire_d1_83),.data_out(wire_d1_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2185(.data_in(wire_d1_84),.data_out(wire_d1_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2186(.data_in(wire_d1_85),.data_out(wire_d1_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2187(.data_in(wire_d1_86),.data_out(wire_d1_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2188(.data_in(wire_d1_87),.data_out(wire_d1_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2189(.data_in(wire_d1_88),.data_out(wire_d1_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2190(.data_in(wire_d1_89),.data_out(wire_d1_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2191(.data_in(wire_d1_90),.data_out(wire_d1_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2192(.data_in(wire_d1_91),.data_out(wire_d1_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2193(.data_in(wire_d1_92),.data_out(wire_d1_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2194(.data_in(wire_d1_93),.data_out(wire_d1_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2195(.data_in(wire_d1_94),.data_out(wire_d1_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2196(.data_in(wire_d1_95),.data_out(wire_d1_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2197(.data_in(wire_d1_96),.data_out(wire_d1_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2198(.data_in(wire_d1_97),.data_out(wire_d1_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2199(.data_in(wire_d1_98),.data_out(wire_d1_99),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21100(.data_in(wire_d1_99),.data_out(wire_d1_100),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21101(.data_in(wire_d1_100),.data_out(wire_d1_101),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21102(.data_in(wire_d1_101),.data_out(wire_d1_102),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21103(.data_in(wire_d1_102),.data_out(wire_d1_103),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21104(.data_in(wire_d1_103),.data_out(wire_d1_104),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21105(.data_in(wire_d1_104),.data_out(wire_d1_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21106(.data_in(wire_d1_105),.data_out(wire_d1_106),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21107(.data_in(wire_d1_106),.data_out(wire_d1_107),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21108(.data_in(wire_d1_107),.data_out(wire_d1_108),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21109(.data_in(wire_d1_108),.data_out(wire_d1_109),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21110(.data_in(wire_d1_109),.data_out(wire_d1_110),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21111(.data_in(wire_d1_110),.data_out(wire_d1_111),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21112(.data_in(wire_d1_111),.data_out(wire_d1_112),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21113(.data_in(wire_d1_112),.data_out(wire_d1_113),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21114(.data_in(wire_d1_113),.data_out(wire_d1_114),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21115(.data_in(wire_d1_114),.data_out(wire_d1_115),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21116(.data_in(wire_d1_115),.data_out(wire_d1_116),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21117(.data_in(wire_d1_116),.data_out(wire_d1_117),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21118(.data_in(wire_d1_117),.data_out(wire_d1_118),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21119(.data_in(wire_d1_118),.data_out(wire_d1_119),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21120(.data_in(wire_d1_119),.data_out(wire_d1_120),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21121(.data_in(wire_d1_120),.data_out(wire_d1_121),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21122(.data_in(wire_d1_121),.data_out(wire_d1_122),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21123(.data_in(wire_d1_122),.data_out(wire_d1_123),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21124(.data_in(wire_d1_123),.data_out(wire_d1_124),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21125(.data_in(wire_d1_124),.data_out(wire_d1_125),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21126(.data_in(wire_d1_125),.data_out(wire_d1_126),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21127(.data_in(wire_d1_126),.data_out(wire_d1_127),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21128(.data_in(wire_d1_127),.data_out(wire_d1_128),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21129(.data_in(wire_d1_128),.data_out(wire_d1_129),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21130(.data_in(wire_d1_129),.data_out(wire_d1_130),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21131(.data_in(wire_d1_130),.data_out(wire_d1_131),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21132(.data_in(wire_d1_131),.data_out(wire_d1_132),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21133(.data_in(wire_d1_132),.data_out(wire_d1_133),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21134(.data_in(wire_d1_133),.data_out(wire_d1_134),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21135(.data_in(wire_d1_134),.data_out(wire_d1_135),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21136(.data_in(wire_d1_135),.data_out(wire_d1_136),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21137(.data_in(wire_d1_136),.data_out(wire_d1_137),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21138(.data_in(wire_d1_137),.data_out(wire_d1_138),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21139(.data_in(wire_d1_138),.data_out(wire_d1_139),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21140(.data_in(wire_d1_139),.data_out(wire_d1_140),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21141(.data_in(wire_d1_140),.data_out(wire_d1_141),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21142(.data_in(wire_d1_141),.data_out(wire_d1_142),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21143(.data_in(wire_d1_142),.data_out(wire_d1_143),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21144(.data_in(wire_d1_143),.data_out(wire_d1_144),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21145(.data_in(wire_d1_144),.data_out(wire_d1_145),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21146(.data_in(wire_d1_145),.data_out(wire_d1_146),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21147(.data_in(wire_d1_146),.data_out(wire_d1_147),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21148(.data_in(wire_d1_147),.data_out(wire_d1_148),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21149(.data_in(wire_d1_148),.data_out(wire_d1_149),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21150(.data_in(wire_d1_149),.data_out(wire_d1_150),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21151(.data_in(wire_d1_150),.data_out(wire_d1_151),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21152(.data_in(wire_d1_151),.data_out(wire_d1_152),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21153(.data_in(wire_d1_152),.data_out(wire_d1_153),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21154(.data_in(wire_d1_153),.data_out(wire_d1_154),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21155(.data_in(wire_d1_154),.data_out(wire_d1_155),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21156(.data_in(wire_d1_155),.data_out(wire_d1_156),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21157(.data_in(wire_d1_156),.data_out(wire_d1_157),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21158(.data_in(wire_d1_157),.data_out(wire_d1_158),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21159(.data_in(wire_d1_158),.data_out(wire_d1_159),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21160(.data_in(wire_d1_159),.data_out(wire_d1_160),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21161(.data_in(wire_d1_160),.data_out(wire_d1_161),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21162(.data_in(wire_d1_161),.data_out(wire_d1_162),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21163(.data_in(wire_d1_162),.data_out(wire_d1_163),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21164(.data_in(wire_d1_163),.data_out(wire_d1_164),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21165(.data_in(wire_d1_164),.data_out(wire_d1_165),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21166(.data_in(wire_d1_165),.data_out(wire_d1_166),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21167(.data_in(wire_d1_166),.data_out(wire_d1_167),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21168(.data_in(wire_d1_167),.data_out(wire_d1_168),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21169(.data_in(wire_d1_168),.data_out(wire_d1_169),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21170(.data_in(wire_d1_169),.data_out(wire_d1_170),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21171(.data_in(wire_d1_170),.data_out(wire_d1_171),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21172(.data_in(wire_d1_171),.data_out(wire_d1_172),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21173(.data_in(wire_d1_172),.data_out(wire_d1_173),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21174(.data_in(wire_d1_173),.data_out(wire_d1_174),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21175(.data_in(wire_d1_174),.data_out(wire_d1_175),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21176(.data_in(wire_d1_175),.data_out(wire_d1_176),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21177(.data_in(wire_d1_176),.data_out(wire_d1_177),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21178(.data_in(wire_d1_177),.data_out(wire_d1_178),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21179(.data_in(wire_d1_178),.data_out(wire_d1_179),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21180(.data_in(wire_d1_179),.data_out(wire_d1_180),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21181(.data_in(wire_d1_180),.data_out(wire_d1_181),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21182(.data_in(wire_d1_181),.data_out(wire_d1_182),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21183(.data_in(wire_d1_182),.data_out(wire_d1_183),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21184(.data_in(wire_d1_183),.data_out(wire_d1_184),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21185(.data_in(wire_d1_184),.data_out(wire_d1_185),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21186(.data_in(wire_d1_185),.data_out(wire_d1_186),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21187(.data_in(wire_d1_186),.data_out(wire_d1_187),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21188(.data_in(wire_d1_187),.data_out(wire_d1_188),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21189(.data_in(wire_d1_188),.data_out(wire_d1_189),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21190(.data_in(wire_d1_189),.data_out(wire_d1_190),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21191(.data_in(wire_d1_190),.data_out(wire_d1_191),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21192(.data_in(wire_d1_191),.data_out(wire_d1_192),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21193(.data_in(wire_d1_192),.data_out(wire_d1_193),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21194(.data_in(wire_d1_193),.data_out(wire_d1_194),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21195(.data_in(wire_d1_194),.data_out(wire_d1_195),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21196(.data_in(wire_d1_195),.data_out(wire_d1_196),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21197(.data_in(wire_d1_196),.data_out(wire_d1_197),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21198(.data_in(wire_d1_197),.data_out(wire_d1_198),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21199(.data_in(wire_d1_198),.data_out(d_out1),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance320(.data_in(d_in2),.data_out(wire_d2_0),.clk(clk),.rst(rst));            //channel 3
	encoder #(.WIDTH(WIDTH)) encoder_instance321(.data_in(wire_d2_0),.data_out(wire_d2_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance322(.data_in(wire_d2_1),.data_out(wire_d2_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323(.data_in(wire_d2_2),.data_out(wire_d2_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance324(.data_in(wire_d2_3),.data_out(wire_d2_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance325(.data_in(wire_d2_4),.data_out(wire_d2_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance326(.data_in(wire_d2_5),.data_out(wire_d2_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance327(.data_in(wire_d2_6),.data_out(wire_d2_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance328(.data_in(wire_d2_7),.data_out(wire_d2_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance329(.data_in(wire_d2_8),.data_out(wire_d2_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3210(.data_in(wire_d2_9),.data_out(wire_d2_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3211(.data_in(wire_d2_10),.data_out(wire_d2_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3212(.data_in(wire_d2_11),.data_out(wire_d2_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3213(.data_in(wire_d2_12),.data_out(wire_d2_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3214(.data_in(wire_d2_13),.data_out(wire_d2_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3215(.data_in(wire_d2_14),.data_out(wire_d2_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3216(.data_in(wire_d2_15),.data_out(wire_d2_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3217(.data_in(wire_d2_16),.data_out(wire_d2_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3218(.data_in(wire_d2_17),.data_out(wire_d2_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3219(.data_in(wire_d2_18),.data_out(wire_d2_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3220(.data_in(wire_d2_19),.data_out(wire_d2_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3221(.data_in(wire_d2_20),.data_out(wire_d2_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3222(.data_in(wire_d2_21),.data_out(wire_d2_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3223(.data_in(wire_d2_22),.data_out(wire_d2_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3224(.data_in(wire_d2_23),.data_out(wire_d2_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3225(.data_in(wire_d2_24),.data_out(wire_d2_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3226(.data_in(wire_d2_25),.data_out(wire_d2_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3227(.data_in(wire_d2_26),.data_out(wire_d2_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3228(.data_in(wire_d2_27),.data_out(wire_d2_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3229(.data_in(wire_d2_28),.data_out(wire_d2_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3230(.data_in(wire_d2_29),.data_out(wire_d2_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3231(.data_in(wire_d2_30),.data_out(wire_d2_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3232(.data_in(wire_d2_31),.data_out(wire_d2_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3233(.data_in(wire_d2_32),.data_out(wire_d2_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3234(.data_in(wire_d2_33),.data_out(wire_d2_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3235(.data_in(wire_d2_34),.data_out(wire_d2_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3236(.data_in(wire_d2_35),.data_out(wire_d2_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3237(.data_in(wire_d2_36),.data_out(wire_d2_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3238(.data_in(wire_d2_37),.data_out(wire_d2_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3239(.data_in(wire_d2_38),.data_out(wire_d2_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3240(.data_in(wire_d2_39),.data_out(wire_d2_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3241(.data_in(wire_d2_40),.data_out(wire_d2_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3242(.data_in(wire_d2_41),.data_out(wire_d2_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3243(.data_in(wire_d2_42),.data_out(wire_d2_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3244(.data_in(wire_d2_43),.data_out(wire_d2_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3245(.data_in(wire_d2_44),.data_out(wire_d2_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3246(.data_in(wire_d2_45),.data_out(wire_d2_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3247(.data_in(wire_d2_46),.data_out(wire_d2_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3248(.data_in(wire_d2_47),.data_out(wire_d2_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3249(.data_in(wire_d2_48),.data_out(wire_d2_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3250(.data_in(wire_d2_49),.data_out(wire_d2_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3251(.data_in(wire_d2_50),.data_out(wire_d2_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3252(.data_in(wire_d2_51),.data_out(wire_d2_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3253(.data_in(wire_d2_52),.data_out(wire_d2_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3254(.data_in(wire_d2_53),.data_out(wire_d2_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3255(.data_in(wire_d2_54),.data_out(wire_d2_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3256(.data_in(wire_d2_55),.data_out(wire_d2_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3257(.data_in(wire_d2_56),.data_out(wire_d2_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3258(.data_in(wire_d2_57),.data_out(wire_d2_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3259(.data_in(wire_d2_58),.data_out(wire_d2_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3260(.data_in(wire_d2_59),.data_out(wire_d2_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3261(.data_in(wire_d2_60),.data_out(wire_d2_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3262(.data_in(wire_d2_61),.data_out(wire_d2_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3263(.data_in(wire_d2_62),.data_out(wire_d2_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3264(.data_in(wire_d2_63),.data_out(wire_d2_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3265(.data_in(wire_d2_64),.data_out(wire_d2_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3266(.data_in(wire_d2_65),.data_out(wire_d2_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3267(.data_in(wire_d2_66),.data_out(wire_d2_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3268(.data_in(wire_d2_67),.data_out(wire_d2_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3269(.data_in(wire_d2_68),.data_out(wire_d2_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3270(.data_in(wire_d2_69),.data_out(wire_d2_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3271(.data_in(wire_d2_70),.data_out(wire_d2_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3272(.data_in(wire_d2_71),.data_out(wire_d2_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3273(.data_in(wire_d2_72),.data_out(wire_d2_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3274(.data_in(wire_d2_73),.data_out(wire_d2_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3275(.data_in(wire_d2_74),.data_out(wire_d2_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3276(.data_in(wire_d2_75),.data_out(wire_d2_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3277(.data_in(wire_d2_76),.data_out(wire_d2_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3278(.data_in(wire_d2_77),.data_out(wire_d2_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3279(.data_in(wire_d2_78),.data_out(wire_d2_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3280(.data_in(wire_d2_79),.data_out(wire_d2_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3281(.data_in(wire_d2_80),.data_out(wire_d2_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3282(.data_in(wire_d2_81),.data_out(wire_d2_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3283(.data_in(wire_d2_82),.data_out(wire_d2_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3284(.data_in(wire_d2_83),.data_out(wire_d2_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3285(.data_in(wire_d2_84),.data_out(wire_d2_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3286(.data_in(wire_d2_85),.data_out(wire_d2_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3287(.data_in(wire_d2_86),.data_out(wire_d2_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3288(.data_in(wire_d2_87),.data_out(wire_d2_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3289(.data_in(wire_d2_88),.data_out(wire_d2_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3290(.data_in(wire_d2_89),.data_out(wire_d2_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3291(.data_in(wire_d2_90),.data_out(wire_d2_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3292(.data_in(wire_d2_91),.data_out(wire_d2_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3293(.data_in(wire_d2_92),.data_out(wire_d2_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3294(.data_in(wire_d2_93),.data_out(wire_d2_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3295(.data_in(wire_d2_94),.data_out(wire_d2_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3296(.data_in(wire_d2_95),.data_out(wire_d2_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3297(.data_in(wire_d2_96),.data_out(wire_d2_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3298(.data_in(wire_d2_97),.data_out(wire_d2_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3299(.data_in(wire_d2_98),.data_out(wire_d2_99),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32100(.data_in(wire_d2_99),.data_out(wire_d2_100),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32101(.data_in(wire_d2_100),.data_out(wire_d2_101),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32102(.data_in(wire_d2_101),.data_out(wire_d2_102),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32103(.data_in(wire_d2_102),.data_out(wire_d2_103),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32104(.data_in(wire_d2_103),.data_out(wire_d2_104),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32105(.data_in(wire_d2_104),.data_out(wire_d2_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32106(.data_in(wire_d2_105),.data_out(wire_d2_106),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32107(.data_in(wire_d2_106),.data_out(wire_d2_107),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32108(.data_in(wire_d2_107),.data_out(wire_d2_108),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32109(.data_in(wire_d2_108),.data_out(wire_d2_109),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32110(.data_in(wire_d2_109),.data_out(wire_d2_110),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32111(.data_in(wire_d2_110),.data_out(wire_d2_111),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32112(.data_in(wire_d2_111),.data_out(wire_d2_112),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32113(.data_in(wire_d2_112),.data_out(wire_d2_113),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32114(.data_in(wire_d2_113),.data_out(wire_d2_114),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32115(.data_in(wire_d2_114),.data_out(wire_d2_115),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32116(.data_in(wire_d2_115),.data_out(wire_d2_116),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32117(.data_in(wire_d2_116),.data_out(wire_d2_117),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32118(.data_in(wire_d2_117),.data_out(wire_d2_118),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32119(.data_in(wire_d2_118),.data_out(wire_d2_119),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32120(.data_in(wire_d2_119),.data_out(wire_d2_120),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32121(.data_in(wire_d2_120),.data_out(wire_d2_121),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32122(.data_in(wire_d2_121),.data_out(wire_d2_122),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32123(.data_in(wire_d2_122),.data_out(wire_d2_123),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32124(.data_in(wire_d2_123),.data_out(wire_d2_124),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32125(.data_in(wire_d2_124),.data_out(wire_d2_125),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32126(.data_in(wire_d2_125),.data_out(wire_d2_126),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32127(.data_in(wire_d2_126),.data_out(wire_d2_127),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32128(.data_in(wire_d2_127),.data_out(wire_d2_128),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32129(.data_in(wire_d2_128),.data_out(wire_d2_129),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32130(.data_in(wire_d2_129),.data_out(wire_d2_130),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32131(.data_in(wire_d2_130),.data_out(wire_d2_131),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32132(.data_in(wire_d2_131),.data_out(wire_d2_132),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32133(.data_in(wire_d2_132),.data_out(wire_d2_133),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32134(.data_in(wire_d2_133),.data_out(wire_d2_134),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32135(.data_in(wire_d2_134),.data_out(wire_d2_135),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32136(.data_in(wire_d2_135),.data_out(wire_d2_136),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32137(.data_in(wire_d2_136),.data_out(wire_d2_137),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32138(.data_in(wire_d2_137),.data_out(wire_d2_138),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32139(.data_in(wire_d2_138),.data_out(wire_d2_139),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32140(.data_in(wire_d2_139),.data_out(wire_d2_140),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32141(.data_in(wire_d2_140),.data_out(wire_d2_141),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32142(.data_in(wire_d2_141),.data_out(wire_d2_142),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32143(.data_in(wire_d2_142),.data_out(wire_d2_143),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32144(.data_in(wire_d2_143),.data_out(wire_d2_144),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32145(.data_in(wire_d2_144),.data_out(wire_d2_145),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32146(.data_in(wire_d2_145),.data_out(wire_d2_146),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32147(.data_in(wire_d2_146),.data_out(wire_d2_147),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32148(.data_in(wire_d2_147),.data_out(wire_d2_148),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32149(.data_in(wire_d2_148),.data_out(wire_d2_149),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32150(.data_in(wire_d2_149),.data_out(wire_d2_150),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32151(.data_in(wire_d2_150),.data_out(wire_d2_151),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32152(.data_in(wire_d2_151),.data_out(wire_d2_152),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32153(.data_in(wire_d2_152),.data_out(wire_d2_153),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32154(.data_in(wire_d2_153),.data_out(wire_d2_154),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32155(.data_in(wire_d2_154),.data_out(wire_d2_155),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32156(.data_in(wire_d2_155),.data_out(wire_d2_156),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32157(.data_in(wire_d2_156),.data_out(wire_d2_157),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32158(.data_in(wire_d2_157),.data_out(wire_d2_158),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32159(.data_in(wire_d2_158),.data_out(wire_d2_159),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32160(.data_in(wire_d2_159),.data_out(wire_d2_160),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32161(.data_in(wire_d2_160),.data_out(wire_d2_161),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32162(.data_in(wire_d2_161),.data_out(wire_d2_162),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32163(.data_in(wire_d2_162),.data_out(wire_d2_163),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32164(.data_in(wire_d2_163),.data_out(wire_d2_164),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32165(.data_in(wire_d2_164),.data_out(wire_d2_165),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32166(.data_in(wire_d2_165),.data_out(wire_d2_166),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32167(.data_in(wire_d2_166),.data_out(wire_d2_167),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32168(.data_in(wire_d2_167),.data_out(wire_d2_168),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32169(.data_in(wire_d2_168),.data_out(wire_d2_169),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32170(.data_in(wire_d2_169),.data_out(wire_d2_170),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32171(.data_in(wire_d2_170),.data_out(wire_d2_171),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32172(.data_in(wire_d2_171),.data_out(wire_d2_172),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32173(.data_in(wire_d2_172),.data_out(wire_d2_173),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32174(.data_in(wire_d2_173),.data_out(wire_d2_174),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32175(.data_in(wire_d2_174),.data_out(wire_d2_175),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32176(.data_in(wire_d2_175),.data_out(wire_d2_176),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32177(.data_in(wire_d2_176),.data_out(wire_d2_177),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32178(.data_in(wire_d2_177),.data_out(wire_d2_178),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32179(.data_in(wire_d2_178),.data_out(wire_d2_179),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32180(.data_in(wire_d2_179),.data_out(wire_d2_180),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32181(.data_in(wire_d2_180),.data_out(wire_d2_181),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32182(.data_in(wire_d2_181),.data_out(wire_d2_182),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32183(.data_in(wire_d2_182),.data_out(wire_d2_183),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32184(.data_in(wire_d2_183),.data_out(wire_d2_184),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32185(.data_in(wire_d2_184),.data_out(wire_d2_185),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32186(.data_in(wire_d2_185),.data_out(wire_d2_186),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32187(.data_in(wire_d2_186),.data_out(wire_d2_187),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32188(.data_in(wire_d2_187),.data_out(wire_d2_188),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32189(.data_in(wire_d2_188),.data_out(wire_d2_189),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32190(.data_in(wire_d2_189),.data_out(wire_d2_190),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32191(.data_in(wire_d2_190),.data_out(wire_d2_191),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32192(.data_in(wire_d2_191),.data_out(wire_d2_192),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32193(.data_in(wire_d2_192),.data_out(wire_d2_193),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32194(.data_in(wire_d2_193),.data_out(wire_d2_194),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32195(.data_in(wire_d2_194),.data_out(wire_d2_195),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32196(.data_in(wire_d2_195),.data_out(wire_d2_196),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32197(.data_in(wire_d2_196),.data_out(wire_d2_197),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32198(.data_in(wire_d2_197),.data_out(wire_d2_198),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32199(.data_in(wire_d2_198),.data_out(d_out2),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance430(.data_in(d_in3),.data_out(wire_d3_0),.clk(clk),.rst(rst));            //channel 4
	encoder #(.WIDTH(WIDTH)) encoder_instance431(.data_in(wire_d3_0),.data_out(wire_d3_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance432(.data_in(wire_d3_1),.data_out(wire_d3_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance433(.data_in(wire_d3_2),.data_out(wire_d3_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434(.data_in(wire_d3_3),.data_out(wire_d3_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance435(.data_in(wire_d3_4),.data_out(wire_d3_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance436(.data_in(wire_d3_5),.data_out(wire_d3_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance437(.data_in(wire_d3_6),.data_out(wire_d3_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance438(.data_in(wire_d3_7),.data_out(wire_d3_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance439(.data_in(wire_d3_8),.data_out(wire_d3_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4310(.data_in(wire_d3_9),.data_out(wire_d3_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4311(.data_in(wire_d3_10),.data_out(wire_d3_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4312(.data_in(wire_d3_11),.data_out(wire_d3_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4313(.data_in(wire_d3_12),.data_out(wire_d3_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4314(.data_in(wire_d3_13),.data_out(wire_d3_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4315(.data_in(wire_d3_14),.data_out(wire_d3_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4316(.data_in(wire_d3_15),.data_out(wire_d3_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4317(.data_in(wire_d3_16),.data_out(wire_d3_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4318(.data_in(wire_d3_17),.data_out(wire_d3_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4319(.data_in(wire_d3_18),.data_out(wire_d3_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4320(.data_in(wire_d3_19),.data_out(wire_d3_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4321(.data_in(wire_d3_20),.data_out(wire_d3_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4322(.data_in(wire_d3_21),.data_out(wire_d3_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4323(.data_in(wire_d3_22),.data_out(wire_d3_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4324(.data_in(wire_d3_23),.data_out(wire_d3_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4325(.data_in(wire_d3_24),.data_out(wire_d3_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4326(.data_in(wire_d3_25),.data_out(wire_d3_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4327(.data_in(wire_d3_26),.data_out(wire_d3_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4328(.data_in(wire_d3_27),.data_out(wire_d3_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4329(.data_in(wire_d3_28),.data_out(wire_d3_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4330(.data_in(wire_d3_29),.data_out(wire_d3_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4331(.data_in(wire_d3_30),.data_out(wire_d3_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4332(.data_in(wire_d3_31),.data_out(wire_d3_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4333(.data_in(wire_d3_32),.data_out(wire_d3_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4334(.data_in(wire_d3_33),.data_out(wire_d3_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4335(.data_in(wire_d3_34),.data_out(wire_d3_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4336(.data_in(wire_d3_35),.data_out(wire_d3_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4337(.data_in(wire_d3_36),.data_out(wire_d3_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4338(.data_in(wire_d3_37),.data_out(wire_d3_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4339(.data_in(wire_d3_38),.data_out(wire_d3_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4340(.data_in(wire_d3_39),.data_out(wire_d3_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4341(.data_in(wire_d3_40),.data_out(wire_d3_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4342(.data_in(wire_d3_41),.data_out(wire_d3_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4343(.data_in(wire_d3_42),.data_out(wire_d3_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4344(.data_in(wire_d3_43),.data_out(wire_d3_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4345(.data_in(wire_d3_44),.data_out(wire_d3_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4346(.data_in(wire_d3_45),.data_out(wire_d3_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4347(.data_in(wire_d3_46),.data_out(wire_d3_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4348(.data_in(wire_d3_47),.data_out(wire_d3_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4349(.data_in(wire_d3_48),.data_out(wire_d3_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4350(.data_in(wire_d3_49),.data_out(wire_d3_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4351(.data_in(wire_d3_50),.data_out(wire_d3_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4352(.data_in(wire_d3_51),.data_out(wire_d3_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4353(.data_in(wire_d3_52),.data_out(wire_d3_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4354(.data_in(wire_d3_53),.data_out(wire_d3_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4355(.data_in(wire_d3_54),.data_out(wire_d3_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4356(.data_in(wire_d3_55),.data_out(wire_d3_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4357(.data_in(wire_d3_56),.data_out(wire_d3_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4358(.data_in(wire_d3_57),.data_out(wire_d3_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4359(.data_in(wire_d3_58),.data_out(wire_d3_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4360(.data_in(wire_d3_59),.data_out(wire_d3_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4361(.data_in(wire_d3_60),.data_out(wire_d3_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4362(.data_in(wire_d3_61),.data_out(wire_d3_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4363(.data_in(wire_d3_62),.data_out(wire_d3_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4364(.data_in(wire_d3_63),.data_out(wire_d3_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4365(.data_in(wire_d3_64),.data_out(wire_d3_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4366(.data_in(wire_d3_65),.data_out(wire_d3_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4367(.data_in(wire_d3_66),.data_out(wire_d3_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4368(.data_in(wire_d3_67),.data_out(wire_d3_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4369(.data_in(wire_d3_68),.data_out(wire_d3_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4370(.data_in(wire_d3_69),.data_out(wire_d3_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4371(.data_in(wire_d3_70),.data_out(wire_d3_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4372(.data_in(wire_d3_71),.data_out(wire_d3_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4373(.data_in(wire_d3_72),.data_out(wire_d3_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4374(.data_in(wire_d3_73),.data_out(wire_d3_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4375(.data_in(wire_d3_74),.data_out(wire_d3_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4376(.data_in(wire_d3_75),.data_out(wire_d3_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4377(.data_in(wire_d3_76),.data_out(wire_d3_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4378(.data_in(wire_d3_77),.data_out(wire_d3_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4379(.data_in(wire_d3_78),.data_out(wire_d3_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4380(.data_in(wire_d3_79),.data_out(wire_d3_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4381(.data_in(wire_d3_80),.data_out(wire_d3_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4382(.data_in(wire_d3_81),.data_out(wire_d3_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4383(.data_in(wire_d3_82),.data_out(wire_d3_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4384(.data_in(wire_d3_83),.data_out(wire_d3_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4385(.data_in(wire_d3_84),.data_out(wire_d3_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4386(.data_in(wire_d3_85),.data_out(wire_d3_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4387(.data_in(wire_d3_86),.data_out(wire_d3_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4388(.data_in(wire_d3_87),.data_out(wire_d3_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4389(.data_in(wire_d3_88),.data_out(wire_d3_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4390(.data_in(wire_d3_89),.data_out(wire_d3_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4391(.data_in(wire_d3_90),.data_out(wire_d3_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4392(.data_in(wire_d3_91),.data_out(wire_d3_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4393(.data_in(wire_d3_92),.data_out(wire_d3_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4394(.data_in(wire_d3_93),.data_out(wire_d3_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4395(.data_in(wire_d3_94),.data_out(wire_d3_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4396(.data_in(wire_d3_95),.data_out(wire_d3_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4397(.data_in(wire_d3_96),.data_out(wire_d3_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4398(.data_in(wire_d3_97),.data_out(wire_d3_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4399(.data_in(wire_d3_98),.data_out(wire_d3_99),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43100(.data_in(wire_d3_99),.data_out(wire_d3_100),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43101(.data_in(wire_d3_100),.data_out(wire_d3_101),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43102(.data_in(wire_d3_101),.data_out(wire_d3_102),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43103(.data_in(wire_d3_102),.data_out(wire_d3_103),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43104(.data_in(wire_d3_103),.data_out(wire_d3_104),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43105(.data_in(wire_d3_104),.data_out(wire_d3_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43106(.data_in(wire_d3_105),.data_out(wire_d3_106),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43107(.data_in(wire_d3_106),.data_out(wire_d3_107),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43108(.data_in(wire_d3_107),.data_out(wire_d3_108),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43109(.data_in(wire_d3_108),.data_out(wire_d3_109),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43110(.data_in(wire_d3_109),.data_out(wire_d3_110),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43111(.data_in(wire_d3_110),.data_out(wire_d3_111),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43112(.data_in(wire_d3_111),.data_out(wire_d3_112),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43113(.data_in(wire_d3_112),.data_out(wire_d3_113),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43114(.data_in(wire_d3_113),.data_out(wire_d3_114),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43115(.data_in(wire_d3_114),.data_out(wire_d3_115),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43116(.data_in(wire_d3_115),.data_out(wire_d3_116),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43117(.data_in(wire_d3_116),.data_out(wire_d3_117),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43118(.data_in(wire_d3_117),.data_out(wire_d3_118),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43119(.data_in(wire_d3_118),.data_out(wire_d3_119),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43120(.data_in(wire_d3_119),.data_out(wire_d3_120),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43121(.data_in(wire_d3_120),.data_out(wire_d3_121),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43122(.data_in(wire_d3_121),.data_out(wire_d3_122),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43123(.data_in(wire_d3_122),.data_out(wire_d3_123),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43124(.data_in(wire_d3_123),.data_out(wire_d3_124),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43125(.data_in(wire_d3_124),.data_out(wire_d3_125),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43126(.data_in(wire_d3_125),.data_out(wire_d3_126),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43127(.data_in(wire_d3_126),.data_out(wire_d3_127),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43128(.data_in(wire_d3_127),.data_out(wire_d3_128),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43129(.data_in(wire_d3_128),.data_out(wire_d3_129),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43130(.data_in(wire_d3_129),.data_out(wire_d3_130),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43131(.data_in(wire_d3_130),.data_out(wire_d3_131),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43132(.data_in(wire_d3_131),.data_out(wire_d3_132),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43133(.data_in(wire_d3_132),.data_out(wire_d3_133),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43134(.data_in(wire_d3_133),.data_out(wire_d3_134),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43135(.data_in(wire_d3_134),.data_out(wire_d3_135),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43136(.data_in(wire_d3_135),.data_out(wire_d3_136),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43137(.data_in(wire_d3_136),.data_out(wire_d3_137),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43138(.data_in(wire_d3_137),.data_out(wire_d3_138),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43139(.data_in(wire_d3_138),.data_out(wire_d3_139),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43140(.data_in(wire_d3_139),.data_out(wire_d3_140),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43141(.data_in(wire_d3_140),.data_out(wire_d3_141),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43142(.data_in(wire_d3_141),.data_out(wire_d3_142),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43143(.data_in(wire_d3_142),.data_out(wire_d3_143),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43144(.data_in(wire_d3_143),.data_out(wire_d3_144),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43145(.data_in(wire_d3_144),.data_out(wire_d3_145),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43146(.data_in(wire_d3_145),.data_out(wire_d3_146),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43147(.data_in(wire_d3_146),.data_out(wire_d3_147),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43148(.data_in(wire_d3_147),.data_out(wire_d3_148),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43149(.data_in(wire_d3_148),.data_out(wire_d3_149),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43150(.data_in(wire_d3_149),.data_out(wire_d3_150),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43151(.data_in(wire_d3_150),.data_out(wire_d3_151),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43152(.data_in(wire_d3_151),.data_out(wire_d3_152),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43153(.data_in(wire_d3_152),.data_out(wire_d3_153),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43154(.data_in(wire_d3_153),.data_out(wire_d3_154),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43155(.data_in(wire_d3_154),.data_out(wire_d3_155),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43156(.data_in(wire_d3_155),.data_out(wire_d3_156),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43157(.data_in(wire_d3_156),.data_out(wire_d3_157),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43158(.data_in(wire_d3_157),.data_out(wire_d3_158),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43159(.data_in(wire_d3_158),.data_out(wire_d3_159),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43160(.data_in(wire_d3_159),.data_out(wire_d3_160),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43161(.data_in(wire_d3_160),.data_out(wire_d3_161),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43162(.data_in(wire_d3_161),.data_out(wire_d3_162),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43163(.data_in(wire_d3_162),.data_out(wire_d3_163),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43164(.data_in(wire_d3_163),.data_out(wire_d3_164),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43165(.data_in(wire_d3_164),.data_out(wire_d3_165),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43166(.data_in(wire_d3_165),.data_out(wire_d3_166),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43167(.data_in(wire_d3_166),.data_out(wire_d3_167),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43168(.data_in(wire_d3_167),.data_out(wire_d3_168),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43169(.data_in(wire_d3_168),.data_out(wire_d3_169),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43170(.data_in(wire_d3_169),.data_out(wire_d3_170),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43171(.data_in(wire_d3_170),.data_out(wire_d3_171),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43172(.data_in(wire_d3_171),.data_out(wire_d3_172),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43173(.data_in(wire_d3_172),.data_out(wire_d3_173),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43174(.data_in(wire_d3_173),.data_out(wire_d3_174),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43175(.data_in(wire_d3_174),.data_out(wire_d3_175),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43176(.data_in(wire_d3_175),.data_out(wire_d3_176),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43177(.data_in(wire_d3_176),.data_out(wire_d3_177),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43178(.data_in(wire_d3_177),.data_out(wire_d3_178),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43179(.data_in(wire_d3_178),.data_out(wire_d3_179),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43180(.data_in(wire_d3_179),.data_out(wire_d3_180),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43181(.data_in(wire_d3_180),.data_out(wire_d3_181),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43182(.data_in(wire_d3_181),.data_out(wire_d3_182),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43183(.data_in(wire_d3_182),.data_out(wire_d3_183),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43184(.data_in(wire_d3_183),.data_out(wire_d3_184),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43185(.data_in(wire_d3_184),.data_out(wire_d3_185),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43186(.data_in(wire_d3_185),.data_out(wire_d3_186),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43187(.data_in(wire_d3_186),.data_out(wire_d3_187),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43188(.data_in(wire_d3_187),.data_out(wire_d3_188),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43189(.data_in(wire_d3_188),.data_out(wire_d3_189),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43190(.data_in(wire_d3_189),.data_out(wire_d3_190),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43191(.data_in(wire_d3_190),.data_out(wire_d3_191),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43192(.data_in(wire_d3_191),.data_out(wire_d3_192),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43193(.data_in(wire_d3_192),.data_out(wire_d3_193),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43194(.data_in(wire_d3_193),.data_out(wire_d3_194),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43195(.data_in(wire_d3_194),.data_out(wire_d3_195),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43196(.data_in(wire_d3_195),.data_out(wire_d3_196),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43197(.data_in(wire_d3_196),.data_out(wire_d3_197),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43198(.data_in(wire_d3_197),.data_out(wire_d3_198),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43199(.data_in(wire_d3_198),.data_out(d_out3),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance540(.data_in(d_in4),.data_out(wire_d4_0),.clk(clk),.rst(rst));            //channel 5
	encoder #(.WIDTH(WIDTH)) encoder_instance541(.data_in(wire_d4_0),.data_out(wire_d4_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance542(.data_in(wire_d4_1),.data_out(wire_d4_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance543(.data_in(wire_d4_2),.data_out(wire_d4_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance544(.data_in(wire_d4_3),.data_out(wire_d4_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545(.data_in(wire_d4_4),.data_out(wire_d4_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance546(.data_in(wire_d4_5),.data_out(wire_d4_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance547(.data_in(wire_d4_6),.data_out(wire_d4_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance548(.data_in(wire_d4_7),.data_out(wire_d4_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance549(.data_in(wire_d4_8),.data_out(wire_d4_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5410(.data_in(wire_d4_9),.data_out(wire_d4_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5411(.data_in(wire_d4_10),.data_out(wire_d4_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5412(.data_in(wire_d4_11),.data_out(wire_d4_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5413(.data_in(wire_d4_12),.data_out(wire_d4_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5414(.data_in(wire_d4_13),.data_out(wire_d4_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5415(.data_in(wire_d4_14),.data_out(wire_d4_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5416(.data_in(wire_d4_15),.data_out(wire_d4_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5417(.data_in(wire_d4_16),.data_out(wire_d4_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5418(.data_in(wire_d4_17),.data_out(wire_d4_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5419(.data_in(wire_d4_18),.data_out(wire_d4_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5420(.data_in(wire_d4_19),.data_out(wire_d4_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5421(.data_in(wire_d4_20),.data_out(wire_d4_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5422(.data_in(wire_d4_21),.data_out(wire_d4_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5423(.data_in(wire_d4_22),.data_out(wire_d4_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5424(.data_in(wire_d4_23),.data_out(wire_d4_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5425(.data_in(wire_d4_24),.data_out(wire_d4_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5426(.data_in(wire_d4_25),.data_out(wire_d4_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5427(.data_in(wire_d4_26),.data_out(wire_d4_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5428(.data_in(wire_d4_27),.data_out(wire_d4_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5429(.data_in(wire_d4_28),.data_out(wire_d4_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5430(.data_in(wire_d4_29),.data_out(wire_d4_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5431(.data_in(wire_d4_30),.data_out(wire_d4_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5432(.data_in(wire_d4_31),.data_out(wire_d4_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5433(.data_in(wire_d4_32),.data_out(wire_d4_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5434(.data_in(wire_d4_33),.data_out(wire_d4_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5435(.data_in(wire_d4_34),.data_out(wire_d4_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5436(.data_in(wire_d4_35),.data_out(wire_d4_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5437(.data_in(wire_d4_36),.data_out(wire_d4_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5438(.data_in(wire_d4_37),.data_out(wire_d4_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5439(.data_in(wire_d4_38),.data_out(wire_d4_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5440(.data_in(wire_d4_39),.data_out(wire_d4_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5441(.data_in(wire_d4_40),.data_out(wire_d4_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5442(.data_in(wire_d4_41),.data_out(wire_d4_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5443(.data_in(wire_d4_42),.data_out(wire_d4_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5444(.data_in(wire_d4_43),.data_out(wire_d4_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5445(.data_in(wire_d4_44),.data_out(wire_d4_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5446(.data_in(wire_d4_45),.data_out(wire_d4_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5447(.data_in(wire_d4_46),.data_out(wire_d4_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5448(.data_in(wire_d4_47),.data_out(wire_d4_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5449(.data_in(wire_d4_48),.data_out(wire_d4_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5450(.data_in(wire_d4_49),.data_out(wire_d4_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5451(.data_in(wire_d4_50),.data_out(wire_d4_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5452(.data_in(wire_d4_51),.data_out(wire_d4_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5453(.data_in(wire_d4_52),.data_out(wire_d4_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5454(.data_in(wire_d4_53),.data_out(wire_d4_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5455(.data_in(wire_d4_54),.data_out(wire_d4_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5456(.data_in(wire_d4_55),.data_out(wire_d4_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5457(.data_in(wire_d4_56),.data_out(wire_d4_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5458(.data_in(wire_d4_57),.data_out(wire_d4_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5459(.data_in(wire_d4_58),.data_out(wire_d4_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5460(.data_in(wire_d4_59),.data_out(wire_d4_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5461(.data_in(wire_d4_60),.data_out(wire_d4_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5462(.data_in(wire_d4_61),.data_out(wire_d4_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5463(.data_in(wire_d4_62),.data_out(wire_d4_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5464(.data_in(wire_d4_63),.data_out(wire_d4_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5465(.data_in(wire_d4_64),.data_out(wire_d4_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5466(.data_in(wire_d4_65),.data_out(wire_d4_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5467(.data_in(wire_d4_66),.data_out(wire_d4_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5468(.data_in(wire_d4_67),.data_out(wire_d4_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5469(.data_in(wire_d4_68),.data_out(wire_d4_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5470(.data_in(wire_d4_69),.data_out(wire_d4_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5471(.data_in(wire_d4_70),.data_out(wire_d4_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5472(.data_in(wire_d4_71),.data_out(wire_d4_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5473(.data_in(wire_d4_72),.data_out(wire_d4_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5474(.data_in(wire_d4_73),.data_out(wire_d4_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5475(.data_in(wire_d4_74),.data_out(wire_d4_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5476(.data_in(wire_d4_75),.data_out(wire_d4_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5477(.data_in(wire_d4_76),.data_out(wire_d4_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5478(.data_in(wire_d4_77),.data_out(wire_d4_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5479(.data_in(wire_d4_78),.data_out(wire_d4_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5480(.data_in(wire_d4_79),.data_out(wire_d4_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5481(.data_in(wire_d4_80),.data_out(wire_d4_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5482(.data_in(wire_d4_81),.data_out(wire_d4_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5483(.data_in(wire_d4_82),.data_out(wire_d4_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5484(.data_in(wire_d4_83),.data_out(wire_d4_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5485(.data_in(wire_d4_84),.data_out(wire_d4_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5486(.data_in(wire_d4_85),.data_out(wire_d4_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5487(.data_in(wire_d4_86),.data_out(wire_d4_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5488(.data_in(wire_d4_87),.data_out(wire_d4_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5489(.data_in(wire_d4_88),.data_out(wire_d4_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5490(.data_in(wire_d4_89),.data_out(wire_d4_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5491(.data_in(wire_d4_90),.data_out(wire_d4_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5492(.data_in(wire_d4_91),.data_out(wire_d4_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5493(.data_in(wire_d4_92),.data_out(wire_d4_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5494(.data_in(wire_d4_93),.data_out(wire_d4_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5495(.data_in(wire_d4_94),.data_out(wire_d4_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5496(.data_in(wire_d4_95),.data_out(wire_d4_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5497(.data_in(wire_d4_96),.data_out(wire_d4_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5498(.data_in(wire_d4_97),.data_out(wire_d4_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5499(.data_in(wire_d4_98),.data_out(wire_d4_99),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54100(.data_in(wire_d4_99),.data_out(wire_d4_100),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54101(.data_in(wire_d4_100),.data_out(wire_d4_101),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54102(.data_in(wire_d4_101),.data_out(wire_d4_102),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54103(.data_in(wire_d4_102),.data_out(wire_d4_103),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54104(.data_in(wire_d4_103),.data_out(wire_d4_104),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54105(.data_in(wire_d4_104),.data_out(wire_d4_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54106(.data_in(wire_d4_105),.data_out(wire_d4_106),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54107(.data_in(wire_d4_106),.data_out(wire_d4_107),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54108(.data_in(wire_d4_107),.data_out(wire_d4_108),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54109(.data_in(wire_d4_108),.data_out(wire_d4_109),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54110(.data_in(wire_d4_109),.data_out(wire_d4_110),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54111(.data_in(wire_d4_110),.data_out(wire_d4_111),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54112(.data_in(wire_d4_111),.data_out(wire_d4_112),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54113(.data_in(wire_d4_112),.data_out(wire_d4_113),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54114(.data_in(wire_d4_113),.data_out(wire_d4_114),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54115(.data_in(wire_d4_114),.data_out(wire_d4_115),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54116(.data_in(wire_d4_115),.data_out(wire_d4_116),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54117(.data_in(wire_d4_116),.data_out(wire_d4_117),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54118(.data_in(wire_d4_117),.data_out(wire_d4_118),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54119(.data_in(wire_d4_118),.data_out(wire_d4_119),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54120(.data_in(wire_d4_119),.data_out(wire_d4_120),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54121(.data_in(wire_d4_120),.data_out(wire_d4_121),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54122(.data_in(wire_d4_121),.data_out(wire_d4_122),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54123(.data_in(wire_d4_122),.data_out(wire_d4_123),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54124(.data_in(wire_d4_123),.data_out(wire_d4_124),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54125(.data_in(wire_d4_124),.data_out(wire_d4_125),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54126(.data_in(wire_d4_125),.data_out(wire_d4_126),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54127(.data_in(wire_d4_126),.data_out(wire_d4_127),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54128(.data_in(wire_d4_127),.data_out(wire_d4_128),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54129(.data_in(wire_d4_128),.data_out(wire_d4_129),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54130(.data_in(wire_d4_129),.data_out(wire_d4_130),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54131(.data_in(wire_d4_130),.data_out(wire_d4_131),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54132(.data_in(wire_d4_131),.data_out(wire_d4_132),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54133(.data_in(wire_d4_132),.data_out(wire_d4_133),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54134(.data_in(wire_d4_133),.data_out(wire_d4_134),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54135(.data_in(wire_d4_134),.data_out(wire_d4_135),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54136(.data_in(wire_d4_135),.data_out(wire_d4_136),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54137(.data_in(wire_d4_136),.data_out(wire_d4_137),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54138(.data_in(wire_d4_137),.data_out(wire_d4_138),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54139(.data_in(wire_d4_138),.data_out(wire_d4_139),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54140(.data_in(wire_d4_139),.data_out(wire_d4_140),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54141(.data_in(wire_d4_140),.data_out(wire_d4_141),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54142(.data_in(wire_d4_141),.data_out(wire_d4_142),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54143(.data_in(wire_d4_142),.data_out(wire_d4_143),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54144(.data_in(wire_d4_143),.data_out(wire_d4_144),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54145(.data_in(wire_d4_144),.data_out(wire_d4_145),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54146(.data_in(wire_d4_145),.data_out(wire_d4_146),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54147(.data_in(wire_d4_146),.data_out(wire_d4_147),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54148(.data_in(wire_d4_147),.data_out(wire_d4_148),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54149(.data_in(wire_d4_148),.data_out(wire_d4_149),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54150(.data_in(wire_d4_149),.data_out(wire_d4_150),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54151(.data_in(wire_d4_150),.data_out(wire_d4_151),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54152(.data_in(wire_d4_151),.data_out(wire_d4_152),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54153(.data_in(wire_d4_152),.data_out(wire_d4_153),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54154(.data_in(wire_d4_153),.data_out(wire_d4_154),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54155(.data_in(wire_d4_154),.data_out(wire_d4_155),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54156(.data_in(wire_d4_155),.data_out(wire_d4_156),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54157(.data_in(wire_d4_156),.data_out(wire_d4_157),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54158(.data_in(wire_d4_157),.data_out(wire_d4_158),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54159(.data_in(wire_d4_158),.data_out(wire_d4_159),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54160(.data_in(wire_d4_159),.data_out(wire_d4_160),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54161(.data_in(wire_d4_160),.data_out(wire_d4_161),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54162(.data_in(wire_d4_161),.data_out(wire_d4_162),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54163(.data_in(wire_d4_162),.data_out(wire_d4_163),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54164(.data_in(wire_d4_163),.data_out(wire_d4_164),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54165(.data_in(wire_d4_164),.data_out(wire_d4_165),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54166(.data_in(wire_d4_165),.data_out(wire_d4_166),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54167(.data_in(wire_d4_166),.data_out(wire_d4_167),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54168(.data_in(wire_d4_167),.data_out(wire_d4_168),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54169(.data_in(wire_d4_168),.data_out(wire_d4_169),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54170(.data_in(wire_d4_169),.data_out(wire_d4_170),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54171(.data_in(wire_d4_170),.data_out(wire_d4_171),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54172(.data_in(wire_d4_171),.data_out(wire_d4_172),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54173(.data_in(wire_d4_172),.data_out(wire_d4_173),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54174(.data_in(wire_d4_173),.data_out(wire_d4_174),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54175(.data_in(wire_d4_174),.data_out(wire_d4_175),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54176(.data_in(wire_d4_175),.data_out(wire_d4_176),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54177(.data_in(wire_d4_176),.data_out(wire_d4_177),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54178(.data_in(wire_d4_177),.data_out(wire_d4_178),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54179(.data_in(wire_d4_178),.data_out(wire_d4_179),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54180(.data_in(wire_d4_179),.data_out(wire_d4_180),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54181(.data_in(wire_d4_180),.data_out(wire_d4_181),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54182(.data_in(wire_d4_181),.data_out(wire_d4_182),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54183(.data_in(wire_d4_182),.data_out(wire_d4_183),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54184(.data_in(wire_d4_183),.data_out(wire_d4_184),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54185(.data_in(wire_d4_184),.data_out(wire_d4_185),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54186(.data_in(wire_d4_185),.data_out(wire_d4_186),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54187(.data_in(wire_d4_186),.data_out(wire_d4_187),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54188(.data_in(wire_d4_187),.data_out(wire_d4_188),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54189(.data_in(wire_d4_188),.data_out(wire_d4_189),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54190(.data_in(wire_d4_189),.data_out(wire_d4_190),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54191(.data_in(wire_d4_190),.data_out(wire_d4_191),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54192(.data_in(wire_d4_191),.data_out(wire_d4_192),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54193(.data_in(wire_d4_192),.data_out(wire_d4_193),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54194(.data_in(wire_d4_193),.data_out(wire_d4_194),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54195(.data_in(wire_d4_194),.data_out(wire_d4_195),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54196(.data_in(wire_d4_195),.data_out(wire_d4_196),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54197(.data_in(wire_d4_196),.data_out(wire_d4_197),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54198(.data_in(wire_d4_197),.data_out(wire_d4_198),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54199(.data_in(wire_d4_198),.data_out(d_out4),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance650(.data_in(d_in5),.data_out(wire_d5_0),.clk(clk),.rst(rst));            //channel 6
	encoder #(.WIDTH(WIDTH)) encoder_instance651(.data_in(wire_d5_0),.data_out(wire_d5_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance652(.data_in(wire_d5_1),.data_out(wire_d5_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance653(.data_in(wire_d5_2),.data_out(wire_d5_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance654(.data_in(wire_d5_3),.data_out(wire_d5_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance655(.data_in(wire_d5_4),.data_out(wire_d5_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656(.data_in(wire_d5_5),.data_out(wire_d5_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance657(.data_in(wire_d5_6),.data_out(wire_d5_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance658(.data_in(wire_d5_7),.data_out(wire_d5_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance659(.data_in(wire_d5_8),.data_out(wire_d5_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6510(.data_in(wire_d5_9),.data_out(wire_d5_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6511(.data_in(wire_d5_10),.data_out(wire_d5_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6512(.data_in(wire_d5_11),.data_out(wire_d5_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6513(.data_in(wire_d5_12),.data_out(wire_d5_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6514(.data_in(wire_d5_13),.data_out(wire_d5_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6515(.data_in(wire_d5_14),.data_out(wire_d5_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6516(.data_in(wire_d5_15),.data_out(wire_d5_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6517(.data_in(wire_d5_16),.data_out(wire_d5_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6518(.data_in(wire_d5_17),.data_out(wire_d5_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6519(.data_in(wire_d5_18),.data_out(wire_d5_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6520(.data_in(wire_d5_19),.data_out(wire_d5_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6521(.data_in(wire_d5_20),.data_out(wire_d5_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6522(.data_in(wire_d5_21),.data_out(wire_d5_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6523(.data_in(wire_d5_22),.data_out(wire_d5_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6524(.data_in(wire_d5_23),.data_out(wire_d5_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6525(.data_in(wire_d5_24),.data_out(wire_d5_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6526(.data_in(wire_d5_25),.data_out(wire_d5_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6527(.data_in(wire_d5_26),.data_out(wire_d5_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6528(.data_in(wire_d5_27),.data_out(wire_d5_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6529(.data_in(wire_d5_28),.data_out(wire_d5_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6530(.data_in(wire_d5_29),.data_out(wire_d5_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6531(.data_in(wire_d5_30),.data_out(wire_d5_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6532(.data_in(wire_d5_31),.data_out(wire_d5_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6533(.data_in(wire_d5_32),.data_out(wire_d5_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6534(.data_in(wire_d5_33),.data_out(wire_d5_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6535(.data_in(wire_d5_34),.data_out(wire_d5_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6536(.data_in(wire_d5_35),.data_out(wire_d5_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6537(.data_in(wire_d5_36),.data_out(wire_d5_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6538(.data_in(wire_d5_37),.data_out(wire_d5_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6539(.data_in(wire_d5_38),.data_out(wire_d5_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6540(.data_in(wire_d5_39),.data_out(wire_d5_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6541(.data_in(wire_d5_40),.data_out(wire_d5_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6542(.data_in(wire_d5_41),.data_out(wire_d5_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6543(.data_in(wire_d5_42),.data_out(wire_d5_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6544(.data_in(wire_d5_43),.data_out(wire_d5_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6545(.data_in(wire_d5_44),.data_out(wire_d5_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6546(.data_in(wire_d5_45),.data_out(wire_d5_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6547(.data_in(wire_d5_46),.data_out(wire_d5_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6548(.data_in(wire_d5_47),.data_out(wire_d5_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6549(.data_in(wire_d5_48),.data_out(wire_d5_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6550(.data_in(wire_d5_49),.data_out(wire_d5_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6551(.data_in(wire_d5_50),.data_out(wire_d5_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6552(.data_in(wire_d5_51),.data_out(wire_d5_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6553(.data_in(wire_d5_52),.data_out(wire_d5_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6554(.data_in(wire_d5_53),.data_out(wire_d5_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6555(.data_in(wire_d5_54),.data_out(wire_d5_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6556(.data_in(wire_d5_55),.data_out(wire_d5_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6557(.data_in(wire_d5_56),.data_out(wire_d5_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6558(.data_in(wire_d5_57),.data_out(wire_d5_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6559(.data_in(wire_d5_58),.data_out(wire_d5_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6560(.data_in(wire_d5_59),.data_out(wire_d5_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6561(.data_in(wire_d5_60),.data_out(wire_d5_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6562(.data_in(wire_d5_61),.data_out(wire_d5_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6563(.data_in(wire_d5_62),.data_out(wire_d5_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6564(.data_in(wire_d5_63),.data_out(wire_d5_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6565(.data_in(wire_d5_64),.data_out(wire_d5_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6566(.data_in(wire_d5_65),.data_out(wire_d5_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6567(.data_in(wire_d5_66),.data_out(wire_d5_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6568(.data_in(wire_d5_67),.data_out(wire_d5_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6569(.data_in(wire_d5_68),.data_out(wire_d5_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6570(.data_in(wire_d5_69),.data_out(wire_d5_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6571(.data_in(wire_d5_70),.data_out(wire_d5_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6572(.data_in(wire_d5_71),.data_out(wire_d5_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6573(.data_in(wire_d5_72),.data_out(wire_d5_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6574(.data_in(wire_d5_73),.data_out(wire_d5_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6575(.data_in(wire_d5_74),.data_out(wire_d5_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6576(.data_in(wire_d5_75),.data_out(wire_d5_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6577(.data_in(wire_d5_76),.data_out(wire_d5_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6578(.data_in(wire_d5_77),.data_out(wire_d5_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6579(.data_in(wire_d5_78),.data_out(wire_d5_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6580(.data_in(wire_d5_79),.data_out(wire_d5_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6581(.data_in(wire_d5_80),.data_out(wire_d5_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6582(.data_in(wire_d5_81),.data_out(wire_d5_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6583(.data_in(wire_d5_82),.data_out(wire_d5_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6584(.data_in(wire_d5_83),.data_out(wire_d5_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6585(.data_in(wire_d5_84),.data_out(wire_d5_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6586(.data_in(wire_d5_85),.data_out(wire_d5_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6587(.data_in(wire_d5_86),.data_out(wire_d5_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6588(.data_in(wire_d5_87),.data_out(wire_d5_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6589(.data_in(wire_d5_88),.data_out(wire_d5_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6590(.data_in(wire_d5_89),.data_out(wire_d5_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6591(.data_in(wire_d5_90),.data_out(wire_d5_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6592(.data_in(wire_d5_91),.data_out(wire_d5_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6593(.data_in(wire_d5_92),.data_out(wire_d5_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6594(.data_in(wire_d5_93),.data_out(wire_d5_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6595(.data_in(wire_d5_94),.data_out(wire_d5_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6596(.data_in(wire_d5_95),.data_out(wire_d5_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6597(.data_in(wire_d5_96),.data_out(wire_d5_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6598(.data_in(wire_d5_97),.data_out(wire_d5_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6599(.data_in(wire_d5_98),.data_out(wire_d5_99),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65100(.data_in(wire_d5_99),.data_out(wire_d5_100),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65101(.data_in(wire_d5_100),.data_out(wire_d5_101),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65102(.data_in(wire_d5_101),.data_out(wire_d5_102),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65103(.data_in(wire_d5_102),.data_out(wire_d5_103),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65104(.data_in(wire_d5_103),.data_out(wire_d5_104),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65105(.data_in(wire_d5_104),.data_out(wire_d5_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65106(.data_in(wire_d5_105),.data_out(wire_d5_106),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65107(.data_in(wire_d5_106),.data_out(wire_d5_107),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65108(.data_in(wire_d5_107),.data_out(wire_d5_108),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65109(.data_in(wire_d5_108),.data_out(wire_d5_109),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65110(.data_in(wire_d5_109),.data_out(wire_d5_110),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65111(.data_in(wire_d5_110),.data_out(wire_d5_111),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65112(.data_in(wire_d5_111),.data_out(wire_d5_112),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65113(.data_in(wire_d5_112),.data_out(wire_d5_113),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65114(.data_in(wire_d5_113),.data_out(wire_d5_114),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65115(.data_in(wire_d5_114),.data_out(wire_d5_115),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65116(.data_in(wire_d5_115),.data_out(wire_d5_116),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65117(.data_in(wire_d5_116),.data_out(wire_d5_117),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65118(.data_in(wire_d5_117),.data_out(wire_d5_118),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65119(.data_in(wire_d5_118),.data_out(wire_d5_119),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65120(.data_in(wire_d5_119),.data_out(wire_d5_120),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65121(.data_in(wire_d5_120),.data_out(wire_d5_121),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65122(.data_in(wire_d5_121),.data_out(wire_d5_122),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65123(.data_in(wire_d5_122),.data_out(wire_d5_123),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65124(.data_in(wire_d5_123),.data_out(wire_d5_124),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65125(.data_in(wire_d5_124),.data_out(wire_d5_125),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65126(.data_in(wire_d5_125),.data_out(wire_d5_126),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65127(.data_in(wire_d5_126),.data_out(wire_d5_127),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65128(.data_in(wire_d5_127),.data_out(wire_d5_128),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65129(.data_in(wire_d5_128),.data_out(wire_d5_129),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65130(.data_in(wire_d5_129),.data_out(wire_d5_130),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65131(.data_in(wire_d5_130),.data_out(wire_d5_131),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65132(.data_in(wire_d5_131),.data_out(wire_d5_132),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65133(.data_in(wire_d5_132),.data_out(wire_d5_133),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65134(.data_in(wire_d5_133),.data_out(wire_d5_134),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65135(.data_in(wire_d5_134),.data_out(wire_d5_135),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65136(.data_in(wire_d5_135),.data_out(wire_d5_136),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65137(.data_in(wire_d5_136),.data_out(wire_d5_137),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65138(.data_in(wire_d5_137),.data_out(wire_d5_138),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65139(.data_in(wire_d5_138),.data_out(wire_d5_139),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65140(.data_in(wire_d5_139),.data_out(wire_d5_140),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65141(.data_in(wire_d5_140),.data_out(wire_d5_141),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65142(.data_in(wire_d5_141),.data_out(wire_d5_142),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65143(.data_in(wire_d5_142),.data_out(wire_d5_143),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65144(.data_in(wire_d5_143),.data_out(wire_d5_144),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65145(.data_in(wire_d5_144),.data_out(wire_d5_145),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65146(.data_in(wire_d5_145),.data_out(wire_d5_146),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65147(.data_in(wire_d5_146),.data_out(wire_d5_147),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65148(.data_in(wire_d5_147),.data_out(wire_d5_148),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65149(.data_in(wire_d5_148),.data_out(wire_d5_149),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65150(.data_in(wire_d5_149),.data_out(wire_d5_150),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65151(.data_in(wire_d5_150),.data_out(wire_d5_151),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65152(.data_in(wire_d5_151),.data_out(wire_d5_152),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65153(.data_in(wire_d5_152),.data_out(wire_d5_153),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65154(.data_in(wire_d5_153),.data_out(wire_d5_154),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65155(.data_in(wire_d5_154),.data_out(wire_d5_155),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65156(.data_in(wire_d5_155),.data_out(wire_d5_156),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65157(.data_in(wire_d5_156),.data_out(wire_d5_157),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65158(.data_in(wire_d5_157),.data_out(wire_d5_158),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65159(.data_in(wire_d5_158),.data_out(wire_d5_159),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65160(.data_in(wire_d5_159),.data_out(wire_d5_160),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65161(.data_in(wire_d5_160),.data_out(wire_d5_161),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65162(.data_in(wire_d5_161),.data_out(wire_d5_162),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65163(.data_in(wire_d5_162),.data_out(wire_d5_163),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65164(.data_in(wire_d5_163),.data_out(wire_d5_164),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65165(.data_in(wire_d5_164),.data_out(wire_d5_165),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65166(.data_in(wire_d5_165),.data_out(wire_d5_166),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65167(.data_in(wire_d5_166),.data_out(wire_d5_167),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65168(.data_in(wire_d5_167),.data_out(wire_d5_168),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65169(.data_in(wire_d5_168),.data_out(wire_d5_169),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65170(.data_in(wire_d5_169),.data_out(wire_d5_170),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65171(.data_in(wire_d5_170),.data_out(wire_d5_171),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65172(.data_in(wire_d5_171),.data_out(wire_d5_172),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65173(.data_in(wire_d5_172),.data_out(wire_d5_173),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65174(.data_in(wire_d5_173),.data_out(wire_d5_174),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65175(.data_in(wire_d5_174),.data_out(wire_d5_175),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65176(.data_in(wire_d5_175),.data_out(wire_d5_176),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65177(.data_in(wire_d5_176),.data_out(wire_d5_177),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65178(.data_in(wire_d5_177),.data_out(wire_d5_178),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65179(.data_in(wire_d5_178),.data_out(wire_d5_179),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65180(.data_in(wire_d5_179),.data_out(wire_d5_180),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65181(.data_in(wire_d5_180),.data_out(wire_d5_181),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65182(.data_in(wire_d5_181),.data_out(wire_d5_182),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65183(.data_in(wire_d5_182),.data_out(wire_d5_183),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65184(.data_in(wire_d5_183),.data_out(wire_d5_184),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65185(.data_in(wire_d5_184),.data_out(wire_d5_185),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65186(.data_in(wire_d5_185),.data_out(wire_d5_186),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65187(.data_in(wire_d5_186),.data_out(wire_d5_187),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65188(.data_in(wire_d5_187),.data_out(wire_d5_188),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65189(.data_in(wire_d5_188),.data_out(wire_d5_189),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65190(.data_in(wire_d5_189),.data_out(wire_d5_190),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65191(.data_in(wire_d5_190),.data_out(wire_d5_191),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65192(.data_in(wire_d5_191),.data_out(wire_d5_192),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65193(.data_in(wire_d5_192),.data_out(wire_d5_193),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65194(.data_in(wire_d5_193),.data_out(wire_d5_194),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65195(.data_in(wire_d5_194),.data_out(wire_d5_195),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65196(.data_in(wire_d5_195),.data_out(wire_d5_196),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65197(.data_in(wire_d5_196),.data_out(wire_d5_197),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65198(.data_in(wire_d5_197),.data_out(wire_d5_198),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65199(.data_in(wire_d5_198),.data_out(d_out5),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance760(.data_in(d_in6),.data_out(wire_d6_0),.clk(clk),.rst(rst));            //channel 7
	encoder #(.WIDTH(WIDTH)) encoder_instance761(.data_in(wire_d6_0),.data_out(wire_d6_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance762(.data_in(wire_d6_1),.data_out(wire_d6_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance763(.data_in(wire_d6_2),.data_out(wire_d6_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance764(.data_in(wire_d6_3),.data_out(wire_d6_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance765(.data_in(wire_d6_4),.data_out(wire_d6_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance766(.data_in(wire_d6_5),.data_out(wire_d6_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767(.data_in(wire_d6_6),.data_out(wire_d6_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance768(.data_in(wire_d6_7),.data_out(wire_d6_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance769(.data_in(wire_d6_8),.data_out(wire_d6_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7610(.data_in(wire_d6_9),.data_out(wire_d6_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7611(.data_in(wire_d6_10),.data_out(wire_d6_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7612(.data_in(wire_d6_11),.data_out(wire_d6_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7613(.data_in(wire_d6_12),.data_out(wire_d6_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7614(.data_in(wire_d6_13),.data_out(wire_d6_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7615(.data_in(wire_d6_14),.data_out(wire_d6_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7616(.data_in(wire_d6_15),.data_out(wire_d6_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7617(.data_in(wire_d6_16),.data_out(wire_d6_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7618(.data_in(wire_d6_17),.data_out(wire_d6_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7619(.data_in(wire_d6_18),.data_out(wire_d6_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7620(.data_in(wire_d6_19),.data_out(wire_d6_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7621(.data_in(wire_d6_20),.data_out(wire_d6_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7622(.data_in(wire_d6_21),.data_out(wire_d6_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7623(.data_in(wire_d6_22),.data_out(wire_d6_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7624(.data_in(wire_d6_23),.data_out(wire_d6_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7625(.data_in(wire_d6_24),.data_out(wire_d6_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7626(.data_in(wire_d6_25),.data_out(wire_d6_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7627(.data_in(wire_d6_26),.data_out(wire_d6_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7628(.data_in(wire_d6_27),.data_out(wire_d6_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7629(.data_in(wire_d6_28),.data_out(wire_d6_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7630(.data_in(wire_d6_29),.data_out(wire_d6_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7631(.data_in(wire_d6_30),.data_out(wire_d6_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7632(.data_in(wire_d6_31),.data_out(wire_d6_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7633(.data_in(wire_d6_32),.data_out(wire_d6_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7634(.data_in(wire_d6_33),.data_out(wire_d6_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7635(.data_in(wire_d6_34),.data_out(wire_d6_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7636(.data_in(wire_d6_35),.data_out(wire_d6_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7637(.data_in(wire_d6_36),.data_out(wire_d6_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7638(.data_in(wire_d6_37),.data_out(wire_d6_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7639(.data_in(wire_d6_38),.data_out(wire_d6_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7640(.data_in(wire_d6_39),.data_out(wire_d6_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7641(.data_in(wire_d6_40),.data_out(wire_d6_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7642(.data_in(wire_d6_41),.data_out(wire_d6_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7643(.data_in(wire_d6_42),.data_out(wire_d6_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7644(.data_in(wire_d6_43),.data_out(wire_d6_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7645(.data_in(wire_d6_44),.data_out(wire_d6_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7646(.data_in(wire_d6_45),.data_out(wire_d6_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7647(.data_in(wire_d6_46),.data_out(wire_d6_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7648(.data_in(wire_d6_47),.data_out(wire_d6_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7649(.data_in(wire_d6_48),.data_out(wire_d6_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7650(.data_in(wire_d6_49),.data_out(wire_d6_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7651(.data_in(wire_d6_50),.data_out(wire_d6_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7652(.data_in(wire_d6_51),.data_out(wire_d6_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7653(.data_in(wire_d6_52),.data_out(wire_d6_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7654(.data_in(wire_d6_53),.data_out(wire_d6_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7655(.data_in(wire_d6_54),.data_out(wire_d6_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7656(.data_in(wire_d6_55),.data_out(wire_d6_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7657(.data_in(wire_d6_56),.data_out(wire_d6_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7658(.data_in(wire_d6_57),.data_out(wire_d6_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7659(.data_in(wire_d6_58),.data_out(wire_d6_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7660(.data_in(wire_d6_59),.data_out(wire_d6_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7661(.data_in(wire_d6_60),.data_out(wire_d6_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7662(.data_in(wire_d6_61),.data_out(wire_d6_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7663(.data_in(wire_d6_62),.data_out(wire_d6_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7664(.data_in(wire_d6_63),.data_out(wire_d6_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7665(.data_in(wire_d6_64),.data_out(wire_d6_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7666(.data_in(wire_d6_65),.data_out(wire_d6_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7667(.data_in(wire_d6_66),.data_out(wire_d6_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7668(.data_in(wire_d6_67),.data_out(wire_d6_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7669(.data_in(wire_d6_68),.data_out(wire_d6_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7670(.data_in(wire_d6_69),.data_out(wire_d6_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7671(.data_in(wire_d6_70),.data_out(wire_d6_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7672(.data_in(wire_d6_71),.data_out(wire_d6_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7673(.data_in(wire_d6_72),.data_out(wire_d6_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7674(.data_in(wire_d6_73),.data_out(wire_d6_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7675(.data_in(wire_d6_74),.data_out(wire_d6_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7676(.data_in(wire_d6_75),.data_out(wire_d6_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7677(.data_in(wire_d6_76),.data_out(wire_d6_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7678(.data_in(wire_d6_77),.data_out(wire_d6_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7679(.data_in(wire_d6_78),.data_out(wire_d6_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7680(.data_in(wire_d6_79),.data_out(wire_d6_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7681(.data_in(wire_d6_80),.data_out(wire_d6_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7682(.data_in(wire_d6_81),.data_out(wire_d6_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7683(.data_in(wire_d6_82),.data_out(wire_d6_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7684(.data_in(wire_d6_83),.data_out(wire_d6_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7685(.data_in(wire_d6_84),.data_out(wire_d6_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7686(.data_in(wire_d6_85),.data_out(wire_d6_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7687(.data_in(wire_d6_86),.data_out(wire_d6_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7688(.data_in(wire_d6_87),.data_out(wire_d6_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7689(.data_in(wire_d6_88),.data_out(wire_d6_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7690(.data_in(wire_d6_89),.data_out(wire_d6_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7691(.data_in(wire_d6_90),.data_out(wire_d6_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7692(.data_in(wire_d6_91),.data_out(wire_d6_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7693(.data_in(wire_d6_92),.data_out(wire_d6_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7694(.data_in(wire_d6_93),.data_out(wire_d6_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7695(.data_in(wire_d6_94),.data_out(wire_d6_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7696(.data_in(wire_d6_95),.data_out(wire_d6_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7697(.data_in(wire_d6_96),.data_out(wire_d6_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7698(.data_in(wire_d6_97),.data_out(wire_d6_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7699(.data_in(wire_d6_98),.data_out(wire_d6_99),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76100(.data_in(wire_d6_99),.data_out(wire_d6_100),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76101(.data_in(wire_d6_100),.data_out(wire_d6_101),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76102(.data_in(wire_d6_101),.data_out(wire_d6_102),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76103(.data_in(wire_d6_102),.data_out(wire_d6_103),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76104(.data_in(wire_d6_103),.data_out(wire_d6_104),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76105(.data_in(wire_d6_104),.data_out(wire_d6_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76106(.data_in(wire_d6_105),.data_out(wire_d6_106),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76107(.data_in(wire_d6_106),.data_out(wire_d6_107),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76108(.data_in(wire_d6_107),.data_out(wire_d6_108),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76109(.data_in(wire_d6_108),.data_out(wire_d6_109),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76110(.data_in(wire_d6_109),.data_out(wire_d6_110),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76111(.data_in(wire_d6_110),.data_out(wire_d6_111),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76112(.data_in(wire_d6_111),.data_out(wire_d6_112),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76113(.data_in(wire_d6_112),.data_out(wire_d6_113),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76114(.data_in(wire_d6_113),.data_out(wire_d6_114),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76115(.data_in(wire_d6_114),.data_out(wire_d6_115),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76116(.data_in(wire_d6_115),.data_out(wire_d6_116),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76117(.data_in(wire_d6_116),.data_out(wire_d6_117),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76118(.data_in(wire_d6_117),.data_out(wire_d6_118),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76119(.data_in(wire_d6_118),.data_out(wire_d6_119),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76120(.data_in(wire_d6_119),.data_out(wire_d6_120),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76121(.data_in(wire_d6_120),.data_out(wire_d6_121),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76122(.data_in(wire_d6_121),.data_out(wire_d6_122),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76123(.data_in(wire_d6_122),.data_out(wire_d6_123),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76124(.data_in(wire_d6_123),.data_out(wire_d6_124),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76125(.data_in(wire_d6_124),.data_out(wire_d6_125),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76126(.data_in(wire_d6_125),.data_out(wire_d6_126),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76127(.data_in(wire_d6_126),.data_out(wire_d6_127),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76128(.data_in(wire_d6_127),.data_out(wire_d6_128),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76129(.data_in(wire_d6_128),.data_out(wire_d6_129),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76130(.data_in(wire_d6_129),.data_out(wire_d6_130),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76131(.data_in(wire_d6_130),.data_out(wire_d6_131),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76132(.data_in(wire_d6_131),.data_out(wire_d6_132),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76133(.data_in(wire_d6_132),.data_out(wire_d6_133),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76134(.data_in(wire_d6_133),.data_out(wire_d6_134),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76135(.data_in(wire_d6_134),.data_out(wire_d6_135),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76136(.data_in(wire_d6_135),.data_out(wire_d6_136),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76137(.data_in(wire_d6_136),.data_out(wire_d6_137),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76138(.data_in(wire_d6_137),.data_out(wire_d6_138),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76139(.data_in(wire_d6_138),.data_out(wire_d6_139),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76140(.data_in(wire_d6_139),.data_out(wire_d6_140),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76141(.data_in(wire_d6_140),.data_out(wire_d6_141),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76142(.data_in(wire_d6_141),.data_out(wire_d6_142),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76143(.data_in(wire_d6_142),.data_out(wire_d6_143),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76144(.data_in(wire_d6_143),.data_out(wire_d6_144),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76145(.data_in(wire_d6_144),.data_out(wire_d6_145),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76146(.data_in(wire_d6_145),.data_out(wire_d6_146),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76147(.data_in(wire_d6_146),.data_out(wire_d6_147),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76148(.data_in(wire_d6_147),.data_out(wire_d6_148),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76149(.data_in(wire_d6_148),.data_out(wire_d6_149),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76150(.data_in(wire_d6_149),.data_out(wire_d6_150),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76151(.data_in(wire_d6_150),.data_out(wire_d6_151),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76152(.data_in(wire_d6_151),.data_out(wire_d6_152),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76153(.data_in(wire_d6_152),.data_out(wire_d6_153),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76154(.data_in(wire_d6_153),.data_out(wire_d6_154),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76155(.data_in(wire_d6_154),.data_out(wire_d6_155),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76156(.data_in(wire_d6_155),.data_out(wire_d6_156),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76157(.data_in(wire_d6_156),.data_out(wire_d6_157),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76158(.data_in(wire_d6_157),.data_out(wire_d6_158),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76159(.data_in(wire_d6_158),.data_out(wire_d6_159),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76160(.data_in(wire_d6_159),.data_out(wire_d6_160),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76161(.data_in(wire_d6_160),.data_out(wire_d6_161),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76162(.data_in(wire_d6_161),.data_out(wire_d6_162),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76163(.data_in(wire_d6_162),.data_out(wire_d6_163),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76164(.data_in(wire_d6_163),.data_out(wire_d6_164),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76165(.data_in(wire_d6_164),.data_out(wire_d6_165),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76166(.data_in(wire_d6_165),.data_out(wire_d6_166),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76167(.data_in(wire_d6_166),.data_out(wire_d6_167),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76168(.data_in(wire_d6_167),.data_out(wire_d6_168),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76169(.data_in(wire_d6_168),.data_out(wire_d6_169),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76170(.data_in(wire_d6_169),.data_out(wire_d6_170),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76171(.data_in(wire_d6_170),.data_out(wire_d6_171),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76172(.data_in(wire_d6_171),.data_out(wire_d6_172),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76173(.data_in(wire_d6_172),.data_out(wire_d6_173),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76174(.data_in(wire_d6_173),.data_out(wire_d6_174),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76175(.data_in(wire_d6_174),.data_out(wire_d6_175),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76176(.data_in(wire_d6_175),.data_out(wire_d6_176),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76177(.data_in(wire_d6_176),.data_out(wire_d6_177),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76178(.data_in(wire_d6_177),.data_out(wire_d6_178),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76179(.data_in(wire_d6_178),.data_out(wire_d6_179),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76180(.data_in(wire_d6_179),.data_out(wire_d6_180),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76181(.data_in(wire_d6_180),.data_out(wire_d6_181),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76182(.data_in(wire_d6_181),.data_out(wire_d6_182),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76183(.data_in(wire_d6_182),.data_out(wire_d6_183),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76184(.data_in(wire_d6_183),.data_out(wire_d6_184),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76185(.data_in(wire_d6_184),.data_out(wire_d6_185),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76186(.data_in(wire_d6_185),.data_out(wire_d6_186),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76187(.data_in(wire_d6_186),.data_out(wire_d6_187),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76188(.data_in(wire_d6_187),.data_out(wire_d6_188),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76189(.data_in(wire_d6_188),.data_out(wire_d6_189),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76190(.data_in(wire_d6_189),.data_out(wire_d6_190),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76191(.data_in(wire_d6_190),.data_out(wire_d6_191),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76192(.data_in(wire_d6_191),.data_out(wire_d6_192),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76193(.data_in(wire_d6_192),.data_out(wire_d6_193),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76194(.data_in(wire_d6_193),.data_out(wire_d6_194),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76195(.data_in(wire_d6_194),.data_out(wire_d6_195),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76196(.data_in(wire_d6_195),.data_out(wire_d6_196),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76197(.data_in(wire_d6_196),.data_out(wire_d6_197),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76198(.data_in(wire_d6_197),.data_out(wire_d6_198),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76199(.data_in(wire_d6_198),.data_out(d_out6),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance870(.data_in(d_in7),.data_out(wire_d7_0),.clk(clk),.rst(rst));            //channel 8
	encoder #(.WIDTH(WIDTH)) encoder_instance871(.data_in(wire_d7_0),.data_out(wire_d7_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance872(.data_in(wire_d7_1),.data_out(wire_d7_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance873(.data_in(wire_d7_2),.data_out(wire_d7_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance874(.data_in(wire_d7_3),.data_out(wire_d7_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance875(.data_in(wire_d7_4),.data_out(wire_d7_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance876(.data_in(wire_d7_5),.data_out(wire_d7_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance877(.data_in(wire_d7_6),.data_out(wire_d7_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878(.data_in(wire_d7_7),.data_out(wire_d7_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance879(.data_in(wire_d7_8),.data_out(wire_d7_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8710(.data_in(wire_d7_9),.data_out(wire_d7_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8711(.data_in(wire_d7_10),.data_out(wire_d7_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8712(.data_in(wire_d7_11),.data_out(wire_d7_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8713(.data_in(wire_d7_12),.data_out(wire_d7_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8714(.data_in(wire_d7_13),.data_out(wire_d7_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8715(.data_in(wire_d7_14),.data_out(wire_d7_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8716(.data_in(wire_d7_15),.data_out(wire_d7_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8717(.data_in(wire_d7_16),.data_out(wire_d7_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8718(.data_in(wire_d7_17),.data_out(wire_d7_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8719(.data_in(wire_d7_18),.data_out(wire_d7_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8720(.data_in(wire_d7_19),.data_out(wire_d7_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8721(.data_in(wire_d7_20),.data_out(wire_d7_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8722(.data_in(wire_d7_21),.data_out(wire_d7_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8723(.data_in(wire_d7_22),.data_out(wire_d7_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8724(.data_in(wire_d7_23),.data_out(wire_d7_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8725(.data_in(wire_d7_24),.data_out(wire_d7_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8726(.data_in(wire_d7_25),.data_out(wire_d7_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8727(.data_in(wire_d7_26),.data_out(wire_d7_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8728(.data_in(wire_d7_27),.data_out(wire_d7_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8729(.data_in(wire_d7_28),.data_out(wire_d7_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8730(.data_in(wire_d7_29),.data_out(wire_d7_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8731(.data_in(wire_d7_30),.data_out(wire_d7_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8732(.data_in(wire_d7_31),.data_out(wire_d7_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8733(.data_in(wire_d7_32),.data_out(wire_d7_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8734(.data_in(wire_d7_33),.data_out(wire_d7_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8735(.data_in(wire_d7_34),.data_out(wire_d7_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8736(.data_in(wire_d7_35),.data_out(wire_d7_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8737(.data_in(wire_d7_36),.data_out(wire_d7_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8738(.data_in(wire_d7_37),.data_out(wire_d7_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8739(.data_in(wire_d7_38),.data_out(wire_d7_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8740(.data_in(wire_d7_39),.data_out(wire_d7_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8741(.data_in(wire_d7_40),.data_out(wire_d7_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8742(.data_in(wire_d7_41),.data_out(wire_d7_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8743(.data_in(wire_d7_42),.data_out(wire_d7_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8744(.data_in(wire_d7_43),.data_out(wire_d7_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8745(.data_in(wire_d7_44),.data_out(wire_d7_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8746(.data_in(wire_d7_45),.data_out(wire_d7_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8747(.data_in(wire_d7_46),.data_out(wire_d7_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8748(.data_in(wire_d7_47),.data_out(wire_d7_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8749(.data_in(wire_d7_48),.data_out(wire_d7_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8750(.data_in(wire_d7_49),.data_out(wire_d7_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8751(.data_in(wire_d7_50),.data_out(wire_d7_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8752(.data_in(wire_d7_51),.data_out(wire_d7_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8753(.data_in(wire_d7_52),.data_out(wire_d7_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8754(.data_in(wire_d7_53),.data_out(wire_d7_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8755(.data_in(wire_d7_54),.data_out(wire_d7_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8756(.data_in(wire_d7_55),.data_out(wire_d7_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8757(.data_in(wire_d7_56),.data_out(wire_d7_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8758(.data_in(wire_d7_57),.data_out(wire_d7_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8759(.data_in(wire_d7_58),.data_out(wire_d7_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8760(.data_in(wire_d7_59),.data_out(wire_d7_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8761(.data_in(wire_d7_60),.data_out(wire_d7_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8762(.data_in(wire_d7_61),.data_out(wire_d7_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8763(.data_in(wire_d7_62),.data_out(wire_d7_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8764(.data_in(wire_d7_63),.data_out(wire_d7_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8765(.data_in(wire_d7_64),.data_out(wire_d7_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8766(.data_in(wire_d7_65),.data_out(wire_d7_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8767(.data_in(wire_d7_66),.data_out(wire_d7_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8768(.data_in(wire_d7_67),.data_out(wire_d7_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8769(.data_in(wire_d7_68),.data_out(wire_d7_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8770(.data_in(wire_d7_69),.data_out(wire_d7_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8771(.data_in(wire_d7_70),.data_out(wire_d7_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8772(.data_in(wire_d7_71),.data_out(wire_d7_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8773(.data_in(wire_d7_72),.data_out(wire_d7_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8774(.data_in(wire_d7_73),.data_out(wire_d7_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8775(.data_in(wire_d7_74),.data_out(wire_d7_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8776(.data_in(wire_d7_75),.data_out(wire_d7_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8777(.data_in(wire_d7_76),.data_out(wire_d7_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8778(.data_in(wire_d7_77),.data_out(wire_d7_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8779(.data_in(wire_d7_78),.data_out(wire_d7_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8780(.data_in(wire_d7_79),.data_out(wire_d7_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8781(.data_in(wire_d7_80),.data_out(wire_d7_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8782(.data_in(wire_d7_81),.data_out(wire_d7_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8783(.data_in(wire_d7_82),.data_out(wire_d7_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8784(.data_in(wire_d7_83),.data_out(wire_d7_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8785(.data_in(wire_d7_84),.data_out(wire_d7_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8786(.data_in(wire_d7_85),.data_out(wire_d7_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8787(.data_in(wire_d7_86),.data_out(wire_d7_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8788(.data_in(wire_d7_87),.data_out(wire_d7_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8789(.data_in(wire_d7_88),.data_out(wire_d7_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8790(.data_in(wire_d7_89),.data_out(wire_d7_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8791(.data_in(wire_d7_90),.data_out(wire_d7_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8792(.data_in(wire_d7_91),.data_out(wire_d7_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8793(.data_in(wire_d7_92),.data_out(wire_d7_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8794(.data_in(wire_d7_93),.data_out(wire_d7_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8795(.data_in(wire_d7_94),.data_out(wire_d7_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8796(.data_in(wire_d7_95),.data_out(wire_d7_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8797(.data_in(wire_d7_96),.data_out(wire_d7_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8798(.data_in(wire_d7_97),.data_out(wire_d7_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8799(.data_in(wire_d7_98),.data_out(wire_d7_99),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87100(.data_in(wire_d7_99),.data_out(wire_d7_100),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87101(.data_in(wire_d7_100),.data_out(wire_d7_101),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87102(.data_in(wire_d7_101),.data_out(wire_d7_102),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87103(.data_in(wire_d7_102),.data_out(wire_d7_103),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87104(.data_in(wire_d7_103),.data_out(wire_d7_104),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87105(.data_in(wire_d7_104),.data_out(wire_d7_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87106(.data_in(wire_d7_105),.data_out(wire_d7_106),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87107(.data_in(wire_d7_106),.data_out(wire_d7_107),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87108(.data_in(wire_d7_107),.data_out(wire_d7_108),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87109(.data_in(wire_d7_108),.data_out(wire_d7_109),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87110(.data_in(wire_d7_109),.data_out(wire_d7_110),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87111(.data_in(wire_d7_110),.data_out(wire_d7_111),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87112(.data_in(wire_d7_111),.data_out(wire_d7_112),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87113(.data_in(wire_d7_112),.data_out(wire_d7_113),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87114(.data_in(wire_d7_113),.data_out(wire_d7_114),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87115(.data_in(wire_d7_114),.data_out(wire_d7_115),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87116(.data_in(wire_d7_115),.data_out(wire_d7_116),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87117(.data_in(wire_d7_116),.data_out(wire_d7_117),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87118(.data_in(wire_d7_117),.data_out(wire_d7_118),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87119(.data_in(wire_d7_118),.data_out(wire_d7_119),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87120(.data_in(wire_d7_119),.data_out(wire_d7_120),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87121(.data_in(wire_d7_120),.data_out(wire_d7_121),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87122(.data_in(wire_d7_121),.data_out(wire_d7_122),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87123(.data_in(wire_d7_122),.data_out(wire_d7_123),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87124(.data_in(wire_d7_123),.data_out(wire_d7_124),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87125(.data_in(wire_d7_124),.data_out(wire_d7_125),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87126(.data_in(wire_d7_125),.data_out(wire_d7_126),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87127(.data_in(wire_d7_126),.data_out(wire_d7_127),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87128(.data_in(wire_d7_127),.data_out(wire_d7_128),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87129(.data_in(wire_d7_128),.data_out(wire_d7_129),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87130(.data_in(wire_d7_129),.data_out(wire_d7_130),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87131(.data_in(wire_d7_130),.data_out(wire_d7_131),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87132(.data_in(wire_d7_131),.data_out(wire_d7_132),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87133(.data_in(wire_d7_132),.data_out(wire_d7_133),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87134(.data_in(wire_d7_133),.data_out(wire_d7_134),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87135(.data_in(wire_d7_134),.data_out(wire_d7_135),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87136(.data_in(wire_d7_135),.data_out(wire_d7_136),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87137(.data_in(wire_d7_136),.data_out(wire_d7_137),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87138(.data_in(wire_d7_137),.data_out(wire_d7_138),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87139(.data_in(wire_d7_138),.data_out(wire_d7_139),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87140(.data_in(wire_d7_139),.data_out(wire_d7_140),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87141(.data_in(wire_d7_140),.data_out(wire_d7_141),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87142(.data_in(wire_d7_141),.data_out(wire_d7_142),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87143(.data_in(wire_d7_142),.data_out(wire_d7_143),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87144(.data_in(wire_d7_143),.data_out(wire_d7_144),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87145(.data_in(wire_d7_144),.data_out(wire_d7_145),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87146(.data_in(wire_d7_145),.data_out(wire_d7_146),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87147(.data_in(wire_d7_146),.data_out(wire_d7_147),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87148(.data_in(wire_d7_147),.data_out(wire_d7_148),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87149(.data_in(wire_d7_148),.data_out(wire_d7_149),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87150(.data_in(wire_d7_149),.data_out(wire_d7_150),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87151(.data_in(wire_d7_150),.data_out(wire_d7_151),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87152(.data_in(wire_d7_151),.data_out(wire_d7_152),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87153(.data_in(wire_d7_152),.data_out(wire_d7_153),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87154(.data_in(wire_d7_153),.data_out(wire_d7_154),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87155(.data_in(wire_d7_154),.data_out(wire_d7_155),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87156(.data_in(wire_d7_155),.data_out(wire_d7_156),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87157(.data_in(wire_d7_156),.data_out(wire_d7_157),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87158(.data_in(wire_d7_157),.data_out(wire_d7_158),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87159(.data_in(wire_d7_158),.data_out(wire_d7_159),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87160(.data_in(wire_d7_159),.data_out(wire_d7_160),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87161(.data_in(wire_d7_160),.data_out(wire_d7_161),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87162(.data_in(wire_d7_161),.data_out(wire_d7_162),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87163(.data_in(wire_d7_162),.data_out(wire_d7_163),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87164(.data_in(wire_d7_163),.data_out(wire_d7_164),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87165(.data_in(wire_d7_164),.data_out(wire_d7_165),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87166(.data_in(wire_d7_165),.data_out(wire_d7_166),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87167(.data_in(wire_d7_166),.data_out(wire_d7_167),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87168(.data_in(wire_d7_167),.data_out(wire_d7_168),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87169(.data_in(wire_d7_168),.data_out(wire_d7_169),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87170(.data_in(wire_d7_169),.data_out(wire_d7_170),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87171(.data_in(wire_d7_170),.data_out(wire_d7_171),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87172(.data_in(wire_d7_171),.data_out(wire_d7_172),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87173(.data_in(wire_d7_172),.data_out(wire_d7_173),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87174(.data_in(wire_d7_173),.data_out(wire_d7_174),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87175(.data_in(wire_d7_174),.data_out(wire_d7_175),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87176(.data_in(wire_d7_175),.data_out(wire_d7_176),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87177(.data_in(wire_d7_176),.data_out(wire_d7_177),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87178(.data_in(wire_d7_177),.data_out(wire_d7_178),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87179(.data_in(wire_d7_178),.data_out(wire_d7_179),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87180(.data_in(wire_d7_179),.data_out(wire_d7_180),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87181(.data_in(wire_d7_180),.data_out(wire_d7_181),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87182(.data_in(wire_d7_181),.data_out(wire_d7_182),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87183(.data_in(wire_d7_182),.data_out(wire_d7_183),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87184(.data_in(wire_d7_183),.data_out(wire_d7_184),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87185(.data_in(wire_d7_184),.data_out(wire_d7_185),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87186(.data_in(wire_d7_185),.data_out(wire_d7_186),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87187(.data_in(wire_d7_186),.data_out(wire_d7_187),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87188(.data_in(wire_d7_187),.data_out(wire_d7_188),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87189(.data_in(wire_d7_188),.data_out(wire_d7_189),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87190(.data_in(wire_d7_189),.data_out(wire_d7_190),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87191(.data_in(wire_d7_190),.data_out(wire_d7_191),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87192(.data_in(wire_d7_191),.data_out(wire_d7_192),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87193(.data_in(wire_d7_192),.data_out(wire_d7_193),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87194(.data_in(wire_d7_193),.data_out(wire_d7_194),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87195(.data_in(wire_d7_194),.data_out(wire_d7_195),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87196(.data_in(wire_d7_195),.data_out(wire_d7_196),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87197(.data_in(wire_d7_196),.data_out(wire_d7_197),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87198(.data_in(wire_d7_197),.data_out(wire_d7_198),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87199(.data_in(wire_d7_198),.data_out(d_out7),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance980(.data_in(d_in8),.data_out(wire_d8_0),.clk(clk),.rst(rst));            //channel 9
	encoder #(.WIDTH(WIDTH)) encoder_instance981(.data_in(wire_d8_0),.data_out(wire_d8_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance982(.data_in(wire_d8_1),.data_out(wire_d8_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance983(.data_in(wire_d8_2),.data_out(wire_d8_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance984(.data_in(wire_d8_3),.data_out(wire_d8_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance985(.data_in(wire_d8_4),.data_out(wire_d8_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance986(.data_in(wire_d8_5),.data_out(wire_d8_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance987(.data_in(wire_d8_6),.data_out(wire_d8_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance988(.data_in(wire_d8_7),.data_out(wire_d8_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance989(.data_in(wire_d8_8),.data_out(wire_d8_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9810(.data_in(wire_d8_9),.data_out(wire_d8_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9811(.data_in(wire_d8_10),.data_out(wire_d8_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9812(.data_in(wire_d8_11),.data_out(wire_d8_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9813(.data_in(wire_d8_12),.data_out(wire_d8_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9814(.data_in(wire_d8_13),.data_out(wire_d8_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9815(.data_in(wire_d8_14),.data_out(wire_d8_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9816(.data_in(wire_d8_15),.data_out(wire_d8_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9817(.data_in(wire_d8_16),.data_out(wire_d8_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9818(.data_in(wire_d8_17),.data_out(wire_d8_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9819(.data_in(wire_d8_18),.data_out(wire_d8_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9820(.data_in(wire_d8_19),.data_out(wire_d8_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9821(.data_in(wire_d8_20),.data_out(wire_d8_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9822(.data_in(wire_d8_21),.data_out(wire_d8_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9823(.data_in(wire_d8_22),.data_out(wire_d8_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9824(.data_in(wire_d8_23),.data_out(wire_d8_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9825(.data_in(wire_d8_24),.data_out(wire_d8_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9826(.data_in(wire_d8_25),.data_out(wire_d8_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9827(.data_in(wire_d8_26),.data_out(wire_d8_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9828(.data_in(wire_d8_27),.data_out(wire_d8_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9829(.data_in(wire_d8_28),.data_out(wire_d8_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9830(.data_in(wire_d8_29),.data_out(wire_d8_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9831(.data_in(wire_d8_30),.data_out(wire_d8_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9832(.data_in(wire_d8_31),.data_out(wire_d8_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9833(.data_in(wire_d8_32),.data_out(wire_d8_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9834(.data_in(wire_d8_33),.data_out(wire_d8_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9835(.data_in(wire_d8_34),.data_out(wire_d8_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9836(.data_in(wire_d8_35),.data_out(wire_d8_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9837(.data_in(wire_d8_36),.data_out(wire_d8_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9838(.data_in(wire_d8_37),.data_out(wire_d8_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9839(.data_in(wire_d8_38),.data_out(wire_d8_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9840(.data_in(wire_d8_39),.data_out(wire_d8_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9841(.data_in(wire_d8_40),.data_out(wire_d8_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9842(.data_in(wire_d8_41),.data_out(wire_d8_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9843(.data_in(wire_d8_42),.data_out(wire_d8_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9844(.data_in(wire_d8_43),.data_out(wire_d8_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9845(.data_in(wire_d8_44),.data_out(wire_d8_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9846(.data_in(wire_d8_45),.data_out(wire_d8_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9847(.data_in(wire_d8_46),.data_out(wire_d8_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9848(.data_in(wire_d8_47),.data_out(wire_d8_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9849(.data_in(wire_d8_48),.data_out(wire_d8_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9850(.data_in(wire_d8_49),.data_out(wire_d8_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9851(.data_in(wire_d8_50),.data_out(wire_d8_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9852(.data_in(wire_d8_51),.data_out(wire_d8_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9853(.data_in(wire_d8_52),.data_out(wire_d8_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9854(.data_in(wire_d8_53),.data_out(wire_d8_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9855(.data_in(wire_d8_54),.data_out(wire_d8_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9856(.data_in(wire_d8_55),.data_out(wire_d8_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9857(.data_in(wire_d8_56),.data_out(wire_d8_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9858(.data_in(wire_d8_57),.data_out(wire_d8_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9859(.data_in(wire_d8_58),.data_out(wire_d8_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9860(.data_in(wire_d8_59),.data_out(wire_d8_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9861(.data_in(wire_d8_60),.data_out(wire_d8_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9862(.data_in(wire_d8_61),.data_out(wire_d8_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9863(.data_in(wire_d8_62),.data_out(wire_d8_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9864(.data_in(wire_d8_63),.data_out(wire_d8_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9865(.data_in(wire_d8_64),.data_out(wire_d8_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9866(.data_in(wire_d8_65),.data_out(wire_d8_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9867(.data_in(wire_d8_66),.data_out(wire_d8_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9868(.data_in(wire_d8_67),.data_out(wire_d8_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9869(.data_in(wire_d8_68),.data_out(wire_d8_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9870(.data_in(wire_d8_69),.data_out(wire_d8_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9871(.data_in(wire_d8_70),.data_out(wire_d8_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9872(.data_in(wire_d8_71),.data_out(wire_d8_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9873(.data_in(wire_d8_72),.data_out(wire_d8_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9874(.data_in(wire_d8_73),.data_out(wire_d8_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9875(.data_in(wire_d8_74),.data_out(wire_d8_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9876(.data_in(wire_d8_75),.data_out(wire_d8_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9877(.data_in(wire_d8_76),.data_out(wire_d8_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9878(.data_in(wire_d8_77),.data_out(wire_d8_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9879(.data_in(wire_d8_78),.data_out(wire_d8_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9880(.data_in(wire_d8_79),.data_out(wire_d8_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9881(.data_in(wire_d8_80),.data_out(wire_d8_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9882(.data_in(wire_d8_81),.data_out(wire_d8_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9883(.data_in(wire_d8_82),.data_out(wire_d8_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9884(.data_in(wire_d8_83),.data_out(wire_d8_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9885(.data_in(wire_d8_84),.data_out(wire_d8_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9886(.data_in(wire_d8_85),.data_out(wire_d8_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9887(.data_in(wire_d8_86),.data_out(wire_d8_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9888(.data_in(wire_d8_87),.data_out(wire_d8_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9889(.data_in(wire_d8_88),.data_out(wire_d8_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9890(.data_in(wire_d8_89),.data_out(wire_d8_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9891(.data_in(wire_d8_90),.data_out(wire_d8_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9892(.data_in(wire_d8_91),.data_out(wire_d8_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9893(.data_in(wire_d8_92),.data_out(wire_d8_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9894(.data_in(wire_d8_93),.data_out(wire_d8_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9895(.data_in(wire_d8_94),.data_out(wire_d8_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9896(.data_in(wire_d8_95),.data_out(wire_d8_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9897(.data_in(wire_d8_96),.data_out(wire_d8_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9898(.data_in(wire_d8_97),.data_out(wire_d8_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9899(.data_in(wire_d8_98),.data_out(wire_d8_99),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98100(.data_in(wire_d8_99),.data_out(wire_d8_100),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98101(.data_in(wire_d8_100),.data_out(wire_d8_101),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98102(.data_in(wire_d8_101),.data_out(wire_d8_102),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98103(.data_in(wire_d8_102),.data_out(wire_d8_103),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98104(.data_in(wire_d8_103),.data_out(wire_d8_104),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98105(.data_in(wire_d8_104),.data_out(wire_d8_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98106(.data_in(wire_d8_105),.data_out(wire_d8_106),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98107(.data_in(wire_d8_106),.data_out(wire_d8_107),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98108(.data_in(wire_d8_107),.data_out(wire_d8_108),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98109(.data_in(wire_d8_108),.data_out(wire_d8_109),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98110(.data_in(wire_d8_109),.data_out(wire_d8_110),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98111(.data_in(wire_d8_110),.data_out(wire_d8_111),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98112(.data_in(wire_d8_111),.data_out(wire_d8_112),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98113(.data_in(wire_d8_112),.data_out(wire_d8_113),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98114(.data_in(wire_d8_113),.data_out(wire_d8_114),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98115(.data_in(wire_d8_114),.data_out(wire_d8_115),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98116(.data_in(wire_d8_115),.data_out(wire_d8_116),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98117(.data_in(wire_d8_116),.data_out(wire_d8_117),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98118(.data_in(wire_d8_117),.data_out(wire_d8_118),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98119(.data_in(wire_d8_118),.data_out(wire_d8_119),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98120(.data_in(wire_d8_119),.data_out(wire_d8_120),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98121(.data_in(wire_d8_120),.data_out(wire_d8_121),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98122(.data_in(wire_d8_121),.data_out(wire_d8_122),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98123(.data_in(wire_d8_122),.data_out(wire_d8_123),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98124(.data_in(wire_d8_123),.data_out(wire_d8_124),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98125(.data_in(wire_d8_124),.data_out(wire_d8_125),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98126(.data_in(wire_d8_125),.data_out(wire_d8_126),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98127(.data_in(wire_d8_126),.data_out(wire_d8_127),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98128(.data_in(wire_d8_127),.data_out(wire_d8_128),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98129(.data_in(wire_d8_128),.data_out(wire_d8_129),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98130(.data_in(wire_d8_129),.data_out(wire_d8_130),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98131(.data_in(wire_d8_130),.data_out(wire_d8_131),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98132(.data_in(wire_d8_131),.data_out(wire_d8_132),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98133(.data_in(wire_d8_132),.data_out(wire_d8_133),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98134(.data_in(wire_d8_133),.data_out(wire_d8_134),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98135(.data_in(wire_d8_134),.data_out(wire_d8_135),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98136(.data_in(wire_d8_135),.data_out(wire_d8_136),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98137(.data_in(wire_d8_136),.data_out(wire_d8_137),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98138(.data_in(wire_d8_137),.data_out(wire_d8_138),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98139(.data_in(wire_d8_138),.data_out(wire_d8_139),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98140(.data_in(wire_d8_139),.data_out(wire_d8_140),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98141(.data_in(wire_d8_140),.data_out(wire_d8_141),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98142(.data_in(wire_d8_141),.data_out(wire_d8_142),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98143(.data_in(wire_d8_142),.data_out(wire_d8_143),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98144(.data_in(wire_d8_143),.data_out(wire_d8_144),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98145(.data_in(wire_d8_144),.data_out(wire_d8_145),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98146(.data_in(wire_d8_145),.data_out(wire_d8_146),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98147(.data_in(wire_d8_146),.data_out(wire_d8_147),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98148(.data_in(wire_d8_147),.data_out(wire_d8_148),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98149(.data_in(wire_d8_148),.data_out(wire_d8_149),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98150(.data_in(wire_d8_149),.data_out(wire_d8_150),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98151(.data_in(wire_d8_150),.data_out(wire_d8_151),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98152(.data_in(wire_d8_151),.data_out(wire_d8_152),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98153(.data_in(wire_d8_152),.data_out(wire_d8_153),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98154(.data_in(wire_d8_153),.data_out(wire_d8_154),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98155(.data_in(wire_d8_154),.data_out(wire_d8_155),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98156(.data_in(wire_d8_155),.data_out(wire_d8_156),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98157(.data_in(wire_d8_156),.data_out(wire_d8_157),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98158(.data_in(wire_d8_157),.data_out(wire_d8_158),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98159(.data_in(wire_d8_158),.data_out(wire_d8_159),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98160(.data_in(wire_d8_159),.data_out(wire_d8_160),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98161(.data_in(wire_d8_160),.data_out(wire_d8_161),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98162(.data_in(wire_d8_161),.data_out(wire_d8_162),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98163(.data_in(wire_d8_162),.data_out(wire_d8_163),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98164(.data_in(wire_d8_163),.data_out(wire_d8_164),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98165(.data_in(wire_d8_164),.data_out(wire_d8_165),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98166(.data_in(wire_d8_165),.data_out(wire_d8_166),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98167(.data_in(wire_d8_166),.data_out(wire_d8_167),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98168(.data_in(wire_d8_167),.data_out(wire_d8_168),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98169(.data_in(wire_d8_168),.data_out(wire_d8_169),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98170(.data_in(wire_d8_169),.data_out(wire_d8_170),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98171(.data_in(wire_d8_170),.data_out(wire_d8_171),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98172(.data_in(wire_d8_171),.data_out(wire_d8_172),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98173(.data_in(wire_d8_172),.data_out(wire_d8_173),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98174(.data_in(wire_d8_173),.data_out(wire_d8_174),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98175(.data_in(wire_d8_174),.data_out(wire_d8_175),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98176(.data_in(wire_d8_175),.data_out(wire_d8_176),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98177(.data_in(wire_d8_176),.data_out(wire_d8_177),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98178(.data_in(wire_d8_177),.data_out(wire_d8_178),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98179(.data_in(wire_d8_178),.data_out(wire_d8_179),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98180(.data_in(wire_d8_179),.data_out(wire_d8_180),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98181(.data_in(wire_d8_180),.data_out(wire_d8_181),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98182(.data_in(wire_d8_181),.data_out(wire_d8_182),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98183(.data_in(wire_d8_182),.data_out(wire_d8_183),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98184(.data_in(wire_d8_183),.data_out(wire_d8_184),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98185(.data_in(wire_d8_184),.data_out(wire_d8_185),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98186(.data_in(wire_d8_185),.data_out(wire_d8_186),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98187(.data_in(wire_d8_186),.data_out(wire_d8_187),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98188(.data_in(wire_d8_187),.data_out(wire_d8_188),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98189(.data_in(wire_d8_188),.data_out(wire_d8_189),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98190(.data_in(wire_d8_189),.data_out(wire_d8_190),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98191(.data_in(wire_d8_190),.data_out(wire_d8_191),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98192(.data_in(wire_d8_191),.data_out(wire_d8_192),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98193(.data_in(wire_d8_192),.data_out(wire_d8_193),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98194(.data_in(wire_d8_193),.data_out(wire_d8_194),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98195(.data_in(wire_d8_194),.data_out(wire_d8_195),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98196(.data_in(wire_d8_195),.data_out(wire_d8_196),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98197(.data_in(wire_d8_196),.data_out(wire_d8_197),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98198(.data_in(wire_d8_197),.data_out(wire_d8_198),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98199(.data_in(wire_d8_198),.data_out(d_out8),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance10090(.data_in(d_in9),.data_out(wire_d9_0),.clk(clk),.rst(rst));            //channel 10
	encoder #(.WIDTH(WIDTH)) encoder_instance10091(.data_in(wire_d9_0),.data_out(wire_d9_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10092(.data_in(wire_d9_1),.data_out(wire_d9_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10093(.data_in(wire_d9_2),.data_out(wire_d9_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10094(.data_in(wire_d9_3),.data_out(wire_d9_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10095(.data_in(wire_d9_4),.data_out(wire_d9_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10096(.data_in(wire_d9_5),.data_out(wire_d9_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10097(.data_in(wire_d9_6),.data_out(wire_d9_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10098(.data_in(wire_d9_7),.data_out(wire_d9_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10099(.data_in(wire_d9_8),.data_out(wire_d9_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100910(.data_in(wire_d9_9),.data_out(wire_d9_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100911(.data_in(wire_d9_10),.data_out(wire_d9_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100912(.data_in(wire_d9_11),.data_out(wire_d9_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100913(.data_in(wire_d9_12),.data_out(wire_d9_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100914(.data_in(wire_d9_13),.data_out(wire_d9_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100915(.data_in(wire_d9_14),.data_out(wire_d9_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100916(.data_in(wire_d9_15),.data_out(wire_d9_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100917(.data_in(wire_d9_16),.data_out(wire_d9_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100918(.data_in(wire_d9_17),.data_out(wire_d9_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100919(.data_in(wire_d9_18),.data_out(wire_d9_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100920(.data_in(wire_d9_19),.data_out(wire_d9_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100921(.data_in(wire_d9_20),.data_out(wire_d9_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100922(.data_in(wire_d9_21),.data_out(wire_d9_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100923(.data_in(wire_d9_22),.data_out(wire_d9_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100924(.data_in(wire_d9_23),.data_out(wire_d9_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100925(.data_in(wire_d9_24),.data_out(wire_d9_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100926(.data_in(wire_d9_25),.data_out(wire_d9_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100927(.data_in(wire_d9_26),.data_out(wire_d9_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100928(.data_in(wire_d9_27),.data_out(wire_d9_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100929(.data_in(wire_d9_28),.data_out(wire_d9_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100930(.data_in(wire_d9_29),.data_out(wire_d9_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100931(.data_in(wire_d9_30),.data_out(wire_d9_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100932(.data_in(wire_d9_31),.data_out(wire_d9_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100933(.data_in(wire_d9_32),.data_out(wire_d9_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100934(.data_in(wire_d9_33),.data_out(wire_d9_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100935(.data_in(wire_d9_34),.data_out(wire_d9_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100936(.data_in(wire_d9_35),.data_out(wire_d9_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100937(.data_in(wire_d9_36),.data_out(wire_d9_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100938(.data_in(wire_d9_37),.data_out(wire_d9_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100939(.data_in(wire_d9_38),.data_out(wire_d9_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100940(.data_in(wire_d9_39),.data_out(wire_d9_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100941(.data_in(wire_d9_40),.data_out(wire_d9_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100942(.data_in(wire_d9_41),.data_out(wire_d9_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100943(.data_in(wire_d9_42),.data_out(wire_d9_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100944(.data_in(wire_d9_43),.data_out(wire_d9_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100945(.data_in(wire_d9_44),.data_out(wire_d9_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100946(.data_in(wire_d9_45),.data_out(wire_d9_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100947(.data_in(wire_d9_46),.data_out(wire_d9_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100948(.data_in(wire_d9_47),.data_out(wire_d9_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100949(.data_in(wire_d9_48),.data_out(wire_d9_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100950(.data_in(wire_d9_49),.data_out(wire_d9_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100951(.data_in(wire_d9_50),.data_out(wire_d9_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100952(.data_in(wire_d9_51),.data_out(wire_d9_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100953(.data_in(wire_d9_52),.data_out(wire_d9_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100954(.data_in(wire_d9_53),.data_out(wire_d9_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100955(.data_in(wire_d9_54),.data_out(wire_d9_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100956(.data_in(wire_d9_55),.data_out(wire_d9_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100957(.data_in(wire_d9_56),.data_out(wire_d9_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100958(.data_in(wire_d9_57),.data_out(wire_d9_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100959(.data_in(wire_d9_58),.data_out(wire_d9_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100960(.data_in(wire_d9_59),.data_out(wire_d9_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100961(.data_in(wire_d9_60),.data_out(wire_d9_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100962(.data_in(wire_d9_61),.data_out(wire_d9_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100963(.data_in(wire_d9_62),.data_out(wire_d9_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100964(.data_in(wire_d9_63),.data_out(wire_d9_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100965(.data_in(wire_d9_64),.data_out(wire_d9_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100966(.data_in(wire_d9_65),.data_out(wire_d9_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100967(.data_in(wire_d9_66),.data_out(wire_d9_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100968(.data_in(wire_d9_67),.data_out(wire_d9_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100969(.data_in(wire_d9_68),.data_out(wire_d9_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100970(.data_in(wire_d9_69),.data_out(wire_d9_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100971(.data_in(wire_d9_70),.data_out(wire_d9_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100972(.data_in(wire_d9_71),.data_out(wire_d9_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100973(.data_in(wire_d9_72),.data_out(wire_d9_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100974(.data_in(wire_d9_73),.data_out(wire_d9_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100975(.data_in(wire_d9_74),.data_out(wire_d9_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100976(.data_in(wire_d9_75),.data_out(wire_d9_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100977(.data_in(wire_d9_76),.data_out(wire_d9_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100978(.data_in(wire_d9_77),.data_out(wire_d9_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100979(.data_in(wire_d9_78),.data_out(wire_d9_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100980(.data_in(wire_d9_79),.data_out(wire_d9_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100981(.data_in(wire_d9_80),.data_out(wire_d9_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100982(.data_in(wire_d9_81),.data_out(wire_d9_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100983(.data_in(wire_d9_82),.data_out(wire_d9_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100984(.data_in(wire_d9_83),.data_out(wire_d9_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100985(.data_in(wire_d9_84),.data_out(wire_d9_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100986(.data_in(wire_d9_85),.data_out(wire_d9_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100987(.data_in(wire_d9_86),.data_out(wire_d9_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100988(.data_in(wire_d9_87),.data_out(wire_d9_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100989(.data_in(wire_d9_88),.data_out(wire_d9_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100990(.data_in(wire_d9_89),.data_out(wire_d9_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100991(.data_in(wire_d9_90),.data_out(wire_d9_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100992(.data_in(wire_d9_91),.data_out(wire_d9_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100993(.data_in(wire_d9_92),.data_out(wire_d9_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100994(.data_in(wire_d9_93),.data_out(wire_d9_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100995(.data_in(wire_d9_94),.data_out(wire_d9_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100996(.data_in(wire_d9_95),.data_out(wire_d9_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100997(.data_in(wire_d9_96),.data_out(wire_d9_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100998(.data_in(wire_d9_97),.data_out(wire_d9_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100999(.data_in(wire_d9_98),.data_out(wire_d9_99),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009100(.data_in(wire_d9_99),.data_out(wire_d9_100),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009101(.data_in(wire_d9_100),.data_out(wire_d9_101),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009102(.data_in(wire_d9_101),.data_out(wire_d9_102),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009103(.data_in(wire_d9_102),.data_out(wire_d9_103),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009104(.data_in(wire_d9_103),.data_out(wire_d9_104),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009105(.data_in(wire_d9_104),.data_out(wire_d9_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009106(.data_in(wire_d9_105),.data_out(wire_d9_106),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009107(.data_in(wire_d9_106),.data_out(wire_d9_107),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009108(.data_in(wire_d9_107),.data_out(wire_d9_108),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009109(.data_in(wire_d9_108),.data_out(wire_d9_109),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009110(.data_in(wire_d9_109),.data_out(wire_d9_110),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009111(.data_in(wire_d9_110),.data_out(wire_d9_111),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009112(.data_in(wire_d9_111),.data_out(wire_d9_112),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009113(.data_in(wire_d9_112),.data_out(wire_d9_113),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009114(.data_in(wire_d9_113),.data_out(wire_d9_114),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009115(.data_in(wire_d9_114),.data_out(wire_d9_115),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009116(.data_in(wire_d9_115),.data_out(wire_d9_116),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009117(.data_in(wire_d9_116),.data_out(wire_d9_117),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009118(.data_in(wire_d9_117),.data_out(wire_d9_118),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009119(.data_in(wire_d9_118),.data_out(wire_d9_119),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009120(.data_in(wire_d9_119),.data_out(wire_d9_120),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009121(.data_in(wire_d9_120),.data_out(wire_d9_121),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009122(.data_in(wire_d9_121),.data_out(wire_d9_122),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009123(.data_in(wire_d9_122),.data_out(wire_d9_123),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009124(.data_in(wire_d9_123),.data_out(wire_d9_124),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009125(.data_in(wire_d9_124),.data_out(wire_d9_125),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009126(.data_in(wire_d9_125),.data_out(wire_d9_126),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009127(.data_in(wire_d9_126),.data_out(wire_d9_127),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009128(.data_in(wire_d9_127),.data_out(wire_d9_128),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009129(.data_in(wire_d9_128),.data_out(wire_d9_129),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009130(.data_in(wire_d9_129),.data_out(wire_d9_130),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009131(.data_in(wire_d9_130),.data_out(wire_d9_131),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009132(.data_in(wire_d9_131),.data_out(wire_d9_132),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009133(.data_in(wire_d9_132),.data_out(wire_d9_133),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009134(.data_in(wire_d9_133),.data_out(wire_d9_134),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009135(.data_in(wire_d9_134),.data_out(wire_d9_135),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009136(.data_in(wire_d9_135),.data_out(wire_d9_136),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009137(.data_in(wire_d9_136),.data_out(wire_d9_137),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009138(.data_in(wire_d9_137),.data_out(wire_d9_138),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009139(.data_in(wire_d9_138),.data_out(wire_d9_139),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009140(.data_in(wire_d9_139),.data_out(wire_d9_140),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009141(.data_in(wire_d9_140),.data_out(wire_d9_141),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009142(.data_in(wire_d9_141),.data_out(wire_d9_142),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009143(.data_in(wire_d9_142),.data_out(wire_d9_143),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009144(.data_in(wire_d9_143),.data_out(wire_d9_144),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009145(.data_in(wire_d9_144),.data_out(wire_d9_145),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009146(.data_in(wire_d9_145),.data_out(wire_d9_146),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009147(.data_in(wire_d9_146),.data_out(wire_d9_147),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009148(.data_in(wire_d9_147),.data_out(wire_d9_148),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009149(.data_in(wire_d9_148),.data_out(wire_d9_149),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009150(.data_in(wire_d9_149),.data_out(wire_d9_150),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009151(.data_in(wire_d9_150),.data_out(wire_d9_151),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009152(.data_in(wire_d9_151),.data_out(wire_d9_152),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009153(.data_in(wire_d9_152),.data_out(wire_d9_153),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009154(.data_in(wire_d9_153),.data_out(wire_d9_154),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009155(.data_in(wire_d9_154),.data_out(wire_d9_155),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009156(.data_in(wire_d9_155),.data_out(wire_d9_156),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009157(.data_in(wire_d9_156),.data_out(wire_d9_157),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009158(.data_in(wire_d9_157),.data_out(wire_d9_158),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009159(.data_in(wire_d9_158),.data_out(wire_d9_159),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009160(.data_in(wire_d9_159),.data_out(wire_d9_160),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009161(.data_in(wire_d9_160),.data_out(wire_d9_161),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009162(.data_in(wire_d9_161),.data_out(wire_d9_162),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009163(.data_in(wire_d9_162),.data_out(wire_d9_163),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009164(.data_in(wire_d9_163),.data_out(wire_d9_164),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009165(.data_in(wire_d9_164),.data_out(wire_d9_165),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009166(.data_in(wire_d9_165),.data_out(wire_d9_166),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009167(.data_in(wire_d9_166),.data_out(wire_d9_167),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009168(.data_in(wire_d9_167),.data_out(wire_d9_168),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009169(.data_in(wire_d9_168),.data_out(wire_d9_169),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009170(.data_in(wire_d9_169),.data_out(wire_d9_170),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009171(.data_in(wire_d9_170),.data_out(wire_d9_171),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009172(.data_in(wire_d9_171),.data_out(wire_d9_172),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009173(.data_in(wire_d9_172),.data_out(wire_d9_173),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009174(.data_in(wire_d9_173),.data_out(wire_d9_174),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009175(.data_in(wire_d9_174),.data_out(wire_d9_175),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009176(.data_in(wire_d9_175),.data_out(wire_d9_176),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009177(.data_in(wire_d9_176),.data_out(wire_d9_177),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009178(.data_in(wire_d9_177),.data_out(wire_d9_178),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009179(.data_in(wire_d9_178),.data_out(wire_d9_179),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009180(.data_in(wire_d9_179),.data_out(wire_d9_180),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009181(.data_in(wire_d9_180),.data_out(wire_d9_181),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009182(.data_in(wire_d9_181),.data_out(wire_d9_182),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009183(.data_in(wire_d9_182),.data_out(wire_d9_183),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009184(.data_in(wire_d9_183),.data_out(wire_d9_184),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009185(.data_in(wire_d9_184),.data_out(wire_d9_185),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009186(.data_in(wire_d9_185),.data_out(wire_d9_186),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009187(.data_in(wire_d9_186),.data_out(wire_d9_187),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009188(.data_in(wire_d9_187),.data_out(wire_d9_188),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009189(.data_in(wire_d9_188),.data_out(wire_d9_189),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009190(.data_in(wire_d9_189),.data_out(wire_d9_190),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009191(.data_in(wire_d9_190),.data_out(wire_d9_191),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009192(.data_in(wire_d9_191),.data_out(wire_d9_192),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009193(.data_in(wire_d9_192),.data_out(wire_d9_193),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009194(.data_in(wire_d9_193),.data_out(wire_d9_194),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009195(.data_in(wire_d9_194),.data_out(wire_d9_195),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009196(.data_in(wire_d9_195),.data_out(wire_d9_196),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009197(.data_in(wire_d9_196),.data_out(wire_d9_197),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009198(.data_in(wire_d9_197),.data_out(wire_d9_198),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009199(.data_in(wire_d9_198),.data_out(d_out9),.clk(clk),.rst(rst));


endmodule