`include "encoder.v"
`include "invertion.v"
`include "large_mux.v"
`include "register.v"
module design39_90_100_top #(parameter WIDTH=32,CHANNEL=90) (clk, rst, in, out);

	localparam OUT_BUS=CHANNEL*WIDTH;
	input clk,rst;
	input [WIDTH-1:0] in;
	output [WIDTH-1:0] out;

	reg [WIDTH-1:0] d_in0;
	reg [WIDTH-1:0] d_in1;
	reg [WIDTH-1:0] d_in2;
	reg [WIDTH-1:0] d_in3;
	reg [WIDTH-1:0] d_in4;
	reg [WIDTH-1:0] d_in5;
	reg [WIDTH-1:0] d_in6;
	reg [WIDTH-1:0] d_in7;
	reg [WIDTH-1:0] d_in8;
	reg [WIDTH-1:0] d_in9;
	reg [WIDTH-1:0] d_in10;
	reg [WIDTH-1:0] d_in11;
	reg [WIDTH-1:0] d_in12;
	reg [WIDTH-1:0] d_in13;
	reg [WIDTH-1:0] d_in14;
	reg [WIDTH-1:0] d_in15;
	reg [WIDTH-1:0] d_in16;
	reg [WIDTH-1:0] d_in17;
	reg [WIDTH-1:0] d_in18;
	reg [WIDTH-1:0] d_in19;
	reg [WIDTH-1:0] d_in20;
	reg [WIDTH-1:0] d_in21;
	reg [WIDTH-1:0] d_in22;
	reg [WIDTH-1:0] d_in23;
	reg [WIDTH-1:0] d_in24;
	reg [WIDTH-1:0] d_in25;
	reg [WIDTH-1:0] d_in26;
	reg [WIDTH-1:0] d_in27;
	reg [WIDTH-1:0] d_in28;
	reg [WIDTH-1:0] d_in29;
	reg [WIDTH-1:0] d_in30;
	reg [WIDTH-1:0] d_in31;
	reg [WIDTH-1:0] d_in32;
	reg [WIDTH-1:0] d_in33;
	reg [WIDTH-1:0] d_in34;
	reg [WIDTH-1:0] d_in35;
	reg [WIDTH-1:0] d_in36;
	reg [WIDTH-1:0] d_in37;
	reg [WIDTH-1:0] d_in38;
	reg [WIDTH-1:0] d_in39;
	reg [WIDTH-1:0] d_in40;
	reg [WIDTH-1:0] d_in41;
	reg [WIDTH-1:0] d_in42;
	reg [WIDTH-1:0] d_in43;
	reg [WIDTH-1:0] d_in44;
	reg [WIDTH-1:0] d_in45;
	reg [WIDTH-1:0] d_in46;
	reg [WIDTH-1:0] d_in47;
	reg [WIDTH-1:0] d_in48;
	reg [WIDTH-1:0] d_in49;
	reg [WIDTH-1:0] d_in50;
	reg [WIDTH-1:0] d_in51;
	reg [WIDTH-1:0] d_in52;
	reg [WIDTH-1:0] d_in53;
	reg [WIDTH-1:0] d_in54;
	reg [WIDTH-1:0] d_in55;
	reg [WIDTH-1:0] d_in56;
	reg [WIDTH-1:0] d_in57;
	reg [WIDTH-1:0] d_in58;
	reg [WIDTH-1:0] d_in59;
	reg [WIDTH-1:0] d_in60;
	reg [WIDTH-1:0] d_in61;
	reg [WIDTH-1:0] d_in62;
	reg [WIDTH-1:0] d_in63;
	reg [WIDTH-1:0] d_in64;
	reg [WIDTH-1:0] d_in65;
	reg [WIDTH-1:0] d_in66;
	reg [WIDTH-1:0] d_in67;
	reg [WIDTH-1:0] d_in68;
	reg [WIDTH-1:0] d_in69;
	reg [WIDTH-1:0] d_in70;
	reg [WIDTH-1:0] d_in71;
	reg [WIDTH-1:0] d_in72;
	reg [WIDTH-1:0] d_in73;
	reg [WIDTH-1:0] d_in74;
	reg [WIDTH-1:0] d_in75;
	reg [WIDTH-1:0] d_in76;
	reg [WIDTH-1:0] d_in77;
	reg [WIDTH-1:0] d_in78;
	reg [WIDTH-1:0] d_in79;
	reg [WIDTH-1:0] d_in80;
	reg [WIDTH-1:0] d_in81;
	reg [WIDTH-1:0] d_in82;
	reg [WIDTH-1:0] d_in83;
	reg [WIDTH-1:0] d_in84;
	reg [WIDTH-1:0] d_in85;
	reg [WIDTH-1:0] d_in86;
	reg [WIDTH-1:0] d_in87;
	reg [WIDTH-1:0] d_in88;
	reg [WIDTH-1:0] d_in89;
	wire [WIDTH-1:0] d_out0;
	wire [WIDTH-1:0] d_out1;
	wire [WIDTH-1:0] d_out2;
	wire [WIDTH-1:0] d_out3;
	wire [WIDTH-1:0] d_out4;
	wire [WIDTH-1:0] d_out5;
	wire [WIDTH-1:0] d_out6;
	wire [WIDTH-1:0] d_out7;
	wire [WIDTH-1:0] d_out8;
	wire [WIDTH-1:0] d_out9;
	wire [WIDTH-1:0] d_out10;
	wire [WIDTH-1:0] d_out11;
	wire [WIDTH-1:0] d_out12;
	wire [WIDTH-1:0] d_out13;
	wire [WIDTH-1:0] d_out14;
	wire [WIDTH-1:0] d_out15;
	wire [WIDTH-1:0] d_out16;
	wire [WIDTH-1:0] d_out17;
	wire [WIDTH-1:0] d_out18;
	wire [WIDTH-1:0] d_out19;
	wire [WIDTH-1:0] d_out20;
	wire [WIDTH-1:0] d_out21;
	wire [WIDTH-1:0] d_out22;
	wire [WIDTH-1:0] d_out23;
	wire [WIDTH-1:0] d_out24;
	wire [WIDTH-1:0] d_out25;
	wire [WIDTH-1:0] d_out26;
	wire [WIDTH-1:0] d_out27;
	wire [WIDTH-1:0] d_out28;
	wire [WIDTH-1:0] d_out29;
	wire [WIDTH-1:0] d_out30;
	wire [WIDTH-1:0] d_out31;
	wire [WIDTH-1:0] d_out32;
	wire [WIDTH-1:0] d_out33;
	wire [WIDTH-1:0] d_out34;
	wire [WIDTH-1:0] d_out35;
	wire [WIDTH-1:0] d_out36;
	wire [WIDTH-1:0] d_out37;
	wire [WIDTH-1:0] d_out38;
	wire [WIDTH-1:0] d_out39;
	wire [WIDTH-1:0] d_out40;
	wire [WIDTH-1:0] d_out41;
	wire [WIDTH-1:0] d_out42;
	wire [WIDTH-1:0] d_out43;
	wire [WIDTH-1:0] d_out44;
	wire [WIDTH-1:0] d_out45;
	wire [WIDTH-1:0] d_out46;
	wire [WIDTH-1:0] d_out47;
	wire [WIDTH-1:0] d_out48;
	wire [WIDTH-1:0] d_out49;
	wire [WIDTH-1:0] d_out50;
	wire [WIDTH-1:0] d_out51;
	wire [WIDTH-1:0] d_out52;
	wire [WIDTH-1:0] d_out53;
	wire [WIDTH-1:0] d_out54;
	wire [WIDTH-1:0] d_out55;
	wire [WIDTH-1:0] d_out56;
	wire [WIDTH-1:0] d_out57;
	wire [WIDTH-1:0] d_out58;
	wire [WIDTH-1:0] d_out59;
	wire [WIDTH-1:0] d_out60;
	wire [WIDTH-1:0] d_out61;
	wire [WIDTH-1:0] d_out62;
	wire [WIDTH-1:0] d_out63;
	wire [WIDTH-1:0] d_out64;
	wire [WIDTH-1:0] d_out65;
	wire [WIDTH-1:0] d_out66;
	wire [WIDTH-1:0] d_out67;
	wire [WIDTH-1:0] d_out68;
	wire [WIDTH-1:0] d_out69;
	wire [WIDTH-1:0] d_out70;
	wire [WIDTH-1:0] d_out71;
	wire [WIDTH-1:0] d_out72;
	wire [WIDTH-1:0] d_out73;
	wire [WIDTH-1:0] d_out74;
	wire [WIDTH-1:0] d_out75;
	wire [WIDTH-1:0] d_out76;
	wire [WIDTH-1:0] d_out77;
	wire [WIDTH-1:0] d_out78;
	wire [WIDTH-1:0] d_out79;
	wire [WIDTH-1:0] d_out80;
	wire [WIDTH-1:0] d_out81;
	wire [WIDTH-1:0] d_out82;
	wire [WIDTH-1:0] d_out83;
	wire [WIDTH-1:0] d_out84;
	wire [WIDTH-1:0] d_out85;
	wire [WIDTH-1:0] d_out86;
	wire [WIDTH-1:0] d_out87;
	wire [WIDTH-1:0] d_out88;
	wire [WIDTH-1:0] d_out89;

	reg [OUT_BUS-1:0] tmp;

	always @ (posedge clk or posedge rst) begin
		if (rst)
			tmp <= 0;
		else
			tmp <= {tmp[OUT_BUS-(WIDTH-1):0],in};
	end

	always @ (posedge clk) begin
		d_in0 <= tmp[WIDTH-1:0];
		d_in1 <= tmp[(WIDTH*2)-1:WIDTH*1];
		d_in2 <= tmp[(WIDTH*3)-1:WIDTH*2];
		d_in3 <= tmp[(WIDTH*4)-1:WIDTH*3];
		d_in4 <= tmp[(WIDTH*5)-1:WIDTH*4];
		d_in5 <= tmp[(WIDTH*6)-1:WIDTH*5];
		d_in6 <= tmp[(WIDTH*7)-1:WIDTH*6];
		d_in7 <= tmp[(WIDTH*8)-1:WIDTH*7];
		d_in8 <= tmp[(WIDTH*9)-1:WIDTH*8];
		d_in9 <= tmp[(WIDTH*10)-1:WIDTH*9];
		d_in10 <= tmp[(WIDTH*11)-1:WIDTH*10];
		d_in11 <= tmp[(WIDTH*12)-1:WIDTH*11];
		d_in12 <= tmp[(WIDTH*13)-1:WIDTH*12];
		d_in13 <= tmp[(WIDTH*14)-1:WIDTH*13];
		d_in14 <= tmp[(WIDTH*15)-1:WIDTH*14];
		d_in15 <= tmp[(WIDTH*16)-1:WIDTH*15];
		d_in16 <= tmp[(WIDTH*17)-1:WIDTH*16];
		d_in17 <= tmp[(WIDTH*18)-1:WIDTH*17];
		d_in18 <= tmp[(WIDTH*19)-1:WIDTH*18];
		d_in19 <= tmp[(WIDTH*20)-1:WIDTH*19];
		d_in20 <= tmp[(WIDTH*21)-1:WIDTH*20];
		d_in21 <= tmp[(WIDTH*22)-1:WIDTH*21];
		d_in22 <= tmp[(WIDTH*23)-1:WIDTH*22];
		d_in23 <= tmp[(WIDTH*24)-1:WIDTH*23];
		d_in24 <= tmp[(WIDTH*25)-1:WIDTH*24];
		d_in25 <= tmp[(WIDTH*26)-1:WIDTH*25];
		d_in26 <= tmp[(WIDTH*27)-1:WIDTH*26];
		d_in27 <= tmp[(WIDTH*28)-1:WIDTH*27];
		d_in28 <= tmp[(WIDTH*29)-1:WIDTH*28];
		d_in29 <= tmp[(WIDTH*30)-1:WIDTH*29];
		d_in30 <= tmp[(WIDTH*31)-1:WIDTH*30];
		d_in31 <= tmp[(WIDTH*32)-1:WIDTH*31];
		d_in32 <= tmp[(WIDTH*33)-1:WIDTH*32];
		d_in33 <= tmp[(WIDTH*34)-1:WIDTH*33];
		d_in34 <= tmp[(WIDTH*35)-1:WIDTH*34];
		d_in35 <= tmp[(WIDTH*36)-1:WIDTH*35];
		d_in36 <= tmp[(WIDTH*37)-1:WIDTH*36];
		d_in37 <= tmp[(WIDTH*38)-1:WIDTH*37];
		d_in38 <= tmp[(WIDTH*39)-1:WIDTH*38];
		d_in39 <= tmp[(WIDTH*40)-1:WIDTH*39];
		d_in40 <= tmp[(WIDTH*41)-1:WIDTH*40];
		d_in41 <= tmp[(WIDTH*42)-1:WIDTH*41];
		d_in42 <= tmp[(WIDTH*43)-1:WIDTH*42];
		d_in43 <= tmp[(WIDTH*44)-1:WIDTH*43];
		d_in44 <= tmp[(WIDTH*45)-1:WIDTH*44];
		d_in45 <= tmp[(WIDTH*46)-1:WIDTH*45];
		d_in46 <= tmp[(WIDTH*47)-1:WIDTH*46];
		d_in47 <= tmp[(WIDTH*48)-1:WIDTH*47];
		d_in48 <= tmp[(WIDTH*49)-1:WIDTH*48];
		d_in49 <= tmp[(WIDTH*50)-1:WIDTH*49];
		d_in50 <= tmp[(WIDTH*51)-1:WIDTH*50];
		d_in51 <= tmp[(WIDTH*52)-1:WIDTH*51];
		d_in52 <= tmp[(WIDTH*53)-1:WIDTH*52];
		d_in53 <= tmp[(WIDTH*54)-1:WIDTH*53];
		d_in54 <= tmp[(WIDTH*55)-1:WIDTH*54];
		d_in55 <= tmp[(WIDTH*56)-1:WIDTH*55];
		d_in56 <= tmp[(WIDTH*57)-1:WIDTH*56];
		d_in57 <= tmp[(WIDTH*58)-1:WIDTH*57];
		d_in58 <= tmp[(WIDTH*59)-1:WIDTH*58];
		d_in59 <= tmp[(WIDTH*60)-1:WIDTH*59];
		d_in60 <= tmp[(WIDTH*61)-1:WIDTH*60];
		d_in61 <= tmp[(WIDTH*62)-1:WIDTH*61];
		d_in62 <= tmp[(WIDTH*63)-1:WIDTH*62];
		d_in63 <= tmp[(WIDTH*64)-1:WIDTH*63];
		d_in64 <= tmp[(WIDTH*65)-1:WIDTH*64];
		d_in65 <= tmp[(WIDTH*66)-1:WIDTH*65];
		d_in66 <= tmp[(WIDTH*67)-1:WIDTH*66];
		d_in67 <= tmp[(WIDTH*68)-1:WIDTH*67];
		d_in68 <= tmp[(WIDTH*69)-1:WIDTH*68];
		d_in69 <= tmp[(WIDTH*70)-1:WIDTH*69];
		d_in70 <= tmp[(WIDTH*71)-1:WIDTH*70];
		d_in71 <= tmp[(WIDTH*72)-1:WIDTH*71];
		d_in72 <= tmp[(WIDTH*73)-1:WIDTH*72];
		d_in73 <= tmp[(WIDTH*74)-1:WIDTH*73];
		d_in74 <= tmp[(WIDTH*75)-1:WIDTH*74];
		d_in75 <= tmp[(WIDTH*76)-1:WIDTH*75];
		d_in76 <= tmp[(WIDTH*77)-1:WIDTH*76];
		d_in77 <= tmp[(WIDTH*78)-1:WIDTH*77];
		d_in78 <= tmp[(WIDTH*79)-1:WIDTH*78];
		d_in79 <= tmp[(WIDTH*80)-1:WIDTH*79];
		d_in80 <= tmp[(WIDTH*81)-1:WIDTH*80];
		d_in81 <= tmp[(WIDTH*82)-1:WIDTH*81];
		d_in82 <= tmp[(WIDTH*83)-1:WIDTH*82];
		d_in83 <= tmp[(WIDTH*84)-1:WIDTH*83];
		d_in84 <= tmp[(WIDTH*85)-1:WIDTH*84];
		d_in85 <= tmp[(WIDTH*86)-1:WIDTH*85];
		d_in86 <= tmp[(WIDTH*87)-1:WIDTH*86];
		d_in87 <= tmp[(WIDTH*88)-1:WIDTH*87];
		d_in88 <= tmp[(WIDTH*89)-1:WIDTH*88];
		d_in89 <= tmp[(WIDTH*90)-1:WIDTH*89];
	end

	design39_90_100 #(.WIDTH(WIDTH)) design39_90_100_inst(.d_in0(d_in0),.d_in1(d_in1),.d_in2(d_in2),.d_in3(d_in3),.d_in4(d_in4),.d_in5(d_in5),.d_in6(d_in6),.d_in7(d_in7),.d_in8(d_in8),.d_in9(d_in9),.d_in10(d_in10),.d_in11(d_in11),.d_in12(d_in12),.d_in13(d_in13),.d_in14(d_in14),.d_in15(d_in15),.d_in16(d_in16),.d_in17(d_in17),.d_in18(d_in18),.d_in19(d_in19),.d_in20(d_in20),.d_in21(d_in21),.d_in22(d_in22),.d_in23(d_in23),.d_in24(d_in24),.d_in25(d_in25),.d_in26(d_in26),.d_in27(d_in27),.d_in28(d_in28),.d_in29(d_in29),.d_in30(d_in30),.d_in31(d_in31),.d_in32(d_in32),.d_in33(d_in33),.d_in34(d_in34),.d_in35(d_in35),.d_in36(d_in36),.d_in37(d_in37),.d_in38(d_in38),.d_in39(d_in39),.d_in40(d_in40),.d_in41(d_in41),.d_in42(d_in42),.d_in43(d_in43),.d_in44(d_in44),.d_in45(d_in45),.d_in46(d_in46),.d_in47(d_in47),.d_in48(d_in48),.d_in49(d_in49),.d_in50(d_in50),.d_in51(d_in51),.d_in52(d_in52),.d_in53(d_in53),.d_in54(d_in54),.d_in55(d_in55),.d_in56(d_in56),.d_in57(d_in57),.d_in58(d_in58),.d_in59(d_in59),.d_in60(d_in60),.d_in61(d_in61),.d_in62(d_in62),.d_in63(d_in63),.d_in64(d_in64),.d_in65(d_in65),.d_in66(d_in66),.d_in67(d_in67),.d_in68(d_in68),.d_in69(d_in69),.d_in70(d_in70),.d_in71(d_in71),.d_in72(d_in72),.d_in73(d_in73),.d_in74(d_in74),.d_in75(d_in75),.d_in76(d_in76),.d_in77(d_in77),.d_in78(d_in78),.d_in79(d_in79),.d_in80(d_in80),.d_in81(d_in81),.d_in82(d_in82),.d_in83(d_in83),.d_in84(d_in84),.d_in85(d_in85),.d_in86(d_in86),.d_in87(d_in87),.d_in88(d_in88),.d_in89(d_in89),.d_out0(d_out0),.d_out1(d_out1),.d_out2(d_out2),.d_out3(d_out3),.d_out4(d_out4),.d_out5(d_out5),.d_out6(d_out6),.d_out7(d_out7),.d_out8(d_out8),.d_out9(d_out9),.d_out10(d_out10),.d_out11(d_out11),.d_out12(d_out12),.d_out13(d_out13),.d_out14(d_out14),.d_out15(d_out15),.d_out16(d_out16),.d_out17(d_out17),.d_out18(d_out18),.d_out19(d_out19),.d_out20(d_out20),.d_out21(d_out21),.d_out22(d_out22),.d_out23(d_out23),.d_out24(d_out24),.d_out25(d_out25),.d_out26(d_out26),.d_out27(d_out27),.d_out28(d_out28),.d_out29(d_out29),.d_out30(d_out30),.d_out31(d_out31),.d_out32(d_out32),.d_out33(d_out33),.d_out34(d_out34),.d_out35(d_out35),.d_out36(d_out36),.d_out37(d_out37),.d_out38(d_out38),.d_out39(d_out39),.d_out40(d_out40),.d_out41(d_out41),.d_out42(d_out42),.d_out43(d_out43),.d_out44(d_out44),.d_out45(d_out45),.d_out46(d_out46),.d_out47(d_out47),.d_out48(d_out48),.d_out49(d_out49),.d_out50(d_out50),.d_out51(d_out51),.d_out52(d_out52),.d_out53(d_out53),.d_out54(d_out54),.d_out55(d_out55),.d_out56(d_out56),.d_out57(d_out57),.d_out58(d_out58),.d_out59(d_out59),.d_out60(d_out60),.d_out61(d_out61),.d_out62(d_out62),.d_out63(d_out63),.d_out64(d_out64),.d_out65(d_out65),.d_out66(d_out66),.d_out67(d_out67),.d_out68(d_out68),.d_out69(d_out69),.d_out70(d_out70),.d_out71(d_out71),.d_out72(d_out72),.d_out73(d_out73),.d_out74(d_out74),.d_out75(d_out75),.d_out76(d_out76),.d_out77(d_out77),.d_out78(d_out78),.d_out79(d_out79),.d_out80(d_out80),.d_out81(d_out81),.d_out82(d_out82),.d_out83(d_out83),.d_out84(d_out84),.d_out85(d_out85),.d_out86(d_out86),.d_out87(d_out87),.d_out88(d_out88),.d_out89(d_out89),.clk(clk),.rst(rst));

	assign out = d_out0^d_out1^d_out2^d_out3^d_out4^d_out5^d_out6^d_out7^d_out8^d_out9^d_out10^d_out11^d_out12^d_out13^d_out14^d_out15^d_out16^d_out17^d_out18^d_out19^d_out20^d_out21^d_out22^d_out23^d_out24^d_out25^d_out26^d_out27^d_out28^d_out29^d_out30^d_out31^d_out32^d_out33^d_out34^d_out35^d_out36^d_out37^d_out38^d_out39^d_out40^d_out41^d_out42^d_out43^d_out44^d_out45^d_out46^d_out47^d_out48^d_out49^d_out50^d_out51^d_out52^d_out53^d_out54^d_out55^d_out56^d_out57^d_out58^d_out59^d_out60^d_out61^d_out62^d_out63^d_out64^d_out65^d_out66^d_out67^d_out68^d_out69^d_out70^d_out71^d_out72^d_out73^d_out74^d_out75^d_out76^d_out77^d_out78^d_out79^d_out80^d_out81^d_out82^d_out83^d_out84^d_out85^d_out86^d_out87^d_out88^d_out89;

endmodule

module design39_90_100 #(parameter WIDTH=32) (d_in0, d_in1, d_in2, d_in3, d_in4, d_in5, d_in6, d_in7, d_in8, d_in9, d_in10, d_in11, d_in12, d_in13, d_in14, d_in15, d_in16, d_in17, d_in18, d_in19, d_in20, d_in21, d_in22, d_in23, d_in24, d_in25, d_in26, d_in27, d_in28, d_in29, d_in30, d_in31, d_in32, d_in33, d_in34, d_in35, d_in36, d_in37, d_in38, d_in39, d_in40, d_in41, d_in42, d_in43, d_in44, d_in45, d_in46, d_in47, d_in48, d_in49, d_in50, d_in51, d_in52, d_in53, d_in54, d_in55, d_in56, d_in57, d_in58, d_in59, d_in60, d_in61, d_in62, d_in63, d_in64, d_in65, d_in66, d_in67, d_in68, d_in69, d_in70, d_in71, d_in72, d_in73, d_in74, d_in75, d_in76, d_in77, d_in78, d_in79, d_in80, d_in81, d_in82, d_in83, d_in84, d_in85, d_in86, d_in87, d_in88, d_in89, d_out0, d_out1, d_out2, d_out3, d_out4, d_out5, d_out6, d_out7, d_out8, d_out9, d_out10, d_out11, d_out12, d_out13, d_out14, d_out15, d_out16, d_out17, d_out18, d_out19, d_out20, d_out21, d_out22, d_out23, d_out24, d_out25, d_out26, d_out27, d_out28, d_out29, d_out30, d_out31, d_out32, d_out33, d_out34, d_out35, d_out36, d_out37, d_out38, d_out39, d_out40, d_out41, d_out42, d_out43, d_out44, d_out45, d_out46, d_out47, d_out48, d_out49, d_out50, d_out51, d_out52, d_out53, d_out54, d_out55, d_out56, d_out57, d_out58, d_out59, d_out60, d_out61, d_out62, d_out63, d_out64, d_out65, d_out66, d_out67, d_out68, d_out69, d_out70, d_out71, d_out72, d_out73, d_out74, d_out75, d_out76, d_out77, d_out78, d_out79, d_out80, d_out81, d_out82, d_out83, d_out84, d_out85, d_out86, d_out87, d_out88, d_out89, clk, rst);
	input clk;
	input rst;
	input [WIDTH-1:0] d_in0; 
	input [WIDTH-1:0] d_in1; 
	input [WIDTH-1:0] d_in2; 
	input [WIDTH-1:0] d_in3; 
	input [WIDTH-1:0] d_in4; 
	input [WIDTH-1:0] d_in5; 
	input [WIDTH-1:0] d_in6; 
	input [WIDTH-1:0] d_in7; 
	input [WIDTH-1:0] d_in8; 
	input [WIDTH-1:0] d_in9; 
	input [WIDTH-1:0] d_in10; 
	input [WIDTH-1:0] d_in11; 
	input [WIDTH-1:0] d_in12; 
	input [WIDTH-1:0] d_in13; 
	input [WIDTH-1:0] d_in14; 
	input [WIDTH-1:0] d_in15; 
	input [WIDTH-1:0] d_in16; 
	input [WIDTH-1:0] d_in17; 
	input [WIDTH-1:0] d_in18; 
	input [WIDTH-1:0] d_in19; 
	input [WIDTH-1:0] d_in20; 
	input [WIDTH-1:0] d_in21; 
	input [WIDTH-1:0] d_in22; 
	input [WIDTH-1:0] d_in23; 
	input [WIDTH-1:0] d_in24; 
	input [WIDTH-1:0] d_in25; 
	input [WIDTH-1:0] d_in26; 
	input [WIDTH-1:0] d_in27; 
	input [WIDTH-1:0] d_in28; 
	input [WIDTH-1:0] d_in29; 
	input [WIDTH-1:0] d_in30; 
	input [WIDTH-1:0] d_in31; 
	input [WIDTH-1:0] d_in32; 
	input [WIDTH-1:0] d_in33; 
	input [WIDTH-1:0] d_in34; 
	input [WIDTH-1:0] d_in35; 
	input [WIDTH-1:0] d_in36; 
	input [WIDTH-1:0] d_in37; 
	input [WIDTH-1:0] d_in38; 
	input [WIDTH-1:0] d_in39; 
	input [WIDTH-1:0] d_in40; 
	input [WIDTH-1:0] d_in41; 
	input [WIDTH-1:0] d_in42; 
	input [WIDTH-1:0] d_in43; 
	input [WIDTH-1:0] d_in44; 
	input [WIDTH-1:0] d_in45; 
	input [WIDTH-1:0] d_in46; 
	input [WIDTH-1:0] d_in47; 
	input [WIDTH-1:0] d_in48; 
	input [WIDTH-1:0] d_in49; 
	input [WIDTH-1:0] d_in50; 
	input [WIDTH-1:0] d_in51; 
	input [WIDTH-1:0] d_in52; 
	input [WIDTH-1:0] d_in53; 
	input [WIDTH-1:0] d_in54; 
	input [WIDTH-1:0] d_in55; 
	input [WIDTH-1:0] d_in56; 
	input [WIDTH-1:0] d_in57; 
	input [WIDTH-1:0] d_in58; 
	input [WIDTH-1:0] d_in59; 
	input [WIDTH-1:0] d_in60; 
	input [WIDTH-1:0] d_in61; 
	input [WIDTH-1:0] d_in62; 
	input [WIDTH-1:0] d_in63; 
	input [WIDTH-1:0] d_in64; 
	input [WIDTH-1:0] d_in65; 
	input [WIDTH-1:0] d_in66; 
	input [WIDTH-1:0] d_in67; 
	input [WIDTH-1:0] d_in68; 
	input [WIDTH-1:0] d_in69; 
	input [WIDTH-1:0] d_in70; 
	input [WIDTH-1:0] d_in71; 
	input [WIDTH-1:0] d_in72; 
	input [WIDTH-1:0] d_in73; 
	input [WIDTH-1:0] d_in74; 
	input [WIDTH-1:0] d_in75; 
	input [WIDTH-1:0] d_in76; 
	input [WIDTH-1:0] d_in77; 
	input [WIDTH-1:0] d_in78; 
	input [WIDTH-1:0] d_in79; 
	input [WIDTH-1:0] d_in80; 
	input [WIDTH-1:0] d_in81; 
	input [WIDTH-1:0] d_in82; 
	input [WIDTH-1:0] d_in83; 
	input [WIDTH-1:0] d_in84; 
	input [WIDTH-1:0] d_in85; 
	input [WIDTH-1:0] d_in86; 
	input [WIDTH-1:0] d_in87; 
	input [WIDTH-1:0] d_in88; 
	input [WIDTH-1:0] d_in89; 
	output [WIDTH-1:0] d_out0; 
	output [WIDTH-1:0] d_out1; 
	output [WIDTH-1:0] d_out2; 
	output [WIDTH-1:0] d_out3; 
	output [WIDTH-1:0] d_out4; 
	output [WIDTH-1:0] d_out5; 
	output [WIDTH-1:0] d_out6; 
	output [WIDTH-1:0] d_out7; 
	output [WIDTH-1:0] d_out8; 
	output [WIDTH-1:0] d_out9; 
	output [WIDTH-1:0] d_out10; 
	output [WIDTH-1:0] d_out11; 
	output [WIDTH-1:0] d_out12; 
	output [WIDTH-1:0] d_out13; 
	output [WIDTH-1:0] d_out14; 
	output [WIDTH-1:0] d_out15; 
	output [WIDTH-1:0] d_out16; 
	output [WIDTH-1:0] d_out17; 
	output [WIDTH-1:0] d_out18; 
	output [WIDTH-1:0] d_out19; 
	output [WIDTH-1:0] d_out20; 
	output [WIDTH-1:0] d_out21; 
	output [WIDTH-1:0] d_out22; 
	output [WIDTH-1:0] d_out23; 
	output [WIDTH-1:0] d_out24; 
	output [WIDTH-1:0] d_out25; 
	output [WIDTH-1:0] d_out26; 
	output [WIDTH-1:0] d_out27; 
	output [WIDTH-1:0] d_out28; 
	output [WIDTH-1:0] d_out29; 
	output [WIDTH-1:0] d_out30; 
	output [WIDTH-1:0] d_out31; 
	output [WIDTH-1:0] d_out32; 
	output [WIDTH-1:0] d_out33; 
	output [WIDTH-1:0] d_out34; 
	output [WIDTH-1:0] d_out35; 
	output [WIDTH-1:0] d_out36; 
	output [WIDTH-1:0] d_out37; 
	output [WIDTH-1:0] d_out38; 
	output [WIDTH-1:0] d_out39; 
	output [WIDTH-1:0] d_out40; 
	output [WIDTH-1:0] d_out41; 
	output [WIDTH-1:0] d_out42; 
	output [WIDTH-1:0] d_out43; 
	output [WIDTH-1:0] d_out44; 
	output [WIDTH-1:0] d_out45; 
	output [WIDTH-1:0] d_out46; 
	output [WIDTH-1:0] d_out47; 
	output [WIDTH-1:0] d_out48; 
	output [WIDTH-1:0] d_out49; 
	output [WIDTH-1:0] d_out50; 
	output [WIDTH-1:0] d_out51; 
	output [WIDTH-1:0] d_out52; 
	output [WIDTH-1:0] d_out53; 
	output [WIDTH-1:0] d_out54; 
	output [WIDTH-1:0] d_out55; 
	output [WIDTH-1:0] d_out56; 
	output [WIDTH-1:0] d_out57; 
	output [WIDTH-1:0] d_out58; 
	output [WIDTH-1:0] d_out59; 
	output [WIDTH-1:0] d_out60; 
	output [WIDTH-1:0] d_out61; 
	output [WIDTH-1:0] d_out62; 
	output [WIDTH-1:0] d_out63; 
	output [WIDTH-1:0] d_out64; 
	output [WIDTH-1:0] d_out65; 
	output [WIDTH-1:0] d_out66; 
	output [WIDTH-1:0] d_out67; 
	output [WIDTH-1:0] d_out68; 
	output [WIDTH-1:0] d_out69; 
	output [WIDTH-1:0] d_out70; 
	output [WIDTH-1:0] d_out71; 
	output [WIDTH-1:0] d_out72; 
	output [WIDTH-1:0] d_out73; 
	output [WIDTH-1:0] d_out74; 
	output [WIDTH-1:0] d_out75; 
	output [WIDTH-1:0] d_out76; 
	output [WIDTH-1:0] d_out77; 
	output [WIDTH-1:0] d_out78; 
	output [WIDTH-1:0] d_out79; 
	output [WIDTH-1:0] d_out80; 
	output [WIDTH-1:0] d_out81; 
	output [WIDTH-1:0] d_out82; 
	output [WIDTH-1:0] d_out83; 
	output [WIDTH-1:0] d_out84; 
	output [WIDTH-1:0] d_out85; 
	output [WIDTH-1:0] d_out86; 
	output [WIDTH-1:0] d_out87; 
	output [WIDTH-1:0] d_out88; 
	output [WIDTH-1:0] d_out89; 

	wire [WIDTH-1:0] wire_d0_0;
	wire [WIDTH-1:0] wire_d0_1;
	wire [WIDTH-1:0] wire_d0_2;
	wire [WIDTH-1:0] wire_d0_3;
	wire [WIDTH-1:0] wire_d0_4;
	wire [WIDTH-1:0] wire_d0_5;
	wire [WIDTH-1:0] wire_d0_6;
	wire [WIDTH-1:0] wire_d0_7;
	wire [WIDTH-1:0] wire_d0_8;
	wire [WIDTH-1:0] wire_d0_9;
	wire [WIDTH-1:0] wire_d0_10;
	wire [WIDTH-1:0] wire_d0_11;
	wire [WIDTH-1:0] wire_d0_12;
	wire [WIDTH-1:0] wire_d0_13;
	wire [WIDTH-1:0] wire_d0_14;
	wire [WIDTH-1:0] wire_d0_15;
	wire [WIDTH-1:0] wire_d0_16;
	wire [WIDTH-1:0] wire_d0_17;
	wire [WIDTH-1:0] wire_d0_18;
	wire [WIDTH-1:0] wire_d0_19;
	wire [WIDTH-1:0] wire_d0_20;
	wire [WIDTH-1:0] wire_d0_21;
	wire [WIDTH-1:0] wire_d0_22;
	wire [WIDTH-1:0] wire_d0_23;
	wire [WIDTH-1:0] wire_d0_24;
	wire [WIDTH-1:0] wire_d0_25;
	wire [WIDTH-1:0] wire_d0_26;
	wire [WIDTH-1:0] wire_d0_27;
	wire [WIDTH-1:0] wire_d0_28;
	wire [WIDTH-1:0] wire_d0_29;
	wire [WIDTH-1:0] wire_d0_30;
	wire [WIDTH-1:0] wire_d0_31;
	wire [WIDTH-1:0] wire_d0_32;
	wire [WIDTH-1:0] wire_d0_33;
	wire [WIDTH-1:0] wire_d0_34;
	wire [WIDTH-1:0] wire_d0_35;
	wire [WIDTH-1:0] wire_d0_36;
	wire [WIDTH-1:0] wire_d0_37;
	wire [WIDTH-1:0] wire_d0_38;
	wire [WIDTH-1:0] wire_d0_39;
	wire [WIDTH-1:0] wire_d0_40;
	wire [WIDTH-1:0] wire_d0_41;
	wire [WIDTH-1:0] wire_d0_42;
	wire [WIDTH-1:0] wire_d0_43;
	wire [WIDTH-1:0] wire_d0_44;
	wire [WIDTH-1:0] wire_d0_45;
	wire [WIDTH-1:0] wire_d0_46;
	wire [WIDTH-1:0] wire_d0_47;
	wire [WIDTH-1:0] wire_d0_48;
	wire [WIDTH-1:0] wire_d0_49;
	wire [WIDTH-1:0] wire_d0_50;
	wire [WIDTH-1:0] wire_d0_51;
	wire [WIDTH-1:0] wire_d0_52;
	wire [WIDTH-1:0] wire_d0_53;
	wire [WIDTH-1:0] wire_d0_54;
	wire [WIDTH-1:0] wire_d0_55;
	wire [WIDTH-1:0] wire_d0_56;
	wire [WIDTH-1:0] wire_d0_57;
	wire [WIDTH-1:0] wire_d0_58;
	wire [WIDTH-1:0] wire_d0_59;
	wire [WIDTH-1:0] wire_d0_60;
	wire [WIDTH-1:0] wire_d0_61;
	wire [WIDTH-1:0] wire_d0_62;
	wire [WIDTH-1:0] wire_d0_63;
	wire [WIDTH-1:0] wire_d0_64;
	wire [WIDTH-1:0] wire_d0_65;
	wire [WIDTH-1:0] wire_d0_66;
	wire [WIDTH-1:0] wire_d0_67;
	wire [WIDTH-1:0] wire_d0_68;
	wire [WIDTH-1:0] wire_d0_69;
	wire [WIDTH-1:0] wire_d0_70;
	wire [WIDTH-1:0] wire_d0_71;
	wire [WIDTH-1:0] wire_d0_72;
	wire [WIDTH-1:0] wire_d0_73;
	wire [WIDTH-1:0] wire_d0_74;
	wire [WIDTH-1:0] wire_d0_75;
	wire [WIDTH-1:0] wire_d0_76;
	wire [WIDTH-1:0] wire_d0_77;
	wire [WIDTH-1:0] wire_d0_78;
	wire [WIDTH-1:0] wire_d0_79;
	wire [WIDTH-1:0] wire_d0_80;
	wire [WIDTH-1:0] wire_d0_81;
	wire [WIDTH-1:0] wire_d0_82;
	wire [WIDTH-1:0] wire_d0_83;
	wire [WIDTH-1:0] wire_d0_84;
	wire [WIDTH-1:0] wire_d0_85;
	wire [WIDTH-1:0] wire_d0_86;
	wire [WIDTH-1:0] wire_d0_87;
	wire [WIDTH-1:0] wire_d0_88;
	wire [WIDTH-1:0] wire_d0_89;
	wire [WIDTH-1:0] wire_d0_90;
	wire [WIDTH-1:0] wire_d0_91;
	wire [WIDTH-1:0] wire_d0_92;
	wire [WIDTH-1:0] wire_d0_93;
	wire [WIDTH-1:0] wire_d0_94;
	wire [WIDTH-1:0] wire_d0_95;
	wire [WIDTH-1:0] wire_d0_96;
	wire [WIDTH-1:0] wire_d0_97;
	wire [WIDTH-1:0] wire_d0_98;
	wire [WIDTH-1:0] wire_d1_0;
	wire [WIDTH-1:0] wire_d1_1;
	wire [WIDTH-1:0] wire_d1_2;
	wire [WIDTH-1:0] wire_d1_3;
	wire [WIDTH-1:0] wire_d1_4;
	wire [WIDTH-1:0] wire_d1_5;
	wire [WIDTH-1:0] wire_d1_6;
	wire [WIDTH-1:0] wire_d1_7;
	wire [WIDTH-1:0] wire_d1_8;
	wire [WIDTH-1:0] wire_d1_9;
	wire [WIDTH-1:0] wire_d1_10;
	wire [WIDTH-1:0] wire_d1_11;
	wire [WIDTH-1:0] wire_d1_12;
	wire [WIDTH-1:0] wire_d1_13;
	wire [WIDTH-1:0] wire_d1_14;
	wire [WIDTH-1:0] wire_d1_15;
	wire [WIDTH-1:0] wire_d1_16;
	wire [WIDTH-1:0] wire_d1_17;
	wire [WIDTH-1:0] wire_d1_18;
	wire [WIDTH-1:0] wire_d1_19;
	wire [WIDTH-1:0] wire_d1_20;
	wire [WIDTH-1:0] wire_d1_21;
	wire [WIDTH-1:0] wire_d1_22;
	wire [WIDTH-1:0] wire_d1_23;
	wire [WIDTH-1:0] wire_d1_24;
	wire [WIDTH-1:0] wire_d1_25;
	wire [WIDTH-1:0] wire_d1_26;
	wire [WIDTH-1:0] wire_d1_27;
	wire [WIDTH-1:0] wire_d1_28;
	wire [WIDTH-1:0] wire_d1_29;
	wire [WIDTH-1:0] wire_d1_30;
	wire [WIDTH-1:0] wire_d1_31;
	wire [WIDTH-1:0] wire_d1_32;
	wire [WIDTH-1:0] wire_d1_33;
	wire [WIDTH-1:0] wire_d1_34;
	wire [WIDTH-1:0] wire_d1_35;
	wire [WIDTH-1:0] wire_d1_36;
	wire [WIDTH-1:0] wire_d1_37;
	wire [WIDTH-1:0] wire_d1_38;
	wire [WIDTH-1:0] wire_d1_39;
	wire [WIDTH-1:0] wire_d1_40;
	wire [WIDTH-1:0] wire_d1_41;
	wire [WIDTH-1:0] wire_d1_42;
	wire [WIDTH-1:0] wire_d1_43;
	wire [WIDTH-1:0] wire_d1_44;
	wire [WIDTH-1:0] wire_d1_45;
	wire [WIDTH-1:0] wire_d1_46;
	wire [WIDTH-1:0] wire_d1_47;
	wire [WIDTH-1:0] wire_d1_48;
	wire [WIDTH-1:0] wire_d1_49;
	wire [WIDTH-1:0] wire_d1_50;
	wire [WIDTH-1:0] wire_d1_51;
	wire [WIDTH-1:0] wire_d1_52;
	wire [WIDTH-1:0] wire_d1_53;
	wire [WIDTH-1:0] wire_d1_54;
	wire [WIDTH-1:0] wire_d1_55;
	wire [WIDTH-1:0] wire_d1_56;
	wire [WIDTH-1:0] wire_d1_57;
	wire [WIDTH-1:0] wire_d1_58;
	wire [WIDTH-1:0] wire_d1_59;
	wire [WIDTH-1:0] wire_d1_60;
	wire [WIDTH-1:0] wire_d1_61;
	wire [WIDTH-1:0] wire_d1_62;
	wire [WIDTH-1:0] wire_d1_63;
	wire [WIDTH-1:0] wire_d1_64;
	wire [WIDTH-1:0] wire_d1_65;
	wire [WIDTH-1:0] wire_d1_66;
	wire [WIDTH-1:0] wire_d1_67;
	wire [WIDTH-1:0] wire_d1_68;
	wire [WIDTH-1:0] wire_d1_69;
	wire [WIDTH-1:0] wire_d1_70;
	wire [WIDTH-1:0] wire_d1_71;
	wire [WIDTH-1:0] wire_d1_72;
	wire [WIDTH-1:0] wire_d1_73;
	wire [WIDTH-1:0] wire_d1_74;
	wire [WIDTH-1:0] wire_d1_75;
	wire [WIDTH-1:0] wire_d1_76;
	wire [WIDTH-1:0] wire_d1_77;
	wire [WIDTH-1:0] wire_d1_78;
	wire [WIDTH-1:0] wire_d1_79;
	wire [WIDTH-1:0] wire_d1_80;
	wire [WIDTH-1:0] wire_d1_81;
	wire [WIDTH-1:0] wire_d1_82;
	wire [WIDTH-1:0] wire_d1_83;
	wire [WIDTH-1:0] wire_d1_84;
	wire [WIDTH-1:0] wire_d1_85;
	wire [WIDTH-1:0] wire_d1_86;
	wire [WIDTH-1:0] wire_d1_87;
	wire [WIDTH-1:0] wire_d1_88;
	wire [WIDTH-1:0] wire_d1_89;
	wire [WIDTH-1:0] wire_d1_90;
	wire [WIDTH-1:0] wire_d1_91;
	wire [WIDTH-1:0] wire_d1_92;
	wire [WIDTH-1:0] wire_d1_93;
	wire [WIDTH-1:0] wire_d1_94;
	wire [WIDTH-1:0] wire_d1_95;
	wire [WIDTH-1:0] wire_d1_96;
	wire [WIDTH-1:0] wire_d1_97;
	wire [WIDTH-1:0] wire_d1_98;
	wire [WIDTH-1:0] wire_d2_0;
	wire [WIDTH-1:0] wire_d2_1;
	wire [WIDTH-1:0] wire_d2_2;
	wire [WIDTH-1:0] wire_d2_3;
	wire [WIDTH-1:0] wire_d2_4;
	wire [WIDTH-1:0] wire_d2_5;
	wire [WIDTH-1:0] wire_d2_6;
	wire [WIDTH-1:0] wire_d2_7;
	wire [WIDTH-1:0] wire_d2_8;
	wire [WIDTH-1:0] wire_d2_9;
	wire [WIDTH-1:0] wire_d2_10;
	wire [WIDTH-1:0] wire_d2_11;
	wire [WIDTH-1:0] wire_d2_12;
	wire [WIDTH-1:0] wire_d2_13;
	wire [WIDTH-1:0] wire_d2_14;
	wire [WIDTH-1:0] wire_d2_15;
	wire [WIDTH-1:0] wire_d2_16;
	wire [WIDTH-1:0] wire_d2_17;
	wire [WIDTH-1:0] wire_d2_18;
	wire [WIDTH-1:0] wire_d2_19;
	wire [WIDTH-1:0] wire_d2_20;
	wire [WIDTH-1:0] wire_d2_21;
	wire [WIDTH-1:0] wire_d2_22;
	wire [WIDTH-1:0] wire_d2_23;
	wire [WIDTH-1:0] wire_d2_24;
	wire [WIDTH-1:0] wire_d2_25;
	wire [WIDTH-1:0] wire_d2_26;
	wire [WIDTH-1:0] wire_d2_27;
	wire [WIDTH-1:0] wire_d2_28;
	wire [WIDTH-1:0] wire_d2_29;
	wire [WIDTH-1:0] wire_d2_30;
	wire [WIDTH-1:0] wire_d2_31;
	wire [WIDTH-1:0] wire_d2_32;
	wire [WIDTH-1:0] wire_d2_33;
	wire [WIDTH-1:0] wire_d2_34;
	wire [WIDTH-1:0] wire_d2_35;
	wire [WIDTH-1:0] wire_d2_36;
	wire [WIDTH-1:0] wire_d2_37;
	wire [WIDTH-1:0] wire_d2_38;
	wire [WIDTH-1:0] wire_d2_39;
	wire [WIDTH-1:0] wire_d2_40;
	wire [WIDTH-1:0] wire_d2_41;
	wire [WIDTH-1:0] wire_d2_42;
	wire [WIDTH-1:0] wire_d2_43;
	wire [WIDTH-1:0] wire_d2_44;
	wire [WIDTH-1:0] wire_d2_45;
	wire [WIDTH-1:0] wire_d2_46;
	wire [WIDTH-1:0] wire_d2_47;
	wire [WIDTH-1:0] wire_d2_48;
	wire [WIDTH-1:0] wire_d2_49;
	wire [WIDTH-1:0] wire_d2_50;
	wire [WIDTH-1:0] wire_d2_51;
	wire [WIDTH-1:0] wire_d2_52;
	wire [WIDTH-1:0] wire_d2_53;
	wire [WIDTH-1:0] wire_d2_54;
	wire [WIDTH-1:0] wire_d2_55;
	wire [WIDTH-1:0] wire_d2_56;
	wire [WIDTH-1:0] wire_d2_57;
	wire [WIDTH-1:0] wire_d2_58;
	wire [WIDTH-1:0] wire_d2_59;
	wire [WIDTH-1:0] wire_d2_60;
	wire [WIDTH-1:0] wire_d2_61;
	wire [WIDTH-1:0] wire_d2_62;
	wire [WIDTH-1:0] wire_d2_63;
	wire [WIDTH-1:0] wire_d2_64;
	wire [WIDTH-1:0] wire_d2_65;
	wire [WIDTH-1:0] wire_d2_66;
	wire [WIDTH-1:0] wire_d2_67;
	wire [WIDTH-1:0] wire_d2_68;
	wire [WIDTH-1:0] wire_d2_69;
	wire [WIDTH-1:0] wire_d2_70;
	wire [WIDTH-1:0] wire_d2_71;
	wire [WIDTH-1:0] wire_d2_72;
	wire [WIDTH-1:0] wire_d2_73;
	wire [WIDTH-1:0] wire_d2_74;
	wire [WIDTH-1:0] wire_d2_75;
	wire [WIDTH-1:0] wire_d2_76;
	wire [WIDTH-1:0] wire_d2_77;
	wire [WIDTH-1:0] wire_d2_78;
	wire [WIDTH-1:0] wire_d2_79;
	wire [WIDTH-1:0] wire_d2_80;
	wire [WIDTH-1:0] wire_d2_81;
	wire [WIDTH-1:0] wire_d2_82;
	wire [WIDTH-1:0] wire_d2_83;
	wire [WIDTH-1:0] wire_d2_84;
	wire [WIDTH-1:0] wire_d2_85;
	wire [WIDTH-1:0] wire_d2_86;
	wire [WIDTH-1:0] wire_d2_87;
	wire [WIDTH-1:0] wire_d2_88;
	wire [WIDTH-1:0] wire_d2_89;
	wire [WIDTH-1:0] wire_d2_90;
	wire [WIDTH-1:0] wire_d2_91;
	wire [WIDTH-1:0] wire_d2_92;
	wire [WIDTH-1:0] wire_d2_93;
	wire [WIDTH-1:0] wire_d2_94;
	wire [WIDTH-1:0] wire_d2_95;
	wire [WIDTH-1:0] wire_d2_96;
	wire [WIDTH-1:0] wire_d2_97;
	wire [WIDTH-1:0] wire_d2_98;
	wire [WIDTH-1:0] wire_d3_0;
	wire [WIDTH-1:0] wire_d3_1;
	wire [WIDTH-1:0] wire_d3_2;
	wire [WIDTH-1:0] wire_d3_3;
	wire [WIDTH-1:0] wire_d3_4;
	wire [WIDTH-1:0] wire_d3_5;
	wire [WIDTH-1:0] wire_d3_6;
	wire [WIDTH-1:0] wire_d3_7;
	wire [WIDTH-1:0] wire_d3_8;
	wire [WIDTH-1:0] wire_d3_9;
	wire [WIDTH-1:0] wire_d3_10;
	wire [WIDTH-1:0] wire_d3_11;
	wire [WIDTH-1:0] wire_d3_12;
	wire [WIDTH-1:0] wire_d3_13;
	wire [WIDTH-1:0] wire_d3_14;
	wire [WIDTH-1:0] wire_d3_15;
	wire [WIDTH-1:0] wire_d3_16;
	wire [WIDTH-1:0] wire_d3_17;
	wire [WIDTH-1:0] wire_d3_18;
	wire [WIDTH-1:0] wire_d3_19;
	wire [WIDTH-1:0] wire_d3_20;
	wire [WIDTH-1:0] wire_d3_21;
	wire [WIDTH-1:0] wire_d3_22;
	wire [WIDTH-1:0] wire_d3_23;
	wire [WIDTH-1:0] wire_d3_24;
	wire [WIDTH-1:0] wire_d3_25;
	wire [WIDTH-1:0] wire_d3_26;
	wire [WIDTH-1:0] wire_d3_27;
	wire [WIDTH-1:0] wire_d3_28;
	wire [WIDTH-1:0] wire_d3_29;
	wire [WIDTH-1:0] wire_d3_30;
	wire [WIDTH-1:0] wire_d3_31;
	wire [WIDTH-1:0] wire_d3_32;
	wire [WIDTH-1:0] wire_d3_33;
	wire [WIDTH-1:0] wire_d3_34;
	wire [WIDTH-1:0] wire_d3_35;
	wire [WIDTH-1:0] wire_d3_36;
	wire [WIDTH-1:0] wire_d3_37;
	wire [WIDTH-1:0] wire_d3_38;
	wire [WIDTH-1:0] wire_d3_39;
	wire [WIDTH-1:0] wire_d3_40;
	wire [WIDTH-1:0] wire_d3_41;
	wire [WIDTH-1:0] wire_d3_42;
	wire [WIDTH-1:0] wire_d3_43;
	wire [WIDTH-1:0] wire_d3_44;
	wire [WIDTH-1:0] wire_d3_45;
	wire [WIDTH-1:0] wire_d3_46;
	wire [WIDTH-1:0] wire_d3_47;
	wire [WIDTH-1:0] wire_d3_48;
	wire [WIDTH-1:0] wire_d3_49;
	wire [WIDTH-1:0] wire_d3_50;
	wire [WIDTH-1:0] wire_d3_51;
	wire [WIDTH-1:0] wire_d3_52;
	wire [WIDTH-1:0] wire_d3_53;
	wire [WIDTH-1:0] wire_d3_54;
	wire [WIDTH-1:0] wire_d3_55;
	wire [WIDTH-1:0] wire_d3_56;
	wire [WIDTH-1:0] wire_d3_57;
	wire [WIDTH-1:0] wire_d3_58;
	wire [WIDTH-1:0] wire_d3_59;
	wire [WIDTH-1:0] wire_d3_60;
	wire [WIDTH-1:0] wire_d3_61;
	wire [WIDTH-1:0] wire_d3_62;
	wire [WIDTH-1:0] wire_d3_63;
	wire [WIDTH-1:0] wire_d3_64;
	wire [WIDTH-1:0] wire_d3_65;
	wire [WIDTH-1:0] wire_d3_66;
	wire [WIDTH-1:0] wire_d3_67;
	wire [WIDTH-1:0] wire_d3_68;
	wire [WIDTH-1:0] wire_d3_69;
	wire [WIDTH-1:0] wire_d3_70;
	wire [WIDTH-1:0] wire_d3_71;
	wire [WIDTH-1:0] wire_d3_72;
	wire [WIDTH-1:0] wire_d3_73;
	wire [WIDTH-1:0] wire_d3_74;
	wire [WIDTH-1:0] wire_d3_75;
	wire [WIDTH-1:0] wire_d3_76;
	wire [WIDTH-1:0] wire_d3_77;
	wire [WIDTH-1:0] wire_d3_78;
	wire [WIDTH-1:0] wire_d3_79;
	wire [WIDTH-1:0] wire_d3_80;
	wire [WIDTH-1:0] wire_d3_81;
	wire [WIDTH-1:0] wire_d3_82;
	wire [WIDTH-1:0] wire_d3_83;
	wire [WIDTH-1:0] wire_d3_84;
	wire [WIDTH-1:0] wire_d3_85;
	wire [WIDTH-1:0] wire_d3_86;
	wire [WIDTH-1:0] wire_d3_87;
	wire [WIDTH-1:0] wire_d3_88;
	wire [WIDTH-1:0] wire_d3_89;
	wire [WIDTH-1:0] wire_d3_90;
	wire [WIDTH-1:0] wire_d3_91;
	wire [WIDTH-1:0] wire_d3_92;
	wire [WIDTH-1:0] wire_d3_93;
	wire [WIDTH-1:0] wire_d3_94;
	wire [WIDTH-1:0] wire_d3_95;
	wire [WIDTH-1:0] wire_d3_96;
	wire [WIDTH-1:0] wire_d3_97;
	wire [WIDTH-1:0] wire_d3_98;
	wire [WIDTH-1:0] wire_d4_0;
	wire [WIDTH-1:0] wire_d4_1;
	wire [WIDTH-1:0] wire_d4_2;
	wire [WIDTH-1:0] wire_d4_3;
	wire [WIDTH-1:0] wire_d4_4;
	wire [WIDTH-1:0] wire_d4_5;
	wire [WIDTH-1:0] wire_d4_6;
	wire [WIDTH-1:0] wire_d4_7;
	wire [WIDTH-1:0] wire_d4_8;
	wire [WIDTH-1:0] wire_d4_9;
	wire [WIDTH-1:0] wire_d4_10;
	wire [WIDTH-1:0] wire_d4_11;
	wire [WIDTH-1:0] wire_d4_12;
	wire [WIDTH-1:0] wire_d4_13;
	wire [WIDTH-1:0] wire_d4_14;
	wire [WIDTH-1:0] wire_d4_15;
	wire [WIDTH-1:0] wire_d4_16;
	wire [WIDTH-1:0] wire_d4_17;
	wire [WIDTH-1:0] wire_d4_18;
	wire [WIDTH-1:0] wire_d4_19;
	wire [WIDTH-1:0] wire_d4_20;
	wire [WIDTH-1:0] wire_d4_21;
	wire [WIDTH-1:0] wire_d4_22;
	wire [WIDTH-1:0] wire_d4_23;
	wire [WIDTH-1:0] wire_d4_24;
	wire [WIDTH-1:0] wire_d4_25;
	wire [WIDTH-1:0] wire_d4_26;
	wire [WIDTH-1:0] wire_d4_27;
	wire [WIDTH-1:0] wire_d4_28;
	wire [WIDTH-1:0] wire_d4_29;
	wire [WIDTH-1:0] wire_d4_30;
	wire [WIDTH-1:0] wire_d4_31;
	wire [WIDTH-1:0] wire_d4_32;
	wire [WIDTH-1:0] wire_d4_33;
	wire [WIDTH-1:0] wire_d4_34;
	wire [WIDTH-1:0] wire_d4_35;
	wire [WIDTH-1:0] wire_d4_36;
	wire [WIDTH-1:0] wire_d4_37;
	wire [WIDTH-1:0] wire_d4_38;
	wire [WIDTH-1:0] wire_d4_39;
	wire [WIDTH-1:0] wire_d4_40;
	wire [WIDTH-1:0] wire_d4_41;
	wire [WIDTH-1:0] wire_d4_42;
	wire [WIDTH-1:0] wire_d4_43;
	wire [WIDTH-1:0] wire_d4_44;
	wire [WIDTH-1:0] wire_d4_45;
	wire [WIDTH-1:0] wire_d4_46;
	wire [WIDTH-1:0] wire_d4_47;
	wire [WIDTH-1:0] wire_d4_48;
	wire [WIDTH-1:0] wire_d4_49;
	wire [WIDTH-1:0] wire_d4_50;
	wire [WIDTH-1:0] wire_d4_51;
	wire [WIDTH-1:0] wire_d4_52;
	wire [WIDTH-1:0] wire_d4_53;
	wire [WIDTH-1:0] wire_d4_54;
	wire [WIDTH-1:0] wire_d4_55;
	wire [WIDTH-1:0] wire_d4_56;
	wire [WIDTH-1:0] wire_d4_57;
	wire [WIDTH-1:0] wire_d4_58;
	wire [WIDTH-1:0] wire_d4_59;
	wire [WIDTH-1:0] wire_d4_60;
	wire [WIDTH-1:0] wire_d4_61;
	wire [WIDTH-1:0] wire_d4_62;
	wire [WIDTH-1:0] wire_d4_63;
	wire [WIDTH-1:0] wire_d4_64;
	wire [WIDTH-1:0] wire_d4_65;
	wire [WIDTH-1:0] wire_d4_66;
	wire [WIDTH-1:0] wire_d4_67;
	wire [WIDTH-1:0] wire_d4_68;
	wire [WIDTH-1:0] wire_d4_69;
	wire [WIDTH-1:0] wire_d4_70;
	wire [WIDTH-1:0] wire_d4_71;
	wire [WIDTH-1:0] wire_d4_72;
	wire [WIDTH-1:0] wire_d4_73;
	wire [WIDTH-1:0] wire_d4_74;
	wire [WIDTH-1:0] wire_d4_75;
	wire [WIDTH-1:0] wire_d4_76;
	wire [WIDTH-1:0] wire_d4_77;
	wire [WIDTH-1:0] wire_d4_78;
	wire [WIDTH-1:0] wire_d4_79;
	wire [WIDTH-1:0] wire_d4_80;
	wire [WIDTH-1:0] wire_d4_81;
	wire [WIDTH-1:0] wire_d4_82;
	wire [WIDTH-1:0] wire_d4_83;
	wire [WIDTH-1:0] wire_d4_84;
	wire [WIDTH-1:0] wire_d4_85;
	wire [WIDTH-1:0] wire_d4_86;
	wire [WIDTH-1:0] wire_d4_87;
	wire [WIDTH-1:0] wire_d4_88;
	wire [WIDTH-1:0] wire_d4_89;
	wire [WIDTH-1:0] wire_d4_90;
	wire [WIDTH-1:0] wire_d4_91;
	wire [WIDTH-1:0] wire_d4_92;
	wire [WIDTH-1:0] wire_d4_93;
	wire [WIDTH-1:0] wire_d4_94;
	wire [WIDTH-1:0] wire_d4_95;
	wire [WIDTH-1:0] wire_d4_96;
	wire [WIDTH-1:0] wire_d4_97;
	wire [WIDTH-1:0] wire_d4_98;
	wire [WIDTH-1:0] wire_d5_0;
	wire [WIDTH-1:0] wire_d5_1;
	wire [WIDTH-1:0] wire_d5_2;
	wire [WIDTH-1:0] wire_d5_3;
	wire [WIDTH-1:0] wire_d5_4;
	wire [WIDTH-1:0] wire_d5_5;
	wire [WIDTH-1:0] wire_d5_6;
	wire [WIDTH-1:0] wire_d5_7;
	wire [WIDTH-1:0] wire_d5_8;
	wire [WIDTH-1:0] wire_d5_9;
	wire [WIDTH-1:0] wire_d5_10;
	wire [WIDTH-1:0] wire_d5_11;
	wire [WIDTH-1:0] wire_d5_12;
	wire [WIDTH-1:0] wire_d5_13;
	wire [WIDTH-1:0] wire_d5_14;
	wire [WIDTH-1:0] wire_d5_15;
	wire [WIDTH-1:0] wire_d5_16;
	wire [WIDTH-1:0] wire_d5_17;
	wire [WIDTH-1:0] wire_d5_18;
	wire [WIDTH-1:0] wire_d5_19;
	wire [WIDTH-1:0] wire_d5_20;
	wire [WIDTH-1:0] wire_d5_21;
	wire [WIDTH-1:0] wire_d5_22;
	wire [WIDTH-1:0] wire_d5_23;
	wire [WIDTH-1:0] wire_d5_24;
	wire [WIDTH-1:0] wire_d5_25;
	wire [WIDTH-1:0] wire_d5_26;
	wire [WIDTH-1:0] wire_d5_27;
	wire [WIDTH-1:0] wire_d5_28;
	wire [WIDTH-1:0] wire_d5_29;
	wire [WIDTH-1:0] wire_d5_30;
	wire [WIDTH-1:0] wire_d5_31;
	wire [WIDTH-1:0] wire_d5_32;
	wire [WIDTH-1:0] wire_d5_33;
	wire [WIDTH-1:0] wire_d5_34;
	wire [WIDTH-1:0] wire_d5_35;
	wire [WIDTH-1:0] wire_d5_36;
	wire [WIDTH-1:0] wire_d5_37;
	wire [WIDTH-1:0] wire_d5_38;
	wire [WIDTH-1:0] wire_d5_39;
	wire [WIDTH-1:0] wire_d5_40;
	wire [WIDTH-1:0] wire_d5_41;
	wire [WIDTH-1:0] wire_d5_42;
	wire [WIDTH-1:0] wire_d5_43;
	wire [WIDTH-1:0] wire_d5_44;
	wire [WIDTH-1:0] wire_d5_45;
	wire [WIDTH-1:0] wire_d5_46;
	wire [WIDTH-1:0] wire_d5_47;
	wire [WIDTH-1:0] wire_d5_48;
	wire [WIDTH-1:0] wire_d5_49;
	wire [WIDTH-1:0] wire_d5_50;
	wire [WIDTH-1:0] wire_d5_51;
	wire [WIDTH-1:0] wire_d5_52;
	wire [WIDTH-1:0] wire_d5_53;
	wire [WIDTH-1:0] wire_d5_54;
	wire [WIDTH-1:0] wire_d5_55;
	wire [WIDTH-1:0] wire_d5_56;
	wire [WIDTH-1:0] wire_d5_57;
	wire [WIDTH-1:0] wire_d5_58;
	wire [WIDTH-1:0] wire_d5_59;
	wire [WIDTH-1:0] wire_d5_60;
	wire [WIDTH-1:0] wire_d5_61;
	wire [WIDTH-1:0] wire_d5_62;
	wire [WIDTH-1:0] wire_d5_63;
	wire [WIDTH-1:0] wire_d5_64;
	wire [WIDTH-1:0] wire_d5_65;
	wire [WIDTH-1:0] wire_d5_66;
	wire [WIDTH-1:0] wire_d5_67;
	wire [WIDTH-1:0] wire_d5_68;
	wire [WIDTH-1:0] wire_d5_69;
	wire [WIDTH-1:0] wire_d5_70;
	wire [WIDTH-1:0] wire_d5_71;
	wire [WIDTH-1:0] wire_d5_72;
	wire [WIDTH-1:0] wire_d5_73;
	wire [WIDTH-1:0] wire_d5_74;
	wire [WIDTH-1:0] wire_d5_75;
	wire [WIDTH-1:0] wire_d5_76;
	wire [WIDTH-1:0] wire_d5_77;
	wire [WIDTH-1:0] wire_d5_78;
	wire [WIDTH-1:0] wire_d5_79;
	wire [WIDTH-1:0] wire_d5_80;
	wire [WIDTH-1:0] wire_d5_81;
	wire [WIDTH-1:0] wire_d5_82;
	wire [WIDTH-1:0] wire_d5_83;
	wire [WIDTH-1:0] wire_d5_84;
	wire [WIDTH-1:0] wire_d5_85;
	wire [WIDTH-1:0] wire_d5_86;
	wire [WIDTH-1:0] wire_d5_87;
	wire [WIDTH-1:0] wire_d5_88;
	wire [WIDTH-1:0] wire_d5_89;
	wire [WIDTH-1:0] wire_d5_90;
	wire [WIDTH-1:0] wire_d5_91;
	wire [WIDTH-1:0] wire_d5_92;
	wire [WIDTH-1:0] wire_d5_93;
	wire [WIDTH-1:0] wire_d5_94;
	wire [WIDTH-1:0] wire_d5_95;
	wire [WIDTH-1:0] wire_d5_96;
	wire [WIDTH-1:0] wire_d5_97;
	wire [WIDTH-1:0] wire_d5_98;
	wire [WIDTH-1:0] wire_d6_0;
	wire [WIDTH-1:0] wire_d6_1;
	wire [WIDTH-1:0] wire_d6_2;
	wire [WIDTH-1:0] wire_d6_3;
	wire [WIDTH-1:0] wire_d6_4;
	wire [WIDTH-1:0] wire_d6_5;
	wire [WIDTH-1:0] wire_d6_6;
	wire [WIDTH-1:0] wire_d6_7;
	wire [WIDTH-1:0] wire_d6_8;
	wire [WIDTH-1:0] wire_d6_9;
	wire [WIDTH-1:0] wire_d6_10;
	wire [WIDTH-1:0] wire_d6_11;
	wire [WIDTH-1:0] wire_d6_12;
	wire [WIDTH-1:0] wire_d6_13;
	wire [WIDTH-1:0] wire_d6_14;
	wire [WIDTH-1:0] wire_d6_15;
	wire [WIDTH-1:0] wire_d6_16;
	wire [WIDTH-1:0] wire_d6_17;
	wire [WIDTH-1:0] wire_d6_18;
	wire [WIDTH-1:0] wire_d6_19;
	wire [WIDTH-1:0] wire_d6_20;
	wire [WIDTH-1:0] wire_d6_21;
	wire [WIDTH-1:0] wire_d6_22;
	wire [WIDTH-1:0] wire_d6_23;
	wire [WIDTH-1:0] wire_d6_24;
	wire [WIDTH-1:0] wire_d6_25;
	wire [WIDTH-1:0] wire_d6_26;
	wire [WIDTH-1:0] wire_d6_27;
	wire [WIDTH-1:0] wire_d6_28;
	wire [WIDTH-1:0] wire_d6_29;
	wire [WIDTH-1:0] wire_d6_30;
	wire [WIDTH-1:0] wire_d6_31;
	wire [WIDTH-1:0] wire_d6_32;
	wire [WIDTH-1:0] wire_d6_33;
	wire [WIDTH-1:0] wire_d6_34;
	wire [WIDTH-1:0] wire_d6_35;
	wire [WIDTH-1:0] wire_d6_36;
	wire [WIDTH-1:0] wire_d6_37;
	wire [WIDTH-1:0] wire_d6_38;
	wire [WIDTH-1:0] wire_d6_39;
	wire [WIDTH-1:0] wire_d6_40;
	wire [WIDTH-1:0] wire_d6_41;
	wire [WIDTH-1:0] wire_d6_42;
	wire [WIDTH-1:0] wire_d6_43;
	wire [WIDTH-1:0] wire_d6_44;
	wire [WIDTH-1:0] wire_d6_45;
	wire [WIDTH-1:0] wire_d6_46;
	wire [WIDTH-1:0] wire_d6_47;
	wire [WIDTH-1:0] wire_d6_48;
	wire [WIDTH-1:0] wire_d6_49;
	wire [WIDTH-1:0] wire_d6_50;
	wire [WIDTH-1:0] wire_d6_51;
	wire [WIDTH-1:0] wire_d6_52;
	wire [WIDTH-1:0] wire_d6_53;
	wire [WIDTH-1:0] wire_d6_54;
	wire [WIDTH-1:0] wire_d6_55;
	wire [WIDTH-1:0] wire_d6_56;
	wire [WIDTH-1:0] wire_d6_57;
	wire [WIDTH-1:0] wire_d6_58;
	wire [WIDTH-1:0] wire_d6_59;
	wire [WIDTH-1:0] wire_d6_60;
	wire [WIDTH-1:0] wire_d6_61;
	wire [WIDTH-1:0] wire_d6_62;
	wire [WIDTH-1:0] wire_d6_63;
	wire [WIDTH-1:0] wire_d6_64;
	wire [WIDTH-1:0] wire_d6_65;
	wire [WIDTH-1:0] wire_d6_66;
	wire [WIDTH-1:0] wire_d6_67;
	wire [WIDTH-1:0] wire_d6_68;
	wire [WIDTH-1:0] wire_d6_69;
	wire [WIDTH-1:0] wire_d6_70;
	wire [WIDTH-1:0] wire_d6_71;
	wire [WIDTH-1:0] wire_d6_72;
	wire [WIDTH-1:0] wire_d6_73;
	wire [WIDTH-1:0] wire_d6_74;
	wire [WIDTH-1:0] wire_d6_75;
	wire [WIDTH-1:0] wire_d6_76;
	wire [WIDTH-1:0] wire_d6_77;
	wire [WIDTH-1:0] wire_d6_78;
	wire [WIDTH-1:0] wire_d6_79;
	wire [WIDTH-1:0] wire_d6_80;
	wire [WIDTH-1:0] wire_d6_81;
	wire [WIDTH-1:0] wire_d6_82;
	wire [WIDTH-1:0] wire_d6_83;
	wire [WIDTH-1:0] wire_d6_84;
	wire [WIDTH-1:0] wire_d6_85;
	wire [WIDTH-1:0] wire_d6_86;
	wire [WIDTH-1:0] wire_d6_87;
	wire [WIDTH-1:0] wire_d6_88;
	wire [WIDTH-1:0] wire_d6_89;
	wire [WIDTH-1:0] wire_d6_90;
	wire [WIDTH-1:0] wire_d6_91;
	wire [WIDTH-1:0] wire_d6_92;
	wire [WIDTH-1:0] wire_d6_93;
	wire [WIDTH-1:0] wire_d6_94;
	wire [WIDTH-1:0] wire_d6_95;
	wire [WIDTH-1:0] wire_d6_96;
	wire [WIDTH-1:0] wire_d6_97;
	wire [WIDTH-1:0] wire_d6_98;
	wire [WIDTH-1:0] wire_d7_0;
	wire [WIDTH-1:0] wire_d7_1;
	wire [WIDTH-1:0] wire_d7_2;
	wire [WIDTH-1:0] wire_d7_3;
	wire [WIDTH-1:0] wire_d7_4;
	wire [WIDTH-1:0] wire_d7_5;
	wire [WIDTH-1:0] wire_d7_6;
	wire [WIDTH-1:0] wire_d7_7;
	wire [WIDTH-1:0] wire_d7_8;
	wire [WIDTH-1:0] wire_d7_9;
	wire [WIDTH-1:0] wire_d7_10;
	wire [WIDTH-1:0] wire_d7_11;
	wire [WIDTH-1:0] wire_d7_12;
	wire [WIDTH-1:0] wire_d7_13;
	wire [WIDTH-1:0] wire_d7_14;
	wire [WIDTH-1:0] wire_d7_15;
	wire [WIDTH-1:0] wire_d7_16;
	wire [WIDTH-1:0] wire_d7_17;
	wire [WIDTH-1:0] wire_d7_18;
	wire [WIDTH-1:0] wire_d7_19;
	wire [WIDTH-1:0] wire_d7_20;
	wire [WIDTH-1:0] wire_d7_21;
	wire [WIDTH-1:0] wire_d7_22;
	wire [WIDTH-1:0] wire_d7_23;
	wire [WIDTH-1:0] wire_d7_24;
	wire [WIDTH-1:0] wire_d7_25;
	wire [WIDTH-1:0] wire_d7_26;
	wire [WIDTH-1:0] wire_d7_27;
	wire [WIDTH-1:0] wire_d7_28;
	wire [WIDTH-1:0] wire_d7_29;
	wire [WIDTH-1:0] wire_d7_30;
	wire [WIDTH-1:0] wire_d7_31;
	wire [WIDTH-1:0] wire_d7_32;
	wire [WIDTH-1:0] wire_d7_33;
	wire [WIDTH-1:0] wire_d7_34;
	wire [WIDTH-1:0] wire_d7_35;
	wire [WIDTH-1:0] wire_d7_36;
	wire [WIDTH-1:0] wire_d7_37;
	wire [WIDTH-1:0] wire_d7_38;
	wire [WIDTH-1:0] wire_d7_39;
	wire [WIDTH-1:0] wire_d7_40;
	wire [WIDTH-1:0] wire_d7_41;
	wire [WIDTH-1:0] wire_d7_42;
	wire [WIDTH-1:0] wire_d7_43;
	wire [WIDTH-1:0] wire_d7_44;
	wire [WIDTH-1:0] wire_d7_45;
	wire [WIDTH-1:0] wire_d7_46;
	wire [WIDTH-1:0] wire_d7_47;
	wire [WIDTH-1:0] wire_d7_48;
	wire [WIDTH-1:0] wire_d7_49;
	wire [WIDTH-1:0] wire_d7_50;
	wire [WIDTH-1:0] wire_d7_51;
	wire [WIDTH-1:0] wire_d7_52;
	wire [WIDTH-1:0] wire_d7_53;
	wire [WIDTH-1:0] wire_d7_54;
	wire [WIDTH-1:0] wire_d7_55;
	wire [WIDTH-1:0] wire_d7_56;
	wire [WIDTH-1:0] wire_d7_57;
	wire [WIDTH-1:0] wire_d7_58;
	wire [WIDTH-1:0] wire_d7_59;
	wire [WIDTH-1:0] wire_d7_60;
	wire [WIDTH-1:0] wire_d7_61;
	wire [WIDTH-1:0] wire_d7_62;
	wire [WIDTH-1:0] wire_d7_63;
	wire [WIDTH-1:0] wire_d7_64;
	wire [WIDTH-1:0] wire_d7_65;
	wire [WIDTH-1:0] wire_d7_66;
	wire [WIDTH-1:0] wire_d7_67;
	wire [WIDTH-1:0] wire_d7_68;
	wire [WIDTH-1:0] wire_d7_69;
	wire [WIDTH-1:0] wire_d7_70;
	wire [WIDTH-1:0] wire_d7_71;
	wire [WIDTH-1:0] wire_d7_72;
	wire [WIDTH-1:0] wire_d7_73;
	wire [WIDTH-1:0] wire_d7_74;
	wire [WIDTH-1:0] wire_d7_75;
	wire [WIDTH-1:0] wire_d7_76;
	wire [WIDTH-1:0] wire_d7_77;
	wire [WIDTH-1:0] wire_d7_78;
	wire [WIDTH-1:0] wire_d7_79;
	wire [WIDTH-1:0] wire_d7_80;
	wire [WIDTH-1:0] wire_d7_81;
	wire [WIDTH-1:0] wire_d7_82;
	wire [WIDTH-1:0] wire_d7_83;
	wire [WIDTH-1:0] wire_d7_84;
	wire [WIDTH-1:0] wire_d7_85;
	wire [WIDTH-1:0] wire_d7_86;
	wire [WIDTH-1:0] wire_d7_87;
	wire [WIDTH-1:0] wire_d7_88;
	wire [WIDTH-1:0] wire_d7_89;
	wire [WIDTH-1:0] wire_d7_90;
	wire [WIDTH-1:0] wire_d7_91;
	wire [WIDTH-1:0] wire_d7_92;
	wire [WIDTH-1:0] wire_d7_93;
	wire [WIDTH-1:0] wire_d7_94;
	wire [WIDTH-1:0] wire_d7_95;
	wire [WIDTH-1:0] wire_d7_96;
	wire [WIDTH-1:0] wire_d7_97;
	wire [WIDTH-1:0] wire_d7_98;
	wire [WIDTH-1:0] wire_d8_0;
	wire [WIDTH-1:0] wire_d8_1;
	wire [WIDTH-1:0] wire_d8_2;
	wire [WIDTH-1:0] wire_d8_3;
	wire [WIDTH-1:0] wire_d8_4;
	wire [WIDTH-1:0] wire_d8_5;
	wire [WIDTH-1:0] wire_d8_6;
	wire [WIDTH-1:0] wire_d8_7;
	wire [WIDTH-1:0] wire_d8_8;
	wire [WIDTH-1:0] wire_d8_9;
	wire [WIDTH-1:0] wire_d8_10;
	wire [WIDTH-1:0] wire_d8_11;
	wire [WIDTH-1:0] wire_d8_12;
	wire [WIDTH-1:0] wire_d8_13;
	wire [WIDTH-1:0] wire_d8_14;
	wire [WIDTH-1:0] wire_d8_15;
	wire [WIDTH-1:0] wire_d8_16;
	wire [WIDTH-1:0] wire_d8_17;
	wire [WIDTH-1:0] wire_d8_18;
	wire [WIDTH-1:0] wire_d8_19;
	wire [WIDTH-1:0] wire_d8_20;
	wire [WIDTH-1:0] wire_d8_21;
	wire [WIDTH-1:0] wire_d8_22;
	wire [WIDTH-1:0] wire_d8_23;
	wire [WIDTH-1:0] wire_d8_24;
	wire [WIDTH-1:0] wire_d8_25;
	wire [WIDTH-1:0] wire_d8_26;
	wire [WIDTH-1:0] wire_d8_27;
	wire [WIDTH-1:0] wire_d8_28;
	wire [WIDTH-1:0] wire_d8_29;
	wire [WIDTH-1:0] wire_d8_30;
	wire [WIDTH-1:0] wire_d8_31;
	wire [WIDTH-1:0] wire_d8_32;
	wire [WIDTH-1:0] wire_d8_33;
	wire [WIDTH-1:0] wire_d8_34;
	wire [WIDTH-1:0] wire_d8_35;
	wire [WIDTH-1:0] wire_d8_36;
	wire [WIDTH-1:0] wire_d8_37;
	wire [WIDTH-1:0] wire_d8_38;
	wire [WIDTH-1:0] wire_d8_39;
	wire [WIDTH-1:0] wire_d8_40;
	wire [WIDTH-1:0] wire_d8_41;
	wire [WIDTH-1:0] wire_d8_42;
	wire [WIDTH-1:0] wire_d8_43;
	wire [WIDTH-1:0] wire_d8_44;
	wire [WIDTH-1:0] wire_d8_45;
	wire [WIDTH-1:0] wire_d8_46;
	wire [WIDTH-1:0] wire_d8_47;
	wire [WIDTH-1:0] wire_d8_48;
	wire [WIDTH-1:0] wire_d8_49;
	wire [WIDTH-1:0] wire_d8_50;
	wire [WIDTH-1:0] wire_d8_51;
	wire [WIDTH-1:0] wire_d8_52;
	wire [WIDTH-1:0] wire_d8_53;
	wire [WIDTH-1:0] wire_d8_54;
	wire [WIDTH-1:0] wire_d8_55;
	wire [WIDTH-1:0] wire_d8_56;
	wire [WIDTH-1:0] wire_d8_57;
	wire [WIDTH-1:0] wire_d8_58;
	wire [WIDTH-1:0] wire_d8_59;
	wire [WIDTH-1:0] wire_d8_60;
	wire [WIDTH-1:0] wire_d8_61;
	wire [WIDTH-1:0] wire_d8_62;
	wire [WIDTH-1:0] wire_d8_63;
	wire [WIDTH-1:0] wire_d8_64;
	wire [WIDTH-1:0] wire_d8_65;
	wire [WIDTH-1:0] wire_d8_66;
	wire [WIDTH-1:0] wire_d8_67;
	wire [WIDTH-1:0] wire_d8_68;
	wire [WIDTH-1:0] wire_d8_69;
	wire [WIDTH-1:0] wire_d8_70;
	wire [WIDTH-1:0] wire_d8_71;
	wire [WIDTH-1:0] wire_d8_72;
	wire [WIDTH-1:0] wire_d8_73;
	wire [WIDTH-1:0] wire_d8_74;
	wire [WIDTH-1:0] wire_d8_75;
	wire [WIDTH-1:0] wire_d8_76;
	wire [WIDTH-1:0] wire_d8_77;
	wire [WIDTH-1:0] wire_d8_78;
	wire [WIDTH-1:0] wire_d8_79;
	wire [WIDTH-1:0] wire_d8_80;
	wire [WIDTH-1:0] wire_d8_81;
	wire [WIDTH-1:0] wire_d8_82;
	wire [WIDTH-1:0] wire_d8_83;
	wire [WIDTH-1:0] wire_d8_84;
	wire [WIDTH-1:0] wire_d8_85;
	wire [WIDTH-1:0] wire_d8_86;
	wire [WIDTH-1:0] wire_d8_87;
	wire [WIDTH-1:0] wire_d8_88;
	wire [WIDTH-1:0] wire_d8_89;
	wire [WIDTH-1:0] wire_d8_90;
	wire [WIDTH-1:0] wire_d8_91;
	wire [WIDTH-1:0] wire_d8_92;
	wire [WIDTH-1:0] wire_d8_93;
	wire [WIDTH-1:0] wire_d8_94;
	wire [WIDTH-1:0] wire_d8_95;
	wire [WIDTH-1:0] wire_d8_96;
	wire [WIDTH-1:0] wire_d8_97;
	wire [WIDTH-1:0] wire_d8_98;
	wire [WIDTH-1:0] wire_d9_0;
	wire [WIDTH-1:0] wire_d9_1;
	wire [WIDTH-1:0] wire_d9_2;
	wire [WIDTH-1:0] wire_d9_3;
	wire [WIDTH-1:0] wire_d9_4;
	wire [WIDTH-1:0] wire_d9_5;
	wire [WIDTH-1:0] wire_d9_6;
	wire [WIDTH-1:0] wire_d9_7;
	wire [WIDTH-1:0] wire_d9_8;
	wire [WIDTH-1:0] wire_d9_9;
	wire [WIDTH-1:0] wire_d9_10;
	wire [WIDTH-1:0] wire_d9_11;
	wire [WIDTH-1:0] wire_d9_12;
	wire [WIDTH-1:0] wire_d9_13;
	wire [WIDTH-1:0] wire_d9_14;
	wire [WIDTH-1:0] wire_d9_15;
	wire [WIDTH-1:0] wire_d9_16;
	wire [WIDTH-1:0] wire_d9_17;
	wire [WIDTH-1:0] wire_d9_18;
	wire [WIDTH-1:0] wire_d9_19;
	wire [WIDTH-1:0] wire_d9_20;
	wire [WIDTH-1:0] wire_d9_21;
	wire [WIDTH-1:0] wire_d9_22;
	wire [WIDTH-1:0] wire_d9_23;
	wire [WIDTH-1:0] wire_d9_24;
	wire [WIDTH-1:0] wire_d9_25;
	wire [WIDTH-1:0] wire_d9_26;
	wire [WIDTH-1:0] wire_d9_27;
	wire [WIDTH-1:0] wire_d9_28;
	wire [WIDTH-1:0] wire_d9_29;
	wire [WIDTH-1:0] wire_d9_30;
	wire [WIDTH-1:0] wire_d9_31;
	wire [WIDTH-1:0] wire_d9_32;
	wire [WIDTH-1:0] wire_d9_33;
	wire [WIDTH-1:0] wire_d9_34;
	wire [WIDTH-1:0] wire_d9_35;
	wire [WIDTH-1:0] wire_d9_36;
	wire [WIDTH-1:0] wire_d9_37;
	wire [WIDTH-1:0] wire_d9_38;
	wire [WIDTH-1:0] wire_d9_39;
	wire [WIDTH-1:0] wire_d9_40;
	wire [WIDTH-1:0] wire_d9_41;
	wire [WIDTH-1:0] wire_d9_42;
	wire [WIDTH-1:0] wire_d9_43;
	wire [WIDTH-1:0] wire_d9_44;
	wire [WIDTH-1:0] wire_d9_45;
	wire [WIDTH-1:0] wire_d9_46;
	wire [WIDTH-1:0] wire_d9_47;
	wire [WIDTH-1:0] wire_d9_48;
	wire [WIDTH-1:0] wire_d9_49;
	wire [WIDTH-1:0] wire_d9_50;
	wire [WIDTH-1:0] wire_d9_51;
	wire [WIDTH-1:0] wire_d9_52;
	wire [WIDTH-1:0] wire_d9_53;
	wire [WIDTH-1:0] wire_d9_54;
	wire [WIDTH-1:0] wire_d9_55;
	wire [WIDTH-1:0] wire_d9_56;
	wire [WIDTH-1:0] wire_d9_57;
	wire [WIDTH-1:0] wire_d9_58;
	wire [WIDTH-1:0] wire_d9_59;
	wire [WIDTH-1:0] wire_d9_60;
	wire [WIDTH-1:0] wire_d9_61;
	wire [WIDTH-1:0] wire_d9_62;
	wire [WIDTH-1:0] wire_d9_63;
	wire [WIDTH-1:0] wire_d9_64;
	wire [WIDTH-1:0] wire_d9_65;
	wire [WIDTH-1:0] wire_d9_66;
	wire [WIDTH-1:0] wire_d9_67;
	wire [WIDTH-1:0] wire_d9_68;
	wire [WIDTH-1:0] wire_d9_69;
	wire [WIDTH-1:0] wire_d9_70;
	wire [WIDTH-1:0] wire_d9_71;
	wire [WIDTH-1:0] wire_d9_72;
	wire [WIDTH-1:0] wire_d9_73;
	wire [WIDTH-1:0] wire_d9_74;
	wire [WIDTH-1:0] wire_d9_75;
	wire [WIDTH-1:0] wire_d9_76;
	wire [WIDTH-1:0] wire_d9_77;
	wire [WIDTH-1:0] wire_d9_78;
	wire [WIDTH-1:0] wire_d9_79;
	wire [WIDTH-1:0] wire_d9_80;
	wire [WIDTH-1:0] wire_d9_81;
	wire [WIDTH-1:0] wire_d9_82;
	wire [WIDTH-1:0] wire_d9_83;
	wire [WIDTH-1:0] wire_d9_84;
	wire [WIDTH-1:0] wire_d9_85;
	wire [WIDTH-1:0] wire_d9_86;
	wire [WIDTH-1:0] wire_d9_87;
	wire [WIDTH-1:0] wire_d9_88;
	wire [WIDTH-1:0] wire_d9_89;
	wire [WIDTH-1:0] wire_d9_90;
	wire [WIDTH-1:0] wire_d9_91;
	wire [WIDTH-1:0] wire_d9_92;
	wire [WIDTH-1:0] wire_d9_93;
	wire [WIDTH-1:0] wire_d9_94;
	wire [WIDTH-1:0] wire_d9_95;
	wire [WIDTH-1:0] wire_d9_96;
	wire [WIDTH-1:0] wire_d9_97;
	wire [WIDTH-1:0] wire_d9_98;
	wire [WIDTH-1:0] wire_d10_0;
	wire [WIDTH-1:0] wire_d10_1;
	wire [WIDTH-1:0] wire_d10_2;
	wire [WIDTH-1:0] wire_d10_3;
	wire [WIDTH-1:0] wire_d10_4;
	wire [WIDTH-1:0] wire_d10_5;
	wire [WIDTH-1:0] wire_d10_6;
	wire [WIDTH-1:0] wire_d10_7;
	wire [WIDTH-1:0] wire_d10_8;
	wire [WIDTH-1:0] wire_d10_9;
	wire [WIDTH-1:0] wire_d10_10;
	wire [WIDTH-1:0] wire_d10_11;
	wire [WIDTH-1:0] wire_d10_12;
	wire [WIDTH-1:0] wire_d10_13;
	wire [WIDTH-1:0] wire_d10_14;
	wire [WIDTH-1:0] wire_d10_15;
	wire [WIDTH-1:0] wire_d10_16;
	wire [WIDTH-1:0] wire_d10_17;
	wire [WIDTH-1:0] wire_d10_18;
	wire [WIDTH-1:0] wire_d10_19;
	wire [WIDTH-1:0] wire_d10_20;
	wire [WIDTH-1:0] wire_d10_21;
	wire [WIDTH-1:0] wire_d10_22;
	wire [WIDTH-1:0] wire_d10_23;
	wire [WIDTH-1:0] wire_d10_24;
	wire [WIDTH-1:0] wire_d10_25;
	wire [WIDTH-1:0] wire_d10_26;
	wire [WIDTH-1:0] wire_d10_27;
	wire [WIDTH-1:0] wire_d10_28;
	wire [WIDTH-1:0] wire_d10_29;
	wire [WIDTH-1:0] wire_d10_30;
	wire [WIDTH-1:0] wire_d10_31;
	wire [WIDTH-1:0] wire_d10_32;
	wire [WIDTH-1:0] wire_d10_33;
	wire [WIDTH-1:0] wire_d10_34;
	wire [WIDTH-1:0] wire_d10_35;
	wire [WIDTH-1:0] wire_d10_36;
	wire [WIDTH-1:0] wire_d10_37;
	wire [WIDTH-1:0] wire_d10_38;
	wire [WIDTH-1:0] wire_d10_39;
	wire [WIDTH-1:0] wire_d10_40;
	wire [WIDTH-1:0] wire_d10_41;
	wire [WIDTH-1:0] wire_d10_42;
	wire [WIDTH-1:0] wire_d10_43;
	wire [WIDTH-1:0] wire_d10_44;
	wire [WIDTH-1:0] wire_d10_45;
	wire [WIDTH-1:0] wire_d10_46;
	wire [WIDTH-1:0] wire_d10_47;
	wire [WIDTH-1:0] wire_d10_48;
	wire [WIDTH-1:0] wire_d10_49;
	wire [WIDTH-1:0] wire_d10_50;
	wire [WIDTH-1:0] wire_d10_51;
	wire [WIDTH-1:0] wire_d10_52;
	wire [WIDTH-1:0] wire_d10_53;
	wire [WIDTH-1:0] wire_d10_54;
	wire [WIDTH-1:0] wire_d10_55;
	wire [WIDTH-1:0] wire_d10_56;
	wire [WIDTH-1:0] wire_d10_57;
	wire [WIDTH-1:0] wire_d10_58;
	wire [WIDTH-1:0] wire_d10_59;
	wire [WIDTH-1:0] wire_d10_60;
	wire [WIDTH-1:0] wire_d10_61;
	wire [WIDTH-1:0] wire_d10_62;
	wire [WIDTH-1:0] wire_d10_63;
	wire [WIDTH-1:0] wire_d10_64;
	wire [WIDTH-1:0] wire_d10_65;
	wire [WIDTH-1:0] wire_d10_66;
	wire [WIDTH-1:0] wire_d10_67;
	wire [WIDTH-1:0] wire_d10_68;
	wire [WIDTH-1:0] wire_d10_69;
	wire [WIDTH-1:0] wire_d10_70;
	wire [WIDTH-1:0] wire_d10_71;
	wire [WIDTH-1:0] wire_d10_72;
	wire [WIDTH-1:0] wire_d10_73;
	wire [WIDTH-1:0] wire_d10_74;
	wire [WIDTH-1:0] wire_d10_75;
	wire [WIDTH-1:0] wire_d10_76;
	wire [WIDTH-1:0] wire_d10_77;
	wire [WIDTH-1:0] wire_d10_78;
	wire [WIDTH-1:0] wire_d10_79;
	wire [WIDTH-1:0] wire_d10_80;
	wire [WIDTH-1:0] wire_d10_81;
	wire [WIDTH-1:0] wire_d10_82;
	wire [WIDTH-1:0] wire_d10_83;
	wire [WIDTH-1:0] wire_d10_84;
	wire [WIDTH-1:0] wire_d10_85;
	wire [WIDTH-1:0] wire_d10_86;
	wire [WIDTH-1:0] wire_d10_87;
	wire [WIDTH-1:0] wire_d10_88;
	wire [WIDTH-1:0] wire_d10_89;
	wire [WIDTH-1:0] wire_d10_90;
	wire [WIDTH-1:0] wire_d10_91;
	wire [WIDTH-1:0] wire_d10_92;
	wire [WIDTH-1:0] wire_d10_93;
	wire [WIDTH-1:0] wire_d10_94;
	wire [WIDTH-1:0] wire_d10_95;
	wire [WIDTH-1:0] wire_d10_96;
	wire [WIDTH-1:0] wire_d10_97;
	wire [WIDTH-1:0] wire_d10_98;
	wire [WIDTH-1:0] wire_d11_0;
	wire [WIDTH-1:0] wire_d11_1;
	wire [WIDTH-1:0] wire_d11_2;
	wire [WIDTH-1:0] wire_d11_3;
	wire [WIDTH-1:0] wire_d11_4;
	wire [WIDTH-1:0] wire_d11_5;
	wire [WIDTH-1:0] wire_d11_6;
	wire [WIDTH-1:0] wire_d11_7;
	wire [WIDTH-1:0] wire_d11_8;
	wire [WIDTH-1:0] wire_d11_9;
	wire [WIDTH-1:0] wire_d11_10;
	wire [WIDTH-1:0] wire_d11_11;
	wire [WIDTH-1:0] wire_d11_12;
	wire [WIDTH-1:0] wire_d11_13;
	wire [WIDTH-1:0] wire_d11_14;
	wire [WIDTH-1:0] wire_d11_15;
	wire [WIDTH-1:0] wire_d11_16;
	wire [WIDTH-1:0] wire_d11_17;
	wire [WIDTH-1:0] wire_d11_18;
	wire [WIDTH-1:0] wire_d11_19;
	wire [WIDTH-1:0] wire_d11_20;
	wire [WIDTH-1:0] wire_d11_21;
	wire [WIDTH-1:0] wire_d11_22;
	wire [WIDTH-1:0] wire_d11_23;
	wire [WIDTH-1:0] wire_d11_24;
	wire [WIDTH-1:0] wire_d11_25;
	wire [WIDTH-1:0] wire_d11_26;
	wire [WIDTH-1:0] wire_d11_27;
	wire [WIDTH-1:0] wire_d11_28;
	wire [WIDTH-1:0] wire_d11_29;
	wire [WIDTH-1:0] wire_d11_30;
	wire [WIDTH-1:0] wire_d11_31;
	wire [WIDTH-1:0] wire_d11_32;
	wire [WIDTH-1:0] wire_d11_33;
	wire [WIDTH-1:0] wire_d11_34;
	wire [WIDTH-1:0] wire_d11_35;
	wire [WIDTH-1:0] wire_d11_36;
	wire [WIDTH-1:0] wire_d11_37;
	wire [WIDTH-1:0] wire_d11_38;
	wire [WIDTH-1:0] wire_d11_39;
	wire [WIDTH-1:0] wire_d11_40;
	wire [WIDTH-1:0] wire_d11_41;
	wire [WIDTH-1:0] wire_d11_42;
	wire [WIDTH-1:0] wire_d11_43;
	wire [WIDTH-1:0] wire_d11_44;
	wire [WIDTH-1:0] wire_d11_45;
	wire [WIDTH-1:0] wire_d11_46;
	wire [WIDTH-1:0] wire_d11_47;
	wire [WIDTH-1:0] wire_d11_48;
	wire [WIDTH-1:0] wire_d11_49;
	wire [WIDTH-1:0] wire_d11_50;
	wire [WIDTH-1:0] wire_d11_51;
	wire [WIDTH-1:0] wire_d11_52;
	wire [WIDTH-1:0] wire_d11_53;
	wire [WIDTH-1:0] wire_d11_54;
	wire [WIDTH-1:0] wire_d11_55;
	wire [WIDTH-1:0] wire_d11_56;
	wire [WIDTH-1:0] wire_d11_57;
	wire [WIDTH-1:0] wire_d11_58;
	wire [WIDTH-1:0] wire_d11_59;
	wire [WIDTH-1:0] wire_d11_60;
	wire [WIDTH-1:0] wire_d11_61;
	wire [WIDTH-1:0] wire_d11_62;
	wire [WIDTH-1:0] wire_d11_63;
	wire [WIDTH-1:0] wire_d11_64;
	wire [WIDTH-1:0] wire_d11_65;
	wire [WIDTH-1:0] wire_d11_66;
	wire [WIDTH-1:0] wire_d11_67;
	wire [WIDTH-1:0] wire_d11_68;
	wire [WIDTH-1:0] wire_d11_69;
	wire [WIDTH-1:0] wire_d11_70;
	wire [WIDTH-1:0] wire_d11_71;
	wire [WIDTH-1:0] wire_d11_72;
	wire [WIDTH-1:0] wire_d11_73;
	wire [WIDTH-1:0] wire_d11_74;
	wire [WIDTH-1:0] wire_d11_75;
	wire [WIDTH-1:0] wire_d11_76;
	wire [WIDTH-1:0] wire_d11_77;
	wire [WIDTH-1:0] wire_d11_78;
	wire [WIDTH-1:0] wire_d11_79;
	wire [WIDTH-1:0] wire_d11_80;
	wire [WIDTH-1:0] wire_d11_81;
	wire [WIDTH-1:0] wire_d11_82;
	wire [WIDTH-1:0] wire_d11_83;
	wire [WIDTH-1:0] wire_d11_84;
	wire [WIDTH-1:0] wire_d11_85;
	wire [WIDTH-1:0] wire_d11_86;
	wire [WIDTH-1:0] wire_d11_87;
	wire [WIDTH-1:0] wire_d11_88;
	wire [WIDTH-1:0] wire_d11_89;
	wire [WIDTH-1:0] wire_d11_90;
	wire [WIDTH-1:0] wire_d11_91;
	wire [WIDTH-1:0] wire_d11_92;
	wire [WIDTH-1:0] wire_d11_93;
	wire [WIDTH-1:0] wire_d11_94;
	wire [WIDTH-1:0] wire_d11_95;
	wire [WIDTH-1:0] wire_d11_96;
	wire [WIDTH-1:0] wire_d11_97;
	wire [WIDTH-1:0] wire_d11_98;
	wire [WIDTH-1:0] wire_d12_0;
	wire [WIDTH-1:0] wire_d12_1;
	wire [WIDTH-1:0] wire_d12_2;
	wire [WIDTH-1:0] wire_d12_3;
	wire [WIDTH-1:0] wire_d12_4;
	wire [WIDTH-1:0] wire_d12_5;
	wire [WIDTH-1:0] wire_d12_6;
	wire [WIDTH-1:0] wire_d12_7;
	wire [WIDTH-1:0] wire_d12_8;
	wire [WIDTH-1:0] wire_d12_9;
	wire [WIDTH-1:0] wire_d12_10;
	wire [WIDTH-1:0] wire_d12_11;
	wire [WIDTH-1:0] wire_d12_12;
	wire [WIDTH-1:0] wire_d12_13;
	wire [WIDTH-1:0] wire_d12_14;
	wire [WIDTH-1:0] wire_d12_15;
	wire [WIDTH-1:0] wire_d12_16;
	wire [WIDTH-1:0] wire_d12_17;
	wire [WIDTH-1:0] wire_d12_18;
	wire [WIDTH-1:0] wire_d12_19;
	wire [WIDTH-1:0] wire_d12_20;
	wire [WIDTH-1:0] wire_d12_21;
	wire [WIDTH-1:0] wire_d12_22;
	wire [WIDTH-1:0] wire_d12_23;
	wire [WIDTH-1:0] wire_d12_24;
	wire [WIDTH-1:0] wire_d12_25;
	wire [WIDTH-1:0] wire_d12_26;
	wire [WIDTH-1:0] wire_d12_27;
	wire [WIDTH-1:0] wire_d12_28;
	wire [WIDTH-1:0] wire_d12_29;
	wire [WIDTH-1:0] wire_d12_30;
	wire [WIDTH-1:0] wire_d12_31;
	wire [WIDTH-1:0] wire_d12_32;
	wire [WIDTH-1:0] wire_d12_33;
	wire [WIDTH-1:0] wire_d12_34;
	wire [WIDTH-1:0] wire_d12_35;
	wire [WIDTH-1:0] wire_d12_36;
	wire [WIDTH-1:0] wire_d12_37;
	wire [WIDTH-1:0] wire_d12_38;
	wire [WIDTH-1:0] wire_d12_39;
	wire [WIDTH-1:0] wire_d12_40;
	wire [WIDTH-1:0] wire_d12_41;
	wire [WIDTH-1:0] wire_d12_42;
	wire [WIDTH-1:0] wire_d12_43;
	wire [WIDTH-1:0] wire_d12_44;
	wire [WIDTH-1:0] wire_d12_45;
	wire [WIDTH-1:0] wire_d12_46;
	wire [WIDTH-1:0] wire_d12_47;
	wire [WIDTH-1:0] wire_d12_48;
	wire [WIDTH-1:0] wire_d12_49;
	wire [WIDTH-1:0] wire_d12_50;
	wire [WIDTH-1:0] wire_d12_51;
	wire [WIDTH-1:0] wire_d12_52;
	wire [WIDTH-1:0] wire_d12_53;
	wire [WIDTH-1:0] wire_d12_54;
	wire [WIDTH-1:0] wire_d12_55;
	wire [WIDTH-1:0] wire_d12_56;
	wire [WIDTH-1:0] wire_d12_57;
	wire [WIDTH-1:0] wire_d12_58;
	wire [WIDTH-1:0] wire_d12_59;
	wire [WIDTH-1:0] wire_d12_60;
	wire [WIDTH-1:0] wire_d12_61;
	wire [WIDTH-1:0] wire_d12_62;
	wire [WIDTH-1:0] wire_d12_63;
	wire [WIDTH-1:0] wire_d12_64;
	wire [WIDTH-1:0] wire_d12_65;
	wire [WIDTH-1:0] wire_d12_66;
	wire [WIDTH-1:0] wire_d12_67;
	wire [WIDTH-1:0] wire_d12_68;
	wire [WIDTH-1:0] wire_d12_69;
	wire [WIDTH-1:0] wire_d12_70;
	wire [WIDTH-1:0] wire_d12_71;
	wire [WIDTH-1:0] wire_d12_72;
	wire [WIDTH-1:0] wire_d12_73;
	wire [WIDTH-1:0] wire_d12_74;
	wire [WIDTH-1:0] wire_d12_75;
	wire [WIDTH-1:0] wire_d12_76;
	wire [WIDTH-1:0] wire_d12_77;
	wire [WIDTH-1:0] wire_d12_78;
	wire [WIDTH-1:0] wire_d12_79;
	wire [WIDTH-1:0] wire_d12_80;
	wire [WIDTH-1:0] wire_d12_81;
	wire [WIDTH-1:0] wire_d12_82;
	wire [WIDTH-1:0] wire_d12_83;
	wire [WIDTH-1:0] wire_d12_84;
	wire [WIDTH-1:0] wire_d12_85;
	wire [WIDTH-1:0] wire_d12_86;
	wire [WIDTH-1:0] wire_d12_87;
	wire [WIDTH-1:0] wire_d12_88;
	wire [WIDTH-1:0] wire_d12_89;
	wire [WIDTH-1:0] wire_d12_90;
	wire [WIDTH-1:0] wire_d12_91;
	wire [WIDTH-1:0] wire_d12_92;
	wire [WIDTH-1:0] wire_d12_93;
	wire [WIDTH-1:0] wire_d12_94;
	wire [WIDTH-1:0] wire_d12_95;
	wire [WIDTH-1:0] wire_d12_96;
	wire [WIDTH-1:0] wire_d12_97;
	wire [WIDTH-1:0] wire_d12_98;
	wire [WIDTH-1:0] wire_d13_0;
	wire [WIDTH-1:0] wire_d13_1;
	wire [WIDTH-1:0] wire_d13_2;
	wire [WIDTH-1:0] wire_d13_3;
	wire [WIDTH-1:0] wire_d13_4;
	wire [WIDTH-1:0] wire_d13_5;
	wire [WIDTH-1:0] wire_d13_6;
	wire [WIDTH-1:0] wire_d13_7;
	wire [WIDTH-1:0] wire_d13_8;
	wire [WIDTH-1:0] wire_d13_9;
	wire [WIDTH-1:0] wire_d13_10;
	wire [WIDTH-1:0] wire_d13_11;
	wire [WIDTH-1:0] wire_d13_12;
	wire [WIDTH-1:0] wire_d13_13;
	wire [WIDTH-1:0] wire_d13_14;
	wire [WIDTH-1:0] wire_d13_15;
	wire [WIDTH-1:0] wire_d13_16;
	wire [WIDTH-1:0] wire_d13_17;
	wire [WIDTH-1:0] wire_d13_18;
	wire [WIDTH-1:0] wire_d13_19;
	wire [WIDTH-1:0] wire_d13_20;
	wire [WIDTH-1:0] wire_d13_21;
	wire [WIDTH-1:0] wire_d13_22;
	wire [WIDTH-1:0] wire_d13_23;
	wire [WIDTH-1:0] wire_d13_24;
	wire [WIDTH-1:0] wire_d13_25;
	wire [WIDTH-1:0] wire_d13_26;
	wire [WIDTH-1:0] wire_d13_27;
	wire [WIDTH-1:0] wire_d13_28;
	wire [WIDTH-1:0] wire_d13_29;
	wire [WIDTH-1:0] wire_d13_30;
	wire [WIDTH-1:0] wire_d13_31;
	wire [WIDTH-1:0] wire_d13_32;
	wire [WIDTH-1:0] wire_d13_33;
	wire [WIDTH-1:0] wire_d13_34;
	wire [WIDTH-1:0] wire_d13_35;
	wire [WIDTH-1:0] wire_d13_36;
	wire [WIDTH-1:0] wire_d13_37;
	wire [WIDTH-1:0] wire_d13_38;
	wire [WIDTH-1:0] wire_d13_39;
	wire [WIDTH-1:0] wire_d13_40;
	wire [WIDTH-1:0] wire_d13_41;
	wire [WIDTH-1:0] wire_d13_42;
	wire [WIDTH-1:0] wire_d13_43;
	wire [WIDTH-1:0] wire_d13_44;
	wire [WIDTH-1:0] wire_d13_45;
	wire [WIDTH-1:0] wire_d13_46;
	wire [WIDTH-1:0] wire_d13_47;
	wire [WIDTH-1:0] wire_d13_48;
	wire [WIDTH-1:0] wire_d13_49;
	wire [WIDTH-1:0] wire_d13_50;
	wire [WIDTH-1:0] wire_d13_51;
	wire [WIDTH-1:0] wire_d13_52;
	wire [WIDTH-1:0] wire_d13_53;
	wire [WIDTH-1:0] wire_d13_54;
	wire [WIDTH-1:0] wire_d13_55;
	wire [WIDTH-1:0] wire_d13_56;
	wire [WIDTH-1:0] wire_d13_57;
	wire [WIDTH-1:0] wire_d13_58;
	wire [WIDTH-1:0] wire_d13_59;
	wire [WIDTH-1:0] wire_d13_60;
	wire [WIDTH-1:0] wire_d13_61;
	wire [WIDTH-1:0] wire_d13_62;
	wire [WIDTH-1:0] wire_d13_63;
	wire [WIDTH-1:0] wire_d13_64;
	wire [WIDTH-1:0] wire_d13_65;
	wire [WIDTH-1:0] wire_d13_66;
	wire [WIDTH-1:0] wire_d13_67;
	wire [WIDTH-1:0] wire_d13_68;
	wire [WIDTH-1:0] wire_d13_69;
	wire [WIDTH-1:0] wire_d13_70;
	wire [WIDTH-1:0] wire_d13_71;
	wire [WIDTH-1:0] wire_d13_72;
	wire [WIDTH-1:0] wire_d13_73;
	wire [WIDTH-1:0] wire_d13_74;
	wire [WIDTH-1:0] wire_d13_75;
	wire [WIDTH-1:0] wire_d13_76;
	wire [WIDTH-1:0] wire_d13_77;
	wire [WIDTH-1:0] wire_d13_78;
	wire [WIDTH-1:0] wire_d13_79;
	wire [WIDTH-1:0] wire_d13_80;
	wire [WIDTH-1:0] wire_d13_81;
	wire [WIDTH-1:0] wire_d13_82;
	wire [WIDTH-1:0] wire_d13_83;
	wire [WIDTH-1:0] wire_d13_84;
	wire [WIDTH-1:0] wire_d13_85;
	wire [WIDTH-1:0] wire_d13_86;
	wire [WIDTH-1:0] wire_d13_87;
	wire [WIDTH-1:0] wire_d13_88;
	wire [WIDTH-1:0] wire_d13_89;
	wire [WIDTH-1:0] wire_d13_90;
	wire [WIDTH-1:0] wire_d13_91;
	wire [WIDTH-1:0] wire_d13_92;
	wire [WIDTH-1:0] wire_d13_93;
	wire [WIDTH-1:0] wire_d13_94;
	wire [WIDTH-1:0] wire_d13_95;
	wire [WIDTH-1:0] wire_d13_96;
	wire [WIDTH-1:0] wire_d13_97;
	wire [WIDTH-1:0] wire_d13_98;
	wire [WIDTH-1:0] wire_d14_0;
	wire [WIDTH-1:0] wire_d14_1;
	wire [WIDTH-1:0] wire_d14_2;
	wire [WIDTH-1:0] wire_d14_3;
	wire [WIDTH-1:0] wire_d14_4;
	wire [WIDTH-1:0] wire_d14_5;
	wire [WIDTH-1:0] wire_d14_6;
	wire [WIDTH-1:0] wire_d14_7;
	wire [WIDTH-1:0] wire_d14_8;
	wire [WIDTH-1:0] wire_d14_9;
	wire [WIDTH-1:0] wire_d14_10;
	wire [WIDTH-1:0] wire_d14_11;
	wire [WIDTH-1:0] wire_d14_12;
	wire [WIDTH-1:0] wire_d14_13;
	wire [WIDTH-1:0] wire_d14_14;
	wire [WIDTH-1:0] wire_d14_15;
	wire [WIDTH-1:0] wire_d14_16;
	wire [WIDTH-1:0] wire_d14_17;
	wire [WIDTH-1:0] wire_d14_18;
	wire [WIDTH-1:0] wire_d14_19;
	wire [WIDTH-1:0] wire_d14_20;
	wire [WIDTH-1:0] wire_d14_21;
	wire [WIDTH-1:0] wire_d14_22;
	wire [WIDTH-1:0] wire_d14_23;
	wire [WIDTH-1:0] wire_d14_24;
	wire [WIDTH-1:0] wire_d14_25;
	wire [WIDTH-1:0] wire_d14_26;
	wire [WIDTH-1:0] wire_d14_27;
	wire [WIDTH-1:0] wire_d14_28;
	wire [WIDTH-1:0] wire_d14_29;
	wire [WIDTH-1:0] wire_d14_30;
	wire [WIDTH-1:0] wire_d14_31;
	wire [WIDTH-1:0] wire_d14_32;
	wire [WIDTH-1:0] wire_d14_33;
	wire [WIDTH-1:0] wire_d14_34;
	wire [WIDTH-1:0] wire_d14_35;
	wire [WIDTH-1:0] wire_d14_36;
	wire [WIDTH-1:0] wire_d14_37;
	wire [WIDTH-1:0] wire_d14_38;
	wire [WIDTH-1:0] wire_d14_39;
	wire [WIDTH-1:0] wire_d14_40;
	wire [WIDTH-1:0] wire_d14_41;
	wire [WIDTH-1:0] wire_d14_42;
	wire [WIDTH-1:0] wire_d14_43;
	wire [WIDTH-1:0] wire_d14_44;
	wire [WIDTH-1:0] wire_d14_45;
	wire [WIDTH-1:0] wire_d14_46;
	wire [WIDTH-1:0] wire_d14_47;
	wire [WIDTH-1:0] wire_d14_48;
	wire [WIDTH-1:0] wire_d14_49;
	wire [WIDTH-1:0] wire_d14_50;
	wire [WIDTH-1:0] wire_d14_51;
	wire [WIDTH-1:0] wire_d14_52;
	wire [WIDTH-1:0] wire_d14_53;
	wire [WIDTH-1:0] wire_d14_54;
	wire [WIDTH-1:0] wire_d14_55;
	wire [WIDTH-1:0] wire_d14_56;
	wire [WIDTH-1:0] wire_d14_57;
	wire [WIDTH-1:0] wire_d14_58;
	wire [WIDTH-1:0] wire_d14_59;
	wire [WIDTH-1:0] wire_d14_60;
	wire [WIDTH-1:0] wire_d14_61;
	wire [WIDTH-1:0] wire_d14_62;
	wire [WIDTH-1:0] wire_d14_63;
	wire [WIDTH-1:0] wire_d14_64;
	wire [WIDTH-1:0] wire_d14_65;
	wire [WIDTH-1:0] wire_d14_66;
	wire [WIDTH-1:0] wire_d14_67;
	wire [WIDTH-1:0] wire_d14_68;
	wire [WIDTH-1:0] wire_d14_69;
	wire [WIDTH-1:0] wire_d14_70;
	wire [WIDTH-1:0] wire_d14_71;
	wire [WIDTH-1:0] wire_d14_72;
	wire [WIDTH-1:0] wire_d14_73;
	wire [WIDTH-1:0] wire_d14_74;
	wire [WIDTH-1:0] wire_d14_75;
	wire [WIDTH-1:0] wire_d14_76;
	wire [WIDTH-1:0] wire_d14_77;
	wire [WIDTH-1:0] wire_d14_78;
	wire [WIDTH-1:0] wire_d14_79;
	wire [WIDTH-1:0] wire_d14_80;
	wire [WIDTH-1:0] wire_d14_81;
	wire [WIDTH-1:0] wire_d14_82;
	wire [WIDTH-1:0] wire_d14_83;
	wire [WIDTH-1:0] wire_d14_84;
	wire [WIDTH-1:0] wire_d14_85;
	wire [WIDTH-1:0] wire_d14_86;
	wire [WIDTH-1:0] wire_d14_87;
	wire [WIDTH-1:0] wire_d14_88;
	wire [WIDTH-1:0] wire_d14_89;
	wire [WIDTH-1:0] wire_d14_90;
	wire [WIDTH-1:0] wire_d14_91;
	wire [WIDTH-1:0] wire_d14_92;
	wire [WIDTH-1:0] wire_d14_93;
	wire [WIDTH-1:0] wire_d14_94;
	wire [WIDTH-1:0] wire_d14_95;
	wire [WIDTH-1:0] wire_d14_96;
	wire [WIDTH-1:0] wire_d14_97;
	wire [WIDTH-1:0] wire_d14_98;
	wire [WIDTH-1:0] wire_d15_0;
	wire [WIDTH-1:0] wire_d15_1;
	wire [WIDTH-1:0] wire_d15_2;
	wire [WIDTH-1:0] wire_d15_3;
	wire [WIDTH-1:0] wire_d15_4;
	wire [WIDTH-1:0] wire_d15_5;
	wire [WIDTH-1:0] wire_d15_6;
	wire [WIDTH-1:0] wire_d15_7;
	wire [WIDTH-1:0] wire_d15_8;
	wire [WIDTH-1:0] wire_d15_9;
	wire [WIDTH-1:0] wire_d15_10;
	wire [WIDTH-1:0] wire_d15_11;
	wire [WIDTH-1:0] wire_d15_12;
	wire [WIDTH-1:0] wire_d15_13;
	wire [WIDTH-1:0] wire_d15_14;
	wire [WIDTH-1:0] wire_d15_15;
	wire [WIDTH-1:0] wire_d15_16;
	wire [WIDTH-1:0] wire_d15_17;
	wire [WIDTH-1:0] wire_d15_18;
	wire [WIDTH-1:0] wire_d15_19;
	wire [WIDTH-1:0] wire_d15_20;
	wire [WIDTH-1:0] wire_d15_21;
	wire [WIDTH-1:0] wire_d15_22;
	wire [WIDTH-1:0] wire_d15_23;
	wire [WIDTH-1:0] wire_d15_24;
	wire [WIDTH-1:0] wire_d15_25;
	wire [WIDTH-1:0] wire_d15_26;
	wire [WIDTH-1:0] wire_d15_27;
	wire [WIDTH-1:0] wire_d15_28;
	wire [WIDTH-1:0] wire_d15_29;
	wire [WIDTH-1:0] wire_d15_30;
	wire [WIDTH-1:0] wire_d15_31;
	wire [WIDTH-1:0] wire_d15_32;
	wire [WIDTH-1:0] wire_d15_33;
	wire [WIDTH-1:0] wire_d15_34;
	wire [WIDTH-1:0] wire_d15_35;
	wire [WIDTH-1:0] wire_d15_36;
	wire [WIDTH-1:0] wire_d15_37;
	wire [WIDTH-1:0] wire_d15_38;
	wire [WIDTH-1:0] wire_d15_39;
	wire [WIDTH-1:0] wire_d15_40;
	wire [WIDTH-1:0] wire_d15_41;
	wire [WIDTH-1:0] wire_d15_42;
	wire [WIDTH-1:0] wire_d15_43;
	wire [WIDTH-1:0] wire_d15_44;
	wire [WIDTH-1:0] wire_d15_45;
	wire [WIDTH-1:0] wire_d15_46;
	wire [WIDTH-1:0] wire_d15_47;
	wire [WIDTH-1:0] wire_d15_48;
	wire [WIDTH-1:0] wire_d15_49;
	wire [WIDTH-1:0] wire_d15_50;
	wire [WIDTH-1:0] wire_d15_51;
	wire [WIDTH-1:0] wire_d15_52;
	wire [WIDTH-1:0] wire_d15_53;
	wire [WIDTH-1:0] wire_d15_54;
	wire [WIDTH-1:0] wire_d15_55;
	wire [WIDTH-1:0] wire_d15_56;
	wire [WIDTH-1:0] wire_d15_57;
	wire [WIDTH-1:0] wire_d15_58;
	wire [WIDTH-1:0] wire_d15_59;
	wire [WIDTH-1:0] wire_d15_60;
	wire [WIDTH-1:0] wire_d15_61;
	wire [WIDTH-1:0] wire_d15_62;
	wire [WIDTH-1:0] wire_d15_63;
	wire [WIDTH-1:0] wire_d15_64;
	wire [WIDTH-1:0] wire_d15_65;
	wire [WIDTH-1:0] wire_d15_66;
	wire [WIDTH-1:0] wire_d15_67;
	wire [WIDTH-1:0] wire_d15_68;
	wire [WIDTH-1:0] wire_d15_69;
	wire [WIDTH-1:0] wire_d15_70;
	wire [WIDTH-1:0] wire_d15_71;
	wire [WIDTH-1:0] wire_d15_72;
	wire [WIDTH-1:0] wire_d15_73;
	wire [WIDTH-1:0] wire_d15_74;
	wire [WIDTH-1:0] wire_d15_75;
	wire [WIDTH-1:0] wire_d15_76;
	wire [WIDTH-1:0] wire_d15_77;
	wire [WIDTH-1:0] wire_d15_78;
	wire [WIDTH-1:0] wire_d15_79;
	wire [WIDTH-1:0] wire_d15_80;
	wire [WIDTH-1:0] wire_d15_81;
	wire [WIDTH-1:0] wire_d15_82;
	wire [WIDTH-1:0] wire_d15_83;
	wire [WIDTH-1:0] wire_d15_84;
	wire [WIDTH-1:0] wire_d15_85;
	wire [WIDTH-1:0] wire_d15_86;
	wire [WIDTH-1:0] wire_d15_87;
	wire [WIDTH-1:0] wire_d15_88;
	wire [WIDTH-1:0] wire_d15_89;
	wire [WIDTH-1:0] wire_d15_90;
	wire [WIDTH-1:0] wire_d15_91;
	wire [WIDTH-1:0] wire_d15_92;
	wire [WIDTH-1:0] wire_d15_93;
	wire [WIDTH-1:0] wire_d15_94;
	wire [WIDTH-1:0] wire_d15_95;
	wire [WIDTH-1:0] wire_d15_96;
	wire [WIDTH-1:0] wire_d15_97;
	wire [WIDTH-1:0] wire_d15_98;
	wire [WIDTH-1:0] wire_d16_0;
	wire [WIDTH-1:0] wire_d16_1;
	wire [WIDTH-1:0] wire_d16_2;
	wire [WIDTH-1:0] wire_d16_3;
	wire [WIDTH-1:0] wire_d16_4;
	wire [WIDTH-1:0] wire_d16_5;
	wire [WIDTH-1:0] wire_d16_6;
	wire [WIDTH-1:0] wire_d16_7;
	wire [WIDTH-1:0] wire_d16_8;
	wire [WIDTH-1:0] wire_d16_9;
	wire [WIDTH-1:0] wire_d16_10;
	wire [WIDTH-1:0] wire_d16_11;
	wire [WIDTH-1:0] wire_d16_12;
	wire [WIDTH-1:0] wire_d16_13;
	wire [WIDTH-1:0] wire_d16_14;
	wire [WIDTH-1:0] wire_d16_15;
	wire [WIDTH-1:0] wire_d16_16;
	wire [WIDTH-1:0] wire_d16_17;
	wire [WIDTH-1:0] wire_d16_18;
	wire [WIDTH-1:0] wire_d16_19;
	wire [WIDTH-1:0] wire_d16_20;
	wire [WIDTH-1:0] wire_d16_21;
	wire [WIDTH-1:0] wire_d16_22;
	wire [WIDTH-1:0] wire_d16_23;
	wire [WIDTH-1:0] wire_d16_24;
	wire [WIDTH-1:0] wire_d16_25;
	wire [WIDTH-1:0] wire_d16_26;
	wire [WIDTH-1:0] wire_d16_27;
	wire [WIDTH-1:0] wire_d16_28;
	wire [WIDTH-1:0] wire_d16_29;
	wire [WIDTH-1:0] wire_d16_30;
	wire [WIDTH-1:0] wire_d16_31;
	wire [WIDTH-1:0] wire_d16_32;
	wire [WIDTH-1:0] wire_d16_33;
	wire [WIDTH-1:0] wire_d16_34;
	wire [WIDTH-1:0] wire_d16_35;
	wire [WIDTH-1:0] wire_d16_36;
	wire [WIDTH-1:0] wire_d16_37;
	wire [WIDTH-1:0] wire_d16_38;
	wire [WIDTH-1:0] wire_d16_39;
	wire [WIDTH-1:0] wire_d16_40;
	wire [WIDTH-1:0] wire_d16_41;
	wire [WIDTH-1:0] wire_d16_42;
	wire [WIDTH-1:0] wire_d16_43;
	wire [WIDTH-1:0] wire_d16_44;
	wire [WIDTH-1:0] wire_d16_45;
	wire [WIDTH-1:0] wire_d16_46;
	wire [WIDTH-1:0] wire_d16_47;
	wire [WIDTH-1:0] wire_d16_48;
	wire [WIDTH-1:0] wire_d16_49;
	wire [WIDTH-1:0] wire_d16_50;
	wire [WIDTH-1:0] wire_d16_51;
	wire [WIDTH-1:0] wire_d16_52;
	wire [WIDTH-1:0] wire_d16_53;
	wire [WIDTH-1:0] wire_d16_54;
	wire [WIDTH-1:0] wire_d16_55;
	wire [WIDTH-1:0] wire_d16_56;
	wire [WIDTH-1:0] wire_d16_57;
	wire [WIDTH-1:0] wire_d16_58;
	wire [WIDTH-1:0] wire_d16_59;
	wire [WIDTH-1:0] wire_d16_60;
	wire [WIDTH-1:0] wire_d16_61;
	wire [WIDTH-1:0] wire_d16_62;
	wire [WIDTH-1:0] wire_d16_63;
	wire [WIDTH-1:0] wire_d16_64;
	wire [WIDTH-1:0] wire_d16_65;
	wire [WIDTH-1:0] wire_d16_66;
	wire [WIDTH-1:0] wire_d16_67;
	wire [WIDTH-1:0] wire_d16_68;
	wire [WIDTH-1:0] wire_d16_69;
	wire [WIDTH-1:0] wire_d16_70;
	wire [WIDTH-1:0] wire_d16_71;
	wire [WIDTH-1:0] wire_d16_72;
	wire [WIDTH-1:0] wire_d16_73;
	wire [WIDTH-1:0] wire_d16_74;
	wire [WIDTH-1:0] wire_d16_75;
	wire [WIDTH-1:0] wire_d16_76;
	wire [WIDTH-1:0] wire_d16_77;
	wire [WIDTH-1:0] wire_d16_78;
	wire [WIDTH-1:0] wire_d16_79;
	wire [WIDTH-1:0] wire_d16_80;
	wire [WIDTH-1:0] wire_d16_81;
	wire [WIDTH-1:0] wire_d16_82;
	wire [WIDTH-1:0] wire_d16_83;
	wire [WIDTH-1:0] wire_d16_84;
	wire [WIDTH-1:0] wire_d16_85;
	wire [WIDTH-1:0] wire_d16_86;
	wire [WIDTH-1:0] wire_d16_87;
	wire [WIDTH-1:0] wire_d16_88;
	wire [WIDTH-1:0] wire_d16_89;
	wire [WIDTH-1:0] wire_d16_90;
	wire [WIDTH-1:0] wire_d16_91;
	wire [WIDTH-1:0] wire_d16_92;
	wire [WIDTH-1:0] wire_d16_93;
	wire [WIDTH-1:0] wire_d16_94;
	wire [WIDTH-1:0] wire_d16_95;
	wire [WIDTH-1:0] wire_d16_96;
	wire [WIDTH-1:0] wire_d16_97;
	wire [WIDTH-1:0] wire_d16_98;
	wire [WIDTH-1:0] wire_d17_0;
	wire [WIDTH-1:0] wire_d17_1;
	wire [WIDTH-1:0] wire_d17_2;
	wire [WIDTH-1:0] wire_d17_3;
	wire [WIDTH-1:0] wire_d17_4;
	wire [WIDTH-1:0] wire_d17_5;
	wire [WIDTH-1:0] wire_d17_6;
	wire [WIDTH-1:0] wire_d17_7;
	wire [WIDTH-1:0] wire_d17_8;
	wire [WIDTH-1:0] wire_d17_9;
	wire [WIDTH-1:0] wire_d17_10;
	wire [WIDTH-1:0] wire_d17_11;
	wire [WIDTH-1:0] wire_d17_12;
	wire [WIDTH-1:0] wire_d17_13;
	wire [WIDTH-1:0] wire_d17_14;
	wire [WIDTH-1:0] wire_d17_15;
	wire [WIDTH-1:0] wire_d17_16;
	wire [WIDTH-1:0] wire_d17_17;
	wire [WIDTH-1:0] wire_d17_18;
	wire [WIDTH-1:0] wire_d17_19;
	wire [WIDTH-1:0] wire_d17_20;
	wire [WIDTH-1:0] wire_d17_21;
	wire [WIDTH-1:0] wire_d17_22;
	wire [WIDTH-1:0] wire_d17_23;
	wire [WIDTH-1:0] wire_d17_24;
	wire [WIDTH-1:0] wire_d17_25;
	wire [WIDTH-1:0] wire_d17_26;
	wire [WIDTH-1:0] wire_d17_27;
	wire [WIDTH-1:0] wire_d17_28;
	wire [WIDTH-1:0] wire_d17_29;
	wire [WIDTH-1:0] wire_d17_30;
	wire [WIDTH-1:0] wire_d17_31;
	wire [WIDTH-1:0] wire_d17_32;
	wire [WIDTH-1:0] wire_d17_33;
	wire [WIDTH-1:0] wire_d17_34;
	wire [WIDTH-1:0] wire_d17_35;
	wire [WIDTH-1:0] wire_d17_36;
	wire [WIDTH-1:0] wire_d17_37;
	wire [WIDTH-1:0] wire_d17_38;
	wire [WIDTH-1:0] wire_d17_39;
	wire [WIDTH-1:0] wire_d17_40;
	wire [WIDTH-1:0] wire_d17_41;
	wire [WIDTH-1:0] wire_d17_42;
	wire [WIDTH-1:0] wire_d17_43;
	wire [WIDTH-1:0] wire_d17_44;
	wire [WIDTH-1:0] wire_d17_45;
	wire [WIDTH-1:0] wire_d17_46;
	wire [WIDTH-1:0] wire_d17_47;
	wire [WIDTH-1:0] wire_d17_48;
	wire [WIDTH-1:0] wire_d17_49;
	wire [WIDTH-1:0] wire_d17_50;
	wire [WIDTH-1:0] wire_d17_51;
	wire [WIDTH-1:0] wire_d17_52;
	wire [WIDTH-1:0] wire_d17_53;
	wire [WIDTH-1:0] wire_d17_54;
	wire [WIDTH-1:0] wire_d17_55;
	wire [WIDTH-1:0] wire_d17_56;
	wire [WIDTH-1:0] wire_d17_57;
	wire [WIDTH-1:0] wire_d17_58;
	wire [WIDTH-1:0] wire_d17_59;
	wire [WIDTH-1:0] wire_d17_60;
	wire [WIDTH-1:0] wire_d17_61;
	wire [WIDTH-1:0] wire_d17_62;
	wire [WIDTH-1:0] wire_d17_63;
	wire [WIDTH-1:0] wire_d17_64;
	wire [WIDTH-1:0] wire_d17_65;
	wire [WIDTH-1:0] wire_d17_66;
	wire [WIDTH-1:0] wire_d17_67;
	wire [WIDTH-1:0] wire_d17_68;
	wire [WIDTH-1:0] wire_d17_69;
	wire [WIDTH-1:0] wire_d17_70;
	wire [WIDTH-1:0] wire_d17_71;
	wire [WIDTH-1:0] wire_d17_72;
	wire [WIDTH-1:0] wire_d17_73;
	wire [WIDTH-1:0] wire_d17_74;
	wire [WIDTH-1:0] wire_d17_75;
	wire [WIDTH-1:0] wire_d17_76;
	wire [WIDTH-1:0] wire_d17_77;
	wire [WIDTH-1:0] wire_d17_78;
	wire [WIDTH-1:0] wire_d17_79;
	wire [WIDTH-1:0] wire_d17_80;
	wire [WIDTH-1:0] wire_d17_81;
	wire [WIDTH-1:0] wire_d17_82;
	wire [WIDTH-1:0] wire_d17_83;
	wire [WIDTH-1:0] wire_d17_84;
	wire [WIDTH-1:0] wire_d17_85;
	wire [WIDTH-1:0] wire_d17_86;
	wire [WIDTH-1:0] wire_d17_87;
	wire [WIDTH-1:0] wire_d17_88;
	wire [WIDTH-1:0] wire_d17_89;
	wire [WIDTH-1:0] wire_d17_90;
	wire [WIDTH-1:0] wire_d17_91;
	wire [WIDTH-1:0] wire_d17_92;
	wire [WIDTH-1:0] wire_d17_93;
	wire [WIDTH-1:0] wire_d17_94;
	wire [WIDTH-1:0] wire_d17_95;
	wire [WIDTH-1:0] wire_d17_96;
	wire [WIDTH-1:0] wire_d17_97;
	wire [WIDTH-1:0] wire_d17_98;
	wire [WIDTH-1:0] wire_d18_0;
	wire [WIDTH-1:0] wire_d18_1;
	wire [WIDTH-1:0] wire_d18_2;
	wire [WIDTH-1:0] wire_d18_3;
	wire [WIDTH-1:0] wire_d18_4;
	wire [WIDTH-1:0] wire_d18_5;
	wire [WIDTH-1:0] wire_d18_6;
	wire [WIDTH-1:0] wire_d18_7;
	wire [WIDTH-1:0] wire_d18_8;
	wire [WIDTH-1:0] wire_d18_9;
	wire [WIDTH-1:0] wire_d18_10;
	wire [WIDTH-1:0] wire_d18_11;
	wire [WIDTH-1:0] wire_d18_12;
	wire [WIDTH-1:0] wire_d18_13;
	wire [WIDTH-1:0] wire_d18_14;
	wire [WIDTH-1:0] wire_d18_15;
	wire [WIDTH-1:0] wire_d18_16;
	wire [WIDTH-1:0] wire_d18_17;
	wire [WIDTH-1:0] wire_d18_18;
	wire [WIDTH-1:0] wire_d18_19;
	wire [WIDTH-1:0] wire_d18_20;
	wire [WIDTH-1:0] wire_d18_21;
	wire [WIDTH-1:0] wire_d18_22;
	wire [WIDTH-1:0] wire_d18_23;
	wire [WIDTH-1:0] wire_d18_24;
	wire [WIDTH-1:0] wire_d18_25;
	wire [WIDTH-1:0] wire_d18_26;
	wire [WIDTH-1:0] wire_d18_27;
	wire [WIDTH-1:0] wire_d18_28;
	wire [WIDTH-1:0] wire_d18_29;
	wire [WIDTH-1:0] wire_d18_30;
	wire [WIDTH-1:0] wire_d18_31;
	wire [WIDTH-1:0] wire_d18_32;
	wire [WIDTH-1:0] wire_d18_33;
	wire [WIDTH-1:0] wire_d18_34;
	wire [WIDTH-1:0] wire_d18_35;
	wire [WIDTH-1:0] wire_d18_36;
	wire [WIDTH-1:0] wire_d18_37;
	wire [WIDTH-1:0] wire_d18_38;
	wire [WIDTH-1:0] wire_d18_39;
	wire [WIDTH-1:0] wire_d18_40;
	wire [WIDTH-1:0] wire_d18_41;
	wire [WIDTH-1:0] wire_d18_42;
	wire [WIDTH-1:0] wire_d18_43;
	wire [WIDTH-1:0] wire_d18_44;
	wire [WIDTH-1:0] wire_d18_45;
	wire [WIDTH-1:0] wire_d18_46;
	wire [WIDTH-1:0] wire_d18_47;
	wire [WIDTH-1:0] wire_d18_48;
	wire [WIDTH-1:0] wire_d18_49;
	wire [WIDTH-1:0] wire_d18_50;
	wire [WIDTH-1:0] wire_d18_51;
	wire [WIDTH-1:0] wire_d18_52;
	wire [WIDTH-1:0] wire_d18_53;
	wire [WIDTH-1:0] wire_d18_54;
	wire [WIDTH-1:0] wire_d18_55;
	wire [WIDTH-1:0] wire_d18_56;
	wire [WIDTH-1:0] wire_d18_57;
	wire [WIDTH-1:0] wire_d18_58;
	wire [WIDTH-1:0] wire_d18_59;
	wire [WIDTH-1:0] wire_d18_60;
	wire [WIDTH-1:0] wire_d18_61;
	wire [WIDTH-1:0] wire_d18_62;
	wire [WIDTH-1:0] wire_d18_63;
	wire [WIDTH-1:0] wire_d18_64;
	wire [WIDTH-1:0] wire_d18_65;
	wire [WIDTH-1:0] wire_d18_66;
	wire [WIDTH-1:0] wire_d18_67;
	wire [WIDTH-1:0] wire_d18_68;
	wire [WIDTH-1:0] wire_d18_69;
	wire [WIDTH-1:0] wire_d18_70;
	wire [WIDTH-1:0] wire_d18_71;
	wire [WIDTH-1:0] wire_d18_72;
	wire [WIDTH-1:0] wire_d18_73;
	wire [WIDTH-1:0] wire_d18_74;
	wire [WIDTH-1:0] wire_d18_75;
	wire [WIDTH-1:0] wire_d18_76;
	wire [WIDTH-1:0] wire_d18_77;
	wire [WIDTH-1:0] wire_d18_78;
	wire [WIDTH-1:0] wire_d18_79;
	wire [WIDTH-1:0] wire_d18_80;
	wire [WIDTH-1:0] wire_d18_81;
	wire [WIDTH-1:0] wire_d18_82;
	wire [WIDTH-1:0] wire_d18_83;
	wire [WIDTH-1:0] wire_d18_84;
	wire [WIDTH-1:0] wire_d18_85;
	wire [WIDTH-1:0] wire_d18_86;
	wire [WIDTH-1:0] wire_d18_87;
	wire [WIDTH-1:0] wire_d18_88;
	wire [WIDTH-1:0] wire_d18_89;
	wire [WIDTH-1:0] wire_d18_90;
	wire [WIDTH-1:0] wire_d18_91;
	wire [WIDTH-1:0] wire_d18_92;
	wire [WIDTH-1:0] wire_d18_93;
	wire [WIDTH-1:0] wire_d18_94;
	wire [WIDTH-1:0] wire_d18_95;
	wire [WIDTH-1:0] wire_d18_96;
	wire [WIDTH-1:0] wire_d18_97;
	wire [WIDTH-1:0] wire_d18_98;
	wire [WIDTH-1:0] wire_d19_0;
	wire [WIDTH-1:0] wire_d19_1;
	wire [WIDTH-1:0] wire_d19_2;
	wire [WIDTH-1:0] wire_d19_3;
	wire [WIDTH-1:0] wire_d19_4;
	wire [WIDTH-1:0] wire_d19_5;
	wire [WIDTH-1:0] wire_d19_6;
	wire [WIDTH-1:0] wire_d19_7;
	wire [WIDTH-1:0] wire_d19_8;
	wire [WIDTH-1:0] wire_d19_9;
	wire [WIDTH-1:0] wire_d19_10;
	wire [WIDTH-1:0] wire_d19_11;
	wire [WIDTH-1:0] wire_d19_12;
	wire [WIDTH-1:0] wire_d19_13;
	wire [WIDTH-1:0] wire_d19_14;
	wire [WIDTH-1:0] wire_d19_15;
	wire [WIDTH-1:0] wire_d19_16;
	wire [WIDTH-1:0] wire_d19_17;
	wire [WIDTH-1:0] wire_d19_18;
	wire [WIDTH-1:0] wire_d19_19;
	wire [WIDTH-1:0] wire_d19_20;
	wire [WIDTH-1:0] wire_d19_21;
	wire [WIDTH-1:0] wire_d19_22;
	wire [WIDTH-1:0] wire_d19_23;
	wire [WIDTH-1:0] wire_d19_24;
	wire [WIDTH-1:0] wire_d19_25;
	wire [WIDTH-1:0] wire_d19_26;
	wire [WIDTH-1:0] wire_d19_27;
	wire [WIDTH-1:0] wire_d19_28;
	wire [WIDTH-1:0] wire_d19_29;
	wire [WIDTH-1:0] wire_d19_30;
	wire [WIDTH-1:0] wire_d19_31;
	wire [WIDTH-1:0] wire_d19_32;
	wire [WIDTH-1:0] wire_d19_33;
	wire [WIDTH-1:0] wire_d19_34;
	wire [WIDTH-1:0] wire_d19_35;
	wire [WIDTH-1:0] wire_d19_36;
	wire [WIDTH-1:0] wire_d19_37;
	wire [WIDTH-1:0] wire_d19_38;
	wire [WIDTH-1:0] wire_d19_39;
	wire [WIDTH-1:0] wire_d19_40;
	wire [WIDTH-1:0] wire_d19_41;
	wire [WIDTH-1:0] wire_d19_42;
	wire [WIDTH-1:0] wire_d19_43;
	wire [WIDTH-1:0] wire_d19_44;
	wire [WIDTH-1:0] wire_d19_45;
	wire [WIDTH-1:0] wire_d19_46;
	wire [WIDTH-1:0] wire_d19_47;
	wire [WIDTH-1:0] wire_d19_48;
	wire [WIDTH-1:0] wire_d19_49;
	wire [WIDTH-1:0] wire_d19_50;
	wire [WIDTH-1:0] wire_d19_51;
	wire [WIDTH-1:0] wire_d19_52;
	wire [WIDTH-1:0] wire_d19_53;
	wire [WIDTH-1:0] wire_d19_54;
	wire [WIDTH-1:0] wire_d19_55;
	wire [WIDTH-1:0] wire_d19_56;
	wire [WIDTH-1:0] wire_d19_57;
	wire [WIDTH-1:0] wire_d19_58;
	wire [WIDTH-1:0] wire_d19_59;
	wire [WIDTH-1:0] wire_d19_60;
	wire [WIDTH-1:0] wire_d19_61;
	wire [WIDTH-1:0] wire_d19_62;
	wire [WIDTH-1:0] wire_d19_63;
	wire [WIDTH-1:0] wire_d19_64;
	wire [WIDTH-1:0] wire_d19_65;
	wire [WIDTH-1:0] wire_d19_66;
	wire [WIDTH-1:0] wire_d19_67;
	wire [WIDTH-1:0] wire_d19_68;
	wire [WIDTH-1:0] wire_d19_69;
	wire [WIDTH-1:0] wire_d19_70;
	wire [WIDTH-1:0] wire_d19_71;
	wire [WIDTH-1:0] wire_d19_72;
	wire [WIDTH-1:0] wire_d19_73;
	wire [WIDTH-1:0] wire_d19_74;
	wire [WIDTH-1:0] wire_d19_75;
	wire [WIDTH-1:0] wire_d19_76;
	wire [WIDTH-1:0] wire_d19_77;
	wire [WIDTH-1:0] wire_d19_78;
	wire [WIDTH-1:0] wire_d19_79;
	wire [WIDTH-1:0] wire_d19_80;
	wire [WIDTH-1:0] wire_d19_81;
	wire [WIDTH-1:0] wire_d19_82;
	wire [WIDTH-1:0] wire_d19_83;
	wire [WIDTH-1:0] wire_d19_84;
	wire [WIDTH-1:0] wire_d19_85;
	wire [WIDTH-1:0] wire_d19_86;
	wire [WIDTH-1:0] wire_d19_87;
	wire [WIDTH-1:0] wire_d19_88;
	wire [WIDTH-1:0] wire_d19_89;
	wire [WIDTH-1:0] wire_d19_90;
	wire [WIDTH-1:0] wire_d19_91;
	wire [WIDTH-1:0] wire_d19_92;
	wire [WIDTH-1:0] wire_d19_93;
	wire [WIDTH-1:0] wire_d19_94;
	wire [WIDTH-1:0] wire_d19_95;
	wire [WIDTH-1:0] wire_d19_96;
	wire [WIDTH-1:0] wire_d19_97;
	wire [WIDTH-1:0] wire_d19_98;
	wire [WIDTH-1:0] wire_d20_0;
	wire [WIDTH-1:0] wire_d20_1;
	wire [WIDTH-1:0] wire_d20_2;
	wire [WIDTH-1:0] wire_d20_3;
	wire [WIDTH-1:0] wire_d20_4;
	wire [WIDTH-1:0] wire_d20_5;
	wire [WIDTH-1:0] wire_d20_6;
	wire [WIDTH-1:0] wire_d20_7;
	wire [WIDTH-1:0] wire_d20_8;
	wire [WIDTH-1:0] wire_d20_9;
	wire [WIDTH-1:0] wire_d20_10;
	wire [WIDTH-1:0] wire_d20_11;
	wire [WIDTH-1:0] wire_d20_12;
	wire [WIDTH-1:0] wire_d20_13;
	wire [WIDTH-1:0] wire_d20_14;
	wire [WIDTH-1:0] wire_d20_15;
	wire [WIDTH-1:0] wire_d20_16;
	wire [WIDTH-1:0] wire_d20_17;
	wire [WIDTH-1:0] wire_d20_18;
	wire [WIDTH-1:0] wire_d20_19;
	wire [WIDTH-1:0] wire_d20_20;
	wire [WIDTH-1:0] wire_d20_21;
	wire [WIDTH-1:0] wire_d20_22;
	wire [WIDTH-1:0] wire_d20_23;
	wire [WIDTH-1:0] wire_d20_24;
	wire [WIDTH-1:0] wire_d20_25;
	wire [WIDTH-1:0] wire_d20_26;
	wire [WIDTH-1:0] wire_d20_27;
	wire [WIDTH-1:0] wire_d20_28;
	wire [WIDTH-1:0] wire_d20_29;
	wire [WIDTH-1:0] wire_d20_30;
	wire [WIDTH-1:0] wire_d20_31;
	wire [WIDTH-1:0] wire_d20_32;
	wire [WIDTH-1:0] wire_d20_33;
	wire [WIDTH-1:0] wire_d20_34;
	wire [WIDTH-1:0] wire_d20_35;
	wire [WIDTH-1:0] wire_d20_36;
	wire [WIDTH-1:0] wire_d20_37;
	wire [WIDTH-1:0] wire_d20_38;
	wire [WIDTH-1:0] wire_d20_39;
	wire [WIDTH-1:0] wire_d20_40;
	wire [WIDTH-1:0] wire_d20_41;
	wire [WIDTH-1:0] wire_d20_42;
	wire [WIDTH-1:0] wire_d20_43;
	wire [WIDTH-1:0] wire_d20_44;
	wire [WIDTH-1:0] wire_d20_45;
	wire [WIDTH-1:0] wire_d20_46;
	wire [WIDTH-1:0] wire_d20_47;
	wire [WIDTH-1:0] wire_d20_48;
	wire [WIDTH-1:0] wire_d20_49;
	wire [WIDTH-1:0] wire_d20_50;
	wire [WIDTH-1:0] wire_d20_51;
	wire [WIDTH-1:0] wire_d20_52;
	wire [WIDTH-1:0] wire_d20_53;
	wire [WIDTH-1:0] wire_d20_54;
	wire [WIDTH-1:0] wire_d20_55;
	wire [WIDTH-1:0] wire_d20_56;
	wire [WIDTH-1:0] wire_d20_57;
	wire [WIDTH-1:0] wire_d20_58;
	wire [WIDTH-1:0] wire_d20_59;
	wire [WIDTH-1:0] wire_d20_60;
	wire [WIDTH-1:0] wire_d20_61;
	wire [WIDTH-1:0] wire_d20_62;
	wire [WIDTH-1:0] wire_d20_63;
	wire [WIDTH-1:0] wire_d20_64;
	wire [WIDTH-1:0] wire_d20_65;
	wire [WIDTH-1:0] wire_d20_66;
	wire [WIDTH-1:0] wire_d20_67;
	wire [WIDTH-1:0] wire_d20_68;
	wire [WIDTH-1:0] wire_d20_69;
	wire [WIDTH-1:0] wire_d20_70;
	wire [WIDTH-1:0] wire_d20_71;
	wire [WIDTH-1:0] wire_d20_72;
	wire [WIDTH-1:0] wire_d20_73;
	wire [WIDTH-1:0] wire_d20_74;
	wire [WIDTH-1:0] wire_d20_75;
	wire [WIDTH-1:0] wire_d20_76;
	wire [WIDTH-1:0] wire_d20_77;
	wire [WIDTH-1:0] wire_d20_78;
	wire [WIDTH-1:0] wire_d20_79;
	wire [WIDTH-1:0] wire_d20_80;
	wire [WIDTH-1:0] wire_d20_81;
	wire [WIDTH-1:0] wire_d20_82;
	wire [WIDTH-1:0] wire_d20_83;
	wire [WIDTH-1:0] wire_d20_84;
	wire [WIDTH-1:0] wire_d20_85;
	wire [WIDTH-1:0] wire_d20_86;
	wire [WIDTH-1:0] wire_d20_87;
	wire [WIDTH-1:0] wire_d20_88;
	wire [WIDTH-1:0] wire_d20_89;
	wire [WIDTH-1:0] wire_d20_90;
	wire [WIDTH-1:0] wire_d20_91;
	wire [WIDTH-1:0] wire_d20_92;
	wire [WIDTH-1:0] wire_d20_93;
	wire [WIDTH-1:0] wire_d20_94;
	wire [WIDTH-1:0] wire_d20_95;
	wire [WIDTH-1:0] wire_d20_96;
	wire [WIDTH-1:0] wire_d20_97;
	wire [WIDTH-1:0] wire_d20_98;
	wire [WIDTH-1:0] wire_d21_0;
	wire [WIDTH-1:0] wire_d21_1;
	wire [WIDTH-1:0] wire_d21_2;
	wire [WIDTH-1:0] wire_d21_3;
	wire [WIDTH-1:0] wire_d21_4;
	wire [WIDTH-1:0] wire_d21_5;
	wire [WIDTH-1:0] wire_d21_6;
	wire [WIDTH-1:0] wire_d21_7;
	wire [WIDTH-1:0] wire_d21_8;
	wire [WIDTH-1:0] wire_d21_9;
	wire [WIDTH-1:0] wire_d21_10;
	wire [WIDTH-1:0] wire_d21_11;
	wire [WIDTH-1:0] wire_d21_12;
	wire [WIDTH-1:0] wire_d21_13;
	wire [WIDTH-1:0] wire_d21_14;
	wire [WIDTH-1:0] wire_d21_15;
	wire [WIDTH-1:0] wire_d21_16;
	wire [WIDTH-1:0] wire_d21_17;
	wire [WIDTH-1:0] wire_d21_18;
	wire [WIDTH-1:0] wire_d21_19;
	wire [WIDTH-1:0] wire_d21_20;
	wire [WIDTH-1:0] wire_d21_21;
	wire [WIDTH-1:0] wire_d21_22;
	wire [WIDTH-1:0] wire_d21_23;
	wire [WIDTH-1:0] wire_d21_24;
	wire [WIDTH-1:0] wire_d21_25;
	wire [WIDTH-1:0] wire_d21_26;
	wire [WIDTH-1:0] wire_d21_27;
	wire [WIDTH-1:0] wire_d21_28;
	wire [WIDTH-1:0] wire_d21_29;
	wire [WIDTH-1:0] wire_d21_30;
	wire [WIDTH-1:0] wire_d21_31;
	wire [WIDTH-1:0] wire_d21_32;
	wire [WIDTH-1:0] wire_d21_33;
	wire [WIDTH-1:0] wire_d21_34;
	wire [WIDTH-1:0] wire_d21_35;
	wire [WIDTH-1:0] wire_d21_36;
	wire [WIDTH-1:0] wire_d21_37;
	wire [WIDTH-1:0] wire_d21_38;
	wire [WIDTH-1:0] wire_d21_39;
	wire [WIDTH-1:0] wire_d21_40;
	wire [WIDTH-1:0] wire_d21_41;
	wire [WIDTH-1:0] wire_d21_42;
	wire [WIDTH-1:0] wire_d21_43;
	wire [WIDTH-1:0] wire_d21_44;
	wire [WIDTH-1:0] wire_d21_45;
	wire [WIDTH-1:0] wire_d21_46;
	wire [WIDTH-1:0] wire_d21_47;
	wire [WIDTH-1:0] wire_d21_48;
	wire [WIDTH-1:0] wire_d21_49;
	wire [WIDTH-1:0] wire_d21_50;
	wire [WIDTH-1:0] wire_d21_51;
	wire [WIDTH-1:0] wire_d21_52;
	wire [WIDTH-1:0] wire_d21_53;
	wire [WIDTH-1:0] wire_d21_54;
	wire [WIDTH-1:0] wire_d21_55;
	wire [WIDTH-1:0] wire_d21_56;
	wire [WIDTH-1:0] wire_d21_57;
	wire [WIDTH-1:0] wire_d21_58;
	wire [WIDTH-1:0] wire_d21_59;
	wire [WIDTH-1:0] wire_d21_60;
	wire [WIDTH-1:0] wire_d21_61;
	wire [WIDTH-1:0] wire_d21_62;
	wire [WIDTH-1:0] wire_d21_63;
	wire [WIDTH-1:0] wire_d21_64;
	wire [WIDTH-1:0] wire_d21_65;
	wire [WIDTH-1:0] wire_d21_66;
	wire [WIDTH-1:0] wire_d21_67;
	wire [WIDTH-1:0] wire_d21_68;
	wire [WIDTH-1:0] wire_d21_69;
	wire [WIDTH-1:0] wire_d21_70;
	wire [WIDTH-1:0] wire_d21_71;
	wire [WIDTH-1:0] wire_d21_72;
	wire [WIDTH-1:0] wire_d21_73;
	wire [WIDTH-1:0] wire_d21_74;
	wire [WIDTH-1:0] wire_d21_75;
	wire [WIDTH-1:0] wire_d21_76;
	wire [WIDTH-1:0] wire_d21_77;
	wire [WIDTH-1:0] wire_d21_78;
	wire [WIDTH-1:0] wire_d21_79;
	wire [WIDTH-1:0] wire_d21_80;
	wire [WIDTH-1:0] wire_d21_81;
	wire [WIDTH-1:0] wire_d21_82;
	wire [WIDTH-1:0] wire_d21_83;
	wire [WIDTH-1:0] wire_d21_84;
	wire [WIDTH-1:0] wire_d21_85;
	wire [WIDTH-1:0] wire_d21_86;
	wire [WIDTH-1:0] wire_d21_87;
	wire [WIDTH-1:0] wire_d21_88;
	wire [WIDTH-1:0] wire_d21_89;
	wire [WIDTH-1:0] wire_d21_90;
	wire [WIDTH-1:0] wire_d21_91;
	wire [WIDTH-1:0] wire_d21_92;
	wire [WIDTH-1:0] wire_d21_93;
	wire [WIDTH-1:0] wire_d21_94;
	wire [WIDTH-1:0] wire_d21_95;
	wire [WIDTH-1:0] wire_d21_96;
	wire [WIDTH-1:0] wire_d21_97;
	wire [WIDTH-1:0] wire_d21_98;
	wire [WIDTH-1:0] wire_d22_0;
	wire [WIDTH-1:0] wire_d22_1;
	wire [WIDTH-1:0] wire_d22_2;
	wire [WIDTH-1:0] wire_d22_3;
	wire [WIDTH-1:0] wire_d22_4;
	wire [WIDTH-1:0] wire_d22_5;
	wire [WIDTH-1:0] wire_d22_6;
	wire [WIDTH-1:0] wire_d22_7;
	wire [WIDTH-1:0] wire_d22_8;
	wire [WIDTH-1:0] wire_d22_9;
	wire [WIDTH-1:0] wire_d22_10;
	wire [WIDTH-1:0] wire_d22_11;
	wire [WIDTH-1:0] wire_d22_12;
	wire [WIDTH-1:0] wire_d22_13;
	wire [WIDTH-1:0] wire_d22_14;
	wire [WIDTH-1:0] wire_d22_15;
	wire [WIDTH-1:0] wire_d22_16;
	wire [WIDTH-1:0] wire_d22_17;
	wire [WIDTH-1:0] wire_d22_18;
	wire [WIDTH-1:0] wire_d22_19;
	wire [WIDTH-1:0] wire_d22_20;
	wire [WIDTH-1:0] wire_d22_21;
	wire [WIDTH-1:0] wire_d22_22;
	wire [WIDTH-1:0] wire_d22_23;
	wire [WIDTH-1:0] wire_d22_24;
	wire [WIDTH-1:0] wire_d22_25;
	wire [WIDTH-1:0] wire_d22_26;
	wire [WIDTH-1:0] wire_d22_27;
	wire [WIDTH-1:0] wire_d22_28;
	wire [WIDTH-1:0] wire_d22_29;
	wire [WIDTH-1:0] wire_d22_30;
	wire [WIDTH-1:0] wire_d22_31;
	wire [WIDTH-1:0] wire_d22_32;
	wire [WIDTH-1:0] wire_d22_33;
	wire [WIDTH-1:0] wire_d22_34;
	wire [WIDTH-1:0] wire_d22_35;
	wire [WIDTH-1:0] wire_d22_36;
	wire [WIDTH-1:0] wire_d22_37;
	wire [WIDTH-1:0] wire_d22_38;
	wire [WIDTH-1:0] wire_d22_39;
	wire [WIDTH-1:0] wire_d22_40;
	wire [WIDTH-1:0] wire_d22_41;
	wire [WIDTH-1:0] wire_d22_42;
	wire [WIDTH-1:0] wire_d22_43;
	wire [WIDTH-1:0] wire_d22_44;
	wire [WIDTH-1:0] wire_d22_45;
	wire [WIDTH-1:0] wire_d22_46;
	wire [WIDTH-1:0] wire_d22_47;
	wire [WIDTH-1:0] wire_d22_48;
	wire [WIDTH-1:0] wire_d22_49;
	wire [WIDTH-1:0] wire_d22_50;
	wire [WIDTH-1:0] wire_d22_51;
	wire [WIDTH-1:0] wire_d22_52;
	wire [WIDTH-1:0] wire_d22_53;
	wire [WIDTH-1:0] wire_d22_54;
	wire [WIDTH-1:0] wire_d22_55;
	wire [WIDTH-1:0] wire_d22_56;
	wire [WIDTH-1:0] wire_d22_57;
	wire [WIDTH-1:0] wire_d22_58;
	wire [WIDTH-1:0] wire_d22_59;
	wire [WIDTH-1:0] wire_d22_60;
	wire [WIDTH-1:0] wire_d22_61;
	wire [WIDTH-1:0] wire_d22_62;
	wire [WIDTH-1:0] wire_d22_63;
	wire [WIDTH-1:0] wire_d22_64;
	wire [WIDTH-1:0] wire_d22_65;
	wire [WIDTH-1:0] wire_d22_66;
	wire [WIDTH-1:0] wire_d22_67;
	wire [WIDTH-1:0] wire_d22_68;
	wire [WIDTH-1:0] wire_d22_69;
	wire [WIDTH-1:0] wire_d22_70;
	wire [WIDTH-1:0] wire_d22_71;
	wire [WIDTH-1:0] wire_d22_72;
	wire [WIDTH-1:0] wire_d22_73;
	wire [WIDTH-1:0] wire_d22_74;
	wire [WIDTH-1:0] wire_d22_75;
	wire [WIDTH-1:0] wire_d22_76;
	wire [WIDTH-1:0] wire_d22_77;
	wire [WIDTH-1:0] wire_d22_78;
	wire [WIDTH-1:0] wire_d22_79;
	wire [WIDTH-1:0] wire_d22_80;
	wire [WIDTH-1:0] wire_d22_81;
	wire [WIDTH-1:0] wire_d22_82;
	wire [WIDTH-1:0] wire_d22_83;
	wire [WIDTH-1:0] wire_d22_84;
	wire [WIDTH-1:0] wire_d22_85;
	wire [WIDTH-1:0] wire_d22_86;
	wire [WIDTH-1:0] wire_d22_87;
	wire [WIDTH-1:0] wire_d22_88;
	wire [WIDTH-1:0] wire_d22_89;
	wire [WIDTH-1:0] wire_d22_90;
	wire [WIDTH-1:0] wire_d22_91;
	wire [WIDTH-1:0] wire_d22_92;
	wire [WIDTH-1:0] wire_d22_93;
	wire [WIDTH-1:0] wire_d22_94;
	wire [WIDTH-1:0] wire_d22_95;
	wire [WIDTH-1:0] wire_d22_96;
	wire [WIDTH-1:0] wire_d22_97;
	wire [WIDTH-1:0] wire_d22_98;
	wire [WIDTH-1:0] wire_d23_0;
	wire [WIDTH-1:0] wire_d23_1;
	wire [WIDTH-1:0] wire_d23_2;
	wire [WIDTH-1:0] wire_d23_3;
	wire [WIDTH-1:0] wire_d23_4;
	wire [WIDTH-1:0] wire_d23_5;
	wire [WIDTH-1:0] wire_d23_6;
	wire [WIDTH-1:0] wire_d23_7;
	wire [WIDTH-1:0] wire_d23_8;
	wire [WIDTH-1:0] wire_d23_9;
	wire [WIDTH-1:0] wire_d23_10;
	wire [WIDTH-1:0] wire_d23_11;
	wire [WIDTH-1:0] wire_d23_12;
	wire [WIDTH-1:0] wire_d23_13;
	wire [WIDTH-1:0] wire_d23_14;
	wire [WIDTH-1:0] wire_d23_15;
	wire [WIDTH-1:0] wire_d23_16;
	wire [WIDTH-1:0] wire_d23_17;
	wire [WIDTH-1:0] wire_d23_18;
	wire [WIDTH-1:0] wire_d23_19;
	wire [WIDTH-1:0] wire_d23_20;
	wire [WIDTH-1:0] wire_d23_21;
	wire [WIDTH-1:0] wire_d23_22;
	wire [WIDTH-1:0] wire_d23_23;
	wire [WIDTH-1:0] wire_d23_24;
	wire [WIDTH-1:0] wire_d23_25;
	wire [WIDTH-1:0] wire_d23_26;
	wire [WIDTH-1:0] wire_d23_27;
	wire [WIDTH-1:0] wire_d23_28;
	wire [WIDTH-1:0] wire_d23_29;
	wire [WIDTH-1:0] wire_d23_30;
	wire [WIDTH-1:0] wire_d23_31;
	wire [WIDTH-1:0] wire_d23_32;
	wire [WIDTH-1:0] wire_d23_33;
	wire [WIDTH-1:0] wire_d23_34;
	wire [WIDTH-1:0] wire_d23_35;
	wire [WIDTH-1:0] wire_d23_36;
	wire [WIDTH-1:0] wire_d23_37;
	wire [WIDTH-1:0] wire_d23_38;
	wire [WIDTH-1:0] wire_d23_39;
	wire [WIDTH-1:0] wire_d23_40;
	wire [WIDTH-1:0] wire_d23_41;
	wire [WIDTH-1:0] wire_d23_42;
	wire [WIDTH-1:0] wire_d23_43;
	wire [WIDTH-1:0] wire_d23_44;
	wire [WIDTH-1:0] wire_d23_45;
	wire [WIDTH-1:0] wire_d23_46;
	wire [WIDTH-1:0] wire_d23_47;
	wire [WIDTH-1:0] wire_d23_48;
	wire [WIDTH-1:0] wire_d23_49;
	wire [WIDTH-1:0] wire_d23_50;
	wire [WIDTH-1:0] wire_d23_51;
	wire [WIDTH-1:0] wire_d23_52;
	wire [WIDTH-1:0] wire_d23_53;
	wire [WIDTH-1:0] wire_d23_54;
	wire [WIDTH-1:0] wire_d23_55;
	wire [WIDTH-1:0] wire_d23_56;
	wire [WIDTH-1:0] wire_d23_57;
	wire [WIDTH-1:0] wire_d23_58;
	wire [WIDTH-1:0] wire_d23_59;
	wire [WIDTH-1:0] wire_d23_60;
	wire [WIDTH-1:0] wire_d23_61;
	wire [WIDTH-1:0] wire_d23_62;
	wire [WIDTH-1:0] wire_d23_63;
	wire [WIDTH-1:0] wire_d23_64;
	wire [WIDTH-1:0] wire_d23_65;
	wire [WIDTH-1:0] wire_d23_66;
	wire [WIDTH-1:0] wire_d23_67;
	wire [WIDTH-1:0] wire_d23_68;
	wire [WIDTH-1:0] wire_d23_69;
	wire [WIDTH-1:0] wire_d23_70;
	wire [WIDTH-1:0] wire_d23_71;
	wire [WIDTH-1:0] wire_d23_72;
	wire [WIDTH-1:0] wire_d23_73;
	wire [WIDTH-1:0] wire_d23_74;
	wire [WIDTH-1:0] wire_d23_75;
	wire [WIDTH-1:0] wire_d23_76;
	wire [WIDTH-1:0] wire_d23_77;
	wire [WIDTH-1:0] wire_d23_78;
	wire [WIDTH-1:0] wire_d23_79;
	wire [WIDTH-1:0] wire_d23_80;
	wire [WIDTH-1:0] wire_d23_81;
	wire [WIDTH-1:0] wire_d23_82;
	wire [WIDTH-1:0] wire_d23_83;
	wire [WIDTH-1:0] wire_d23_84;
	wire [WIDTH-1:0] wire_d23_85;
	wire [WIDTH-1:0] wire_d23_86;
	wire [WIDTH-1:0] wire_d23_87;
	wire [WIDTH-1:0] wire_d23_88;
	wire [WIDTH-1:0] wire_d23_89;
	wire [WIDTH-1:0] wire_d23_90;
	wire [WIDTH-1:0] wire_d23_91;
	wire [WIDTH-1:0] wire_d23_92;
	wire [WIDTH-1:0] wire_d23_93;
	wire [WIDTH-1:0] wire_d23_94;
	wire [WIDTH-1:0] wire_d23_95;
	wire [WIDTH-1:0] wire_d23_96;
	wire [WIDTH-1:0] wire_d23_97;
	wire [WIDTH-1:0] wire_d23_98;
	wire [WIDTH-1:0] wire_d24_0;
	wire [WIDTH-1:0] wire_d24_1;
	wire [WIDTH-1:0] wire_d24_2;
	wire [WIDTH-1:0] wire_d24_3;
	wire [WIDTH-1:0] wire_d24_4;
	wire [WIDTH-1:0] wire_d24_5;
	wire [WIDTH-1:0] wire_d24_6;
	wire [WIDTH-1:0] wire_d24_7;
	wire [WIDTH-1:0] wire_d24_8;
	wire [WIDTH-1:0] wire_d24_9;
	wire [WIDTH-1:0] wire_d24_10;
	wire [WIDTH-1:0] wire_d24_11;
	wire [WIDTH-1:0] wire_d24_12;
	wire [WIDTH-1:0] wire_d24_13;
	wire [WIDTH-1:0] wire_d24_14;
	wire [WIDTH-1:0] wire_d24_15;
	wire [WIDTH-1:0] wire_d24_16;
	wire [WIDTH-1:0] wire_d24_17;
	wire [WIDTH-1:0] wire_d24_18;
	wire [WIDTH-1:0] wire_d24_19;
	wire [WIDTH-1:0] wire_d24_20;
	wire [WIDTH-1:0] wire_d24_21;
	wire [WIDTH-1:0] wire_d24_22;
	wire [WIDTH-1:0] wire_d24_23;
	wire [WIDTH-1:0] wire_d24_24;
	wire [WIDTH-1:0] wire_d24_25;
	wire [WIDTH-1:0] wire_d24_26;
	wire [WIDTH-1:0] wire_d24_27;
	wire [WIDTH-1:0] wire_d24_28;
	wire [WIDTH-1:0] wire_d24_29;
	wire [WIDTH-1:0] wire_d24_30;
	wire [WIDTH-1:0] wire_d24_31;
	wire [WIDTH-1:0] wire_d24_32;
	wire [WIDTH-1:0] wire_d24_33;
	wire [WIDTH-1:0] wire_d24_34;
	wire [WIDTH-1:0] wire_d24_35;
	wire [WIDTH-1:0] wire_d24_36;
	wire [WIDTH-1:0] wire_d24_37;
	wire [WIDTH-1:0] wire_d24_38;
	wire [WIDTH-1:0] wire_d24_39;
	wire [WIDTH-1:0] wire_d24_40;
	wire [WIDTH-1:0] wire_d24_41;
	wire [WIDTH-1:0] wire_d24_42;
	wire [WIDTH-1:0] wire_d24_43;
	wire [WIDTH-1:0] wire_d24_44;
	wire [WIDTH-1:0] wire_d24_45;
	wire [WIDTH-1:0] wire_d24_46;
	wire [WIDTH-1:0] wire_d24_47;
	wire [WIDTH-1:0] wire_d24_48;
	wire [WIDTH-1:0] wire_d24_49;
	wire [WIDTH-1:0] wire_d24_50;
	wire [WIDTH-1:0] wire_d24_51;
	wire [WIDTH-1:0] wire_d24_52;
	wire [WIDTH-1:0] wire_d24_53;
	wire [WIDTH-1:0] wire_d24_54;
	wire [WIDTH-1:0] wire_d24_55;
	wire [WIDTH-1:0] wire_d24_56;
	wire [WIDTH-1:0] wire_d24_57;
	wire [WIDTH-1:0] wire_d24_58;
	wire [WIDTH-1:0] wire_d24_59;
	wire [WIDTH-1:0] wire_d24_60;
	wire [WIDTH-1:0] wire_d24_61;
	wire [WIDTH-1:0] wire_d24_62;
	wire [WIDTH-1:0] wire_d24_63;
	wire [WIDTH-1:0] wire_d24_64;
	wire [WIDTH-1:0] wire_d24_65;
	wire [WIDTH-1:0] wire_d24_66;
	wire [WIDTH-1:0] wire_d24_67;
	wire [WIDTH-1:0] wire_d24_68;
	wire [WIDTH-1:0] wire_d24_69;
	wire [WIDTH-1:0] wire_d24_70;
	wire [WIDTH-1:0] wire_d24_71;
	wire [WIDTH-1:0] wire_d24_72;
	wire [WIDTH-1:0] wire_d24_73;
	wire [WIDTH-1:0] wire_d24_74;
	wire [WIDTH-1:0] wire_d24_75;
	wire [WIDTH-1:0] wire_d24_76;
	wire [WIDTH-1:0] wire_d24_77;
	wire [WIDTH-1:0] wire_d24_78;
	wire [WIDTH-1:0] wire_d24_79;
	wire [WIDTH-1:0] wire_d24_80;
	wire [WIDTH-1:0] wire_d24_81;
	wire [WIDTH-1:0] wire_d24_82;
	wire [WIDTH-1:0] wire_d24_83;
	wire [WIDTH-1:0] wire_d24_84;
	wire [WIDTH-1:0] wire_d24_85;
	wire [WIDTH-1:0] wire_d24_86;
	wire [WIDTH-1:0] wire_d24_87;
	wire [WIDTH-1:0] wire_d24_88;
	wire [WIDTH-1:0] wire_d24_89;
	wire [WIDTH-1:0] wire_d24_90;
	wire [WIDTH-1:0] wire_d24_91;
	wire [WIDTH-1:0] wire_d24_92;
	wire [WIDTH-1:0] wire_d24_93;
	wire [WIDTH-1:0] wire_d24_94;
	wire [WIDTH-1:0] wire_d24_95;
	wire [WIDTH-1:0] wire_d24_96;
	wire [WIDTH-1:0] wire_d24_97;
	wire [WIDTH-1:0] wire_d24_98;
	wire [WIDTH-1:0] wire_d25_0;
	wire [WIDTH-1:0] wire_d25_1;
	wire [WIDTH-1:0] wire_d25_2;
	wire [WIDTH-1:0] wire_d25_3;
	wire [WIDTH-1:0] wire_d25_4;
	wire [WIDTH-1:0] wire_d25_5;
	wire [WIDTH-1:0] wire_d25_6;
	wire [WIDTH-1:0] wire_d25_7;
	wire [WIDTH-1:0] wire_d25_8;
	wire [WIDTH-1:0] wire_d25_9;
	wire [WIDTH-1:0] wire_d25_10;
	wire [WIDTH-1:0] wire_d25_11;
	wire [WIDTH-1:0] wire_d25_12;
	wire [WIDTH-1:0] wire_d25_13;
	wire [WIDTH-1:0] wire_d25_14;
	wire [WIDTH-1:0] wire_d25_15;
	wire [WIDTH-1:0] wire_d25_16;
	wire [WIDTH-1:0] wire_d25_17;
	wire [WIDTH-1:0] wire_d25_18;
	wire [WIDTH-1:0] wire_d25_19;
	wire [WIDTH-1:0] wire_d25_20;
	wire [WIDTH-1:0] wire_d25_21;
	wire [WIDTH-1:0] wire_d25_22;
	wire [WIDTH-1:0] wire_d25_23;
	wire [WIDTH-1:0] wire_d25_24;
	wire [WIDTH-1:0] wire_d25_25;
	wire [WIDTH-1:0] wire_d25_26;
	wire [WIDTH-1:0] wire_d25_27;
	wire [WIDTH-1:0] wire_d25_28;
	wire [WIDTH-1:0] wire_d25_29;
	wire [WIDTH-1:0] wire_d25_30;
	wire [WIDTH-1:0] wire_d25_31;
	wire [WIDTH-1:0] wire_d25_32;
	wire [WIDTH-1:0] wire_d25_33;
	wire [WIDTH-1:0] wire_d25_34;
	wire [WIDTH-1:0] wire_d25_35;
	wire [WIDTH-1:0] wire_d25_36;
	wire [WIDTH-1:0] wire_d25_37;
	wire [WIDTH-1:0] wire_d25_38;
	wire [WIDTH-1:0] wire_d25_39;
	wire [WIDTH-1:0] wire_d25_40;
	wire [WIDTH-1:0] wire_d25_41;
	wire [WIDTH-1:0] wire_d25_42;
	wire [WIDTH-1:0] wire_d25_43;
	wire [WIDTH-1:0] wire_d25_44;
	wire [WIDTH-1:0] wire_d25_45;
	wire [WIDTH-1:0] wire_d25_46;
	wire [WIDTH-1:0] wire_d25_47;
	wire [WIDTH-1:0] wire_d25_48;
	wire [WIDTH-1:0] wire_d25_49;
	wire [WIDTH-1:0] wire_d25_50;
	wire [WIDTH-1:0] wire_d25_51;
	wire [WIDTH-1:0] wire_d25_52;
	wire [WIDTH-1:0] wire_d25_53;
	wire [WIDTH-1:0] wire_d25_54;
	wire [WIDTH-1:0] wire_d25_55;
	wire [WIDTH-1:0] wire_d25_56;
	wire [WIDTH-1:0] wire_d25_57;
	wire [WIDTH-1:0] wire_d25_58;
	wire [WIDTH-1:0] wire_d25_59;
	wire [WIDTH-1:0] wire_d25_60;
	wire [WIDTH-1:0] wire_d25_61;
	wire [WIDTH-1:0] wire_d25_62;
	wire [WIDTH-1:0] wire_d25_63;
	wire [WIDTH-1:0] wire_d25_64;
	wire [WIDTH-1:0] wire_d25_65;
	wire [WIDTH-1:0] wire_d25_66;
	wire [WIDTH-1:0] wire_d25_67;
	wire [WIDTH-1:0] wire_d25_68;
	wire [WIDTH-1:0] wire_d25_69;
	wire [WIDTH-1:0] wire_d25_70;
	wire [WIDTH-1:0] wire_d25_71;
	wire [WIDTH-1:0] wire_d25_72;
	wire [WIDTH-1:0] wire_d25_73;
	wire [WIDTH-1:0] wire_d25_74;
	wire [WIDTH-1:0] wire_d25_75;
	wire [WIDTH-1:0] wire_d25_76;
	wire [WIDTH-1:0] wire_d25_77;
	wire [WIDTH-1:0] wire_d25_78;
	wire [WIDTH-1:0] wire_d25_79;
	wire [WIDTH-1:0] wire_d25_80;
	wire [WIDTH-1:0] wire_d25_81;
	wire [WIDTH-1:0] wire_d25_82;
	wire [WIDTH-1:0] wire_d25_83;
	wire [WIDTH-1:0] wire_d25_84;
	wire [WIDTH-1:0] wire_d25_85;
	wire [WIDTH-1:0] wire_d25_86;
	wire [WIDTH-1:0] wire_d25_87;
	wire [WIDTH-1:0] wire_d25_88;
	wire [WIDTH-1:0] wire_d25_89;
	wire [WIDTH-1:0] wire_d25_90;
	wire [WIDTH-1:0] wire_d25_91;
	wire [WIDTH-1:0] wire_d25_92;
	wire [WIDTH-1:0] wire_d25_93;
	wire [WIDTH-1:0] wire_d25_94;
	wire [WIDTH-1:0] wire_d25_95;
	wire [WIDTH-1:0] wire_d25_96;
	wire [WIDTH-1:0] wire_d25_97;
	wire [WIDTH-1:0] wire_d25_98;
	wire [WIDTH-1:0] wire_d26_0;
	wire [WIDTH-1:0] wire_d26_1;
	wire [WIDTH-1:0] wire_d26_2;
	wire [WIDTH-1:0] wire_d26_3;
	wire [WIDTH-1:0] wire_d26_4;
	wire [WIDTH-1:0] wire_d26_5;
	wire [WIDTH-1:0] wire_d26_6;
	wire [WIDTH-1:0] wire_d26_7;
	wire [WIDTH-1:0] wire_d26_8;
	wire [WIDTH-1:0] wire_d26_9;
	wire [WIDTH-1:0] wire_d26_10;
	wire [WIDTH-1:0] wire_d26_11;
	wire [WIDTH-1:0] wire_d26_12;
	wire [WIDTH-1:0] wire_d26_13;
	wire [WIDTH-1:0] wire_d26_14;
	wire [WIDTH-1:0] wire_d26_15;
	wire [WIDTH-1:0] wire_d26_16;
	wire [WIDTH-1:0] wire_d26_17;
	wire [WIDTH-1:0] wire_d26_18;
	wire [WIDTH-1:0] wire_d26_19;
	wire [WIDTH-1:0] wire_d26_20;
	wire [WIDTH-1:0] wire_d26_21;
	wire [WIDTH-1:0] wire_d26_22;
	wire [WIDTH-1:0] wire_d26_23;
	wire [WIDTH-1:0] wire_d26_24;
	wire [WIDTH-1:0] wire_d26_25;
	wire [WIDTH-1:0] wire_d26_26;
	wire [WIDTH-1:0] wire_d26_27;
	wire [WIDTH-1:0] wire_d26_28;
	wire [WIDTH-1:0] wire_d26_29;
	wire [WIDTH-1:0] wire_d26_30;
	wire [WIDTH-1:0] wire_d26_31;
	wire [WIDTH-1:0] wire_d26_32;
	wire [WIDTH-1:0] wire_d26_33;
	wire [WIDTH-1:0] wire_d26_34;
	wire [WIDTH-1:0] wire_d26_35;
	wire [WIDTH-1:0] wire_d26_36;
	wire [WIDTH-1:0] wire_d26_37;
	wire [WIDTH-1:0] wire_d26_38;
	wire [WIDTH-1:0] wire_d26_39;
	wire [WIDTH-1:0] wire_d26_40;
	wire [WIDTH-1:0] wire_d26_41;
	wire [WIDTH-1:0] wire_d26_42;
	wire [WIDTH-1:0] wire_d26_43;
	wire [WIDTH-1:0] wire_d26_44;
	wire [WIDTH-1:0] wire_d26_45;
	wire [WIDTH-1:0] wire_d26_46;
	wire [WIDTH-1:0] wire_d26_47;
	wire [WIDTH-1:0] wire_d26_48;
	wire [WIDTH-1:0] wire_d26_49;
	wire [WIDTH-1:0] wire_d26_50;
	wire [WIDTH-1:0] wire_d26_51;
	wire [WIDTH-1:0] wire_d26_52;
	wire [WIDTH-1:0] wire_d26_53;
	wire [WIDTH-1:0] wire_d26_54;
	wire [WIDTH-1:0] wire_d26_55;
	wire [WIDTH-1:0] wire_d26_56;
	wire [WIDTH-1:0] wire_d26_57;
	wire [WIDTH-1:0] wire_d26_58;
	wire [WIDTH-1:0] wire_d26_59;
	wire [WIDTH-1:0] wire_d26_60;
	wire [WIDTH-1:0] wire_d26_61;
	wire [WIDTH-1:0] wire_d26_62;
	wire [WIDTH-1:0] wire_d26_63;
	wire [WIDTH-1:0] wire_d26_64;
	wire [WIDTH-1:0] wire_d26_65;
	wire [WIDTH-1:0] wire_d26_66;
	wire [WIDTH-1:0] wire_d26_67;
	wire [WIDTH-1:0] wire_d26_68;
	wire [WIDTH-1:0] wire_d26_69;
	wire [WIDTH-1:0] wire_d26_70;
	wire [WIDTH-1:0] wire_d26_71;
	wire [WIDTH-1:0] wire_d26_72;
	wire [WIDTH-1:0] wire_d26_73;
	wire [WIDTH-1:0] wire_d26_74;
	wire [WIDTH-1:0] wire_d26_75;
	wire [WIDTH-1:0] wire_d26_76;
	wire [WIDTH-1:0] wire_d26_77;
	wire [WIDTH-1:0] wire_d26_78;
	wire [WIDTH-1:0] wire_d26_79;
	wire [WIDTH-1:0] wire_d26_80;
	wire [WIDTH-1:0] wire_d26_81;
	wire [WIDTH-1:0] wire_d26_82;
	wire [WIDTH-1:0] wire_d26_83;
	wire [WIDTH-1:0] wire_d26_84;
	wire [WIDTH-1:0] wire_d26_85;
	wire [WIDTH-1:0] wire_d26_86;
	wire [WIDTH-1:0] wire_d26_87;
	wire [WIDTH-1:0] wire_d26_88;
	wire [WIDTH-1:0] wire_d26_89;
	wire [WIDTH-1:0] wire_d26_90;
	wire [WIDTH-1:0] wire_d26_91;
	wire [WIDTH-1:0] wire_d26_92;
	wire [WIDTH-1:0] wire_d26_93;
	wire [WIDTH-1:0] wire_d26_94;
	wire [WIDTH-1:0] wire_d26_95;
	wire [WIDTH-1:0] wire_d26_96;
	wire [WIDTH-1:0] wire_d26_97;
	wire [WIDTH-1:0] wire_d26_98;
	wire [WIDTH-1:0] wire_d27_0;
	wire [WIDTH-1:0] wire_d27_1;
	wire [WIDTH-1:0] wire_d27_2;
	wire [WIDTH-1:0] wire_d27_3;
	wire [WIDTH-1:0] wire_d27_4;
	wire [WIDTH-1:0] wire_d27_5;
	wire [WIDTH-1:0] wire_d27_6;
	wire [WIDTH-1:0] wire_d27_7;
	wire [WIDTH-1:0] wire_d27_8;
	wire [WIDTH-1:0] wire_d27_9;
	wire [WIDTH-1:0] wire_d27_10;
	wire [WIDTH-1:0] wire_d27_11;
	wire [WIDTH-1:0] wire_d27_12;
	wire [WIDTH-1:0] wire_d27_13;
	wire [WIDTH-1:0] wire_d27_14;
	wire [WIDTH-1:0] wire_d27_15;
	wire [WIDTH-1:0] wire_d27_16;
	wire [WIDTH-1:0] wire_d27_17;
	wire [WIDTH-1:0] wire_d27_18;
	wire [WIDTH-1:0] wire_d27_19;
	wire [WIDTH-1:0] wire_d27_20;
	wire [WIDTH-1:0] wire_d27_21;
	wire [WIDTH-1:0] wire_d27_22;
	wire [WIDTH-1:0] wire_d27_23;
	wire [WIDTH-1:0] wire_d27_24;
	wire [WIDTH-1:0] wire_d27_25;
	wire [WIDTH-1:0] wire_d27_26;
	wire [WIDTH-1:0] wire_d27_27;
	wire [WIDTH-1:0] wire_d27_28;
	wire [WIDTH-1:0] wire_d27_29;
	wire [WIDTH-1:0] wire_d27_30;
	wire [WIDTH-1:0] wire_d27_31;
	wire [WIDTH-1:0] wire_d27_32;
	wire [WIDTH-1:0] wire_d27_33;
	wire [WIDTH-1:0] wire_d27_34;
	wire [WIDTH-1:0] wire_d27_35;
	wire [WIDTH-1:0] wire_d27_36;
	wire [WIDTH-1:0] wire_d27_37;
	wire [WIDTH-1:0] wire_d27_38;
	wire [WIDTH-1:0] wire_d27_39;
	wire [WIDTH-1:0] wire_d27_40;
	wire [WIDTH-1:0] wire_d27_41;
	wire [WIDTH-1:0] wire_d27_42;
	wire [WIDTH-1:0] wire_d27_43;
	wire [WIDTH-1:0] wire_d27_44;
	wire [WIDTH-1:0] wire_d27_45;
	wire [WIDTH-1:0] wire_d27_46;
	wire [WIDTH-1:0] wire_d27_47;
	wire [WIDTH-1:0] wire_d27_48;
	wire [WIDTH-1:0] wire_d27_49;
	wire [WIDTH-1:0] wire_d27_50;
	wire [WIDTH-1:0] wire_d27_51;
	wire [WIDTH-1:0] wire_d27_52;
	wire [WIDTH-1:0] wire_d27_53;
	wire [WIDTH-1:0] wire_d27_54;
	wire [WIDTH-1:0] wire_d27_55;
	wire [WIDTH-1:0] wire_d27_56;
	wire [WIDTH-1:0] wire_d27_57;
	wire [WIDTH-1:0] wire_d27_58;
	wire [WIDTH-1:0] wire_d27_59;
	wire [WIDTH-1:0] wire_d27_60;
	wire [WIDTH-1:0] wire_d27_61;
	wire [WIDTH-1:0] wire_d27_62;
	wire [WIDTH-1:0] wire_d27_63;
	wire [WIDTH-1:0] wire_d27_64;
	wire [WIDTH-1:0] wire_d27_65;
	wire [WIDTH-1:0] wire_d27_66;
	wire [WIDTH-1:0] wire_d27_67;
	wire [WIDTH-1:0] wire_d27_68;
	wire [WIDTH-1:0] wire_d27_69;
	wire [WIDTH-1:0] wire_d27_70;
	wire [WIDTH-1:0] wire_d27_71;
	wire [WIDTH-1:0] wire_d27_72;
	wire [WIDTH-1:0] wire_d27_73;
	wire [WIDTH-1:0] wire_d27_74;
	wire [WIDTH-1:0] wire_d27_75;
	wire [WIDTH-1:0] wire_d27_76;
	wire [WIDTH-1:0] wire_d27_77;
	wire [WIDTH-1:0] wire_d27_78;
	wire [WIDTH-1:0] wire_d27_79;
	wire [WIDTH-1:0] wire_d27_80;
	wire [WIDTH-1:0] wire_d27_81;
	wire [WIDTH-1:0] wire_d27_82;
	wire [WIDTH-1:0] wire_d27_83;
	wire [WIDTH-1:0] wire_d27_84;
	wire [WIDTH-1:0] wire_d27_85;
	wire [WIDTH-1:0] wire_d27_86;
	wire [WIDTH-1:0] wire_d27_87;
	wire [WIDTH-1:0] wire_d27_88;
	wire [WIDTH-1:0] wire_d27_89;
	wire [WIDTH-1:0] wire_d27_90;
	wire [WIDTH-1:0] wire_d27_91;
	wire [WIDTH-1:0] wire_d27_92;
	wire [WIDTH-1:0] wire_d27_93;
	wire [WIDTH-1:0] wire_d27_94;
	wire [WIDTH-1:0] wire_d27_95;
	wire [WIDTH-1:0] wire_d27_96;
	wire [WIDTH-1:0] wire_d27_97;
	wire [WIDTH-1:0] wire_d27_98;
	wire [WIDTH-1:0] wire_d28_0;
	wire [WIDTH-1:0] wire_d28_1;
	wire [WIDTH-1:0] wire_d28_2;
	wire [WIDTH-1:0] wire_d28_3;
	wire [WIDTH-1:0] wire_d28_4;
	wire [WIDTH-1:0] wire_d28_5;
	wire [WIDTH-1:0] wire_d28_6;
	wire [WIDTH-1:0] wire_d28_7;
	wire [WIDTH-1:0] wire_d28_8;
	wire [WIDTH-1:0] wire_d28_9;
	wire [WIDTH-1:0] wire_d28_10;
	wire [WIDTH-1:0] wire_d28_11;
	wire [WIDTH-1:0] wire_d28_12;
	wire [WIDTH-1:0] wire_d28_13;
	wire [WIDTH-1:0] wire_d28_14;
	wire [WIDTH-1:0] wire_d28_15;
	wire [WIDTH-1:0] wire_d28_16;
	wire [WIDTH-1:0] wire_d28_17;
	wire [WIDTH-1:0] wire_d28_18;
	wire [WIDTH-1:0] wire_d28_19;
	wire [WIDTH-1:0] wire_d28_20;
	wire [WIDTH-1:0] wire_d28_21;
	wire [WIDTH-1:0] wire_d28_22;
	wire [WIDTH-1:0] wire_d28_23;
	wire [WIDTH-1:0] wire_d28_24;
	wire [WIDTH-1:0] wire_d28_25;
	wire [WIDTH-1:0] wire_d28_26;
	wire [WIDTH-1:0] wire_d28_27;
	wire [WIDTH-1:0] wire_d28_28;
	wire [WIDTH-1:0] wire_d28_29;
	wire [WIDTH-1:0] wire_d28_30;
	wire [WIDTH-1:0] wire_d28_31;
	wire [WIDTH-1:0] wire_d28_32;
	wire [WIDTH-1:0] wire_d28_33;
	wire [WIDTH-1:0] wire_d28_34;
	wire [WIDTH-1:0] wire_d28_35;
	wire [WIDTH-1:0] wire_d28_36;
	wire [WIDTH-1:0] wire_d28_37;
	wire [WIDTH-1:0] wire_d28_38;
	wire [WIDTH-1:0] wire_d28_39;
	wire [WIDTH-1:0] wire_d28_40;
	wire [WIDTH-1:0] wire_d28_41;
	wire [WIDTH-1:0] wire_d28_42;
	wire [WIDTH-1:0] wire_d28_43;
	wire [WIDTH-1:0] wire_d28_44;
	wire [WIDTH-1:0] wire_d28_45;
	wire [WIDTH-1:0] wire_d28_46;
	wire [WIDTH-1:0] wire_d28_47;
	wire [WIDTH-1:0] wire_d28_48;
	wire [WIDTH-1:0] wire_d28_49;
	wire [WIDTH-1:0] wire_d28_50;
	wire [WIDTH-1:0] wire_d28_51;
	wire [WIDTH-1:0] wire_d28_52;
	wire [WIDTH-1:0] wire_d28_53;
	wire [WIDTH-1:0] wire_d28_54;
	wire [WIDTH-1:0] wire_d28_55;
	wire [WIDTH-1:0] wire_d28_56;
	wire [WIDTH-1:0] wire_d28_57;
	wire [WIDTH-1:0] wire_d28_58;
	wire [WIDTH-1:0] wire_d28_59;
	wire [WIDTH-1:0] wire_d28_60;
	wire [WIDTH-1:0] wire_d28_61;
	wire [WIDTH-1:0] wire_d28_62;
	wire [WIDTH-1:0] wire_d28_63;
	wire [WIDTH-1:0] wire_d28_64;
	wire [WIDTH-1:0] wire_d28_65;
	wire [WIDTH-1:0] wire_d28_66;
	wire [WIDTH-1:0] wire_d28_67;
	wire [WIDTH-1:0] wire_d28_68;
	wire [WIDTH-1:0] wire_d28_69;
	wire [WIDTH-1:0] wire_d28_70;
	wire [WIDTH-1:0] wire_d28_71;
	wire [WIDTH-1:0] wire_d28_72;
	wire [WIDTH-1:0] wire_d28_73;
	wire [WIDTH-1:0] wire_d28_74;
	wire [WIDTH-1:0] wire_d28_75;
	wire [WIDTH-1:0] wire_d28_76;
	wire [WIDTH-1:0] wire_d28_77;
	wire [WIDTH-1:0] wire_d28_78;
	wire [WIDTH-1:0] wire_d28_79;
	wire [WIDTH-1:0] wire_d28_80;
	wire [WIDTH-1:0] wire_d28_81;
	wire [WIDTH-1:0] wire_d28_82;
	wire [WIDTH-1:0] wire_d28_83;
	wire [WIDTH-1:0] wire_d28_84;
	wire [WIDTH-1:0] wire_d28_85;
	wire [WIDTH-1:0] wire_d28_86;
	wire [WIDTH-1:0] wire_d28_87;
	wire [WIDTH-1:0] wire_d28_88;
	wire [WIDTH-1:0] wire_d28_89;
	wire [WIDTH-1:0] wire_d28_90;
	wire [WIDTH-1:0] wire_d28_91;
	wire [WIDTH-1:0] wire_d28_92;
	wire [WIDTH-1:0] wire_d28_93;
	wire [WIDTH-1:0] wire_d28_94;
	wire [WIDTH-1:0] wire_d28_95;
	wire [WIDTH-1:0] wire_d28_96;
	wire [WIDTH-1:0] wire_d28_97;
	wire [WIDTH-1:0] wire_d28_98;
	wire [WIDTH-1:0] wire_d29_0;
	wire [WIDTH-1:0] wire_d29_1;
	wire [WIDTH-1:0] wire_d29_2;
	wire [WIDTH-1:0] wire_d29_3;
	wire [WIDTH-1:0] wire_d29_4;
	wire [WIDTH-1:0] wire_d29_5;
	wire [WIDTH-1:0] wire_d29_6;
	wire [WIDTH-1:0] wire_d29_7;
	wire [WIDTH-1:0] wire_d29_8;
	wire [WIDTH-1:0] wire_d29_9;
	wire [WIDTH-1:0] wire_d29_10;
	wire [WIDTH-1:0] wire_d29_11;
	wire [WIDTH-1:0] wire_d29_12;
	wire [WIDTH-1:0] wire_d29_13;
	wire [WIDTH-1:0] wire_d29_14;
	wire [WIDTH-1:0] wire_d29_15;
	wire [WIDTH-1:0] wire_d29_16;
	wire [WIDTH-1:0] wire_d29_17;
	wire [WIDTH-1:0] wire_d29_18;
	wire [WIDTH-1:0] wire_d29_19;
	wire [WIDTH-1:0] wire_d29_20;
	wire [WIDTH-1:0] wire_d29_21;
	wire [WIDTH-1:0] wire_d29_22;
	wire [WIDTH-1:0] wire_d29_23;
	wire [WIDTH-1:0] wire_d29_24;
	wire [WIDTH-1:0] wire_d29_25;
	wire [WIDTH-1:0] wire_d29_26;
	wire [WIDTH-1:0] wire_d29_27;
	wire [WIDTH-1:0] wire_d29_28;
	wire [WIDTH-1:0] wire_d29_29;
	wire [WIDTH-1:0] wire_d29_30;
	wire [WIDTH-1:0] wire_d29_31;
	wire [WIDTH-1:0] wire_d29_32;
	wire [WIDTH-1:0] wire_d29_33;
	wire [WIDTH-1:0] wire_d29_34;
	wire [WIDTH-1:0] wire_d29_35;
	wire [WIDTH-1:0] wire_d29_36;
	wire [WIDTH-1:0] wire_d29_37;
	wire [WIDTH-1:0] wire_d29_38;
	wire [WIDTH-1:0] wire_d29_39;
	wire [WIDTH-1:0] wire_d29_40;
	wire [WIDTH-1:0] wire_d29_41;
	wire [WIDTH-1:0] wire_d29_42;
	wire [WIDTH-1:0] wire_d29_43;
	wire [WIDTH-1:0] wire_d29_44;
	wire [WIDTH-1:0] wire_d29_45;
	wire [WIDTH-1:0] wire_d29_46;
	wire [WIDTH-1:0] wire_d29_47;
	wire [WIDTH-1:0] wire_d29_48;
	wire [WIDTH-1:0] wire_d29_49;
	wire [WIDTH-1:0] wire_d29_50;
	wire [WIDTH-1:0] wire_d29_51;
	wire [WIDTH-1:0] wire_d29_52;
	wire [WIDTH-1:0] wire_d29_53;
	wire [WIDTH-1:0] wire_d29_54;
	wire [WIDTH-1:0] wire_d29_55;
	wire [WIDTH-1:0] wire_d29_56;
	wire [WIDTH-1:0] wire_d29_57;
	wire [WIDTH-1:0] wire_d29_58;
	wire [WIDTH-1:0] wire_d29_59;
	wire [WIDTH-1:0] wire_d29_60;
	wire [WIDTH-1:0] wire_d29_61;
	wire [WIDTH-1:0] wire_d29_62;
	wire [WIDTH-1:0] wire_d29_63;
	wire [WIDTH-1:0] wire_d29_64;
	wire [WIDTH-1:0] wire_d29_65;
	wire [WIDTH-1:0] wire_d29_66;
	wire [WIDTH-1:0] wire_d29_67;
	wire [WIDTH-1:0] wire_d29_68;
	wire [WIDTH-1:0] wire_d29_69;
	wire [WIDTH-1:0] wire_d29_70;
	wire [WIDTH-1:0] wire_d29_71;
	wire [WIDTH-1:0] wire_d29_72;
	wire [WIDTH-1:0] wire_d29_73;
	wire [WIDTH-1:0] wire_d29_74;
	wire [WIDTH-1:0] wire_d29_75;
	wire [WIDTH-1:0] wire_d29_76;
	wire [WIDTH-1:0] wire_d29_77;
	wire [WIDTH-1:0] wire_d29_78;
	wire [WIDTH-1:0] wire_d29_79;
	wire [WIDTH-1:0] wire_d29_80;
	wire [WIDTH-1:0] wire_d29_81;
	wire [WIDTH-1:0] wire_d29_82;
	wire [WIDTH-1:0] wire_d29_83;
	wire [WIDTH-1:0] wire_d29_84;
	wire [WIDTH-1:0] wire_d29_85;
	wire [WIDTH-1:0] wire_d29_86;
	wire [WIDTH-1:0] wire_d29_87;
	wire [WIDTH-1:0] wire_d29_88;
	wire [WIDTH-1:0] wire_d29_89;
	wire [WIDTH-1:0] wire_d29_90;
	wire [WIDTH-1:0] wire_d29_91;
	wire [WIDTH-1:0] wire_d29_92;
	wire [WIDTH-1:0] wire_d29_93;
	wire [WIDTH-1:0] wire_d29_94;
	wire [WIDTH-1:0] wire_d29_95;
	wire [WIDTH-1:0] wire_d29_96;
	wire [WIDTH-1:0] wire_d29_97;
	wire [WIDTH-1:0] wire_d29_98;
	wire [WIDTH-1:0] wire_d30_0;
	wire [WIDTH-1:0] wire_d30_1;
	wire [WIDTH-1:0] wire_d30_2;
	wire [WIDTH-1:0] wire_d30_3;
	wire [WIDTH-1:0] wire_d30_4;
	wire [WIDTH-1:0] wire_d30_5;
	wire [WIDTH-1:0] wire_d30_6;
	wire [WIDTH-1:0] wire_d30_7;
	wire [WIDTH-1:0] wire_d30_8;
	wire [WIDTH-1:0] wire_d30_9;
	wire [WIDTH-1:0] wire_d30_10;
	wire [WIDTH-1:0] wire_d30_11;
	wire [WIDTH-1:0] wire_d30_12;
	wire [WIDTH-1:0] wire_d30_13;
	wire [WIDTH-1:0] wire_d30_14;
	wire [WIDTH-1:0] wire_d30_15;
	wire [WIDTH-1:0] wire_d30_16;
	wire [WIDTH-1:0] wire_d30_17;
	wire [WIDTH-1:0] wire_d30_18;
	wire [WIDTH-1:0] wire_d30_19;
	wire [WIDTH-1:0] wire_d30_20;
	wire [WIDTH-1:0] wire_d30_21;
	wire [WIDTH-1:0] wire_d30_22;
	wire [WIDTH-1:0] wire_d30_23;
	wire [WIDTH-1:0] wire_d30_24;
	wire [WIDTH-1:0] wire_d30_25;
	wire [WIDTH-1:0] wire_d30_26;
	wire [WIDTH-1:0] wire_d30_27;
	wire [WIDTH-1:0] wire_d30_28;
	wire [WIDTH-1:0] wire_d30_29;
	wire [WIDTH-1:0] wire_d30_30;
	wire [WIDTH-1:0] wire_d30_31;
	wire [WIDTH-1:0] wire_d30_32;
	wire [WIDTH-1:0] wire_d30_33;
	wire [WIDTH-1:0] wire_d30_34;
	wire [WIDTH-1:0] wire_d30_35;
	wire [WIDTH-1:0] wire_d30_36;
	wire [WIDTH-1:0] wire_d30_37;
	wire [WIDTH-1:0] wire_d30_38;
	wire [WIDTH-1:0] wire_d30_39;
	wire [WIDTH-1:0] wire_d30_40;
	wire [WIDTH-1:0] wire_d30_41;
	wire [WIDTH-1:0] wire_d30_42;
	wire [WIDTH-1:0] wire_d30_43;
	wire [WIDTH-1:0] wire_d30_44;
	wire [WIDTH-1:0] wire_d30_45;
	wire [WIDTH-1:0] wire_d30_46;
	wire [WIDTH-1:0] wire_d30_47;
	wire [WIDTH-1:0] wire_d30_48;
	wire [WIDTH-1:0] wire_d30_49;
	wire [WIDTH-1:0] wire_d30_50;
	wire [WIDTH-1:0] wire_d30_51;
	wire [WIDTH-1:0] wire_d30_52;
	wire [WIDTH-1:0] wire_d30_53;
	wire [WIDTH-1:0] wire_d30_54;
	wire [WIDTH-1:0] wire_d30_55;
	wire [WIDTH-1:0] wire_d30_56;
	wire [WIDTH-1:0] wire_d30_57;
	wire [WIDTH-1:0] wire_d30_58;
	wire [WIDTH-1:0] wire_d30_59;
	wire [WIDTH-1:0] wire_d30_60;
	wire [WIDTH-1:0] wire_d30_61;
	wire [WIDTH-1:0] wire_d30_62;
	wire [WIDTH-1:0] wire_d30_63;
	wire [WIDTH-1:0] wire_d30_64;
	wire [WIDTH-1:0] wire_d30_65;
	wire [WIDTH-1:0] wire_d30_66;
	wire [WIDTH-1:0] wire_d30_67;
	wire [WIDTH-1:0] wire_d30_68;
	wire [WIDTH-1:0] wire_d30_69;
	wire [WIDTH-1:0] wire_d30_70;
	wire [WIDTH-1:0] wire_d30_71;
	wire [WIDTH-1:0] wire_d30_72;
	wire [WIDTH-1:0] wire_d30_73;
	wire [WIDTH-1:0] wire_d30_74;
	wire [WIDTH-1:0] wire_d30_75;
	wire [WIDTH-1:0] wire_d30_76;
	wire [WIDTH-1:0] wire_d30_77;
	wire [WIDTH-1:0] wire_d30_78;
	wire [WIDTH-1:0] wire_d30_79;
	wire [WIDTH-1:0] wire_d30_80;
	wire [WIDTH-1:0] wire_d30_81;
	wire [WIDTH-1:0] wire_d30_82;
	wire [WIDTH-1:0] wire_d30_83;
	wire [WIDTH-1:0] wire_d30_84;
	wire [WIDTH-1:0] wire_d30_85;
	wire [WIDTH-1:0] wire_d30_86;
	wire [WIDTH-1:0] wire_d30_87;
	wire [WIDTH-1:0] wire_d30_88;
	wire [WIDTH-1:0] wire_d30_89;
	wire [WIDTH-1:0] wire_d30_90;
	wire [WIDTH-1:0] wire_d30_91;
	wire [WIDTH-1:0] wire_d30_92;
	wire [WIDTH-1:0] wire_d30_93;
	wire [WIDTH-1:0] wire_d30_94;
	wire [WIDTH-1:0] wire_d30_95;
	wire [WIDTH-1:0] wire_d30_96;
	wire [WIDTH-1:0] wire_d30_97;
	wire [WIDTH-1:0] wire_d30_98;
	wire [WIDTH-1:0] wire_d31_0;
	wire [WIDTH-1:0] wire_d31_1;
	wire [WIDTH-1:0] wire_d31_2;
	wire [WIDTH-1:0] wire_d31_3;
	wire [WIDTH-1:0] wire_d31_4;
	wire [WIDTH-1:0] wire_d31_5;
	wire [WIDTH-1:0] wire_d31_6;
	wire [WIDTH-1:0] wire_d31_7;
	wire [WIDTH-1:0] wire_d31_8;
	wire [WIDTH-1:0] wire_d31_9;
	wire [WIDTH-1:0] wire_d31_10;
	wire [WIDTH-1:0] wire_d31_11;
	wire [WIDTH-1:0] wire_d31_12;
	wire [WIDTH-1:0] wire_d31_13;
	wire [WIDTH-1:0] wire_d31_14;
	wire [WIDTH-1:0] wire_d31_15;
	wire [WIDTH-1:0] wire_d31_16;
	wire [WIDTH-1:0] wire_d31_17;
	wire [WIDTH-1:0] wire_d31_18;
	wire [WIDTH-1:0] wire_d31_19;
	wire [WIDTH-1:0] wire_d31_20;
	wire [WIDTH-1:0] wire_d31_21;
	wire [WIDTH-1:0] wire_d31_22;
	wire [WIDTH-1:0] wire_d31_23;
	wire [WIDTH-1:0] wire_d31_24;
	wire [WIDTH-1:0] wire_d31_25;
	wire [WIDTH-1:0] wire_d31_26;
	wire [WIDTH-1:0] wire_d31_27;
	wire [WIDTH-1:0] wire_d31_28;
	wire [WIDTH-1:0] wire_d31_29;
	wire [WIDTH-1:0] wire_d31_30;
	wire [WIDTH-1:0] wire_d31_31;
	wire [WIDTH-1:0] wire_d31_32;
	wire [WIDTH-1:0] wire_d31_33;
	wire [WIDTH-1:0] wire_d31_34;
	wire [WIDTH-1:0] wire_d31_35;
	wire [WIDTH-1:0] wire_d31_36;
	wire [WIDTH-1:0] wire_d31_37;
	wire [WIDTH-1:0] wire_d31_38;
	wire [WIDTH-1:0] wire_d31_39;
	wire [WIDTH-1:0] wire_d31_40;
	wire [WIDTH-1:0] wire_d31_41;
	wire [WIDTH-1:0] wire_d31_42;
	wire [WIDTH-1:0] wire_d31_43;
	wire [WIDTH-1:0] wire_d31_44;
	wire [WIDTH-1:0] wire_d31_45;
	wire [WIDTH-1:0] wire_d31_46;
	wire [WIDTH-1:0] wire_d31_47;
	wire [WIDTH-1:0] wire_d31_48;
	wire [WIDTH-1:0] wire_d31_49;
	wire [WIDTH-1:0] wire_d31_50;
	wire [WIDTH-1:0] wire_d31_51;
	wire [WIDTH-1:0] wire_d31_52;
	wire [WIDTH-1:0] wire_d31_53;
	wire [WIDTH-1:0] wire_d31_54;
	wire [WIDTH-1:0] wire_d31_55;
	wire [WIDTH-1:0] wire_d31_56;
	wire [WIDTH-1:0] wire_d31_57;
	wire [WIDTH-1:0] wire_d31_58;
	wire [WIDTH-1:0] wire_d31_59;
	wire [WIDTH-1:0] wire_d31_60;
	wire [WIDTH-1:0] wire_d31_61;
	wire [WIDTH-1:0] wire_d31_62;
	wire [WIDTH-1:0] wire_d31_63;
	wire [WIDTH-1:0] wire_d31_64;
	wire [WIDTH-1:0] wire_d31_65;
	wire [WIDTH-1:0] wire_d31_66;
	wire [WIDTH-1:0] wire_d31_67;
	wire [WIDTH-1:0] wire_d31_68;
	wire [WIDTH-1:0] wire_d31_69;
	wire [WIDTH-1:0] wire_d31_70;
	wire [WIDTH-1:0] wire_d31_71;
	wire [WIDTH-1:0] wire_d31_72;
	wire [WIDTH-1:0] wire_d31_73;
	wire [WIDTH-1:0] wire_d31_74;
	wire [WIDTH-1:0] wire_d31_75;
	wire [WIDTH-1:0] wire_d31_76;
	wire [WIDTH-1:0] wire_d31_77;
	wire [WIDTH-1:0] wire_d31_78;
	wire [WIDTH-1:0] wire_d31_79;
	wire [WIDTH-1:0] wire_d31_80;
	wire [WIDTH-1:0] wire_d31_81;
	wire [WIDTH-1:0] wire_d31_82;
	wire [WIDTH-1:0] wire_d31_83;
	wire [WIDTH-1:0] wire_d31_84;
	wire [WIDTH-1:0] wire_d31_85;
	wire [WIDTH-1:0] wire_d31_86;
	wire [WIDTH-1:0] wire_d31_87;
	wire [WIDTH-1:0] wire_d31_88;
	wire [WIDTH-1:0] wire_d31_89;
	wire [WIDTH-1:0] wire_d31_90;
	wire [WIDTH-1:0] wire_d31_91;
	wire [WIDTH-1:0] wire_d31_92;
	wire [WIDTH-1:0] wire_d31_93;
	wire [WIDTH-1:0] wire_d31_94;
	wire [WIDTH-1:0] wire_d31_95;
	wire [WIDTH-1:0] wire_d31_96;
	wire [WIDTH-1:0] wire_d31_97;
	wire [WIDTH-1:0] wire_d31_98;
	wire [WIDTH-1:0] wire_d32_0;
	wire [WIDTH-1:0] wire_d32_1;
	wire [WIDTH-1:0] wire_d32_2;
	wire [WIDTH-1:0] wire_d32_3;
	wire [WIDTH-1:0] wire_d32_4;
	wire [WIDTH-1:0] wire_d32_5;
	wire [WIDTH-1:0] wire_d32_6;
	wire [WIDTH-1:0] wire_d32_7;
	wire [WIDTH-1:0] wire_d32_8;
	wire [WIDTH-1:0] wire_d32_9;
	wire [WIDTH-1:0] wire_d32_10;
	wire [WIDTH-1:0] wire_d32_11;
	wire [WIDTH-1:0] wire_d32_12;
	wire [WIDTH-1:0] wire_d32_13;
	wire [WIDTH-1:0] wire_d32_14;
	wire [WIDTH-1:0] wire_d32_15;
	wire [WIDTH-1:0] wire_d32_16;
	wire [WIDTH-1:0] wire_d32_17;
	wire [WIDTH-1:0] wire_d32_18;
	wire [WIDTH-1:0] wire_d32_19;
	wire [WIDTH-1:0] wire_d32_20;
	wire [WIDTH-1:0] wire_d32_21;
	wire [WIDTH-1:0] wire_d32_22;
	wire [WIDTH-1:0] wire_d32_23;
	wire [WIDTH-1:0] wire_d32_24;
	wire [WIDTH-1:0] wire_d32_25;
	wire [WIDTH-1:0] wire_d32_26;
	wire [WIDTH-1:0] wire_d32_27;
	wire [WIDTH-1:0] wire_d32_28;
	wire [WIDTH-1:0] wire_d32_29;
	wire [WIDTH-1:0] wire_d32_30;
	wire [WIDTH-1:0] wire_d32_31;
	wire [WIDTH-1:0] wire_d32_32;
	wire [WIDTH-1:0] wire_d32_33;
	wire [WIDTH-1:0] wire_d32_34;
	wire [WIDTH-1:0] wire_d32_35;
	wire [WIDTH-1:0] wire_d32_36;
	wire [WIDTH-1:0] wire_d32_37;
	wire [WIDTH-1:0] wire_d32_38;
	wire [WIDTH-1:0] wire_d32_39;
	wire [WIDTH-1:0] wire_d32_40;
	wire [WIDTH-1:0] wire_d32_41;
	wire [WIDTH-1:0] wire_d32_42;
	wire [WIDTH-1:0] wire_d32_43;
	wire [WIDTH-1:0] wire_d32_44;
	wire [WIDTH-1:0] wire_d32_45;
	wire [WIDTH-1:0] wire_d32_46;
	wire [WIDTH-1:0] wire_d32_47;
	wire [WIDTH-1:0] wire_d32_48;
	wire [WIDTH-1:0] wire_d32_49;
	wire [WIDTH-1:0] wire_d32_50;
	wire [WIDTH-1:0] wire_d32_51;
	wire [WIDTH-1:0] wire_d32_52;
	wire [WIDTH-1:0] wire_d32_53;
	wire [WIDTH-1:0] wire_d32_54;
	wire [WIDTH-1:0] wire_d32_55;
	wire [WIDTH-1:0] wire_d32_56;
	wire [WIDTH-1:0] wire_d32_57;
	wire [WIDTH-1:0] wire_d32_58;
	wire [WIDTH-1:0] wire_d32_59;
	wire [WIDTH-1:0] wire_d32_60;
	wire [WIDTH-1:0] wire_d32_61;
	wire [WIDTH-1:0] wire_d32_62;
	wire [WIDTH-1:0] wire_d32_63;
	wire [WIDTH-1:0] wire_d32_64;
	wire [WIDTH-1:0] wire_d32_65;
	wire [WIDTH-1:0] wire_d32_66;
	wire [WIDTH-1:0] wire_d32_67;
	wire [WIDTH-1:0] wire_d32_68;
	wire [WIDTH-1:0] wire_d32_69;
	wire [WIDTH-1:0] wire_d32_70;
	wire [WIDTH-1:0] wire_d32_71;
	wire [WIDTH-1:0] wire_d32_72;
	wire [WIDTH-1:0] wire_d32_73;
	wire [WIDTH-1:0] wire_d32_74;
	wire [WIDTH-1:0] wire_d32_75;
	wire [WIDTH-1:0] wire_d32_76;
	wire [WIDTH-1:0] wire_d32_77;
	wire [WIDTH-1:0] wire_d32_78;
	wire [WIDTH-1:0] wire_d32_79;
	wire [WIDTH-1:0] wire_d32_80;
	wire [WIDTH-1:0] wire_d32_81;
	wire [WIDTH-1:0] wire_d32_82;
	wire [WIDTH-1:0] wire_d32_83;
	wire [WIDTH-1:0] wire_d32_84;
	wire [WIDTH-1:0] wire_d32_85;
	wire [WIDTH-1:0] wire_d32_86;
	wire [WIDTH-1:0] wire_d32_87;
	wire [WIDTH-1:0] wire_d32_88;
	wire [WIDTH-1:0] wire_d32_89;
	wire [WIDTH-1:0] wire_d32_90;
	wire [WIDTH-1:0] wire_d32_91;
	wire [WIDTH-1:0] wire_d32_92;
	wire [WIDTH-1:0] wire_d32_93;
	wire [WIDTH-1:0] wire_d32_94;
	wire [WIDTH-1:0] wire_d32_95;
	wire [WIDTH-1:0] wire_d32_96;
	wire [WIDTH-1:0] wire_d32_97;
	wire [WIDTH-1:0] wire_d32_98;
	wire [WIDTH-1:0] wire_d33_0;
	wire [WIDTH-1:0] wire_d33_1;
	wire [WIDTH-1:0] wire_d33_2;
	wire [WIDTH-1:0] wire_d33_3;
	wire [WIDTH-1:0] wire_d33_4;
	wire [WIDTH-1:0] wire_d33_5;
	wire [WIDTH-1:0] wire_d33_6;
	wire [WIDTH-1:0] wire_d33_7;
	wire [WIDTH-1:0] wire_d33_8;
	wire [WIDTH-1:0] wire_d33_9;
	wire [WIDTH-1:0] wire_d33_10;
	wire [WIDTH-1:0] wire_d33_11;
	wire [WIDTH-1:0] wire_d33_12;
	wire [WIDTH-1:0] wire_d33_13;
	wire [WIDTH-1:0] wire_d33_14;
	wire [WIDTH-1:0] wire_d33_15;
	wire [WIDTH-1:0] wire_d33_16;
	wire [WIDTH-1:0] wire_d33_17;
	wire [WIDTH-1:0] wire_d33_18;
	wire [WIDTH-1:0] wire_d33_19;
	wire [WIDTH-1:0] wire_d33_20;
	wire [WIDTH-1:0] wire_d33_21;
	wire [WIDTH-1:0] wire_d33_22;
	wire [WIDTH-1:0] wire_d33_23;
	wire [WIDTH-1:0] wire_d33_24;
	wire [WIDTH-1:0] wire_d33_25;
	wire [WIDTH-1:0] wire_d33_26;
	wire [WIDTH-1:0] wire_d33_27;
	wire [WIDTH-1:0] wire_d33_28;
	wire [WIDTH-1:0] wire_d33_29;
	wire [WIDTH-1:0] wire_d33_30;
	wire [WIDTH-1:0] wire_d33_31;
	wire [WIDTH-1:0] wire_d33_32;
	wire [WIDTH-1:0] wire_d33_33;
	wire [WIDTH-1:0] wire_d33_34;
	wire [WIDTH-1:0] wire_d33_35;
	wire [WIDTH-1:0] wire_d33_36;
	wire [WIDTH-1:0] wire_d33_37;
	wire [WIDTH-1:0] wire_d33_38;
	wire [WIDTH-1:0] wire_d33_39;
	wire [WIDTH-1:0] wire_d33_40;
	wire [WIDTH-1:0] wire_d33_41;
	wire [WIDTH-1:0] wire_d33_42;
	wire [WIDTH-1:0] wire_d33_43;
	wire [WIDTH-1:0] wire_d33_44;
	wire [WIDTH-1:0] wire_d33_45;
	wire [WIDTH-1:0] wire_d33_46;
	wire [WIDTH-1:0] wire_d33_47;
	wire [WIDTH-1:0] wire_d33_48;
	wire [WIDTH-1:0] wire_d33_49;
	wire [WIDTH-1:0] wire_d33_50;
	wire [WIDTH-1:0] wire_d33_51;
	wire [WIDTH-1:0] wire_d33_52;
	wire [WIDTH-1:0] wire_d33_53;
	wire [WIDTH-1:0] wire_d33_54;
	wire [WIDTH-1:0] wire_d33_55;
	wire [WIDTH-1:0] wire_d33_56;
	wire [WIDTH-1:0] wire_d33_57;
	wire [WIDTH-1:0] wire_d33_58;
	wire [WIDTH-1:0] wire_d33_59;
	wire [WIDTH-1:0] wire_d33_60;
	wire [WIDTH-1:0] wire_d33_61;
	wire [WIDTH-1:0] wire_d33_62;
	wire [WIDTH-1:0] wire_d33_63;
	wire [WIDTH-1:0] wire_d33_64;
	wire [WIDTH-1:0] wire_d33_65;
	wire [WIDTH-1:0] wire_d33_66;
	wire [WIDTH-1:0] wire_d33_67;
	wire [WIDTH-1:0] wire_d33_68;
	wire [WIDTH-1:0] wire_d33_69;
	wire [WIDTH-1:0] wire_d33_70;
	wire [WIDTH-1:0] wire_d33_71;
	wire [WIDTH-1:0] wire_d33_72;
	wire [WIDTH-1:0] wire_d33_73;
	wire [WIDTH-1:0] wire_d33_74;
	wire [WIDTH-1:0] wire_d33_75;
	wire [WIDTH-1:0] wire_d33_76;
	wire [WIDTH-1:0] wire_d33_77;
	wire [WIDTH-1:0] wire_d33_78;
	wire [WIDTH-1:0] wire_d33_79;
	wire [WIDTH-1:0] wire_d33_80;
	wire [WIDTH-1:0] wire_d33_81;
	wire [WIDTH-1:0] wire_d33_82;
	wire [WIDTH-1:0] wire_d33_83;
	wire [WIDTH-1:0] wire_d33_84;
	wire [WIDTH-1:0] wire_d33_85;
	wire [WIDTH-1:0] wire_d33_86;
	wire [WIDTH-1:0] wire_d33_87;
	wire [WIDTH-1:0] wire_d33_88;
	wire [WIDTH-1:0] wire_d33_89;
	wire [WIDTH-1:0] wire_d33_90;
	wire [WIDTH-1:0] wire_d33_91;
	wire [WIDTH-1:0] wire_d33_92;
	wire [WIDTH-1:0] wire_d33_93;
	wire [WIDTH-1:0] wire_d33_94;
	wire [WIDTH-1:0] wire_d33_95;
	wire [WIDTH-1:0] wire_d33_96;
	wire [WIDTH-1:0] wire_d33_97;
	wire [WIDTH-1:0] wire_d33_98;
	wire [WIDTH-1:0] wire_d34_0;
	wire [WIDTH-1:0] wire_d34_1;
	wire [WIDTH-1:0] wire_d34_2;
	wire [WIDTH-1:0] wire_d34_3;
	wire [WIDTH-1:0] wire_d34_4;
	wire [WIDTH-1:0] wire_d34_5;
	wire [WIDTH-1:0] wire_d34_6;
	wire [WIDTH-1:0] wire_d34_7;
	wire [WIDTH-1:0] wire_d34_8;
	wire [WIDTH-1:0] wire_d34_9;
	wire [WIDTH-1:0] wire_d34_10;
	wire [WIDTH-1:0] wire_d34_11;
	wire [WIDTH-1:0] wire_d34_12;
	wire [WIDTH-1:0] wire_d34_13;
	wire [WIDTH-1:0] wire_d34_14;
	wire [WIDTH-1:0] wire_d34_15;
	wire [WIDTH-1:0] wire_d34_16;
	wire [WIDTH-1:0] wire_d34_17;
	wire [WIDTH-1:0] wire_d34_18;
	wire [WIDTH-1:0] wire_d34_19;
	wire [WIDTH-1:0] wire_d34_20;
	wire [WIDTH-1:0] wire_d34_21;
	wire [WIDTH-1:0] wire_d34_22;
	wire [WIDTH-1:0] wire_d34_23;
	wire [WIDTH-1:0] wire_d34_24;
	wire [WIDTH-1:0] wire_d34_25;
	wire [WIDTH-1:0] wire_d34_26;
	wire [WIDTH-1:0] wire_d34_27;
	wire [WIDTH-1:0] wire_d34_28;
	wire [WIDTH-1:0] wire_d34_29;
	wire [WIDTH-1:0] wire_d34_30;
	wire [WIDTH-1:0] wire_d34_31;
	wire [WIDTH-1:0] wire_d34_32;
	wire [WIDTH-1:0] wire_d34_33;
	wire [WIDTH-1:0] wire_d34_34;
	wire [WIDTH-1:0] wire_d34_35;
	wire [WIDTH-1:0] wire_d34_36;
	wire [WIDTH-1:0] wire_d34_37;
	wire [WIDTH-1:0] wire_d34_38;
	wire [WIDTH-1:0] wire_d34_39;
	wire [WIDTH-1:0] wire_d34_40;
	wire [WIDTH-1:0] wire_d34_41;
	wire [WIDTH-1:0] wire_d34_42;
	wire [WIDTH-1:0] wire_d34_43;
	wire [WIDTH-1:0] wire_d34_44;
	wire [WIDTH-1:0] wire_d34_45;
	wire [WIDTH-1:0] wire_d34_46;
	wire [WIDTH-1:0] wire_d34_47;
	wire [WIDTH-1:0] wire_d34_48;
	wire [WIDTH-1:0] wire_d34_49;
	wire [WIDTH-1:0] wire_d34_50;
	wire [WIDTH-1:0] wire_d34_51;
	wire [WIDTH-1:0] wire_d34_52;
	wire [WIDTH-1:0] wire_d34_53;
	wire [WIDTH-1:0] wire_d34_54;
	wire [WIDTH-1:0] wire_d34_55;
	wire [WIDTH-1:0] wire_d34_56;
	wire [WIDTH-1:0] wire_d34_57;
	wire [WIDTH-1:0] wire_d34_58;
	wire [WIDTH-1:0] wire_d34_59;
	wire [WIDTH-1:0] wire_d34_60;
	wire [WIDTH-1:0] wire_d34_61;
	wire [WIDTH-1:0] wire_d34_62;
	wire [WIDTH-1:0] wire_d34_63;
	wire [WIDTH-1:0] wire_d34_64;
	wire [WIDTH-1:0] wire_d34_65;
	wire [WIDTH-1:0] wire_d34_66;
	wire [WIDTH-1:0] wire_d34_67;
	wire [WIDTH-1:0] wire_d34_68;
	wire [WIDTH-1:0] wire_d34_69;
	wire [WIDTH-1:0] wire_d34_70;
	wire [WIDTH-1:0] wire_d34_71;
	wire [WIDTH-1:0] wire_d34_72;
	wire [WIDTH-1:0] wire_d34_73;
	wire [WIDTH-1:0] wire_d34_74;
	wire [WIDTH-1:0] wire_d34_75;
	wire [WIDTH-1:0] wire_d34_76;
	wire [WIDTH-1:0] wire_d34_77;
	wire [WIDTH-1:0] wire_d34_78;
	wire [WIDTH-1:0] wire_d34_79;
	wire [WIDTH-1:0] wire_d34_80;
	wire [WIDTH-1:0] wire_d34_81;
	wire [WIDTH-1:0] wire_d34_82;
	wire [WIDTH-1:0] wire_d34_83;
	wire [WIDTH-1:0] wire_d34_84;
	wire [WIDTH-1:0] wire_d34_85;
	wire [WIDTH-1:0] wire_d34_86;
	wire [WIDTH-1:0] wire_d34_87;
	wire [WIDTH-1:0] wire_d34_88;
	wire [WIDTH-1:0] wire_d34_89;
	wire [WIDTH-1:0] wire_d34_90;
	wire [WIDTH-1:0] wire_d34_91;
	wire [WIDTH-1:0] wire_d34_92;
	wire [WIDTH-1:0] wire_d34_93;
	wire [WIDTH-1:0] wire_d34_94;
	wire [WIDTH-1:0] wire_d34_95;
	wire [WIDTH-1:0] wire_d34_96;
	wire [WIDTH-1:0] wire_d34_97;
	wire [WIDTH-1:0] wire_d34_98;
	wire [WIDTH-1:0] wire_d35_0;
	wire [WIDTH-1:0] wire_d35_1;
	wire [WIDTH-1:0] wire_d35_2;
	wire [WIDTH-1:0] wire_d35_3;
	wire [WIDTH-1:0] wire_d35_4;
	wire [WIDTH-1:0] wire_d35_5;
	wire [WIDTH-1:0] wire_d35_6;
	wire [WIDTH-1:0] wire_d35_7;
	wire [WIDTH-1:0] wire_d35_8;
	wire [WIDTH-1:0] wire_d35_9;
	wire [WIDTH-1:0] wire_d35_10;
	wire [WIDTH-1:0] wire_d35_11;
	wire [WIDTH-1:0] wire_d35_12;
	wire [WIDTH-1:0] wire_d35_13;
	wire [WIDTH-1:0] wire_d35_14;
	wire [WIDTH-1:0] wire_d35_15;
	wire [WIDTH-1:0] wire_d35_16;
	wire [WIDTH-1:0] wire_d35_17;
	wire [WIDTH-1:0] wire_d35_18;
	wire [WIDTH-1:0] wire_d35_19;
	wire [WIDTH-1:0] wire_d35_20;
	wire [WIDTH-1:0] wire_d35_21;
	wire [WIDTH-1:0] wire_d35_22;
	wire [WIDTH-1:0] wire_d35_23;
	wire [WIDTH-1:0] wire_d35_24;
	wire [WIDTH-1:0] wire_d35_25;
	wire [WIDTH-1:0] wire_d35_26;
	wire [WIDTH-1:0] wire_d35_27;
	wire [WIDTH-1:0] wire_d35_28;
	wire [WIDTH-1:0] wire_d35_29;
	wire [WIDTH-1:0] wire_d35_30;
	wire [WIDTH-1:0] wire_d35_31;
	wire [WIDTH-1:0] wire_d35_32;
	wire [WIDTH-1:0] wire_d35_33;
	wire [WIDTH-1:0] wire_d35_34;
	wire [WIDTH-1:0] wire_d35_35;
	wire [WIDTH-1:0] wire_d35_36;
	wire [WIDTH-1:0] wire_d35_37;
	wire [WIDTH-1:0] wire_d35_38;
	wire [WIDTH-1:0] wire_d35_39;
	wire [WIDTH-1:0] wire_d35_40;
	wire [WIDTH-1:0] wire_d35_41;
	wire [WIDTH-1:0] wire_d35_42;
	wire [WIDTH-1:0] wire_d35_43;
	wire [WIDTH-1:0] wire_d35_44;
	wire [WIDTH-1:0] wire_d35_45;
	wire [WIDTH-1:0] wire_d35_46;
	wire [WIDTH-1:0] wire_d35_47;
	wire [WIDTH-1:0] wire_d35_48;
	wire [WIDTH-1:0] wire_d35_49;
	wire [WIDTH-1:0] wire_d35_50;
	wire [WIDTH-1:0] wire_d35_51;
	wire [WIDTH-1:0] wire_d35_52;
	wire [WIDTH-1:0] wire_d35_53;
	wire [WIDTH-1:0] wire_d35_54;
	wire [WIDTH-1:0] wire_d35_55;
	wire [WIDTH-1:0] wire_d35_56;
	wire [WIDTH-1:0] wire_d35_57;
	wire [WIDTH-1:0] wire_d35_58;
	wire [WIDTH-1:0] wire_d35_59;
	wire [WIDTH-1:0] wire_d35_60;
	wire [WIDTH-1:0] wire_d35_61;
	wire [WIDTH-1:0] wire_d35_62;
	wire [WIDTH-1:0] wire_d35_63;
	wire [WIDTH-1:0] wire_d35_64;
	wire [WIDTH-1:0] wire_d35_65;
	wire [WIDTH-1:0] wire_d35_66;
	wire [WIDTH-1:0] wire_d35_67;
	wire [WIDTH-1:0] wire_d35_68;
	wire [WIDTH-1:0] wire_d35_69;
	wire [WIDTH-1:0] wire_d35_70;
	wire [WIDTH-1:0] wire_d35_71;
	wire [WIDTH-1:0] wire_d35_72;
	wire [WIDTH-1:0] wire_d35_73;
	wire [WIDTH-1:0] wire_d35_74;
	wire [WIDTH-1:0] wire_d35_75;
	wire [WIDTH-1:0] wire_d35_76;
	wire [WIDTH-1:0] wire_d35_77;
	wire [WIDTH-1:0] wire_d35_78;
	wire [WIDTH-1:0] wire_d35_79;
	wire [WIDTH-1:0] wire_d35_80;
	wire [WIDTH-1:0] wire_d35_81;
	wire [WIDTH-1:0] wire_d35_82;
	wire [WIDTH-1:0] wire_d35_83;
	wire [WIDTH-1:0] wire_d35_84;
	wire [WIDTH-1:0] wire_d35_85;
	wire [WIDTH-1:0] wire_d35_86;
	wire [WIDTH-1:0] wire_d35_87;
	wire [WIDTH-1:0] wire_d35_88;
	wire [WIDTH-1:0] wire_d35_89;
	wire [WIDTH-1:0] wire_d35_90;
	wire [WIDTH-1:0] wire_d35_91;
	wire [WIDTH-1:0] wire_d35_92;
	wire [WIDTH-1:0] wire_d35_93;
	wire [WIDTH-1:0] wire_d35_94;
	wire [WIDTH-1:0] wire_d35_95;
	wire [WIDTH-1:0] wire_d35_96;
	wire [WIDTH-1:0] wire_d35_97;
	wire [WIDTH-1:0] wire_d35_98;
	wire [WIDTH-1:0] wire_d36_0;
	wire [WIDTH-1:0] wire_d36_1;
	wire [WIDTH-1:0] wire_d36_2;
	wire [WIDTH-1:0] wire_d36_3;
	wire [WIDTH-1:0] wire_d36_4;
	wire [WIDTH-1:0] wire_d36_5;
	wire [WIDTH-1:0] wire_d36_6;
	wire [WIDTH-1:0] wire_d36_7;
	wire [WIDTH-1:0] wire_d36_8;
	wire [WIDTH-1:0] wire_d36_9;
	wire [WIDTH-1:0] wire_d36_10;
	wire [WIDTH-1:0] wire_d36_11;
	wire [WIDTH-1:0] wire_d36_12;
	wire [WIDTH-1:0] wire_d36_13;
	wire [WIDTH-1:0] wire_d36_14;
	wire [WIDTH-1:0] wire_d36_15;
	wire [WIDTH-1:0] wire_d36_16;
	wire [WIDTH-1:0] wire_d36_17;
	wire [WIDTH-1:0] wire_d36_18;
	wire [WIDTH-1:0] wire_d36_19;
	wire [WIDTH-1:0] wire_d36_20;
	wire [WIDTH-1:0] wire_d36_21;
	wire [WIDTH-1:0] wire_d36_22;
	wire [WIDTH-1:0] wire_d36_23;
	wire [WIDTH-1:0] wire_d36_24;
	wire [WIDTH-1:0] wire_d36_25;
	wire [WIDTH-1:0] wire_d36_26;
	wire [WIDTH-1:0] wire_d36_27;
	wire [WIDTH-1:0] wire_d36_28;
	wire [WIDTH-1:0] wire_d36_29;
	wire [WIDTH-1:0] wire_d36_30;
	wire [WIDTH-1:0] wire_d36_31;
	wire [WIDTH-1:0] wire_d36_32;
	wire [WIDTH-1:0] wire_d36_33;
	wire [WIDTH-1:0] wire_d36_34;
	wire [WIDTH-1:0] wire_d36_35;
	wire [WIDTH-1:0] wire_d36_36;
	wire [WIDTH-1:0] wire_d36_37;
	wire [WIDTH-1:0] wire_d36_38;
	wire [WIDTH-1:0] wire_d36_39;
	wire [WIDTH-1:0] wire_d36_40;
	wire [WIDTH-1:0] wire_d36_41;
	wire [WIDTH-1:0] wire_d36_42;
	wire [WIDTH-1:0] wire_d36_43;
	wire [WIDTH-1:0] wire_d36_44;
	wire [WIDTH-1:0] wire_d36_45;
	wire [WIDTH-1:0] wire_d36_46;
	wire [WIDTH-1:0] wire_d36_47;
	wire [WIDTH-1:0] wire_d36_48;
	wire [WIDTH-1:0] wire_d36_49;
	wire [WIDTH-1:0] wire_d36_50;
	wire [WIDTH-1:0] wire_d36_51;
	wire [WIDTH-1:0] wire_d36_52;
	wire [WIDTH-1:0] wire_d36_53;
	wire [WIDTH-1:0] wire_d36_54;
	wire [WIDTH-1:0] wire_d36_55;
	wire [WIDTH-1:0] wire_d36_56;
	wire [WIDTH-1:0] wire_d36_57;
	wire [WIDTH-1:0] wire_d36_58;
	wire [WIDTH-1:0] wire_d36_59;
	wire [WIDTH-1:0] wire_d36_60;
	wire [WIDTH-1:0] wire_d36_61;
	wire [WIDTH-1:0] wire_d36_62;
	wire [WIDTH-1:0] wire_d36_63;
	wire [WIDTH-1:0] wire_d36_64;
	wire [WIDTH-1:0] wire_d36_65;
	wire [WIDTH-1:0] wire_d36_66;
	wire [WIDTH-1:0] wire_d36_67;
	wire [WIDTH-1:0] wire_d36_68;
	wire [WIDTH-1:0] wire_d36_69;
	wire [WIDTH-1:0] wire_d36_70;
	wire [WIDTH-1:0] wire_d36_71;
	wire [WIDTH-1:0] wire_d36_72;
	wire [WIDTH-1:0] wire_d36_73;
	wire [WIDTH-1:0] wire_d36_74;
	wire [WIDTH-1:0] wire_d36_75;
	wire [WIDTH-1:0] wire_d36_76;
	wire [WIDTH-1:0] wire_d36_77;
	wire [WIDTH-1:0] wire_d36_78;
	wire [WIDTH-1:0] wire_d36_79;
	wire [WIDTH-1:0] wire_d36_80;
	wire [WIDTH-1:0] wire_d36_81;
	wire [WIDTH-1:0] wire_d36_82;
	wire [WIDTH-1:0] wire_d36_83;
	wire [WIDTH-1:0] wire_d36_84;
	wire [WIDTH-1:0] wire_d36_85;
	wire [WIDTH-1:0] wire_d36_86;
	wire [WIDTH-1:0] wire_d36_87;
	wire [WIDTH-1:0] wire_d36_88;
	wire [WIDTH-1:0] wire_d36_89;
	wire [WIDTH-1:0] wire_d36_90;
	wire [WIDTH-1:0] wire_d36_91;
	wire [WIDTH-1:0] wire_d36_92;
	wire [WIDTH-1:0] wire_d36_93;
	wire [WIDTH-1:0] wire_d36_94;
	wire [WIDTH-1:0] wire_d36_95;
	wire [WIDTH-1:0] wire_d36_96;
	wire [WIDTH-1:0] wire_d36_97;
	wire [WIDTH-1:0] wire_d36_98;
	wire [WIDTH-1:0] wire_d37_0;
	wire [WIDTH-1:0] wire_d37_1;
	wire [WIDTH-1:0] wire_d37_2;
	wire [WIDTH-1:0] wire_d37_3;
	wire [WIDTH-1:0] wire_d37_4;
	wire [WIDTH-1:0] wire_d37_5;
	wire [WIDTH-1:0] wire_d37_6;
	wire [WIDTH-1:0] wire_d37_7;
	wire [WIDTH-1:0] wire_d37_8;
	wire [WIDTH-1:0] wire_d37_9;
	wire [WIDTH-1:0] wire_d37_10;
	wire [WIDTH-1:0] wire_d37_11;
	wire [WIDTH-1:0] wire_d37_12;
	wire [WIDTH-1:0] wire_d37_13;
	wire [WIDTH-1:0] wire_d37_14;
	wire [WIDTH-1:0] wire_d37_15;
	wire [WIDTH-1:0] wire_d37_16;
	wire [WIDTH-1:0] wire_d37_17;
	wire [WIDTH-1:0] wire_d37_18;
	wire [WIDTH-1:0] wire_d37_19;
	wire [WIDTH-1:0] wire_d37_20;
	wire [WIDTH-1:0] wire_d37_21;
	wire [WIDTH-1:0] wire_d37_22;
	wire [WIDTH-1:0] wire_d37_23;
	wire [WIDTH-1:0] wire_d37_24;
	wire [WIDTH-1:0] wire_d37_25;
	wire [WIDTH-1:0] wire_d37_26;
	wire [WIDTH-1:0] wire_d37_27;
	wire [WIDTH-1:0] wire_d37_28;
	wire [WIDTH-1:0] wire_d37_29;
	wire [WIDTH-1:0] wire_d37_30;
	wire [WIDTH-1:0] wire_d37_31;
	wire [WIDTH-1:0] wire_d37_32;
	wire [WIDTH-1:0] wire_d37_33;
	wire [WIDTH-1:0] wire_d37_34;
	wire [WIDTH-1:0] wire_d37_35;
	wire [WIDTH-1:0] wire_d37_36;
	wire [WIDTH-1:0] wire_d37_37;
	wire [WIDTH-1:0] wire_d37_38;
	wire [WIDTH-1:0] wire_d37_39;
	wire [WIDTH-1:0] wire_d37_40;
	wire [WIDTH-1:0] wire_d37_41;
	wire [WIDTH-1:0] wire_d37_42;
	wire [WIDTH-1:0] wire_d37_43;
	wire [WIDTH-1:0] wire_d37_44;
	wire [WIDTH-1:0] wire_d37_45;
	wire [WIDTH-1:0] wire_d37_46;
	wire [WIDTH-1:0] wire_d37_47;
	wire [WIDTH-1:0] wire_d37_48;
	wire [WIDTH-1:0] wire_d37_49;
	wire [WIDTH-1:0] wire_d37_50;
	wire [WIDTH-1:0] wire_d37_51;
	wire [WIDTH-1:0] wire_d37_52;
	wire [WIDTH-1:0] wire_d37_53;
	wire [WIDTH-1:0] wire_d37_54;
	wire [WIDTH-1:0] wire_d37_55;
	wire [WIDTH-1:0] wire_d37_56;
	wire [WIDTH-1:0] wire_d37_57;
	wire [WIDTH-1:0] wire_d37_58;
	wire [WIDTH-1:0] wire_d37_59;
	wire [WIDTH-1:0] wire_d37_60;
	wire [WIDTH-1:0] wire_d37_61;
	wire [WIDTH-1:0] wire_d37_62;
	wire [WIDTH-1:0] wire_d37_63;
	wire [WIDTH-1:0] wire_d37_64;
	wire [WIDTH-1:0] wire_d37_65;
	wire [WIDTH-1:0] wire_d37_66;
	wire [WIDTH-1:0] wire_d37_67;
	wire [WIDTH-1:0] wire_d37_68;
	wire [WIDTH-1:0] wire_d37_69;
	wire [WIDTH-1:0] wire_d37_70;
	wire [WIDTH-1:0] wire_d37_71;
	wire [WIDTH-1:0] wire_d37_72;
	wire [WIDTH-1:0] wire_d37_73;
	wire [WIDTH-1:0] wire_d37_74;
	wire [WIDTH-1:0] wire_d37_75;
	wire [WIDTH-1:0] wire_d37_76;
	wire [WIDTH-1:0] wire_d37_77;
	wire [WIDTH-1:0] wire_d37_78;
	wire [WIDTH-1:0] wire_d37_79;
	wire [WIDTH-1:0] wire_d37_80;
	wire [WIDTH-1:0] wire_d37_81;
	wire [WIDTH-1:0] wire_d37_82;
	wire [WIDTH-1:0] wire_d37_83;
	wire [WIDTH-1:0] wire_d37_84;
	wire [WIDTH-1:0] wire_d37_85;
	wire [WIDTH-1:0] wire_d37_86;
	wire [WIDTH-1:0] wire_d37_87;
	wire [WIDTH-1:0] wire_d37_88;
	wire [WIDTH-1:0] wire_d37_89;
	wire [WIDTH-1:0] wire_d37_90;
	wire [WIDTH-1:0] wire_d37_91;
	wire [WIDTH-1:0] wire_d37_92;
	wire [WIDTH-1:0] wire_d37_93;
	wire [WIDTH-1:0] wire_d37_94;
	wire [WIDTH-1:0] wire_d37_95;
	wire [WIDTH-1:0] wire_d37_96;
	wire [WIDTH-1:0] wire_d37_97;
	wire [WIDTH-1:0] wire_d37_98;
	wire [WIDTH-1:0] wire_d38_0;
	wire [WIDTH-1:0] wire_d38_1;
	wire [WIDTH-1:0] wire_d38_2;
	wire [WIDTH-1:0] wire_d38_3;
	wire [WIDTH-1:0] wire_d38_4;
	wire [WIDTH-1:0] wire_d38_5;
	wire [WIDTH-1:0] wire_d38_6;
	wire [WIDTH-1:0] wire_d38_7;
	wire [WIDTH-1:0] wire_d38_8;
	wire [WIDTH-1:0] wire_d38_9;
	wire [WIDTH-1:0] wire_d38_10;
	wire [WIDTH-1:0] wire_d38_11;
	wire [WIDTH-1:0] wire_d38_12;
	wire [WIDTH-1:0] wire_d38_13;
	wire [WIDTH-1:0] wire_d38_14;
	wire [WIDTH-1:0] wire_d38_15;
	wire [WIDTH-1:0] wire_d38_16;
	wire [WIDTH-1:0] wire_d38_17;
	wire [WIDTH-1:0] wire_d38_18;
	wire [WIDTH-1:0] wire_d38_19;
	wire [WIDTH-1:0] wire_d38_20;
	wire [WIDTH-1:0] wire_d38_21;
	wire [WIDTH-1:0] wire_d38_22;
	wire [WIDTH-1:0] wire_d38_23;
	wire [WIDTH-1:0] wire_d38_24;
	wire [WIDTH-1:0] wire_d38_25;
	wire [WIDTH-1:0] wire_d38_26;
	wire [WIDTH-1:0] wire_d38_27;
	wire [WIDTH-1:0] wire_d38_28;
	wire [WIDTH-1:0] wire_d38_29;
	wire [WIDTH-1:0] wire_d38_30;
	wire [WIDTH-1:0] wire_d38_31;
	wire [WIDTH-1:0] wire_d38_32;
	wire [WIDTH-1:0] wire_d38_33;
	wire [WIDTH-1:0] wire_d38_34;
	wire [WIDTH-1:0] wire_d38_35;
	wire [WIDTH-1:0] wire_d38_36;
	wire [WIDTH-1:0] wire_d38_37;
	wire [WIDTH-1:0] wire_d38_38;
	wire [WIDTH-1:0] wire_d38_39;
	wire [WIDTH-1:0] wire_d38_40;
	wire [WIDTH-1:0] wire_d38_41;
	wire [WIDTH-1:0] wire_d38_42;
	wire [WIDTH-1:0] wire_d38_43;
	wire [WIDTH-1:0] wire_d38_44;
	wire [WIDTH-1:0] wire_d38_45;
	wire [WIDTH-1:0] wire_d38_46;
	wire [WIDTH-1:0] wire_d38_47;
	wire [WIDTH-1:0] wire_d38_48;
	wire [WIDTH-1:0] wire_d38_49;
	wire [WIDTH-1:0] wire_d38_50;
	wire [WIDTH-1:0] wire_d38_51;
	wire [WIDTH-1:0] wire_d38_52;
	wire [WIDTH-1:0] wire_d38_53;
	wire [WIDTH-1:0] wire_d38_54;
	wire [WIDTH-1:0] wire_d38_55;
	wire [WIDTH-1:0] wire_d38_56;
	wire [WIDTH-1:0] wire_d38_57;
	wire [WIDTH-1:0] wire_d38_58;
	wire [WIDTH-1:0] wire_d38_59;
	wire [WIDTH-1:0] wire_d38_60;
	wire [WIDTH-1:0] wire_d38_61;
	wire [WIDTH-1:0] wire_d38_62;
	wire [WIDTH-1:0] wire_d38_63;
	wire [WIDTH-1:0] wire_d38_64;
	wire [WIDTH-1:0] wire_d38_65;
	wire [WIDTH-1:0] wire_d38_66;
	wire [WIDTH-1:0] wire_d38_67;
	wire [WIDTH-1:0] wire_d38_68;
	wire [WIDTH-1:0] wire_d38_69;
	wire [WIDTH-1:0] wire_d38_70;
	wire [WIDTH-1:0] wire_d38_71;
	wire [WIDTH-1:0] wire_d38_72;
	wire [WIDTH-1:0] wire_d38_73;
	wire [WIDTH-1:0] wire_d38_74;
	wire [WIDTH-1:0] wire_d38_75;
	wire [WIDTH-1:0] wire_d38_76;
	wire [WIDTH-1:0] wire_d38_77;
	wire [WIDTH-1:0] wire_d38_78;
	wire [WIDTH-1:0] wire_d38_79;
	wire [WIDTH-1:0] wire_d38_80;
	wire [WIDTH-1:0] wire_d38_81;
	wire [WIDTH-1:0] wire_d38_82;
	wire [WIDTH-1:0] wire_d38_83;
	wire [WIDTH-1:0] wire_d38_84;
	wire [WIDTH-1:0] wire_d38_85;
	wire [WIDTH-1:0] wire_d38_86;
	wire [WIDTH-1:0] wire_d38_87;
	wire [WIDTH-1:0] wire_d38_88;
	wire [WIDTH-1:0] wire_d38_89;
	wire [WIDTH-1:0] wire_d38_90;
	wire [WIDTH-1:0] wire_d38_91;
	wire [WIDTH-1:0] wire_d38_92;
	wire [WIDTH-1:0] wire_d38_93;
	wire [WIDTH-1:0] wire_d38_94;
	wire [WIDTH-1:0] wire_d38_95;
	wire [WIDTH-1:0] wire_d38_96;
	wire [WIDTH-1:0] wire_d38_97;
	wire [WIDTH-1:0] wire_d38_98;
	wire [WIDTH-1:0] wire_d39_0;
	wire [WIDTH-1:0] wire_d39_1;
	wire [WIDTH-1:0] wire_d39_2;
	wire [WIDTH-1:0] wire_d39_3;
	wire [WIDTH-1:0] wire_d39_4;
	wire [WIDTH-1:0] wire_d39_5;
	wire [WIDTH-1:0] wire_d39_6;
	wire [WIDTH-1:0] wire_d39_7;
	wire [WIDTH-1:0] wire_d39_8;
	wire [WIDTH-1:0] wire_d39_9;
	wire [WIDTH-1:0] wire_d39_10;
	wire [WIDTH-1:0] wire_d39_11;
	wire [WIDTH-1:0] wire_d39_12;
	wire [WIDTH-1:0] wire_d39_13;
	wire [WIDTH-1:0] wire_d39_14;
	wire [WIDTH-1:0] wire_d39_15;
	wire [WIDTH-1:0] wire_d39_16;
	wire [WIDTH-1:0] wire_d39_17;
	wire [WIDTH-1:0] wire_d39_18;
	wire [WIDTH-1:0] wire_d39_19;
	wire [WIDTH-1:0] wire_d39_20;
	wire [WIDTH-1:0] wire_d39_21;
	wire [WIDTH-1:0] wire_d39_22;
	wire [WIDTH-1:0] wire_d39_23;
	wire [WIDTH-1:0] wire_d39_24;
	wire [WIDTH-1:0] wire_d39_25;
	wire [WIDTH-1:0] wire_d39_26;
	wire [WIDTH-1:0] wire_d39_27;
	wire [WIDTH-1:0] wire_d39_28;
	wire [WIDTH-1:0] wire_d39_29;
	wire [WIDTH-1:0] wire_d39_30;
	wire [WIDTH-1:0] wire_d39_31;
	wire [WIDTH-1:0] wire_d39_32;
	wire [WIDTH-1:0] wire_d39_33;
	wire [WIDTH-1:0] wire_d39_34;
	wire [WIDTH-1:0] wire_d39_35;
	wire [WIDTH-1:0] wire_d39_36;
	wire [WIDTH-1:0] wire_d39_37;
	wire [WIDTH-1:0] wire_d39_38;
	wire [WIDTH-1:0] wire_d39_39;
	wire [WIDTH-1:0] wire_d39_40;
	wire [WIDTH-1:0] wire_d39_41;
	wire [WIDTH-1:0] wire_d39_42;
	wire [WIDTH-1:0] wire_d39_43;
	wire [WIDTH-1:0] wire_d39_44;
	wire [WIDTH-1:0] wire_d39_45;
	wire [WIDTH-1:0] wire_d39_46;
	wire [WIDTH-1:0] wire_d39_47;
	wire [WIDTH-1:0] wire_d39_48;
	wire [WIDTH-1:0] wire_d39_49;
	wire [WIDTH-1:0] wire_d39_50;
	wire [WIDTH-1:0] wire_d39_51;
	wire [WIDTH-1:0] wire_d39_52;
	wire [WIDTH-1:0] wire_d39_53;
	wire [WIDTH-1:0] wire_d39_54;
	wire [WIDTH-1:0] wire_d39_55;
	wire [WIDTH-1:0] wire_d39_56;
	wire [WIDTH-1:0] wire_d39_57;
	wire [WIDTH-1:0] wire_d39_58;
	wire [WIDTH-1:0] wire_d39_59;
	wire [WIDTH-1:0] wire_d39_60;
	wire [WIDTH-1:0] wire_d39_61;
	wire [WIDTH-1:0] wire_d39_62;
	wire [WIDTH-1:0] wire_d39_63;
	wire [WIDTH-1:0] wire_d39_64;
	wire [WIDTH-1:0] wire_d39_65;
	wire [WIDTH-1:0] wire_d39_66;
	wire [WIDTH-1:0] wire_d39_67;
	wire [WIDTH-1:0] wire_d39_68;
	wire [WIDTH-1:0] wire_d39_69;
	wire [WIDTH-1:0] wire_d39_70;
	wire [WIDTH-1:0] wire_d39_71;
	wire [WIDTH-1:0] wire_d39_72;
	wire [WIDTH-1:0] wire_d39_73;
	wire [WIDTH-1:0] wire_d39_74;
	wire [WIDTH-1:0] wire_d39_75;
	wire [WIDTH-1:0] wire_d39_76;
	wire [WIDTH-1:0] wire_d39_77;
	wire [WIDTH-1:0] wire_d39_78;
	wire [WIDTH-1:0] wire_d39_79;
	wire [WIDTH-1:0] wire_d39_80;
	wire [WIDTH-1:0] wire_d39_81;
	wire [WIDTH-1:0] wire_d39_82;
	wire [WIDTH-1:0] wire_d39_83;
	wire [WIDTH-1:0] wire_d39_84;
	wire [WIDTH-1:0] wire_d39_85;
	wire [WIDTH-1:0] wire_d39_86;
	wire [WIDTH-1:0] wire_d39_87;
	wire [WIDTH-1:0] wire_d39_88;
	wire [WIDTH-1:0] wire_d39_89;
	wire [WIDTH-1:0] wire_d39_90;
	wire [WIDTH-1:0] wire_d39_91;
	wire [WIDTH-1:0] wire_d39_92;
	wire [WIDTH-1:0] wire_d39_93;
	wire [WIDTH-1:0] wire_d39_94;
	wire [WIDTH-1:0] wire_d39_95;
	wire [WIDTH-1:0] wire_d39_96;
	wire [WIDTH-1:0] wire_d39_97;
	wire [WIDTH-1:0] wire_d39_98;
	wire [WIDTH-1:0] wire_d40_0;
	wire [WIDTH-1:0] wire_d40_1;
	wire [WIDTH-1:0] wire_d40_2;
	wire [WIDTH-1:0] wire_d40_3;
	wire [WIDTH-1:0] wire_d40_4;
	wire [WIDTH-1:0] wire_d40_5;
	wire [WIDTH-1:0] wire_d40_6;
	wire [WIDTH-1:0] wire_d40_7;
	wire [WIDTH-1:0] wire_d40_8;
	wire [WIDTH-1:0] wire_d40_9;
	wire [WIDTH-1:0] wire_d40_10;
	wire [WIDTH-1:0] wire_d40_11;
	wire [WIDTH-1:0] wire_d40_12;
	wire [WIDTH-1:0] wire_d40_13;
	wire [WIDTH-1:0] wire_d40_14;
	wire [WIDTH-1:0] wire_d40_15;
	wire [WIDTH-1:0] wire_d40_16;
	wire [WIDTH-1:0] wire_d40_17;
	wire [WIDTH-1:0] wire_d40_18;
	wire [WIDTH-1:0] wire_d40_19;
	wire [WIDTH-1:0] wire_d40_20;
	wire [WIDTH-1:0] wire_d40_21;
	wire [WIDTH-1:0] wire_d40_22;
	wire [WIDTH-1:0] wire_d40_23;
	wire [WIDTH-1:0] wire_d40_24;
	wire [WIDTH-1:0] wire_d40_25;
	wire [WIDTH-1:0] wire_d40_26;
	wire [WIDTH-1:0] wire_d40_27;
	wire [WIDTH-1:0] wire_d40_28;
	wire [WIDTH-1:0] wire_d40_29;
	wire [WIDTH-1:0] wire_d40_30;
	wire [WIDTH-1:0] wire_d40_31;
	wire [WIDTH-1:0] wire_d40_32;
	wire [WIDTH-1:0] wire_d40_33;
	wire [WIDTH-1:0] wire_d40_34;
	wire [WIDTH-1:0] wire_d40_35;
	wire [WIDTH-1:0] wire_d40_36;
	wire [WIDTH-1:0] wire_d40_37;
	wire [WIDTH-1:0] wire_d40_38;
	wire [WIDTH-1:0] wire_d40_39;
	wire [WIDTH-1:0] wire_d40_40;
	wire [WIDTH-1:0] wire_d40_41;
	wire [WIDTH-1:0] wire_d40_42;
	wire [WIDTH-1:0] wire_d40_43;
	wire [WIDTH-1:0] wire_d40_44;
	wire [WIDTH-1:0] wire_d40_45;
	wire [WIDTH-1:0] wire_d40_46;
	wire [WIDTH-1:0] wire_d40_47;
	wire [WIDTH-1:0] wire_d40_48;
	wire [WIDTH-1:0] wire_d40_49;
	wire [WIDTH-1:0] wire_d40_50;
	wire [WIDTH-1:0] wire_d40_51;
	wire [WIDTH-1:0] wire_d40_52;
	wire [WIDTH-1:0] wire_d40_53;
	wire [WIDTH-1:0] wire_d40_54;
	wire [WIDTH-1:0] wire_d40_55;
	wire [WIDTH-1:0] wire_d40_56;
	wire [WIDTH-1:0] wire_d40_57;
	wire [WIDTH-1:0] wire_d40_58;
	wire [WIDTH-1:0] wire_d40_59;
	wire [WIDTH-1:0] wire_d40_60;
	wire [WIDTH-1:0] wire_d40_61;
	wire [WIDTH-1:0] wire_d40_62;
	wire [WIDTH-1:0] wire_d40_63;
	wire [WIDTH-1:0] wire_d40_64;
	wire [WIDTH-1:0] wire_d40_65;
	wire [WIDTH-1:0] wire_d40_66;
	wire [WIDTH-1:0] wire_d40_67;
	wire [WIDTH-1:0] wire_d40_68;
	wire [WIDTH-1:0] wire_d40_69;
	wire [WIDTH-1:0] wire_d40_70;
	wire [WIDTH-1:0] wire_d40_71;
	wire [WIDTH-1:0] wire_d40_72;
	wire [WIDTH-1:0] wire_d40_73;
	wire [WIDTH-1:0] wire_d40_74;
	wire [WIDTH-1:0] wire_d40_75;
	wire [WIDTH-1:0] wire_d40_76;
	wire [WIDTH-1:0] wire_d40_77;
	wire [WIDTH-1:0] wire_d40_78;
	wire [WIDTH-1:0] wire_d40_79;
	wire [WIDTH-1:0] wire_d40_80;
	wire [WIDTH-1:0] wire_d40_81;
	wire [WIDTH-1:0] wire_d40_82;
	wire [WIDTH-1:0] wire_d40_83;
	wire [WIDTH-1:0] wire_d40_84;
	wire [WIDTH-1:0] wire_d40_85;
	wire [WIDTH-1:0] wire_d40_86;
	wire [WIDTH-1:0] wire_d40_87;
	wire [WIDTH-1:0] wire_d40_88;
	wire [WIDTH-1:0] wire_d40_89;
	wire [WIDTH-1:0] wire_d40_90;
	wire [WIDTH-1:0] wire_d40_91;
	wire [WIDTH-1:0] wire_d40_92;
	wire [WIDTH-1:0] wire_d40_93;
	wire [WIDTH-1:0] wire_d40_94;
	wire [WIDTH-1:0] wire_d40_95;
	wire [WIDTH-1:0] wire_d40_96;
	wire [WIDTH-1:0] wire_d40_97;
	wire [WIDTH-1:0] wire_d40_98;
	wire [WIDTH-1:0] wire_d41_0;
	wire [WIDTH-1:0] wire_d41_1;
	wire [WIDTH-1:0] wire_d41_2;
	wire [WIDTH-1:0] wire_d41_3;
	wire [WIDTH-1:0] wire_d41_4;
	wire [WIDTH-1:0] wire_d41_5;
	wire [WIDTH-1:0] wire_d41_6;
	wire [WIDTH-1:0] wire_d41_7;
	wire [WIDTH-1:0] wire_d41_8;
	wire [WIDTH-1:0] wire_d41_9;
	wire [WIDTH-1:0] wire_d41_10;
	wire [WIDTH-1:0] wire_d41_11;
	wire [WIDTH-1:0] wire_d41_12;
	wire [WIDTH-1:0] wire_d41_13;
	wire [WIDTH-1:0] wire_d41_14;
	wire [WIDTH-1:0] wire_d41_15;
	wire [WIDTH-1:0] wire_d41_16;
	wire [WIDTH-1:0] wire_d41_17;
	wire [WIDTH-1:0] wire_d41_18;
	wire [WIDTH-1:0] wire_d41_19;
	wire [WIDTH-1:0] wire_d41_20;
	wire [WIDTH-1:0] wire_d41_21;
	wire [WIDTH-1:0] wire_d41_22;
	wire [WIDTH-1:0] wire_d41_23;
	wire [WIDTH-1:0] wire_d41_24;
	wire [WIDTH-1:0] wire_d41_25;
	wire [WIDTH-1:0] wire_d41_26;
	wire [WIDTH-1:0] wire_d41_27;
	wire [WIDTH-1:0] wire_d41_28;
	wire [WIDTH-1:0] wire_d41_29;
	wire [WIDTH-1:0] wire_d41_30;
	wire [WIDTH-1:0] wire_d41_31;
	wire [WIDTH-1:0] wire_d41_32;
	wire [WIDTH-1:0] wire_d41_33;
	wire [WIDTH-1:0] wire_d41_34;
	wire [WIDTH-1:0] wire_d41_35;
	wire [WIDTH-1:0] wire_d41_36;
	wire [WIDTH-1:0] wire_d41_37;
	wire [WIDTH-1:0] wire_d41_38;
	wire [WIDTH-1:0] wire_d41_39;
	wire [WIDTH-1:0] wire_d41_40;
	wire [WIDTH-1:0] wire_d41_41;
	wire [WIDTH-1:0] wire_d41_42;
	wire [WIDTH-1:0] wire_d41_43;
	wire [WIDTH-1:0] wire_d41_44;
	wire [WIDTH-1:0] wire_d41_45;
	wire [WIDTH-1:0] wire_d41_46;
	wire [WIDTH-1:0] wire_d41_47;
	wire [WIDTH-1:0] wire_d41_48;
	wire [WIDTH-1:0] wire_d41_49;
	wire [WIDTH-1:0] wire_d41_50;
	wire [WIDTH-1:0] wire_d41_51;
	wire [WIDTH-1:0] wire_d41_52;
	wire [WIDTH-1:0] wire_d41_53;
	wire [WIDTH-1:0] wire_d41_54;
	wire [WIDTH-1:0] wire_d41_55;
	wire [WIDTH-1:0] wire_d41_56;
	wire [WIDTH-1:0] wire_d41_57;
	wire [WIDTH-1:0] wire_d41_58;
	wire [WIDTH-1:0] wire_d41_59;
	wire [WIDTH-1:0] wire_d41_60;
	wire [WIDTH-1:0] wire_d41_61;
	wire [WIDTH-1:0] wire_d41_62;
	wire [WIDTH-1:0] wire_d41_63;
	wire [WIDTH-1:0] wire_d41_64;
	wire [WIDTH-1:0] wire_d41_65;
	wire [WIDTH-1:0] wire_d41_66;
	wire [WIDTH-1:0] wire_d41_67;
	wire [WIDTH-1:0] wire_d41_68;
	wire [WIDTH-1:0] wire_d41_69;
	wire [WIDTH-1:0] wire_d41_70;
	wire [WIDTH-1:0] wire_d41_71;
	wire [WIDTH-1:0] wire_d41_72;
	wire [WIDTH-1:0] wire_d41_73;
	wire [WIDTH-1:0] wire_d41_74;
	wire [WIDTH-1:0] wire_d41_75;
	wire [WIDTH-1:0] wire_d41_76;
	wire [WIDTH-1:0] wire_d41_77;
	wire [WIDTH-1:0] wire_d41_78;
	wire [WIDTH-1:0] wire_d41_79;
	wire [WIDTH-1:0] wire_d41_80;
	wire [WIDTH-1:0] wire_d41_81;
	wire [WIDTH-1:0] wire_d41_82;
	wire [WIDTH-1:0] wire_d41_83;
	wire [WIDTH-1:0] wire_d41_84;
	wire [WIDTH-1:0] wire_d41_85;
	wire [WIDTH-1:0] wire_d41_86;
	wire [WIDTH-1:0] wire_d41_87;
	wire [WIDTH-1:0] wire_d41_88;
	wire [WIDTH-1:0] wire_d41_89;
	wire [WIDTH-1:0] wire_d41_90;
	wire [WIDTH-1:0] wire_d41_91;
	wire [WIDTH-1:0] wire_d41_92;
	wire [WIDTH-1:0] wire_d41_93;
	wire [WIDTH-1:0] wire_d41_94;
	wire [WIDTH-1:0] wire_d41_95;
	wire [WIDTH-1:0] wire_d41_96;
	wire [WIDTH-1:0] wire_d41_97;
	wire [WIDTH-1:0] wire_d41_98;
	wire [WIDTH-1:0] wire_d42_0;
	wire [WIDTH-1:0] wire_d42_1;
	wire [WIDTH-1:0] wire_d42_2;
	wire [WIDTH-1:0] wire_d42_3;
	wire [WIDTH-1:0] wire_d42_4;
	wire [WIDTH-1:0] wire_d42_5;
	wire [WIDTH-1:0] wire_d42_6;
	wire [WIDTH-1:0] wire_d42_7;
	wire [WIDTH-1:0] wire_d42_8;
	wire [WIDTH-1:0] wire_d42_9;
	wire [WIDTH-1:0] wire_d42_10;
	wire [WIDTH-1:0] wire_d42_11;
	wire [WIDTH-1:0] wire_d42_12;
	wire [WIDTH-1:0] wire_d42_13;
	wire [WIDTH-1:0] wire_d42_14;
	wire [WIDTH-1:0] wire_d42_15;
	wire [WIDTH-1:0] wire_d42_16;
	wire [WIDTH-1:0] wire_d42_17;
	wire [WIDTH-1:0] wire_d42_18;
	wire [WIDTH-1:0] wire_d42_19;
	wire [WIDTH-1:0] wire_d42_20;
	wire [WIDTH-1:0] wire_d42_21;
	wire [WIDTH-1:0] wire_d42_22;
	wire [WIDTH-1:0] wire_d42_23;
	wire [WIDTH-1:0] wire_d42_24;
	wire [WIDTH-1:0] wire_d42_25;
	wire [WIDTH-1:0] wire_d42_26;
	wire [WIDTH-1:0] wire_d42_27;
	wire [WIDTH-1:0] wire_d42_28;
	wire [WIDTH-1:0] wire_d42_29;
	wire [WIDTH-1:0] wire_d42_30;
	wire [WIDTH-1:0] wire_d42_31;
	wire [WIDTH-1:0] wire_d42_32;
	wire [WIDTH-1:0] wire_d42_33;
	wire [WIDTH-1:0] wire_d42_34;
	wire [WIDTH-1:0] wire_d42_35;
	wire [WIDTH-1:0] wire_d42_36;
	wire [WIDTH-1:0] wire_d42_37;
	wire [WIDTH-1:0] wire_d42_38;
	wire [WIDTH-1:0] wire_d42_39;
	wire [WIDTH-1:0] wire_d42_40;
	wire [WIDTH-1:0] wire_d42_41;
	wire [WIDTH-1:0] wire_d42_42;
	wire [WIDTH-1:0] wire_d42_43;
	wire [WIDTH-1:0] wire_d42_44;
	wire [WIDTH-1:0] wire_d42_45;
	wire [WIDTH-1:0] wire_d42_46;
	wire [WIDTH-1:0] wire_d42_47;
	wire [WIDTH-1:0] wire_d42_48;
	wire [WIDTH-1:0] wire_d42_49;
	wire [WIDTH-1:0] wire_d42_50;
	wire [WIDTH-1:0] wire_d42_51;
	wire [WIDTH-1:0] wire_d42_52;
	wire [WIDTH-1:0] wire_d42_53;
	wire [WIDTH-1:0] wire_d42_54;
	wire [WIDTH-1:0] wire_d42_55;
	wire [WIDTH-1:0] wire_d42_56;
	wire [WIDTH-1:0] wire_d42_57;
	wire [WIDTH-1:0] wire_d42_58;
	wire [WIDTH-1:0] wire_d42_59;
	wire [WIDTH-1:0] wire_d42_60;
	wire [WIDTH-1:0] wire_d42_61;
	wire [WIDTH-1:0] wire_d42_62;
	wire [WIDTH-1:0] wire_d42_63;
	wire [WIDTH-1:0] wire_d42_64;
	wire [WIDTH-1:0] wire_d42_65;
	wire [WIDTH-1:0] wire_d42_66;
	wire [WIDTH-1:0] wire_d42_67;
	wire [WIDTH-1:0] wire_d42_68;
	wire [WIDTH-1:0] wire_d42_69;
	wire [WIDTH-1:0] wire_d42_70;
	wire [WIDTH-1:0] wire_d42_71;
	wire [WIDTH-1:0] wire_d42_72;
	wire [WIDTH-1:0] wire_d42_73;
	wire [WIDTH-1:0] wire_d42_74;
	wire [WIDTH-1:0] wire_d42_75;
	wire [WIDTH-1:0] wire_d42_76;
	wire [WIDTH-1:0] wire_d42_77;
	wire [WIDTH-1:0] wire_d42_78;
	wire [WIDTH-1:0] wire_d42_79;
	wire [WIDTH-1:0] wire_d42_80;
	wire [WIDTH-1:0] wire_d42_81;
	wire [WIDTH-1:0] wire_d42_82;
	wire [WIDTH-1:0] wire_d42_83;
	wire [WIDTH-1:0] wire_d42_84;
	wire [WIDTH-1:0] wire_d42_85;
	wire [WIDTH-1:0] wire_d42_86;
	wire [WIDTH-1:0] wire_d42_87;
	wire [WIDTH-1:0] wire_d42_88;
	wire [WIDTH-1:0] wire_d42_89;
	wire [WIDTH-1:0] wire_d42_90;
	wire [WIDTH-1:0] wire_d42_91;
	wire [WIDTH-1:0] wire_d42_92;
	wire [WIDTH-1:0] wire_d42_93;
	wire [WIDTH-1:0] wire_d42_94;
	wire [WIDTH-1:0] wire_d42_95;
	wire [WIDTH-1:0] wire_d42_96;
	wire [WIDTH-1:0] wire_d42_97;
	wire [WIDTH-1:0] wire_d42_98;
	wire [WIDTH-1:0] wire_d43_0;
	wire [WIDTH-1:0] wire_d43_1;
	wire [WIDTH-1:0] wire_d43_2;
	wire [WIDTH-1:0] wire_d43_3;
	wire [WIDTH-1:0] wire_d43_4;
	wire [WIDTH-1:0] wire_d43_5;
	wire [WIDTH-1:0] wire_d43_6;
	wire [WIDTH-1:0] wire_d43_7;
	wire [WIDTH-1:0] wire_d43_8;
	wire [WIDTH-1:0] wire_d43_9;
	wire [WIDTH-1:0] wire_d43_10;
	wire [WIDTH-1:0] wire_d43_11;
	wire [WIDTH-1:0] wire_d43_12;
	wire [WIDTH-1:0] wire_d43_13;
	wire [WIDTH-1:0] wire_d43_14;
	wire [WIDTH-1:0] wire_d43_15;
	wire [WIDTH-1:0] wire_d43_16;
	wire [WIDTH-1:0] wire_d43_17;
	wire [WIDTH-1:0] wire_d43_18;
	wire [WIDTH-1:0] wire_d43_19;
	wire [WIDTH-1:0] wire_d43_20;
	wire [WIDTH-1:0] wire_d43_21;
	wire [WIDTH-1:0] wire_d43_22;
	wire [WIDTH-1:0] wire_d43_23;
	wire [WIDTH-1:0] wire_d43_24;
	wire [WIDTH-1:0] wire_d43_25;
	wire [WIDTH-1:0] wire_d43_26;
	wire [WIDTH-1:0] wire_d43_27;
	wire [WIDTH-1:0] wire_d43_28;
	wire [WIDTH-1:0] wire_d43_29;
	wire [WIDTH-1:0] wire_d43_30;
	wire [WIDTH-1:0] wire_d43_31;
	wire [WIDTH-1:0] wire_d43_32;
	wire [WIDTH-1:0] wire_d43_33;
	wire [WIDTH-1:0] wire_d43_34;
	wire [WIDTH-1:0] wire_d43_35;
	wire [WIDTH-1:0] wire_d43_36;
	wire [WIDTH-1:0] wire_d43_37;
	wire [WIDTH-1:0] wire_d43_38;
	wire [WIDTH-1:0] wire_d43_39;
	wire [WIDTH-1:0] wire_d43_40;
	wire [WIDTH-1:0] wire_d43_41;
	wire [WIDTH-1:0] wire_d43_42;
	wire [WIDTH-1:0] wire_d43_43;
	wire [WIDTH-1:0] wire_d43_44;
	wire [WIDTH-1:0] wire_d43_45;
	wire [WIDTH-1:0] wire_d43_46;
	wire [WIDTH-1:0] wire_d43_47;
	wire [WIDTH-1:0] wire_d43_48;
	wire [WIDTH-1:0] wire_d43_49;
	wire [WIDTH-1:0] wire_d43_50;
	wire [WIDTH-1:0] wire_d43_51;
	wire [WIDTH-1:0] wire_d43_52;
	wire [WIDTH-1:0] wire_d43_53;
	wire [WIDTH-1:0] wire_d43_54;
	wire [WIDTH-1:0] wire_d43_55;
	wire [WIDTH-1:0] wire_d43_56;
	wire [WIDTH-1:0] wire_d43_57;
	wire [WIDTH-1:0] wire_d43_58;
	wire [WIDTH-1:0] wire_d43_59;
	wire [WIDTH-1:0] wire_d43_60;
	wire [WIDTH-1:0] wire_d43_61;
	wire [WIDTH-1:0] wire_d43_62;
	wire [WIDTH-1:0] wire_d43_63;
	wire [WIDTH-1:0] wire_d43_64;
	wire [WIDTH-1:0] wire_d43_65;
	wire [WIDTH-1:0] wire_d43_66;
	wire [WIDTH-1:0] wire_d43_67;
	wire [WIDTH-1:0] wire_d43_68;
	wire [WIDTH-1:0] wire_d43_69;
	wire [WIDTH-1:0] wire_d43_70;
	wire [WIDTH-1:0] wire_d43_71;
	wire [WIDTH-1:0] wire_d43_72;
	wire [WIDTH-1:0] wire_d43_73;
	wire [WIDTH-1:0] wire_d43_74;
	wire [WIDTH-1:0] wire_d43_75;
	wire [WIDTH-1:0] wire_d43_76;
	wire [WIDTH-1:0] wire_d43_77;
	wire [WIDTH-1:0] wire_d43_78;
	wire [WIDTH-1:0] wire_d43_79;
	wire [WIDTH-1:0] wire_d43_80;
	wire [WIDTH-1:0] wire_d43_81;
	wire [WIDTH-1:0] wire_d43_82;
	wire [WIDTH-1:0] wire_d43_83;
	wire [WIDTH-1:0] wire_d43_84;
	wire [WIDTH-1:0] wire_d43_85;
	wire [WIDTH-1:0] wire_d43_86;
	wire [WIDTH-1:0] wire_d43_87;
	wire [WIDTH-1:0] wire_d43_88;
	wire [WIDTH-1:0] wire_d43_89;
	wire [WIDTH-1:0] wire_d43_90;
	wire [WIDTH-1:0] wire_d43_91;
	wire [WIDTH-1:0] wire_d43_92;
	wire [WIDTH-1:0] wire_d43_93;
	wire [WIDTH-1:0] wire_d43_94;
	wire [WIDTH-1:0] wire_d43_95;
	wire [WIDTH-1:0] wire_d43_96;
	wire [WIDTH-1:0] wire_d43_97;
	wire [WIDTH-1:0] wire_d43_98;
	wire [WIDTH-1:0] wire_d44_0;
	wire [WIDTH-1:0] wire_d44_1;
	wire [WIDTH-1:0] wire_d44_2;
	wire [WIDTH-1:0] wire_d44_3;
	wire [WIDTH-1:0] wire_d44_4;
	wire [WIDTH-1:0] wire_d44_5;
	wire [WIDTH-1:0] wire_d44_6;
	wire [WIDTH-1:0] wire_d44_7;
	wire [WIDTH-1:0] wire_d44_8;
	wire [WIDTH-1:0] wire_d44_9;
	wire [WIDTH-1:0] wire_d44_10;
	wire [WIDTH-1:0] wire_d44_11;
	wire [WIDTH-1:0] wire_d44_12;
	wire [WIDTH-1:0] wire_d44_13;
	wire [WIDTH-1:0] wire_d44_14;
	wire [WIDTH-1:0] wire_d44_15;
	wire [WIDTH-1:0] wire_d44_16;
	wire [WIDTH-1:0] wire_d44_17;
	wire [WIDTH-1:0] wire_d44_18;
	wire [WIDTH-1:0] wire_d44_19;
	wire [WIDTH-1:0] wire_d44_20;
	wire [WIDTH-1:0] wire_d44_21;
	wire [WIDTH-1:0] wire_d44_22;
	wire [WIDTH-1:0] wire_d44_23;
	wire [WIDTH-1:0] wire_d44_24;
	wire [WIDTH-1:0] wire_d44_25;
	wire [WIDTH-1:0] wire_d44_26;
	wire [WIDTH-1:0] wire_d44_27;
	wire [WIDTH-1:0] wire_d44_28;
	wire [WIDTH-1:0] wire_d44_29;
	wire [WIDTH-1:0] wire_d44_30;
	wire [WIDTH-1:0] wire_d44_31;
	wire [WIDTH-1:0] wire_d44_32;
	wire [WIDTH-1:0] wire_d44_33;
	wire [WIDTH-1:0] wire_d44_34;
	wire [WIDTH-1:0] wire_d44_35;
	wire [WIDTH-1:0] wire_d44_36;
	wire [WIDTH-1:0] wire_d44_37;
	wire [WIDTH-1:0] wire_d44_38;
	wire [WIDTH-1:0] wire_d44_39;
	wire [WIDTH-1:0] wire_d44_40;
	wire [WIDTH-1:0] wire_d44_41;
	wire [WIDTH-1:0] wire_d44_42;
	wire [WIDTH-1:0] wire_d44_43;
	wire [WIDTH-1:0] wire_d44_44;
	wire [WIDTH-1:0] wire_d44_45;
	wire [WIDTH-1:0] wire_d44_46;
	wire [WIDTH-1:0] wire_d44_47;
	wire [WIDTH-1:0] wire_d44_48;
	wire [WIDTH-1:0] wire_d44_49;
	wire [WIDTH-1:0] wire_d44_50;
	wire [WIDTH-1:0] wire_d44_51;
	wire [WIDTH-1:0] wire_d44_52;
	wire [WIDTH-1:0] wire_d44_53;
	wire [WIDTH-1:0] wire_d44_54;
	wire [WIDTH-1:0] wire_d44_55;
	wire [WIDTH-1:0] wire_d44_56;
	wire [WIDTH-1:0] wire_d44_57;
	wire [WIDTH-1:0] wire_d44_58;
	wire [WIDTH-1:0] wire_d44_59;
	wire [WIDTH-1:0] wire_d44_60;
	wire [WIDTH-1:0] wire_d44_61;
	wire [WIDTH-1:0] wire_d44_62;
	wire [WIDTH-1:0] wire_d44_63;
	wire [WIDTH-1:0] wire_d44_64;
	wire [WIDTH-1:0] wire_d44_65;
	wire [WIDTH-1:0] wire_d44_66;
	wire [WIDTH-1:0] wire_d44_67;
	wire [WIDTH-1:0] wire_d44_68;
	wire [WIDTH-1:0] wire_d44_69;
	wire [WIDTH-1:0] wire_d44_70;
	wire [WIDTH-1:0] wire_d44_71;
	wire [WIDTH-1:0] wire_d44_72;
	wire [WIDTH-1:0] wire_d44_73;
	wire [WIDTH-1:0] wire_d44_74;
	wire [WIDTH-1:0] wire_d44_75;
	wire [WIDTH-1:0] wire_d44_76;
	wire [WIDTH-1:0] wire_d44_77;
	wire [WIDTH-1:0] wire_d44_78;
	wire [WIDTH-1:0] wire_d44_79;
	wire [WIDTH-1:0] wire_d44_80;
	wire [WIDTH-1:0] wire_d44_81;
	wire [WIDTH-1:0] wire_d44_82;
	wire [WIDTH-1:0] wire_d44_83;
	wire [WIDTH-1:0] wire_d44_84;
	wire [WIDTH-1:0] wire_d44_85;
	wire [WIDTH-1:0] wire_d44_86;
	wire [WIDTH-1:0] wire_d44_87;
	wire [WIDTH-1:0] wire_d44_88;
	wire [WIDTH-1:0] wire_d44_89;
	wire [WIDTH-1:0] wire_d44_90;
	wire [WIDTH-1:0] wire_d44_91;
	wire [WIDTH-1:0] wire_d44_92;
	wire [WIDTH-1:0] wire_d44_93;
	wire [WIDTH-1:0] wire_d44_94;
	wire [WIDTH-1:0] wire_d44_95;
	wire [WIDTH-1:0] wire_d44_96;
	wire [WIDTH-1:0] wire_d44_97;
	wire [WIDTH-1:0] wire_d44_98;
	wire [WIDTH-1:0] wire_d45_0;
	wire [WIDTH-1:0] wire_d45_1;
	wire [WIDTH-1:0] wire_d45_2;
	wire [WIDTH-1:0] wire_d45_3;
	wire [WIDTH-1:0] wire_d45_4;
	wire [WIDTH-1:0] wire_d45_5;
	wire [WIDTH-1:0] wire_d45_6;
	wire [WIDTH-1:0] wire_d45_7;
	wire [WIDTH-1:0] wire_d45_8;
	wire [WIDTH-1:0] wire_d45_9;
	wire [WIDTH-1:0] wire_d45_10;
	wire [WIDTH-1:0] wire_d45_11;
	wire [WIDTH-1:0] wire_d45_12;
	wire [WIDTH-1:0] wire_d45_13;
	wire [WIDTH-1:0] wire_d45_14;
	wire [WIDTH-1:0] wire_d45_15;
	wire [WIDTH-1:0] wire_d45_16;
	wire [WIDTH-1:0] wire_d45_17;
	wire [WIDTH-1:0] wire_d45_18;
	wire [WIDTH-1:0] wire_d45_19;
	wire [WIDTH-1:0] wire_d45_20;
	wire [WIDTH-1:0] wire_d45_21;
	wire [WIDTH-1:0] wire_d45_22;
	wire [WIDTH-1:0] wire_d45_23;
	wire [WIDTH-1:0] wire_d45_24;
	wire [WIDTH-1:0] wire_d45_25;
	wire [WIDTH-1:0] wire_d45_26;
	wire [WIDTH-1:0] wire_d45_27;
	wire [WIDTH-1:0] wire_d45_28;
	wire [WIDTH-1:0] wire_d45_29;
	wire [WIDTH-1:0] wire_d45_30;
	wire [WIDTH-1:0] wire_d45_31;
	wire [WIDTH-1:0] wire_d45_32;
	wire [WIDTH-1:0] wire_d45_33;
	wire [WIDTH-1:0] wire_d45_34;
	wire [WIDTH-1:0] wire_d45_35;
	wire [WIDTH-1:0] wire_d45_36;
	wire [WIDTH-1:0] wire_d45_37;
	wire [WIDTH-1:0] wire_d45_38;
	wire [WIDTH-1:0] wire_d45_39;
	wire [WIDTH-1:0] wire_d45_40;
	wire [WIDTH-1:0] wire_d45_41;
	wire [WIDTH-1:0] wire_d45_42;
	wire [WIDTH-1:0] wire_d45_43;
	wire [WIDTH-1:0] wire_d45_44;
	wire [WIDTH-1:0] wire_d45_45;
	wire [WIDTH-1:0] wire_d45_46;
	wire [WIDTH-1:0] wire_d45_47;
	wire [WIDTH-1:0] wire_d45_48;
	wire [WIDTH-1:0] wire_d45_49;
	wire [WIDTH-1:0] wire_d45_50;
	wire [WIDTH-1:0] wire_d45_51;
	wire [WIDTH-1:0] wire_d45_52;
	wire [WIDTH-1:0] wire_d45_53;
	wire [WIDTH-1:0] wire_d45_54;
	wire [WIDTH-1:0] wire_d45_55;
	wire [WIDTH-1:0] wire_d45_56;
	wire [WIDTH-1:0] wire_d45_57;
	wire [WIDTH-1:0] wire_d45_58;
	wire [WIDTH-1:0] wire_d45_59;
	wire [WIDTH-1:0] wire_d45_60;
	wire [WIDTH-1:0] wire_d45_61;
	wire [WIDTH-1:0] wire_d45_62;
	wire [WIDTH-1:0] wire_d45_63;
	wire [WIDTH-1:0] wire_d45_64;
	wire [WIDTH-1:0] wire_d45_65;
	wire [WIDTH-1:0] wire_d45_66;
	wire [WIDTH-1:0] wire_d45_67;
	wire [WIDTH-1:0] wire_d45_68;
	wire [WIDTH-1:0] wire_d45_69;
	wire [WIDTH-1:0] wire_d45_70;
	wire [WIDTH-1:0] wire_d45_71;
	wire [WIDTH-1:0] wire_d45_72;
	wire [WIDTH-1:0] wire_d45_73;
	wire [WIDTH-1:0] wire_d45_74;
	wire [WIDTH-1:0] wire_d45_75;
	wire [WIDTH-1:0] wire_d45_76;
	wire [WIDTH-1:0] wire_d45_77;
	wire [WIDTH-1:0] wire_d45_78;
	wire [WIDTH-1:0] wire_d45_79;
	wire [WIDTH-1:0] wire_d45_80;
	wire [WIDTH-1:0] wire_d45_81;
	wire [WIDTH-1:0] wire_d45_82;
	wire [WIDTH-1:0] wire_d45_83;
	wire [WIDTH-1:0] wire_d45_84;
	wire [WIDTH-1:0] wire_d45_85;
	wire [WIDTH-1:0] wire_d45_86;
	wire [WIDTH-1:0] wire_d45_87;
	wire [WIDTH-1:0] wire_d45_88;
	wire [WIDTH-1:0] wire_d45_89;
	wire [WIDTH-1:0] wire_d45_90;
	wire [WIDTH-1:0] wire_d45_91;
	wire [WIDTH-1:0] wire_d45_92;
	wire [WIDTH-1:0] wire_d45_93;
	wire [WIDTH-1:0] wire_d45_94;
	wire [WIDTH-1:0] wire_d45_95;
	wire [WIDTH-1:0] wire_d45_96;
	wire [WIDTH-1:0] wire_d45_97;
	wire [WIDTH-1:0] wire_d45_98;
	wire [WIDTH-1:0] wire_d46_0;
	wire [WIDTH-1:0] wire_d46_1;
	wire [WIDTH-1:0] wire_d46_2;
	wire [WIDTH-1:0] wire_d46_3;
	wire [WIDTH-1:0] wire_d46_4;
	wire [WIDTH-1:0] wire_d46_5;
	wire [WIDTH-1:0] wire_d46_6;
	wire [WIDTH-1:0] wire_d46_7;
	wire [WIDTH-1:0] wire_d46_8;
	wire [WIDTH-1:0] wire_d46_9;
	wire [WIDTH-1:0] wire_d46_10;
	wire [WIDTH-1:0] wire_d46_11;
	wire [WIDTH-1:0] wire_d46_12;
	wire [WIDTH-1:0] wire_d46_13;
	wire [WIDTH-1:0] wire_d46_14;
	wire [WIDTH-1:0] wire_d46_15;
	wire [WIDTH-1:0] wire_d46_16;
	wire [WIDTH-1:0] wire_d46_17;
	wire [WIDTH-1:0] wire_d46_18;
	wire [WIDTH-1:0] wire_d46_19;
	wire [WIDTH-1:0] wire_d46_20;
	wire [WIDTH-1:0] wire_d46_21;
	wire [WIDTH-1:0] wire_d46_22;
	wire [WIDTH-1:0] wire_d46_23;
	wire [WIDTH-1:0] wire_d46_24;
	wire [WIDTH-1:0] wire_d46_25;
	wire [WIDTH-1:0] wire_d46_26;
	wire [WIDTH-1:0] wire_d46_27;
	wire [WIDTH-1:0] wire_d46_28;
	wire [WIDTH-1:0] wire_d46_29;
	wire [WIDTH-1:0] wire_d46_30;
	wire [WIDTH-1:0] wire_d46_31;
	wire [WIDTH-1:0] wire_d46_32;
	wire [WIDTH-1:0] wire_d46_33;
	wire [WIDTH-1:0] wire_d46_34;
	wire [WIDTH-1:0] wire_d46_35;
	wire [WIDTH-1:0] wire_d46_36;
	wire [WIDTH-1:0] wire_d46_37;
	wire [WIDTH-1:0] wire_d46_38;
	wire [WIDTH-1:0] wire_d46_39;
	wire [WIDTH-1:0] wire_d46_40;
	wire [WIDTH-1:0] wire_d46_41;
	wire [WIDTH-1:0] wire_d46_42;
	wire [WIDTH-1:0] wire_d46_43;
	wire [WIDTH-1:0] wire_d46_44;
	wire [WIDTH-1:0] wire_d46_45;
	wire [WIDTH-1:0] wire_d46_46;
	wire [WIDTH-1:0] wire_d46_47;
	wire [WIDTH-1:0] wire_d46_48;
	wire [WIDTH-1:0] wire_d46_49;
	wire [WIDTH-1:0] wire_d46_50;
	wire [WIDTH-1:0] wire_d46_51;
	wire [WIDTH-1:0] wire_d46_52;
	wire [WIDTH-1:0] wire_d46_53;
	wire [WIDTH-1:0] wire_d46_54;
	wire [WIDTH-1:0] wire_d46_55;
	wire [WIDTH-1:0] wire_d46_56;
	wire [WIDTH-1:0] wire_d46_57;
	wire [WIDTH-1:0] wire_d46_58;
	wire [WIDTH-1:0] wire_d46_59;
	wire [WIDTH-1:0] wire_d46_60;
	wire [WIDTH-1:0] wire_d46_61;
	wire [WIDTH-1:0] wire_d46_62;
	wire [WIDTH-1:0] wire_d46_63;
	wire [WIDTH-1:0] wire_d46_64;
	wire [WIDTH-1:0] wire_d46_65;
	wire [WIDTH-1:0] wire_d46_66;
	wire [WIDTH-1:0] wire_d46_67;
	wire [WIDTH-1:0] wire_d46_68;
	wire [WIDTH-1:0] wire_d46_69;
	wire [WIDTH-1:0] wire_d46_70;
	wire [WIDTH-1:0] wire_d46_71;
	wire [WIDTH-1:0] wire_d46_72;
	wire [WIDTH-1:0] wire_d46_73;
	wire [WIDTH-1:0] wire_d46_74;
	wire [WIDTH-1:0] wire_d46_75;
	wire [WIDTH-1:0] wire_d46_76;
	wire [WIDTH-1:0] wire_d46_77;
	wire [WIDTH-1:0] wire_d46_78;
	wire [WIDTH-1:0] wire_d46_79;
	wire [WIDTH-1:0] wire_d46_80;
	wire [WIDTH-1:0] wire_d46_81;
	wire [WIDTH-1:0] wire_d46_82;
	wire [WIDTH-1:0] wire_d46_83;
	wire [WIDTH-1:0] wire_d46_84;
	wire [WIDTH-1:0] wire_d46_85;
	wire [WIDTH-1:0] wire_d46_86;
	wire [WIDTH-1:0] wire_d46_87;
	wire [WIDTH-1:0] wire_d46_88;
	wire [WIDTH-1:0] wire_d46_89;
	wire [WIDTH-1:0] wire_d46_90;
	wire [WIDTH-1:0] wire_d46_91;
	wire [WIDTH-1:0] wire_d46_92;
	wire [WIDTH-1:0] wire_d46_93;
	wire [WIDTH-1:0] wire_d46_94;
	wire [WIDTH-1:0] wire_d46_95;
	wire [WIDTH-1:0] wire_d46_96;
	wire [WIDTH-1:0] wire_d46_97;
	wire [WIDTH-1:0] wire_d46_98;
	wire [WIDTH-1:0] wire_d47_0;
	wire [WIDTH-1:0] wire_d47_1;
	wire [WIDTH-1:0] wire_d47_2;
	wire [WIDTH-1:0] wire_d47_3;
	wire [WIDTH-1:0] wire_d47_4;
	wire [WIDTH-1:0] wire_d47_5;
	wire [WIDTH-1:0] wire_d47_6;
	wire [WIDTH-1:0] wire_d47_7;
	wire [WIDTH-1:0] wire_d47_8;
	wire [WIDTH-1:0] wire_d47_9;
	wire [WIDTH-1:0] wire_d47_10;
	wire [WIDTH-1:0] wire_d47_11;
	wire [WIDTH-1:0] wire_d47_12;
	wire [WIDTH-1:0] wire_d47_13;
	wire [WIDTH-1:0] wire_d47_14;
	wire [WIDTH-1:0] wire_d47_15;
	wire [WIDTH-1:0] wire_d47_16;
	wire [WIDTH-1:0] wire_d47_17;
	wire [WIDTH-1:0] wire_d47_18;
	wire [WIDTH-1:0] wire_d47_19;
	wire [WIDTH-1:0] wire_d47_20;
	wire [WIDTH-1:0] wire_d47_21;
	wire [WIDTH-1:0] wire_d47_22;
	wire [WIDTH-1:0] wire_d47_23;
	wire [WIDTH-1:0] wire_d47_24;
	wire [WIDTH-1:0] wire_d47_25;
	wire [WIDTH-1:0] wire_d47_26;
	wire [WIDTH-1:0] wire_d47_27;
	wire [WIDTH-1:0] wire_d47_28;
	wire [WIDTH-1:0] wire_d47_29;
	wire [WIDTH-1:0] wire_d47_30;
	wire [WIDTH-1:0] wire_d47_31;
	wire [WIDTH-1:0] wire_d47_32;
	wire [WIDTH-1:0] wire_d47_33;
	wire [WIDTH-1:0] wire_d47_34;
	wire [WIDTH-1:0] wire_d47_35;
	wire [WIDTH-1:0] wire_d47_36;
	wire [WIDTH-1:0] wire_d47_37;
	wire [WIDTH-1:0] wire_d47_38;
	wire [WIDTH-1:0] wire_d47_39;
	wire [WIDTH-1:0] wire_d47_40;
	wire [WIDTH-1:0] wire_d47_41;
	wire [WIDTH-1:0] wire_d47_42;
	wire [WIDTH-1:0] wire_d47_43;
	wire [WIDTH-1:0] wire_d47_44;
	wire [WIDTH-1:0] wire_d47_45;
	wire [WIDTH-1:0] wire_d47_46;
	wire [WIDTH-1:0] wire_d47_47;
	wire [WIDTH-1:0] wire_d47_48;
	wire [WIDTH-1:0] wire_d47_49;
	wire [WIDTH-1:0] wire_d47_50;
	wire [WIDTH-1:0] wire_d47_51;
	wire [WIDTH-1:0] wire_d47_52;
	wire [WIDTH-1:0] wire_d47_53;
	wire [WIDTH-1:0] wire_d47_54;
	wire [WIDTH-1:0] wire_d47_55;
	wire [WIDTH-1:0] wire_d47_56;
	wire [WIDTH-1:0] wire_d47_57;
	wire [WIDTH-1:0] wire_d47_58;
	wire [WIDTH-1:0] wire_d47_59;
	wire [WIDTH-1:0] wire_d47_60;
	wire [WIDTH-1:0] wire_d47_61;
	wire [WIDTH-1:0] wire_d47_62;
	wire [WIDTH-1:0] wire_d47_63;
	wire [WIDTH-1:0] wire_d47_64;
	wire [WIDTH-1:0] wire_d47_65;
	wire [WIDTH-1:0] wire_d47_66;
	wire [WIDTH-1:0] wire_d47_67;
	wire [WIDTH-1:0] wire_d47_68;
	wire [WIDTH-1:0] wire_d47_69;
	wire [WIDTH-1:0] wire_d47_70;
	wire [WIDTH-1:0] wire_d47_71;
	wire [WIDTH-1:0] wire_d47_72;
	wire [WIDTH-1:0] wire_d47_73;
	wire [WIDTH-1:0] wire_d47_74;
	wire [WIDTH-1:0] wire_d47_75;
	wire [WIDTH-1:0] wire_d47_76;
	wire [WIDTH-1:0] wire_d47_77;
	wire [WIDTH-1:0] wire_d47_78;
	wire [WIDTH-1:0] wire_d47_79;
	wire [WIDTH-1:0] wire_d47_80;
	wire [WIDTH-1:0] wire_d47_81;
	wire [WIDTH-1:0] wire_d47_82;
	wire [WIDTH-1:0] wire_d47_83;
	wire [WIDTH-1:0] wire_d47_84;
	wire [WIDTH-1:0] wire_d47_85;
	wire [WIDTH-1:0] wire_d47_86;
	wire [WIDTH-1:0] wire_d47_87;
	wire [WIDTH-1:0] wire_d47_88;
	wire [WIDTH-1:0] wire_d47_89;
	wire [WIDTH-1:0] wire_d47_90;
	wire [WIDTH-1:0] wire_d47_91;
	wire [WIDTH-1:0] wire_d47_92;
	wire [WIDTH-1:0] wire_d47_93;
	wire [WIDTH-1:0] wire_d47_94;
	wire [WIDTH-1:0] wire_d47_95;
	wire [WIDTH-1:0] wire_d47_96;
	wire [WIDTH-1:0] wire_d47_97;
	wire [WIDTH-1:0] wire_d47_98;
	wire [WIDTH-1:0] wire_d48_0;
	wire [WIDTH-1:0] wire_d48_1;
	wire [WIDTH-1:0] wire_d48_2;
	wire [WIDTH-1:0] wire_d48_3;
	wire [WIDTH-1:0] wire_d48_4;
	wire [WIDTH-1:0] wire_d48_5;
	wire [WIDTH-1:0] wire_d48_6;
	wire [WIDTH-1:0] wire_d48_7;
	wire [WIDTH-1:0] wire_d48_8;
	wire [WIDTH-1:0] wire_d48_9;
	wire [WIDTH-1:0] wire_d48_10;
	wire [WIDTH-1:0] wire_d48_11;
	wire [WIDTH-1:0] wire_d48_12;
	wire [WIDTH-1:0] wire_d48_13;
	wire [WIDTH-1:0] wire_d48_14;
	wire [WIDTH-1:0] wire_d48_15;
	wire [WIDTH-1:0] wire_d48_16;
	wire [WIDTH-1:0] wire_d48_17;
	wire [WIDTH-1:0] wire_d48_18;
	wire [WIDTH-1:0] wire_d48_19;
	wire [WIDTH-1:0] wire_d48_20;
	wire [WIDTH-1:0] wire_d48_21;
	wire [WIDTH-1:0] wire_d48_22;
	wire [WIDTH-1:0] wire_d48_23;
	wire [WIDTH-1:0] wire_d48_24;
	wire [WIDTH-1:0] wire_d48_25;
	wire [WIDTH-1:0] wire_d48_26;
	wire [WIDTH-1:0] wire_d48_27;
	wire [WIDTH-1:0] wire_d48_28;
	wire [WIDTH-1:0] wire_d48_29;
	wire [WIDTH-1:0] wire_d48_30;
	wire [WIDTH-1:0] wire_d48_31;
	wire [WIDTH-1:0] wire_d48_32;
	wire [WIDTH-1:0] wire_d48_33;
	wire [WIDTH-1:0] wire_d48_34;
	wire [WIDTH-1:0] wire_d48_35;
	wire [WIDTH-1:0] wire_d48_36;
	wire [WIDTH-1:0] wire_d48_37;
	wire [WIDTH-1:0] wire_d48_38;
	wire [WIDTH-1:0] wire_d48_39;
	wire [WIDTH-1:0] wire_d48_40;
	wire [WIDTH-1:0] wire_d48_41;
	wire [WIDTH-1:0] wire_d48_42;
	wire [WIDTH-1:0] wire_d48_43;
	wire [WIDTH-1:0] wire_d48_44;
	wire [WIDTH-1:0] wire_d48_45;
	wire [WIDTH-1:0] wire_d48_46;
	wire [WIDTH-1:0] wire_d48_47;
	wire [WIDTH-1:0] wire_d48_48;
	wire [WIDTH-1:0] wire_d48_49;
	wire [WIDTH-1:0] wire_d48_50;
	wire [WIDTH-1:0] wire_d48_51;
	wire [WIDTH-1:0] wire_d48_52;
	wire [WIDTH-1:0] wire_d48_53;
	wire [WIDTH-1:0] wire_d48_54;
	wire [WIDTH-1:0] wire_d48_55;
	wire [WIDTH-1:0] wire_d48_56;
	wire [WIDTH-1:0] wire_d48_57;
	wire [WIDTH-1:0] wire_d48_58;
	wire [WIDTH-1:0] wire_d48_59;
	wire [WIDTH-1:0] wire_d48_60;
	wire [WIDTH-1:0] wire_d48_61;
	wire [WIDTH-1:0] wire_d48_62;
	wire [WIDTH-1:0] wire_d48_63;
	wire [WIDTH-1:0] wire_d48_64;
	wire [WIDTH-1:0] wire_d48_65;
	wire [WIDTH-1:0] wire_d48_66;
	wire [WIDTH-1:0] wire_d48_67;
	wire [WIDTH-1:0] wire_d48_68;
	wire [WIDTH-1:0] wire_d48_69;
	wire [WIDTH-1:0] wire_d48_70;
	wire [WIDTH-1:0] wire_d48_71;
	wire [WIDTH-1:0] wire_d48_72;
	wire [WIDTH-1:0] wire_d48_73;
	wire [WIDTH-1:0] wire_d48_74;
	wire [WIDTH-1:0] wire_d48_75;
	wire [WIDTH-1:0] wire_d48_76;
	wire [WIDTH-1:0] wire_d48_77;
	wire [WIDTH-1:0] wire_d48_78;
	wire [WIDTH-1:0] wire_d48_79;
	wire [WIDTH-1:0] wire_d48_80;
	wire [WIDTH-1:0] wire_d48_81;
	wire [WIDTH-1:0] wire_d48_82;
	wire [WIDTH-1:0] wire_d48_83;
	wire [WIDTH-1:0] wire_d48_84;
	wire [WIDTH-1:0] wire_d48_85;
	wire [WIDTH-1:0] wire_d48_86;
	wire [WIDTH-1:0] wire_d48_87;
	wire [WIDTH-1:0] wire_d48_88;
	wire [WIDTH-1:0] wire_d48_89;
	wire [WIDTH-1:0] wire_d48_90;
	wire [WIDTH-1:0] wire_d48_91;
	wire [WIDTH-1:0] wire_d48_92;
	wire [WIDTH-1:0] wire_d48_93;
	wire [WIDTH-1:0] wire_d48_94;
	wire [WIDTH-1:0] wire_d48_95;
	wire [WIDTH-1:0] wire_d48_96;
	wire [WIDTH-1:0] wire_d48_97;
	wire [WIDTH-1:0] wire_d48_98;
	wire [WIDTH-1:0] wire_d49_0;
	wire [WIDTH-1:0] wire_d49_1;
	wire [WIDTH-1:0] wire_d49_2;
	wire [WIDTH-1:0] wire_d49_3;
	wire [WIDTH-1:0] wire_d49_4;
	wire [WIDTH-1:0] wire_d49_5;
	wire [WIDTH-1:0] wire_d49_6;
	wire [WIDTH-1:0] wire_d49_7;
	wire [WIDTH-1:0] wire_d49_8;
	wire [WIDTH-1:0] wire_d49_9;
	wire [WIDTH-1:0] wire_d49_10;
	wire [WIDTH-1:0] wire_d49_11;
	wire [WIDTH-1:0] wire_d49_12;
	wire [WIDTH-1:0] wire_d49_13;
	wire [WIDTH-1:0] wire_d49_14;
	wire [WIDTH-1:0] wire_d49_15;
	wire [WIDTH-1:0] wire_d49_16;
	wire [WIDTH-1:0] wire_d49_17;
	wire [WIDTH-1:0] wire_d49_18;
	wire [WIDTH-1:0] wire_d49_19;
	wire [WIDTH-1:0] wire_d49_20;
	wire [WIDTH-1:0] wire_d49_21;
	wire [WIDTH-1:0] wire_d49_22;
	wire [WIDTH-1:0] wire_d49_23;
	wire [WIDTH-1:0] wire_d49_24;
	wire [WIDTH-1:0] wire_d49_25;
	wire [WIDTH-1:0] wire_d49_26;
	wire [WIDTH-1:0] wire_d49_27;
	wire [WIDTH-1:0] wire_d49_28;
	wire [WIDTH-1:0] wire_d49_29;
	wire [WIDTH-1:0] wire_d49_30;
	wire [WIDTH-1:0] wire_d49_31;
	wire [WIDTH-1:0] wire_d49_32;
	wire [WIDTH-1:0] wire_d49_33;
	wire [WIDTH-1:0] wire_d49_34;
	wire [WIDTH-1:0] wire_d49_35;
	wire [WIDTH-1:0] wire_d49_36;
	wire [WIDTH-1:0] wire_d49_37;
	wire [WIDTH-1:0] wire_d49_38;
	wire [WIDTH-1:0] wire_d49_39;
	wire [WIDTH-1:0] wire_d49_40;
	wire [WIDTH-1:0] wire_d49_41;
	wire [WIDTH-1:0] wire_d49_42;
	wire [WIDTH-1:0] wire_d49_43;
	wire [WIDTH-1:0] wire_d49_44;
	wire [WIDTH-1:0] wire_d49_45;
	wire [WIDTH-1:0] wire_d49_46;
	wire [WIDTH-1:0] wire_d49_47;
	wire [WIDTH-1:0] wire_d49_48;
	wire [WIDTH-1:0] wire_d49_49;
	wire [WIDTH-1:0] wire_d49_50;
	wire [WIDTH-1:0] wire_d49_51;
	wire [WIDTH-1:0] wire_d49_52;
	wire [WIDTH-1:0] wire_d49_53;
	wire [WIDTH-1:0] wire_d49_54;
	wire [WIDTH-1:0] wire_d49_55;
	wire [WIDTH-1:0] wire_d49_56;
	wire [WIDTH-1:0] wire_d49_57;
	wire [WIDTH-1:0] wire_d49_58;
	wire [WIDTH-1:0] wire_d49_59;
	wire [WIDTH-1:0] wire_d49_60;
	wire [WIDTH-1:0] wire_d49_61;
	wire [WIDTH-1:0] wire_d49_62;
	wire [WIDTH-1:0] wire_d49_63;
	wire [WIDTH-1:0] wire_d49_64;
	wire [WIDTH-1:0] wire_d49_65;
	wire [WIDTH-1:0] wire_d49_66;
	wire [WIDTH-1:0] wire_d49_67;
	wire [WIDTH-1:0] wire_d49_68;
	wire [WIDTH-1:0] wire_d49_69;
	wire [WIDTH-1:0] wire_d49_70;
	wire [WIDTH-1:0] wire_d49_71;
	wire [WIDTH-1:0] wire_d49_72;
	wire [WIDTH-1:0] wire_d49_73;
	wire [WIDTH-1:0] wire_d49_74;
	wire [WIDTH-1:0] wire_d49_75;
	wire [WIDTH-1:0] wire_d49_76;
	wire [WIDTH-1:0] wire_d49_77;
	wire [WIDTH-1:0] wire_d49_78;
	wire [WIDTH-1:0] wire_d49_79;
	wire [WIDTH-1:0] wire_d49_80;
	wire [WIDTH-1:0] wire_d49_81;
	wire [WIDTH-1:0] wire_d49_82;
	wire [WIDTH-1:0] wire_d49_83;
	wire [WIDTH-1:0] wire_d49_84;
	wire [WIDTH-1:0] wire_d49_85;
	wire [WIDTH-1:0] wire_d49_86;
	wire [WIDTH-1:0] wire_d49_87;
	wire [WIDTH-1:0] wire_d49_88;
	wire [WIDTH-1:0] wire_d49_89;
	wire [WIDTH-1:0] wire_d49_90;
	wire [WIDTH-1:0] wire_d49_91;
	wire [WIDTH-1:0] wire_d49_92;
	wire [WIDTH-1:0] wire_d49_93;
	wire [WIDTH-1:0] wire_d49_94;
	wire [WIDTH-1:0] wire_d49_95;
	wire [WIDTH-1:0] wire_d49_96;
	wire [WIDTH-1:0] wire_d49_97;
	wire [WIDTH-1:0] wire_d49_98;
	wire [WIDTH-1:0] wire_d50_0;
	wire [WIDTH-1:0] wire_d50_1;
	wire [WIDTH-1:0] wire_d50_2;
	wire [WIDTH-1:0] wire_d50_3;
	wire [WIDTH-1:0] wire_d50_4;
	wire [WIDTH-1:0] wire_d50_5;
	wire [WIDTH-1:0] wire_d50_6;
	wire [WIDTH-1:0] wire_d50_7;
	wire [WIDTH-1:0] wire_d50_8;
	wire [WIDTH-1:0] wire_d50_9;
	wire [WIDTH-1:0] wire_d50_10;
	wire [WIDTH-1:0] wire_d50_11;
	wire [WIDTH-1:0] wire_d50_12;
	wire [WIDTH-1:0] wire_d50_13;
	wire [WIDTH-1:0] wire_d50_14;
	wire [WIDTH-1:0] wire_d50_15;
	wire [WIDTH-1:0] wire_d50_16;
	wire [WIDTH-1:0] wire_d50_17;
	wire [WIDTH-1:0] wire_d50_18;
	wire [WIDTH-1:0] wire_d50_19;
	wire [WIDTH-1:0] wire_d50_20;
	wire [WIDTH-1:0] wire_d50_21;
	wire [WIDTH-1:0] wire_d50_22;
	wire [WIDTH-1:0] wire_d50_23;
	wire [WIDTH-1:0] wire_d50_24;
	wire [WIDTH-1:0] wire_d50_25;
	wire [WIDTH-1:0] wire_d50_26;
	wire [WIDTH-1:0] wire_d50_27;
	wire [WIDTH-1:0] wire_d50_28;
	wire [WIDTH-1:0] wire_d50_29;
	wire [WIDTH-1:0] wire_d50_30;
	wire [WIDTH-1:0] wire_d50_31;
	wire [WIDTH-1:0] wire_d50_32;
	wire [WIDTH-1:0] wire_d50_33;
	wire [WIDTH-1:0] wire_d50_34;
	wire [WIDTH-1:0] wire_d50_35;
	wire [WIDTH-1:0] wire_d50_36;
	wire [WIDTH-1:0] wire_d50_37;
	wire [WIDTH-1:0] wire_d50_38;
	wire [WIDTH-1:0] wire_d50_39;
	wire [WIDTH-1:0] wire_d50_40;
	wire [WIDTH-1:0] wire_d50_41;
	wire [WIDTH-1:0] wire_d50_42;
	wire [WIDTH-1:0] wire_d50_43;
	wire [WIDTH-1:0] wire_d50_44;
	wire [WIDTH-1:0] wire_d50_45;
	wire [WIDTH-1:0] wire_d50_46;
	wire [WIDTH-1:0] wire_d50_47;
	wire [WIDTH-1:0] wire_d50_48;
	wire [WIDTH-1:0] wire_d50_49;
	wire [WIDTH-1:0] wire_d50_50;
	wire [WIDTH-1:0] wire_d50_51;
	wire [WIDTH-1:0] wire_d50_52;
	wire [WIDTH-1:0] wire_d50_53;
	wire [WIDTH-1:0] wire_d50_54;
	wire [WIDTH-1:0] wire_d50_55;
	wire [WIDTH-1:0] wire_d50_56;
	wire [WIDTH-1:0] wire_d50_57;
	wire [WIDTH-1:0] wire_d50_58;
	wire [WIDTH-1:0] wire_d50_59;
	wire [WIDTH-1:0] wire_d50_60;
	wire [WIDTH-1:0] wire_d50_61;
	wire [WIDTH-1:0] wire_d50_62;
	wire [WIDTH-1:0] wire_d50_63;
	wire [WIDTH-1:0] wire_d50_64;
	wire [WIDTH-1:0] wire_d50_65;
	wire [WIDTH-1:0] wire_d50_66;
	wire [WIDTH-1:0] wire_d50_67;
	wire [WIDTH-1:0] wire_d50_68;
	wire [WIDTH-1:0] wire_d50_69;
	wire [WIDTH-1:0] wire_d50_70;
	wire [WIDTH-1:0] wire_d50_71;
	wire [WIDTH-1:0] wire_d50_72;
	wire [WIDTH-1:0] wire_d50_73;
	wire [WIDTH-1:0] wire_d50_74;
	wire [WIDTH-1:0] wire_d50_75;
	wire [WIDTH-1:0] wire_d50_76;
	wire [WIDTH-1:0] wire_d50_77;
	wire [WIDTH-1:0] wire_d50_78;
	wire [WIDTH-1:0] wire_d50_79;
	wire [WIDTH-1:0] wire_d50_80;
	wire [WIDTH-1:0] wire_d50_81;
	wire [WIDTH-1:0] wire_d50_82;
	wire [WIDTH-1:0] wire_d50_83;
	wire [WIDTH-1:0] wire_d50_84;
	wire [WIDTH-1:0] wire_d50_85;
	wire [WIDTH-1:0] wire_d50_86;
	wire [WIDTH-1:0] wire_d50_87;
	wire [WIDTH-1:0] wire_d50_88;
	wire [WIDTH-1:0] wire_d50_89;
	wire [WIDTH-1:0] wire_d50_90;
	wire [WIDTH-1:0] wire_d50_91;
	wire [WIDTH-1:0] wire_d50_92;
	wire [WIDTH-1:0] wire_d50_93;
	wire [WIDTH-1:0] wire_d50_94;
	wire [WIDTH-1:0] wire_d50_95;
	wire [WIDTH-1:0] wire_d50_96;
	wire [WIDTH-1:0] wire_d50_97;
	wire [WIDTH-1:0] wire_d50_98;
	wire [WIDTH-1:0] wire_d51_0;
	wire [WIDTH-1:0] wire_d51_1;
	wire [WIDTH-1:0] wire_d51_2;
	wire [WIDTH-1:0] wire_d51_3;
	wire [WIDTH-1:0] wire_d51_4;
	wire [WIDTH-1:0] wire_d51_5;
	wire [WIDTH-1:0] wire_d51_6;
	wire [WIDTH-1:0] wire_d51_7;
	wire [WIDTH-1:0] wire_d51_8;
	wire [WIDTH-1:0] wire_d51_9;
	wire [WIDTH-1:0] wire_d51_10;
	wire [WIDTH-1:0] wire_d51_11;
	wire [WIDTH-1:0] wire_d51_12;
	wire [WIDTH-1:0] wire_d51_13;
	wire [WIDTH-1:0] wire_d51_14;
	wire [WIDTH-1:0] wire_d51_15;
	wire [WIDTH-1:0] wire_d51_16;
	wire [WIDTH-1:0] wire_d51_17;
	wire [WIDTH-1:0] wire_d51_18;
	wire [WIDTH-1:0] wire_d51_19;
	wire [WIDTH-1:0] wire_d51_20;
	wire [WIDTH-1:0] wire_d51_21;
	wire [WIDTH-1:0] wire_d51_22;
	wire [WIDTH-1:0] wire_d51_23;
	wire [WIDTH-1:0] wire_d51_24;
	wire [WIDTH-1:0] wire_d51_25;
	wire [WIDTH-1:0] wire_d51_26;
	wire [WIDTH-1:0] wire_d51_27;
	wire [WIDTH-1:0] wire_d51_28;
	wire [WIDTH-1:0] wire_d51_29;
	wire [WIDTH-1:0] wire_d51_30;
	wire [WIDTH-1:0] wire_d51_31;
	wire [WIDTH-1:0] wire_d51_32;
	wire [WIDTH-1:0] wire_d51_33;
	wire [WIDTH-1:0] wire_d51_34;
	wire [WIDTH-1:0] wire_d51_35;
	wire [WIDTH-1:0] wire_d51_36;
	wire [WIDTH-1:0] wire_d51_37;
	wire [WIDTH-1:0] wire_d51_38;
	wire [WIDTH-1:0] wire_d51_39;
	wire [WIDTH-1:0] wire_d51_40;
	wire [WIDTH-1:0] wire_d51_41;
	wire [WIDTH-1:0] wire_d51_42;
	wire [WIDTH-1:0] wire_d51_43;
	wire [WIDTH-1:0] wire_d51_44;
	wire [WIDTH-1:0] wire_d51_45;
	wire [WIDTH-1:0] wire_d51_46;
	wire [WIDTH-1:0] wire_d51_47;
	wire [WIDTH-1:0] wire_d51_48;
	wire [WIDTH-1:0] wire_d51_49;
	wire [WIDTH-1:0] wire_d51_50;
	wire [WIDTH-1:0] wire_d51_51;
	wire [WIDTH-1:0] wire_d51_52;
	wire [WIDTH-1:0] wire_d51_53;
	wire [WIDTH-1:0] wire_d51_54;
	wire [WIDTH-1:0] wire_d51_55;
	wire [WIDTH-1:0] wire_d51_56;
	wire [WIDTH-1:0] wire_d51_57;
	wire [WIDTH-1:0] wire_d51_58;
	wire [WIDTH-1:0] wire_d51_59;
	wire [WIDTH-1:0] wire_d51_60;
	wire [WIDTH-1:0] wire_d51_61;
	wire [WIDTH-1:0] wire_d51_62;
	wire [WIDTH-1:0] wire_d51_63;
	wire [WIDTH-1:0] wire_d51_64;
	wire [WIDTH-1:0] wire_d51_65;
	wire [WIDTH-1:0] wire_d51_66;
	wire [WIDTH-1:0] wire_d51_67;
	wire [WIDTH-1:0] wire_d51_68;
	wire [WIDTH-1:0] wire_d51_69;
	wire [WIDTH-1:0] wire_d51_70;
	wire [WIDTH-1:0] wire_d51_71;
	wire [WIDTH-1:0] wire_d51_72;
	wire [WIDTH-1:0] wire_d51_73;
	wire [WIDTH-1:0] wire_d51_74;
	wire [WIDTH-1:0] wire_d51_75;
	wire [WIDTH-1:0] wire_d51_76;
	wire [WIDTH-1:0] wire_d51_77;
	wire [WIDTH-1:0] wire_d51_78;
	wire [WIDTH-1:0] wire_d51_79;
	wire [WIDTH-1:0] wire_d51_80;
	wire [WIDTH-1:0] wire_d51_81;
	wire [WIDTH-1:0] wire_d51_82;
	wire [WIDTH-1:0] wire_d51_83;
	wire [WIDTH-1:0] wire_d51_84;
	wire [WIDTH-1:0] wire_d51_85;
	wire [WIDTH-1:0] wire_d51_86;
	wire [WIDTH-1:0] wire_d51_87;
	wire [WIDTH-1:0] wire_d51_88;
	wire [WIDTH-1:0] wire_d51_89;
	wire [WIDTH-1:0] wire_d51_90;
	wire [WIDTH-1:0] wire_d51_91;
	wire [WIDTH-1:0] wire_d51_92;
	wire [WIDTH-1:0] wire_d51_93;
	wire [WIDTH-1:0] wire_d51_94;
	wire [WIDTH-1:0] wire_d51_95;
	wire [WIDTH-1:0] wire_d51_96;
	wire [WIDTH-1:0] wire_d51_97;
	wire [WIDTH-1:0] wire_d51_98;
	wire [WIDTH-1:0] wire_d52_0;
	wire [WIDTH-1:0] wire_d52_1;
	wire [WIDTH-1:0] wire_d52_2;
	wire [WIDTH-1:0] wire_d52_3;
	wire [WIDTH-1:0] wire_d52_4;
	wire [WIDTH-1:0] wire_d52_5;
	wire [WIDTH-1:0] wire_d52_6;
	wire [WIDTH-1:0] wire_d52_7;
	wire [WIDTH-1:0] wire_d52_8;
	wire [WIDTH-1:0] wire_d52_9;
	wire [WIDTH-1:0] wire_d52_10;
	wire [WIDTH-1:0] wire_d52_11;
	wire [WIDTH-1:0] wire_d52_12;
	wire [WIDTH-1:0] wire_d52_13;
	wire [WIDTH-1:0] wire_d52_14;
	wire [WIDTH-1:0] wire_d52_15;
	wire [WIDTH-1:0] wire_d52_16;
	wire [WIDTH-1:0] wire_d52_17;
	wire [WIDTH-1:0] wire_d52_18;
	wire [WIDTH-1:0] wire_d52_19;
	wire [WIDTH-1:0] wire_d52_20;
	wire [WIDTH-1:0] wire_d52_21;
	wire [WIDTH-1:0] wire_d52_22;
	wire [WIDTH-1:0] wire_d52_23;
	wire [WIDTH-1:0] wire_d52_24;
	wire [WIDTH-1:0] wire_d52_25;
	wire [WIDTH-1:0] wire_d52_26;
	wire [WIDTH-1:0] wire_d52_27;
	wire [WIDTH-1:0] wire_d52_28;
	wire [WIDTH-1:0] wire_d52_29;
	wire [WIDTH-1:0] wire_d52_30;
	wire [WIDTH-1:0] wire_d52_31;
	wire [WIDTH-1:0] wire_d52_32;
	wire [WIDTH-1:0] wire_d52_33;
	wire [WIDTH-1:0] wire_d52_34;
	wire [WIDTH-1:0] wire_d52_35;
	wire [WIDTH-1:0] wire_d52_36;
	wire [WIDTH-1:0] wire_d52_37;
	wire [WIDTH-1:0] wire_d52_38;
	wire [WIDTH-1:0] wire_d52_39;
	wire [WIDTH-1:0] wire_d52_40;
	wire [WIDTH-1:0] wire_d52_41;
	wire [WIDTH-1:0] wire_d52_42;
	wire [WIDTH-1:0] wire_d52_43;
	wire [WIDTH-1:0] wire_d52_44;
	wire [WIDTH-1:0] wire_d52_45;
	wire [WIDTH-1:0] wire_d52_46;
	wire [WIDTH-1:0] wire_d52_47;
	wire [WIDTH-1:0] wire_d52_48;
	wire [WIDTH-1:0] wire_d52_49;
	wire [WIDTH-1:0] wire_d52_50;
	wire [WIDTH-1:0] wire_d52_51;
	wire [WIDTH-1:0] wire_d52_52;
	wire [WIDTH-1:0] wire_d52_53;
	wire [WIDTH-1:0] wire_d52_54;
	wire [WIDTH-1:0] wire_d52_55;
	wire [WIDTH-1:0] wire_d52_56;
	wire [WIDTH-1:0] wire_d52_57;
	wire [WIDTH-1:0] wire_d52_58;
	wire [WIDTH-1:0] wire_d52_59;
	wire [WIDTH-1:0] wire_d52_60;
	wire [WIDTH-1:0] wire_d52_61;
	wire [WIDTH-1:0] wire_d52_62;
	wire [WIDTH-1:0] wire_d52_63;
	wire [WIDTH-1:0] wire_d52_64;
	wire [WIDTH-1:0] wire_d52_65;
	wire [WIDTH-1:0] wire_d52_66;
	wire [WIDTH-1:0] wire_d52_67;
	wire [WIDTH-1:0] wire_d52_68;
	wire [WIDTH-1:0] wire_d52_69;
	wire [WIDTH-1:0] wire_d52_70;
	wire [WIDTH-1:0] wire_d52_71;
	wire [WIDTH-1:0] wire_d52_72;
	wire [WIDTH-1:0] wire_d52_73;
	wire [WIDTH-1:0] wire_d52_74;
	wire [WIDTH-1:0] wire_d52_75;
	wire [WIDTH-1:0] wire_d52_76;
	wire [WIDTH-1:0] wire_d52_77;
	wire [WIDTH-1:0] wire_d52_78;
	wire [WIDTH-1:0] wire_d52_79;
	wire [WIDTH-1:0] wire_d52_80;
	wire [WIDTH-1:0] wire_d52_81;
	wire [WIDTH-1:0] wire_d52_82;
	wire [WIDTH-1:0] wire_d52_83;
	wire [WIDTH-1:0] wire_d52_84;
	wire [WIDTH-1:0] wire_d52_85;
	wire [WIDTH-1:0] wire_d52_86;
	wire [WIDTH-1:0] wire_d52_87;
	wire [WIDTH-1:0] wire_d52_88;
	wire [WIDTH-1:0] wire_d52_89;
	wire [WIDTH-1:0] wire_d52_90;
	wire [WIDTH-1:0] wire_d52_91;
	wire [WIDTH-1:0] wire_d52_92;
	wire [WIDTH-1:0] wire_d52_93;
	wire [WIDTH-1:0] wire_d52_94;
	wire [WIDTH-1:0] wire_d52_95;
	wire [WIDTH-1:0] wire_d52_96;
	wire [WIDTH-1:0] wire_d52_97;
	wire [WIDTH-1:0] wire_d52_98;
	wire [WIDTH-1:0] wire_d53_0;
	wire [WIDTH-1:0] wire_d53_1;
	wire [WIDTH-1:0] wire_d53_2;
	wire [WIDTH-1:0] wire_d53_3;
	wire [WIDTH-1:0] wire_d53_4;
	wire [WIDTH-1:0] wire_d53_5;
	wire [WIDTH-1:0] wire_d53_6;
	wire [WIDTH-1:0] wire_d53_7;
	wire [WIDTH-1:0] wire_d53_8;
	wire [WIDTH-1:0] wire_d53_9;
	wire [WIDTH-1:0] wire_d53_10;
	wire [WIDTH-1:0] wire_d53_11;
	wire [WIDTH-1:0] wire_d53_12;
	wire [WIDTH-1:0] wire_d53_13;
	wire [WIDTH-1:0] wire_d53_14;
	wire [WIDTH-1:0] wire_d53_15;
	wire [WIDTH-1:0] wire_d53_16;
	wire [WIDTH-1:0] wire_d53_17;
	wire [WIDTH-1:0] wire_d53_18;
	wire [WIDTH-1:0] wire_d53_19;
	wire [WIDTH-1:0] wire_d53_20;
	wire [WIDTH-1:0] wire_d53_21;
	wire [WIDTH-1:0] wire_d53_22;
	wire [WIDTH-1:0] wire_d53_23;
	wire [WIDTH-1:0] wire_d53_24;
	wire [WIDTH-1:0] wire_d53_25;
	wire [WIDTH-1:0] wire_d53_26;
	wire [WIDTH-1:0] wire_d53_27;
	wire [WIDTH-1:0] wire_d53_28;
	wire [WIDTH-1:0] wire_d53_29;
	wire [WIDTH-1:0] wire_d53_30;
	wire [WIDTH-1:0] wire_d53_31;
	wire [WIDTH-1:0] wire_d53_32;
	wire [WIDTH-1:0] wire_d53_33;
	wire [WIDTH-1:0] wire_d53_34;
	wire [WIDTH-1:0] wire_d53_35;
	wire [WIDTH-1:0] wire_d53_36;
	wire [WIDTH-1:0] wire_d53_37;
	wire [WIDTH-1:0] wire_d53_38;
	wire [WIDTH-1:0] wire_d53_39;
	wire [WIDTH-1:0] wire_d53_40;
	wire [WIDTH-1:0] wire_d53_41;
	wire [WIDTH-1:0] wire_d53_42;
	wire [WIDTH-1:0] wire_d53_43;
	wire [WIDTH-1:0] wire_d53_44;
	wire [WIDTH-1:0] wire_d53_45;
	wire [WIDTH-1:0] wire_d53_46;
	wire [WIDTH-1:0] wire_d53_47;
	wire [WIDTH-1:0] wire_d53_48;
	wire [WIDTH-1:0] wire_d53_49;
	wire [WIDTH-1:0] wire_d53_50;
	wire [WIDTH-1:0] wire_d53_51;
	wire [WIDTH-1:0] wire_d53_52;
	wire [WIDTH-1:0] wire_d53_53;
	wire [WIDTH-1:0] wire_d53_54;
	wire [WIDTH-1:0] wire_d53_55;
	wire [WIDTH-1:0] wire_d53_56;
	wire [WIDTH-1:0] wire_d53_57;
	wire [WIDTH-1:0] wire_d53_58;
	wire [WIDTH-1:0] wire_d53_59;
	wire [WIDTH-1:0] wire_d53_60;
	wire [WIDTH-1:0] wire_d53_61;
	wire [WIDTH-1:0] wire_d53_62;
	wire [WIDTH-1:0] wire_d53_63;
	wire [WIDTH-1:0] wire_d53_64;
	wire [WIDTH-1:0] wire_d53_65;
	wire [WIDTH-1:0] wire_d53_66;
	wire [WIDTH-1:0] wire_d53_67;
	wire [WIDTH-1:0] wire_d53_68;
	wire [WIDTH-1:0] wire_d53_69;
	wire [WIDTH-1:0] wire_d53_70;
	wire [WIDTH-1:0] wire_d53_71;
	wire [WIDTH-1:0] wire_d53_72;
	wire [WIDTH-1:0] wire_d53_73;
	wire [WIDTH-1:0] wire_d53_74;
	wire [WIDTH-1:0] wire_d53_75;
	wire [WIDTH-1:0] wire_d53_76;
	wire [WIDTH-1:0] wire_d53_77;
	wire [WIDTH-1:0] wire_d53_78;
	wire [WIDTH-1:0] wire_d53_79;
	wire [WIDTH-1:0] wire_d53_80;
	wire [WIDTH-1:0] wire_d53_81;
	wire [WIDTH-1:0] wire_d53_82;
	wire [WIDTH-1:0] wire_d53_83;
	wire [WIDTH-1:0] wire_d53_84;
	wire [WIDTH-1:0] wire_d53_85;
	wire [WIDTH-1:0] wire_d53_86;
	wire [WIDTH-1:0] wire_d53_87;
	wire [WIDTH-1:0] wire_d53_88;
	wire [WIDTH-1:0] wire_d53_89;
	wire [WIDTH-1:0] wire_d53_90;
	wire [WIDTH-1:0] wire_d53_91;
	wire [WIDTH-1:0] wire_d53_92;
	wire [WIDTH-1:0] wire_d53_93;
	wire [WIDTH-1:0] wire_d53_94;
	wire [WIDTH-1:0] wire_d53_95;
	wire [WIDTH-1:0] wire_d53_96;
	wire [WIDTH-1:0] wire_d53_97;
	wire [WIDTH-1:0] wire_d53_98;
	wire [WIDTH-1:0] wire_d54_0;
	wire [WIDTH-1:0] wire_d54_1;
	wire [WIDTH-1:0] wire_d54_2;
	wire [WIDTH-1:0] wire_d54_3;
	wire [WIDTH-1:0] wire_d54_4;
	wire [WIDTH-1:0] wire_d54_5;
	wire [WIDTH-1:0] wire_d54_6;
	wire [WIDTH-1:0] wire_d54_7;
	wire [WIDTH-1:0] wire_d54_8;
	wire [WIDTH-1:0] wire_d54_9;
	wire [WIDTH-1:0] wire_d54_10;
	wire [WIDTH-1:0] wire_d54_11;
	wire [WIDTH-1:0] wire_d54_12;
	wire [WIDTH-1:0] wire_d54_13;
	wire [WIDTH-1:0] wire_d54_14;
	wire [WIDTH-1:0] wire_d54_15;
	wire [WIDTH-1:0] wire_d54_16;
	wire [WIDTH-1:0] wire_d54_17;
	wire [WIDTH-1:0] wire_d54_18;
	wire [WIDTH-1:0] wire_d54_19;
	wire [WIDTH-1:0] wire_d54_20;
	wire [WIDTH-1:0] wire_d54_21;
	wire [WIDTH-1:0] wire_d54_22;
	wire [WIDTH-1:0] wire_d54_23;
	wire [WIDTH-1:0] wire_d54_24;
	wire [WIDTH-1:0] wire_d54_25;
	wire [WIDTH-1:0] wire_d54_26;
	wire [WIDTH-1:0] wire_d54_27;
	wire [WIDTH-1:0] wire_d54_28;
	wire [WIDTH-1:0] wire_d54_29;
	wire [WIDTH-1:0] wire_d54_30;
	wire [WIDTH-1:0] wire_d54_31;
	wire [WIDTH-1:0] wire_d54_32;
	wire [WIDTH-1:0] wire_d54_33;
	wire [WIDTH-1:0] wire_d54_34;
	wire [WIDTH-1:0] wire_d54_35;
	wire [WIDTH-1:0] wire_d54_36;
	wire [WIDTH-1:0] wire_d54_37;
	wire [WIDTH-1:0] wire_d54_38;
	wire [WIDTH-1:0] wire_d54_39;
	wire [WIDTH-1:0] wire_d54_40;
	wire [WIDTH-1:0] wire_d54_41;
	wire [WIDTH-1:0] wire_d54_42;
	wire [WIDTH-1:0] wire_d54_43;
	wire [WIDTH-1:0] wire_d54_44;
	wire [WIDTH-1:0] wire_d54_45;
	wire [WIDTH-1:0] wire_d54_46;
	wire [WIDTH-1:0] wire_d54_47;
	wire [WIDTH-1:0] wire_d54_48;
	wire [WIDTH-1:0] wire_d54_49;
	wire [WIDTH-1:0] wire_d54_50;
	wire [WIDTH-1:0] wire_d54_51;
	wire [WIDTH-1:0] wire_d54_52;
	wire [WIDTH-1:0] wire_d54_53;
	wire [WIDTH-1:0] wire_d54_54;
	wire [WIDTH-1:0] wire_d54_55;
	wire [WIDTH-1:0] wire_d54_56;
	wire [WIDTH-1:0] wire_d54_57;
	wire [WIDTH-1:0] wire_d54_58;
	wire [WIDTH-1:0] wire_d54_59;
	wire [WIDTH-1:0] wire_d54_60;
	wire [WIDTH-1:0] wire_d54_61;
	wire [WIDTH-1:0] wire_d54_62;
	wire [WIDTH-1:0] wire_d54_63;
	wire [WIDTH-1:0] wire_d54_64;
	wire [WIDTH-1:0] wire_d54_65;
	wire [WIDTH-1:0] wire_d54_66;
	wire [WIDTH-1:0] wire_d54_67;
	wire [WIDTH-1:0] wire_d54_68;
	wire [WIDTH-1:0] wire_d54_69;
	wire [WIDTH-1:0] wire_d54_70;
	wire [WIDTH-1:0] wire_d54_71;
	wire [WIDTH-1:0] wire_d54_72;
	wire [WIDTH-1:0] wire_d54_73;
	wire [WIDTH-1:0] wire_d54_74;
	wire [WIDTH-1:0] wire_d54_75;
	wire [WIDTH-1:0] wire_d54_76;
	wire [WIDTH-1:0] wire_d54_77;
	wire [WIDTH-1:0] wire_d54_78;
	wire [WIDTH-1:0] wire_d54_79;
	wire [WIDTH-1:0] wire_d54_80;
	wire [WIDTH-1:0] wire_d54_81;
	wire [WIDTH-1:0] wire_d54_82;
	wire [WIDTH-1:0] wire_d54_83;
	wire [WIDTH-1:0] wire_d54_84;
	wire [WIDTH-1:0] wire_d54_85;
	wire [WIDTH-1:0] wire_d54_86;
	wire [WIDTH-1:0] wire_d54_87;
	wire [WIDTH-1:0] wire_d54_88;
	wire [WIDTH-1:0] wire_d54_89;
	wire [WIDTH-1:0] wire_d54_90;
	wire [WIDTH-1:0] wire_d54_91;
	wire [WIDTH-1:0] wire_d54_92;
	wire [WIDTH-1:0] wire_d54_93;
	wire [WIDTH-1:0] wire_d54_94;
	wire [WIDTH-1:0] wire_d54_95;
	wire [WIDTH-1:0] wire_d54_96;
	wire [WIDTH-1:0] wire_d54_97;
	wire [WIDTH-1:0] wire_d54_98;
	wire [WIDTH-1:0] wire_d55_0;
	wire [WIDTH-1:0] wire_d55_1;
	wire [WIDTH-1:0] wire_d55_2;
	wire [WIDTH-1:0] wire_d55_3;
	wire [WIDTH-1:0] wire_d55_4;
	wire [WIDTH-1:0] wire_d55_5;
	wire [WIDTH-1:0] wire_d55_6;
	wire [WIDTH-1:0] wire_d55_7;
	wire [WIDTH-1:0] wire_d55_8;
	wire [WIDTH-1:0] wire_d55_9;
	wire [WIDTH-1:0] wire_d55_10;
	wire [WIDTH-1:0] wire_d55_11;
	wire [WIDTH-1:0] wire_d55_12;
	wire [WIDTH-1:0] wire_d55_13;
	wire [WIDTH-1:0] wire_d55_14;
	wire [WIDTH-1:0] wire_d55_15;
	wire [WIDTH-1:0] wire_d55_16;
	wire [WIDTH-1:0] wire_d55_17;
	wire [WIDTH-1:0] wire_d55_18;
	wire [WIDTH-1:0] wire_d55_19;
	wire [WIDTH-1:0] wire_d55_20;
	wire [WIDTH-1:0] wire_d55_21;
	wire [WIDTH-1:0] wire_d55_22;
	wire [WIDTH-1:0] wire_d55_23;
	wire [WIDTH-1:0] wire_d55_24;
	wire [WIDTH-1:0] wire_d55_25;
	wire [WIDTH-1:0] wire_d55_26;
	wire [WIDTH-1:0] wire_d55_27;
	wire [WIDTH-1:0] wire_d55_28;
	wire [WIDTH-1:0] wire_d55_29;
	wire [WIDTH-1:0] wire_d55_30;
	wire [WIDTH-1:0] wire_d55_31;
	wire [WIDTH-1:0] wire_d55_32;
	wire [WIDTH-1:0] wire_d55_33;
	wire [WIDTH-1:0] wire_d55_34;
	wire [WIDTH-1:0] wire_d55_35;
	wire [WIDTH-1:0] wire_d55_36;
	wire [WIDTH-1:0] wire_d55_37;
	wire [WIDTH-1:0] wire_d55_38;
	wire [WIDTH-1:0] wire_d55_39;
	wire [WIDTH-1:0] wire_d55_40;
	wire [WIDTH-1:0] wire_d55_41;
	wire [WIDTH-1:0] wire_d55_42;
	wire [WIDTH-1:0] wire_d55_43;
	wire [WIDTH-1:0] wire_d55_44;
	wire [WIDTH-1:0] wire_d55_45;
	wire [WIDTH-1:0] wire_d55_46;
	wire [WIDTH-1:0] wire_d55_47;
	wire [WIDTH-1:0] wire_d55_48;
	wire [WIDTH-1:0] wire_d55_49;
	wire [WIDTH-1:0] wire_d55_50;
	wire [WIDTH-1:0] wire_d55_51;
	wire [WIDTH-1:0] wire_d55_52;
	wire [WIDTH-1:0] wire_d55_53;
	wire [WIDTH-1:0] wire_d55_54;
	wire [WIDTH-1:0] wire_d55_55;
	wire [WIDTH-1:0] wire_d55_56;
	wire [WIDTH-1:0] wire_d55_57;
	wire [WIDTH-1:0] wire_d55_58;
	wire [WIDTH-1:0] wire_d55_59;
	wire [WIDTH-1:0] wire_d55_60;
	wire [WIDTH-1:0] wire_d55_61;
	wire [WIDTH-1:0] wire_d55_62;
	wire [WIDTH-1:0] wire_d55_63;
	wire [WIDTH-1:0] wire_d55_64;
	wire [WIDTH-1:0] wire_d55_65;
	wire [WIDTH-1:0] wire_d55_66;
	wire [WIDTH-1:0] wire_d55_67;
	wire [WIDTH-1:0] wire_d55_68;
	wire [WIDTH-1:0] wire_d55_69;
	wire [WIDTH-1:0] wire_d55_70;
	wire [WIDTH-1:0] wire_d55_71;
	wire [WIDTH-1:0] wire_d55_72;
	wire [WIDTH-1:0] wire_d55_73;
	wire [WIDTH-1:0] wire_d55_74;
	wire [WIDTH-1:0] wire_d55_75;
	wire [WIDTH-1:0] wire_d55_76;
	wire [WIDTH-1:0] wire_d55_77;
	wire [WIDTH-1:0] wire_d55_78;
	wire [WIDTH-1:0] wire_d55_79;
	wire [WIDTH-1:0] wire_d55_80;
	wire [WIDTH-1:0] wire_d55_81;
	wire [WIDTH-1:0] wire_d55_82;
	wire [WIDTH-1:0] wire_d55_83;
	wire [WIDTH-1:0] wire_d55_84;
	wire [WIDTH-1:0] wire_d55_85;
	wire [WIDTH-1:0] wire_d55_86;
	wire [WIDTH-1:0] wire_d55_87;
	wire [WIDTH-1:0] wire_d55_88;
	wire [WIDTH-1:0] wire_d55_89;
	wire [WIDTH-1:0] wire_d55_90;
	wire [WIDTH-1:0] wire_d55_91;
	wire [WIDTH-1:0] wire_d55_92;
	wire [WIDTH-1:0] wire_d55_93;
	wire [WIDTH-1:0] wire_d55_94;
	wire [WIDTH-1:0] wire_d55_95;
	wire [WIDTH-1:0] wire_d55_96;
	wire [WIDTH-1:0] wire_d55_97;
	wire [WIDTH-1:0] wire_d55_98;
	wire [WIDTH-1:0] wire_d56_0;
	wire [WIDTH-1:0] wire_d56_1;
	wire [WIDTH-1:0] wire_d56_2;
	wire [WIDTH-1:0] wire_d56_3;
	wire [WIDTH-1:0] wire_d56_4;
	wire [WIDTH-1:0] wire_d56_5;
	wire [WIDTH-1:0] wire_d56_6;
	wire [WIDTH-1:0] wire_d56_7;
	wire [WIDTH-1:0] wire_d56_8;
	wire [WIDTH-1:0] wire_d56_9;
	wire [WIDTH-1:0] wire_d56_10;
	wire [WIDTH-1:0] wire_d56_11;
	wire [WIDTH-1:0] wire_d56_12;
	wire [WIDTH-1:0] wire_d56_13;
	wire [WIDTH-1:0] wire_d56_14;
	wire [WIDTH-1:0] wire_d56_15;
	wire [WIDTH-1:0] wire_d56_16;
	wire [WIDTH-1:0] wire_d56_17;
	wire [WIDTH-1:0] wire_d56_18;
	wire [WIDTH-1:0] wire_d56_19;
	wire [WIDTH-1:0] wire_d56_20;
	wire [WIDTH-1:0] wire_d56_21;
	wire [WIDTH-1:0] wire_d56_22;
	wire [WIDTH-1:0] wire_d56_23;
	wire [WIDTH-1:0] wire_d56_24;
	wire [WIDTH-1:0] wire_d56_25;
	wire [WIDTH-1:0] wire_d56_26;
	wire [WIDTH-1:0] wire_d56_27;
	wire [WIDTH-1:0] wire_d56_28;
	wire [WIDTH-1:0] wire_d56_29;
	wire [WIDTH-1:0] wire_d56_30;
	wire [WIDTH-1:0] wire_d56_31;
	wire [WIDTH-1:0] wire_d56_32;
	wire [WIDTH-1:0] wire_d56_33;
	wire [WIDTH-1:0] wire_d56_34;
	wire [WIDTH-1:0] wire_d56_35;
	wire [WIDTH-1:0] wire_d56_36;
	wire [WIDTH-1:0] wire_d56_37;
	wire [WIDTH-1:0] wire_d56_38;
	wire [WIDTH-1:0] wire_d56_39;
	wire [WIDTH-1:0] wire_d56_40;
	wire [WIDTH-1:0] wire_d56_41;
	wire [WIDTH-1:0] wire_d56_42;
	wire [WIDTH-1:0] wire_d56_43;
	wire [WIDTH-1:0] wire_d56_44;
	wire [WIDTH-1:0] wire_d56_45;
	wire [WIDTH-1:0] wire_d56_46;
	wire [WIDTH-1:0] wire_d56_47;
	wire [WIDTH-1:0] wire_d56_48;
	wire [WIDTH-1:0] wire_d56_49;
	wire [WIDTH-1:0] wire_d56_50;
	wire [WIDTH-1:0] wire_d56_51;
	wire [WIDTH-1:0] wire_d56_52;
	wire [WIDTH-1:0] wire_d56_53;
	wire [WIDTH-1:0] wire_d56_54;
	wire [WIDTH-1:0] wire_d56_55;
	wire [WIDTH-1:0] wire_d56_56;
	wire [WIDTH-1:0] wire_d56_57;
	wire [WIDTH-1:0] wire_d56_58;
	wire [WIDTH-1:0] wire_d56_59;
	wire [WIDTH-1:0] wire_d56_60;
	wire [WIDTH-1:0] wire_d56_61;
	wire [WIDTH-1:0] wire_d56_62;
	wire [WIDTH-1:0] wire_d56_63;
	wire [WIDTH-1:0] wire_d56_64;
	wire [WIDTH-1:0] wire_d56_65;
	wire [WIDTH-1:0] wire_d56_66;
	wire [WIDTH-1:0] wire_d56_67;
	wire [WIDTH-1:0] wire_d56_68;
	wire [WIDTH-1:0] wire_d56_69;
	wire [WIDTH-1:0] wire_d56_70;
	wire [WIDTH-1:0] wire_d56_71;
	wire [WIDTH-1:0] wire_d56_72;
	wire [WIDTH-1:0] wire_d56_73;
	wire [WIDTH-1:0] wire_d56_74;
	wire [WIDTH-1:0] wire_d56_75;
	wire [WIDTH-1:0] wire_d56_76;
	wire [WIDTH-1:0] wire_d56_77;
	wire [WIDTH-1:0] wire_d56_78;
	wire [WIDTH-1:0] wire_d56_79;
	wire [WIDTH-1:0] wire_d56_80;
	wire [WIDTH-1:0] wire_d56_81;
	wire [WIDTH-1:0] wire_d56_82;
	wire [WIDTH-1:0] wire_d56_83;
	wire [WIDTH-1:0] wire_d56_84;
	wire [WIDTH-1:0] wire_d56_85;
	wire [WIDTH-1:0] wire_d56_86;
	wire [WIDTH-1:0] wire_d56_87;
	wire [WIDTH-1:0] wire_d56_88;
	wire [WIDTH-1:0] wire_d56_89;
	wire [WIDTH-1:0] wire_d56_90;
	wire [WIDTH-1:0] wire_d56_91;
	wire [WIDTH-1:0] wire_d56_92;
	wire [WIDTH-1:0] wire_d56_93;
	wire [WIDTH-1:0] wire_d56_94;
	wire [WIDTH-1:0] wire_d56_95;
	wire [WIDTH-1:0] wire_d56_96;
	wire [WIDTH-1:0] wire_d56_97;
	wire [WIDTH-1:0] wire_d56_98;
	wire [WIDTH-1:0] wire_d57_0;
	wire [WIDTH-1:0] wire_d57_1;
	wire [WIDTH-1:0] wire_d57_2;
	wire [WIDTH-1:0] wire_d57_3;
	wire [WIDTH-1:0] wire_d57_4;
	wire [WIDTH-1:0] wire_d57_5;
	wire [WIDTH-1:0] wire_d57_6;
	wire [WIDTH-1:0] wire_d57_7;
	wire [WIDTH-1:0] wire_d57_8;
	wire [WIDTH-1:0] wire_d57_9;
	wire [WIDTH-1:0] wire_d57_10;
	wire [WIDTH-1:0] wire_d57_11;
	wire [WIDTH-1:0] wire_d57_12;
	wire [WIDTH-1:0] wire_d57_13;
	wire [WIDTH-1:0] wire_d57_14;
	wire [WIDTH-1:0] wire_d57_15;
	wire [WIDTH-1:0] wire_d57_16;
	wire [WIDTH-1:0] wire_d57_17;
	wire [WIDTH-1:0] wire_d57_18;
	wire [WIDTH-1:0] wire_d57_19;
	wire [WIDTH-1:0] wire_d57_20;
	wire [WIDTH-1:0] wire_d57_21;
	wire [WIDTH-1:0] wire_d57_22;
	wire [WIDTH-1:0] wire_d57_23;
	wire [WIDTH-1:0] wire_d57_24;
	wire [WIDTH-1:0] wire_d57_25;
	wire [WIDTH-1:0] wire_d57_26;
	wire [WIDTH-1:0] wire_d57_27;
	wire [WIDTH-1:0] wire_d57_28;
	wire [WIDTH-1:0] wire_d57_29;
	wire [WIDTH-1:0] wire_d57_30;
	wire [WIDTH-1:0] wire_d57_31;
	wire [WIDTH-1:0] wire_d57_32;
	wire [WIDTH-1:0] wire_d57_33;
	wire [WIDTH-1:0] wire_d57_34;
	wire [WIDTH-1:0] wire_d57_35;
	wire [WIDTH-1:0] wire_d57_36;
	wire [WIDTH-1:0] wire_d57_37;
	wire [WIDTH-1:0] wire_d57_38;
	wire [WIDTH-1:0] wire_d57_39;
	wire [WIDTH-1:0] wire_d57_40;
	wire [WIDTH-1:0] wire_d57_41;
	wire [WIDTH-1:0] wire_d57_42;
	wire [WIDTH-1:0] wire_d57_43;
	wire [WIDTH-1:0] wire_d57_44;
	wire [WIDTH-1:0] wire_d57_45;
	wire [WIDTH-1:0] wire_d57_46;
	wire [WIDTH-1:0] wire_d57_47;
	wire [WIDTH-1:0] wire_d57_48;
	wire [WIDTH-1:0] wire_d57_49;
	wire [WIDTH-1:0] wire_d57_50;
	wire [WIDTH-1:0] wire_d57_51;
	wire [WIDTH-1:0] wire_d57_52;
	wire [WIDTH-1:0] wire_d57_53;
	wire [WIDTH-1:0] wire_d57_54;
	wire [WIDTH-1:0] wire_d57_55;
	wire [WIDTH-1:0] wire_d57_56;
	wire [WIDTH-1:0] wire_d57_57;
	wire [WIDTH-1:0] wire_d57_58;
	wire [WIDTH-1:0] wire_d57_59;
	wire [WIDTH-1:0] wire_d57_60;
	wire [WIDTH-1:0] wire_d57_61;
	wire [WIDTH-1:0] wire_d57_62;
	wire [WIDTH-1:0] wire_d57_63;
	wire [WIDTH-1:0] wire_d57_64;
	wire [WIDTH-1:0] wire_d57_65;
	wire [WIDTH-1:0] wire_d57_66;
	wire [WIDTH-1:0] wire_d57_67;
	wire [WIDTH-1:0] wire_d57_68;
	wire [WIDTH-1:0] wire_d57_69;
	wire [WIDTH-1:0] wire_d57_70;
	wire [WIDTH-1:0] wire_d57_71;
	wire [WIDTH-1:0] wire_d57_72;
	wire [WIDTH-1:0] wire_d57_73;
	wire [WIDTH-1:0] wire_d57_74;
	wire [WIDTH-1:0] wire_d57_75;
	wire [WIDTH-1:0] wire_d57_76;
	wire [WIDTH-1:0] wire_d57_77;
	wire [WIDTH-1:0] wire_d57_78;
	wire [WIDTH-1:0] wire_d57_79;
	wire [WIDTH-1:0] wire_d57_80;
	wire [WIDTH-1:0] wire_d57_81;
	wire [WIDTH-1:0] wire_d57_82;
	wire [WIDTH-1:0] wire_d57_83;
	wire [WIDTH-1:0] wire_d57_84;
	wire [WIDTH-1:0] wire_d57_85;
	wire [WIDTH-1:0] wire_d57_86;
	wire [WIDTH-1:0] wire_d57_87;
	wire [WIDTH-1:0] wire_d57_88;
	wire [WIDTH-1:0] wire_d57_89;
	wire [WIDTH-1:0] wire_d57_90;
	wire [WIDTH-1:0] wire_d57_91;
	wire [WIDTH-1:0] wire_d57_92;
	wire [WIDTH-1:0] wire_d57_93;
	wire [WIDTH-1:0] wire_d57_94;
	wire [WIDTH-1:0] wire_d57_95;
	wire [WIDTH-1:0] wire_d57_96;
	wire [WIDTH-1:0] wire_d57_97;
	wire [WIDTH-1:0] wire_d57_98;
	wire [WIDTH-1:0] wire_d58_0;
	wire [WIDTH-1:0] wire_d58_1;
	wire [WIDTH-1:0] wire_d58_2;
	wire [WIDTH-1:0] wire_d58_3;
	wire [WIDTH-1:0] wire_d58_4;
	wire [WIDTH-1:0] wire_d58_5;
	wire [WIDTH-1:0] wire_d58_6;
	wire [WIDTH-1:0] wire_d58_7;
	wire [WIDTH-1:0] wire_d58_8;
	wire [WIDTH-1:0] wire_d58_9;
	wire [WIDTH-1:0] wire_d58_10;
	wire [WIDTH-1:0] wire_d58_11;
	wire [WIDTH-1:0] wire_d58_12;
	wire [WIDTH-1:0] wire_d58_13;
	wire [WIDTH-1:0] wire_d58_14;
	wire [WIDTH-1:0] wire_d58_15;
	wire [WIDTH-1:0] wire_d58_16;
	wire [WIDTH-1:0] wire_d58_17;
	wire [WIDTH-1:0] wire_d58_18;
	wire [WIDTH-1:0] wire_d58_19;
	wire [WIDTH-1:0] wire_d58_20;
	wire [WIDTH-1:0] wire_d58_21;
	wire [WIDTH-1:0] wire_d58_22;
	wire [WIDTH-1:0] wire_d58_23;
	wire [WIDTH-1:0] wire_d58_24;
	wire [WIDTH-1:0] wire_d58_25;
	wire [WIDTH-1:0] wire_d58_26;
	wire [WIDTH-1:0] wire_d58_27;
	wire [WIDTH-1:0] wire_d58_28;
	wire [WIDTH-1:0] wire_d58_29;
	wire [WIDTH-1:0] wire_d58_30;
	wire [WIDTH-1:0] wire_d58_31;
	wire [WIDTH-1:0] wire_d58_32;
	wire [WIDTH-1:0] wire_d58_33;
	wire [WIDTH-1:0] wire_d58_34;
	wire [WIDTH-1:0] wire_d58_35;
	wire [WIDTH-1:0] wire_d58_36;
	wire [WIDTH-1:0] wire_d58_37;
	wire [WIDTH-1:0] wire_d58_38;
	wire [WIDTH-1:0] wire_d58_39;
	wire [WIDTH-1:0] wire_d58_40;
	wire [WIDTH-1:0] wire_d58_41;
	wire [WIDTH-1:0] wire_d58_42;
	wire [WIDTH-1:0] wire_d58_43;
	wire [WIDTH-1:0] wire_d58_44;
	wire [WIDTH-1:0] wire_d58_45;
	wire [WIDTH-1:0] wire_d58_46;
	wire [WIDTH-1:0] wire_d58_47;
	wire [WIDTH-1:0] wire_d58_48;
	wire [WIDTH-1:0] wire_d58_49;
	wire [WIDTH-1:0] wire_d58_50;
	wire [WIDTH-1:0] wire_d58_51;
	wire [WIDTH-1:0] wire_d58_52;
	wire [WIDTH-1:0] wire_d58_53;
	wire [WIDTH-1:0] wire_d58_54;
	wire [WIDTH-1:0] wire_d58_55;
	wire [WIDTH-1:0] wire_d58_56;
	wire [WIDTH-1:0] wire_d58_57;
	wire [WIDTH-1:0] wire_d58_58;
	wire [WIDTH-1:0] wire_d58_59;
	wire [WIDTH-1:0] wire_d58_60;
	wire [WIDTH-1:0] wire_d58_61;
	wire [WIDTH-1:0] wire_d58_62;
	wire [WIDTH-1:0] wire_d58_63;
	wire [WIDTH-1:0] wire_d58_64;
	wire [WIDTH-1:0] wire_d58_65;
	wire [WIDTH-1:0] wire_d58_66;
	wire [WIDTH-1:0] wire_d58_67;
	wire [WIDTH-1:0] wire_d58_68;
	wire [WIDTH-1:0] wire_d58_69;
	wire [WIDTH-1:0] wire_d58_70;
	wire [WIDTH-1:0] wire_d58_71;
	wire [WIDTH-1:0] wire_d58_72;
	wire [WIDTH-1:0] wire_d58_73;
	wire [WIDTH-1:0] wire_d58_74;
	wire [WIDTH-1:0] wire_d58_75;
	wire [WIDTH-1:0] wire_d58_76;
	wire [WIDTH-1:0] wire_d58_77;
	wire [WIDTH-1:0] wire_d58_78;
	wire [WIDTH-1:0] wire_d58_79;
	wire [WIDTH-1:0] wire_d58_80;
	wire [WIDTH-1:0] wire_d58_81;
	wire [WIDTH-1:0] wire_d58_82;
	wire [WIDTH-1:0] wire_d58_83;
	wire [WIDTH-1:0] wire_d58_84;
	wire [WIDTH-1:0] wire_d58_85;
	wire [WIDTH-1:0] wire_d58_86;
	wire [WIDTH-1:0] wire_d58_87;
	wire [WIDTH-1:0] wire_d58_88;
	wire [WIDTH-1:0] wire_d58_89;
	wire [WIDTH-1:0] wire_d58_90;
	wire [WIDTH-1:0] wire_d58_91;
	wire [WIDTH-1:0] wire_d58_92;
	wire [WIDTH-1:0] wire_d58_93;
	wire [WIDTH-1:0] wire_d58_94;
	wire [WIDTH-1:0] wire_d58_95;
	wire [WIDTH-1:0] wire_d58_96;
	wire [WIDTH-1:0] wire_d58_97;
	wire [WIDTH-1:0] wire_d58_98;
	wire [WIDTH-1:0] wire_d59_0;
	wire [WIDTH-1:0] wire_d59_1;
	wire [WIDTH-1:0] wire_d59_2;
	wire [WIDTH-1:0] wire_d59_3;
	wire [WIDTH-1:0] wire_d59_4;
	wire [WIDTH-1:0] wire_d59_5;
	wire [WIDTH-1:0] wire_d59_6;
	wire [WIDTH-1:0] wire_d59_7;
	wire [WIDTH-1:0] wire_d59_8;
	wire [WIDTH-1:0] wire_d59_9;
	wire [WIDTH-1:0] wire_d59_10;
	wire [WIDTH-1:0] wire_d59_11;
	wire [WIDTH-1:0] wire_d59_12;
	wire [WIDTH-1:0] wire_d59_13;
	wire [WIDTH-1:0] wire_d59_14;
	wire [WIDTH-1:0] wire_d59_15;
	wire [WIDTH-1:0] wire_d59_16;
	wire [WIDTH-1:0] wire_d59_17;
	wire [WIDTH-1:0] wire_d59_18;
	wire [WIDTH-1:0] wire_d59_19;
	wire [WIDTH-1:0] wire_d59_20;
	wire [WIDTH-1:0] wire_d59_21;
	wire [WIDTH-1:0] wire_d59_22;
	wire [WIDTH-1:0] wire_d59_23;
	wire [WIDTH-1:0] wire_d59_24;
	wire [WIDTH-1:0] wire_d59_25;
	wire [WIDTH-1:0] wire_d59_26;
	wire [WIDTH-1:0] wire_d59_27;
	wire [WIDTH-1:0] wire_d59_28;
	wire [WIDTH-1:0] wire_d59_29;
	wire [WIDTH-1:0] wire_d59_30;
	wire [WIDTH-1:0] wire_d59_31;
	wire [WIDTH-1:0] wire_d59_32;
	wire [WIDTH-1:0] wire_d59_33;
	wire [WIDTH-1:0] wire_d59_34;
	wire [WIDTH-1:0] wire_d59_35;
	wire [WIDTH-1:0] wire_d59_36;
	wire [WIDTH-1:0] wire_d59_37;
	wire [WIDTH-1:0] wire_d59_38;
	wire [WIDTH-1:0] wire_d59_39;
	wire [WIDTH-1:0] wire_d59_40;
	wire [WIDTH-1:0] wire_d59_41;
	wire [WIDTH-1:0] wire_d59_42;
	wire [WIDTH-1:0] wire_d59_43;
	wire [WIDTH-1:0] wire_d59_44;
	wire [WIDTH-1:0] wire_d59_45;
	wire [WIDTH-1:0] wire_d59_46;
	wire [WIDTH-1:0] wire_d59_47;
	wire [WIDTH-1:0] wire_d59_48;
	wire [WIDTH-1:0] wire_d59_49;
	wire [WIDTH-1:0] wire_d59_50;
	wire [WIDTH-1:0] wire_d59_51;
	wire [WIDTH-1:0] wire_d59_52;
	wire [WIDTH-1:0] wire_d59_53;
	wire [WIDTH-1:0] wire_d59_54;
	wire [WIDTH-1:0] wire_d59_55;
	wire [WIDTH-1:0] wire_d59_56;
	wire [WIDTH-1:0] wire_d59_57;
	wire [WIDTH-1:0] wire_d59_58;
	wire [WIDTH-1:0] wire_d59_59;
	wire [WIDTH-1:0] wire_d59_60;
	wire [WIDTH-1:0] wire_d59_61;
	wire [WIDTH-1:0] wire_d59_62;
	wire [WIDTH-1:0] wire_d59_63;
	wire [WIDTH-1:0] wire_d59_64;
	wire [WIDTH-1:0] wire_d59_65;
	wire [WIDTH-1:0] wire_d59_66;
	wire [WIDTH-1:0] wire_d59_67;
	wire [WIDTH-1:0] wire_d59_68;
	wire [WIDTH-1:0] wire_d59_69;
	wire [WIDTH-1:0] wire_d59_70;
	wire [WIDTH-1:0] wire_d59_71;
	wire [WIDTH-1:0] wire_d59_72;
	wire [WIDTH-1:0] wire_d59_73;
	wire [WIDTH-1:0] wire_d59_74;
	wire [WIDTH-1:0] wire_d59_75;
	wire [WIDTH-1:0] wire_d59_76;
	wire [WIDTH-1:0] wire_d59_77;
	wire [WIDTH-1:0] wire_d59_78;
	wire [WIDTH-1:0] wire_d59_79;
	wire [WIDTH-1:0] wire_d59_80;
	wire [WIDTH-1:0] wire_d59_81;
	wire [WIDTH-1:0] wire_d59_82;
	wire [WIDTH-1:0] wire_d59_83;
	wire [WIDTH-1:0] wire_d59_84;
	wire [WIDTH-1:0] wire_d59_85;
	wire [WIDTH-1:0] wire_d59_86;
	wire [WIDTH-1:0] wire_d59_87;
	wire [WIDTH-1:0] wire_d59_88;
	wire [WIDTH-1:0] wire_d59_89;
	wire [WIDTH-1:0] wire_d59_90;
	wire [WIDTH-1:0] wire_d59_91;
	wire [WIDTH-1:0] wire_d59_92;
	wire [WIDTH-1:0] wire_d59_93;
	wire [WIDTH-1:0] wire_d59_94;
	wire [WIDTH-1:0] wire_d59_95;
	wire [WIDTH-1:0] wire_d59_96;
	wire [WIDTH-1:0] wire_d59_97;
	wire [WIDTH-1:0] wire_d59_98;
	wire [WIDTH-1:0] wire_d60_0;
	wire [WIDTH-1:0] wire_d60_1;
	wire [WIDTH-1:0] wire_d60_2;
	wire [WIDTH-1:0] wire_d60_3;
	wire [WIDTH-1:0] wire_d60_4;
	wire [WIDTH-1:0] wire_d60_5;
	wire [WIDTH-1:0] wire_d60_6;
	wire [WIDTH-1:0] wire_d60_7;
	wire [WIDTH-1:0] wire_d60_8;
	wire [WIDTH-1:0] wire_d60_9;
	wire [WIDTH-1:0] wire_d60_10;
	wire [WIDTH-1:0] wire_d60_11;
	wire [WIDTH-1:0] wire_d60_12;
	wire [WIDTH-1:0] wire_d60_13;
	wire [WIDTH-1:0] wire_d60_14;
	wire [WIDTH-1:0] wire_d60_15;
	wire [WIDTH-1:0] wire_d60_16;
	wire [WIDTH-1:0] wire_d60_17;
	wire [WIDTH-1:0] wire_d60_18;
	wire [WIDTH-1:0] wire_d60_19;
	wire [WIDTH-1:0] wire_d60_20;
	wire [WIDTH-1:0] wire_d60_21;
	wire [WIDTH-1:0] wire_d60_22;
	wire [WIDTH-1:0] wire_d60_23;
	wire [WIDTH-1:0] wire_d60_24;
	wire [WIDTH-1:0] wire_d60_25;
	wire [WIDTH-1:0] wire_d60_26;
	wire [WIDTH-1:0] wire_d60_27;
	wire [WIDTH-1:0] wire_d60_28;
	wire [WIDTH-1:0] wire_d60_29;
	wire [WIDTH-1:0] wire_d60_30;
	wire [WIDTH-1:0] wire_d60_31;
	wire [WIDTH-1:0] wire_d60_32;
	wire [WIDTH-1:0] wire_d60_33;
	wire [WIDTH-1:0] wire_d60_34;
	wire [WIDTH-1:0] wire_d60_35;
	wire [WIDTH-1:0] wire_d60_36;
	wire [WIDTH-1:0] wire_d60_37;
	wire [WIDTH-1:0] wire_d60_38;
	wire [WIDTH-1:0] wire_d60_39;
	wire [WIDTH-1:0] wire_d60_40;
	wire [WIDTH-1:0] wire_d60_41;
	wire [WIDTH-1:0] wire_d60_42;
	wire [WIDTH-1:0] wire_d60_43;
	wire [WIDTH-1:0] wire_d60_44;
	wire [WIDTH-1:0] wire_d60_45;
	wire [WIDTH-1:0] wire_d60_46;
	wire [WIDTH-1:0] wire_d60_47;
	wire [WIDTH-1:0] wire_d60_48;
	wire [WIDTH-1:0] wire_d60_49;
	wire [WIDTH-1:0] wire_d60_50;
	wire [WIDTH-1:0] wire_d60_51;
	wire [WIDTH-1:0] wire_d60_52;
	wire [WIDTH-1:0] wire_d60_53;
	wire [WIDTH-1:0] wire_d60_54;
	wire [WIDTH-1:0] wire_d60_55;
	wire [WIDTH-1:0] wire_d60_56;
	wire [WIDTH-1:0] wire_d60_57;
	wire [WIDTH-1:0] wire_d60_58;
	wire [WIDTH-1:0] wire_d60_59;
	wire [WIDTH-1:0] wire_d60_60;
	wire [WIDTH-1:0] wire_d60_61;
	wire [WIDTH-1:0] wire_d60_62;
	wire [WIDTH-1:0] wire_d60_63;
	wire [WIDTH-1:0] wire_d60_64;
	wire [WIDTH-1:0] wire_d60_65;
	wire [WIDTH-1:0] wire_d60_66;
	wire [WIDTH-1:0] wire_d60_67;
	wire [WIDTH-1:0] wire_d60_68;
	wire [WIDTH-1:0] wire_d60_69;
	wire [WIDTH-1:0] wire_d60_70;
	wire [WIDTH-1:0] wire_d60_71;
	wire [WIDTH-1:0] wire_d60_72;
	wire [WIDTH-1:0] wire_d60_73;
	wire [WIDTH-1:0] wire_d60_74;
	wire [WIDTH-1:0] wire_d60_75;
	wire [WIDTH-1:0] wire_d60_76;
	wire [WIDTH-1:0] wire_d60_77;
	wire [WIDTH-1:0] wire_d60_78;
	wire [WIDTH-1:0] wire_d60_79;
	wire [WIDTH-1:0] wire_d60_80;
	wire [WIDTH-1:0] wire_d60_81;
	wire [WIDTH-1:0] wire_d60_82;
	wire [WIDTH-1:0] wire_d60_83;
	wire [WIDTH-1:0] wire_d60_84;
	wire [WIDTH-1:0] wire_d60_85;
	wire [WIDTH-1:0] wire_d60_86;
	wire [WIDTH-1:0] wire_d60_87;
	wire [WIDTH-1:0] wire_d60_88;
	wire [WIDTH-1:0] wire_d60_89;
	wire [WIDTH-1:0] wire_d60_90;
	wire [WIDTH-1:0] wire_d60_91;
	wire [WIDTH-1:0] wire_d60_92;
	wire [WIDTH-1:0] wire_d60_93;
	wire [WIDTH-1:0] wire_d60_94;
	wire [WIDTH-1:0] wire_d60_95;
	wire [WIDTH-1:0] wire_d60_96;
	wire [WIDTH-1:0] wire_d60_97;
	wire [WIDTH-1:0] wire_d60_98;
	wire [WIDTH-1:0] wire_d61_0;
	wire [WIDTH-1:0] wire_d61_1;
	wire [WIDTH-1:0] wire_d61_2;
	wire [WIDTH-1:0] wire_d61_3;
	wire [WIDTH-1:0] wire_d61_4;
	wire [WIDTH-1:0] wire_d61_5;
	wire [WIDTH-1:0] wire_d61_6;
	wire [WIDTH-1:0] wire_d61_7;
	wire [WIDTH-1:0] wire_d61_8;
	wire [WIDTH-1:0] wire_d61_9;
	wire [WIDTH-1:0] wire_d61_10;
	wire [WIDTH-1:0] wire_d61_11;
	wire [WIDTH-1:0] wire_d61_12;
	wire [WIDTH-1:0] wire_d61_13;
	wire [WIDTH-1:0] wire_d61_14;
	wire [WIDTH-1:0] wire_d61_15;
	wire [WIDTH-1:0] wire_d61_16;
	wire [WIDTH-1:0] wire_d61_17;
	wire [WIDTH-1:0] wire_d61_18;
	wire [WIDTH-1:0] wire_d61_19;
	wire [WIDTH-1:0] wire_d61_20;
	wire [WIDTH-1:0] wire_d61_21;
	wire [WIDTH-1:0] wire_d61_22;
	wire [WIDTH-1:0] wire_d61_23;
	wire [WIDTH-1:0] wire_d61_24;
	wire [WIDTH-1:0] wire_d61_25;
	wire [WIDTH-1:0] wire_d61_26;
	wire [WIDTH-1:0] wire_d61_27;
	wire [WIDTH-1:0] wire_d61_28;
	wire [WIDTH-1:0] wire_d61_29;
	wire [WIDTH-1:0] wire_d61_30;
	wire [WIDTH-1:0] wire_d61_31;
	wire [WIDTH-1:0] wire_d61_32;
	wire [WIDTH-1:0] wire_d61_33;
	wire [WIDTH-1:0] wire_d61_34;
	wire [WIDTH-1:0] wire_d61_35;
	wire [WIDTH-1:0] wire_d61_36;
	wire [WIDTH-1:0] wire_d61_37;
	wire [WIDTH-1:0] wire_d61_38;
	wire [WIDTH-1:0] wire_d61_39;
	wire [WIDTH-1:0] wire_d61_40;
	wire [WIDTH-1:0] wire_d61_41;
	wire [WIDTH-1:0] wire_d61_42;
	wire [WIDTH-1:0] wire_d61_43;
	wire [WIDTH-1:0] wire_d61_44;
	wire [WIDTH-1:0] wire_d61_45;
	wire [WIDTH-1:0] wire_d61_46;
	wire [WIDTH-1:0] wire_d61_47;
	wire [WIDTH-1:0] wire_d61_48;
	wire [WIDTH-1:0] wire_d61_49;
	wire [WIDTH-1:0] wire_d61_50;
	wire [WIDTH-1:0] wire_d61_51;
	wire [WIDTH-1:0] wire_d61_52;
	wire [WIDTH-1:0] wire_d61_53;
	wire [WIDTH-1:0] wire_d61_54;
	wire [WIDTH-1:0] wire_d61_55;
	wire [WIDTH-1:0] wire_d61_56;
	wire [WIDTH-1:0] wire_d61_57;
	wire [WIDTH-1:0] wire_d61_58;
	wire [WIDTH-1:0] wire_d61_59;
	wire [WIDTH-1:0] wire_d61_60;
	wire [WIDTH-1:0] wire_d61_61;
	wire [WIDTH-1:0] wire_d61_62;
	wire [WIDTH-1:0] wire_d61_63;
	wire [WIDTH-1:0] wire_d61_64;
	wire [WIDTH-1:0] wire_d61_65;
	wire [WIDTH-1:0] wire_d61_66;
	wire [WIDTH-1:0] wire_d61_67;
	wire [WIDTH-1:0] wire_d61_68;
	wire [WIDTH-1:0] wire_d61_69;
	wire [WIDTH-1:0] wire_d61_70;
	wire [WIDTH-1:0] wire_d61_71;
	wire [WIDTH-1:0] wire_d61_72;
	wire [WIDTH-1:0] wire_d61_73;
	wire [WIDTH-1:0] wire_d61_74;
	wire [WIDTH-1:0] wire_d61_75;
	wire [WIDTH-1:0] wire_d61_76;
	wire [WIDTH-1:0] wire_d61_77;
	wire [WIDTH-1:0] wire_d61_78;
	wire [WIDTH-1:0] wire_d61_79;
	wire [WIDTH-1:0] wire_d61_80;
	wire [WIDTH-1:0] wire_d61_81;
	wire [WIDTH-1:0] wire_d61_82;
	wire [WIDTH-1:0] wire_d61_83;
	wire [WIDTH-1:0] wire_d61_84;
	wire [WIDTH-1:0] wire_d61_85;
	wire [WIDTH-1:0] wire_d61_86;
	wire [WIDTH-1:0] wire_d61_87;
	wire [WIDTH-1:0] wire_d61_88;
	wire [WIDTH-1:0] wire_d61_89;
	wire [WIDTH-1:0] wire_d61_90;
	wire [WIDTH-1:0] wire_d61_91;
	wire [WIDTH-1:0] wire_d61_92;
	wire [WIDTH-1:0] wire_d61_93;
	wire [WIDTH-1:0] wire_d61_94;
	wire [WIDTH-1:0] wire_d61_95;
	wire [WIDTH-1:0] wire_d61_96;
	wire [WIDTH-1:0] wire_d61_97;
	wire [WIDTH-1:0] wire_d61_98;
	wire [WIDTH-1:0] wire_d62_0;
	wire [WIDTH-1:0] wire_d62_1;
	wire [WIDTH-1:0] wire_d62_2;
	wire [WIDTH-1:0] wire_d62_3;
	wire [WIDTH-1:0] wire_d62_4;
	wire [WIDTH-1:0] wire_d62_5;
	wire [WIDTH-1:0] wire_d62_6;
	wire [WIDTH-1:0] wire_d62_7;
	wire [WIDTH-1:0] wire_d62_8;
	wire [WIDTH-1:0] wire_d62_9;
	wire [WIDTH-1:0] wire_d62_10;
	wire [WIDTH-1:0] wire_d62_11;
	wire [WIDTH-1:0] wire_d62_12;
	wire [WIDTH-1:0] wire_d62_13;
	wire [WIDTH-1:0] wire_d62_14;
	wire [WIDTH-1:0] wire_d62_15;
	wire [WIDTH-1:0] wire_d62_16;
	wire [WIDTH-1:0] wire_d62_17;
	wire [WIDTH-1:0] wire_d62_18;
	wire [WIDTH-1:0] wire_d62_19;
	wire [WIDTH-1:0] wire_d62_20;
	wire [WIDTH-1:0] wire_d62_21;
	wire [WIDTH-1:0] wire_d62_22;
	wire [WIDTH-1:0] wire_d62_23;
	wire [WIDTH-1:0] wire_d62_24;
	wire [WIDTH-1:0] wire_d62_25;
	wire [WIDTH-1:0] wire_d62_26;
	wire [WIDTH-1:0] wire_d62_27;
	wire [WIDTH-1:0] wire_d62_28;
	wire [WIDTH-1:0] wire_d62_29;
	wire [WIDTH-1:0] wire_d62_30;
	wire [WIDTH-1:0] wire_d62_31;
	wire [WIDTH-1:0] wire_d62_32;
	wire [WIDTH-1:0] wire_d62_33;
	wire [WIDTH-1:0] wire_d62_34;
	wire [WIDTH-1:0] wire_d62_35;
	wire [WIDTH-1:0] wire_d62_36;
	wire [WIDTH-1:0] wire_d62_37;
	wire [WIDTH-1:0] wire_d62_38;
	wire [WIDTH-1:0] wire_d62_39;
	wire [WIDTH-1:0] wire_d62_40;
	wire [WIDTH-1:0] wire_d62_41;
	wire [WIDTH-1:0] wire_d62_42;
	wire [WIDTH-1:0] wire_d62_43;
	wire [WIDTH-1:0] wire_d62_44;
	wire [WIDTH-1:0] wire_d62_45;
	wire [WIDTH-1:0] wire_d62_46;
	wire [WIDTH-1:0] wire_d62_47;
	wire [WIDTH-1:0] wire_d62_48;
	wire [WIDTH-1:0] wire_d62_49;
	wire [WIDTH-1:0] wire_d62_50;
	wire [WIDTH-1:0] wire_d62_51;
	wire [WIDTH-1:0] wire_d62_52;
	wire [WIDTH-1:0] wire_d62_53;
	wire [WIDTH-1:0] wire_d62_54;
	wire [WIDTH-1:0] wire_d62_55;
	wire [WIDTH-1:0] wire_d62_56;
	wire [WIDTH-1:0] wire_d62_57;
	wire [WIDTH-1:0] wire_d62_58;
	wire [WIDTH-1:0] wire_d62_59;
	wire [WIDTH-1:0] wire_d62_60;
	wire [WIDTH-1:0] wire_d62_61;
	wire [WIDTH-1:0] wire_d62_62;
	wire [WIDTH-1:0] wire_d62_63;
	wire [WIDTH-1:0] wire_d62_64;
	wire [WIDTH-1:0] wire_d62_65;
	wire [WIDTH-1:0] wire_d62_66;
	wire [WIDTH-1:0] wire_d62_67;
	wire [WIDTH-1:0] wire_d62_68;
	wire [WIDTH-1:0] wire_d62_69;
	wire [WIDTH-1:0] wire_d62_70;
	wire [WIDTH-1:0] wire_d62_71;
	wire [WIDTH-1:0] wire_d62_72;
	wire [WIDTH-1:0] wire_d62_73;
	wire [WIDTH-1:0] wire_d62_74;
	wire [WIDTH-1:0] wire_d62_75;
	wire [WIDTH-1:0] wire_d62_76;
	wire [WIDTH-1:0] wire_d62_77;
	wire [WIDTH-1:0] wire_d62_78;
	wire [WIDTH-1:0] wire_d62_79;
	wire [WIDTH-1:0] wire_d62_80;
	wire [WIDTH-1:0] wire_d62_81;
	wire [WIDTH-1:0] wire_d62_82;
	wire [WIDTH-1:0] wire_d62_83;
	wire [WIDTH-1:0] wire_d62_84;
	wire [WIDTH-1:0] wire_d62_85;
	wire [WIDTH-1:0] wire_d62_86;
	wire [WIDTH-1:0] wire_d62_87;
	wire [WIDTH-1:0] wire_d62_88;
	wire [WIDTH-1:0] wire_d62_89;
	wire [WIDTH-1:0] wire_d62_90;
	wire [WIDTH-1:0] wire_d62_91;
	wire [WIDTH-1:0] wire_d62_92;
	wire [WIDTH-1:0] wire_d62_93;
	wire [WIDTH-1:0] wire_d62_94;
	wire [WIDTH-1:0] wire_d62_95;
	wire [WIDTH-1:0] wire_d62_96;
	wire [WIDTH-1:0] wire_d62_97;
	wire [WIDTH-1:0] wire_d62_98;
	wire [WIDTH-1:0] wire_d63_0;
	wire [WIDTH-1:0] wire_d63_1;
	wire [WIDTH-1:0] wire_d63_2;
	wire [WIDTH-1:0] wire_d63_3;
	wire [WIDTH-1:0] wire_d63_4;
	wire [WIDTH-1:0] wire_d63_5;
	wire [WIDTH-1:0] wire_d63_6;
	wire [WIDTH-1:0] wire_d63_7;
	wire [WIDTH-1:0] wire_d63_8;
	wire [WIDTH-1:0] wire_d63_9;
	wire [WIDTH-1:0] wire_d63_10;
	wire [WIDTH-1:0] wire_d63_11;
	wire [WIDTH-1:0] wire_d63_12;
	wire [WIDTH-1:0] wire_d63_13;
	wire [WIDTH-1:0] wire_d63_14;
	wire [WIDTH-1:0] wire_d63_15;
	wire [WIDTH-1:0] wire_d63_16;
	wire [WIDTH-1:0] wire_d63_17;
	wire [WIDTH-1:0] wire_d63_18;
	wire [WIDTH-1:0] wire_d63_19;
	wire [WIDTH-1:0] wire_d63_20;
	wire [WIDTH-1:0] wire_d63_21;
	wire [WIDTH-1:0] wire_d63_22;
	wire [WIDTH-1:0] wire_d63_23;
	wire [WIDTH-1:0] wire_d63_24;
	wire [WIDTH-1:0] wire_d63_25;
	wire [WIDTH-1:0] wire_d63_26;
	wire [WIDTH-1:0] wire_d63_27;
	wire [WIDTH-1:0] wire_d63_28;
	wire [WIDTH-1:0] wire_d63_29;
	wire [WIDTH-1:0] wire_d63_30;
	wire [WIDTH-1:0] wire_d63_31;
	wire [WIDTH-1:0] wire_d63_32;
	wire [WIDTH-1:0] wire_d63_33;
	wire [WIDTH-1:0] wire_d63_34;
	wire [WIDTH-1:0] wire_d63_35;
	wire [WIDTH-1:0] wire_d63_36;
	wire [WIDTH-1:0] wire_d63_37;
	wire [WIDTH-1:0] wire_d63_38;
	wire [WIDTH-1:0] wire_d63_39;
	wire [WIDTH-1:0] wire_d63_40;
	wire [WIDTH-1:0] wire_d63_41;
	wire [WIDTH-1:0] wire_d63_42;
	wire [WIDTH-1:0] wire_d63_43;
	wire [WIDTH-1:0] wire_d63_44;
	wire [WIDTH-1:0] wire_d63_45;
	wire [WIDTH-1:0] wire_d63_46;
	wire [WIDTH-1:0] wire_d63_47;
	wire [WIDTH-1:0] wire_d63_48;
	wire [WIDTH-1:0] wire_d63_49;
	wire [WIDTH-1:0] wire_d63_50;
	wire [WIDTH-1:0] wire_d63_51;
	wire [WIDTH-1:0] wire_d63_52;
	wire [WIDTH-1:0] wire_d63_53;
	wire [WIDTH-1:0] wire_d63_54;
	wire [WIDTH-1:0] wire_d63_55;
	wire [WIDTH-1:0] wire_d63_56;
	wire [WIDTH-1:0] wire_d63_57;
	wire [WIDTH-1:0] wire_d63_58;
	wire [WIDTH-1:0] wire_d63_59;
	wire [WIDTH-1:0] wire_d63_60;
	wire [WIDTH-1:0] wire_d63_61;
	wire [WIDTH-1:0] wire_d63_62;
	wire [WIDTH-1:0] wire_d63_63;
	wire [WIDTH-1:0] wire_d63_64;
	wire [WIDTH-1:0] wire_d63_65;
	wire [WIDTH-1:0] wire_d63_66;
	wire [WIDTH-1:0] wire_d63_67;
	wire [WIDTH-1:0] wire_d63_68;
	wire [WIDTH-1:0] wire_d63_69;
	wire [WIDTH-1:0] wire_d63_70;
	wire [WIDTH-1:0] wire_d63_71;
	wire [WIDTH-1:0] wire_d63_72;
	wire [WIDTH-1:0] wire_d63_73;
	wire [WIDTH-1:0] wire_d63_74;
	wire [WIDTH-1:0] wire_d63_75;
	wire [WIDTH-1:0] wire_d63_76;
	wire [WIDTH-1:0] wire_d63_77;
	wire [WIDTH-1:0] wire_d63_78;
	wire [WIDTH-1:0] wire_d63_79;
	wire [WIDTH-1:0] wire_d63_80;
	wire [WIDTH-1:0] wire_d63_81;
	wire [WIDTH-1:0] wire_d63_82;
	wire [WIDTH-1:0] wire_d63_83;
	wire [WIDTH-1:0] wire_d63_84;
	wire [WIDTH-1:0] wire_d63_85;
	wire [WIDTH-1:0] wire_d63_86;
	wire [WIDTH-1:0] wire_d63_87;
	wire [WIDTH-1:0] wire_d63_88;
	wire [WIDTH-1:0] wire_d63_89;
	wire [WIDTH-1:0] wire_d63_90;
	wire [WIDTH-1:0] wire_d63_91;
	wire [WIDTH-1:0] wire_d63_92;
	wire [WIDTH-1:0] wire_d63_93;
	wire [WIDTH-1:0] wire_d63_94;
	wire [WIDTH-1:0] wire_d63_95;
	wire [WIDTH-1:0] wire_d63_96;
	wire [WIDTH-1:0] wire_d63_97;
	wire [WIDTH-1:0] wire_d63_98;
	wire [WIDTH-1:0] wire_d64_0;
	wire [WIDTH-1:0] wire_d64_1;
	wire [WIDTH-1:0] wire_d64_2;
	wire [WIDTH-1:0] wire_d64_3;
	wire [WIDTH-1:0] wire_d64_4;
	wire [WIDTH-1:0] wire_d64_5;
	wire [WIDTH-1:0] wire_d64_6;
	wire [WIDTH-1:0] wire_d64_7;
	wire [WIDTH-1:0] wire_d64_8;
	wire [WIDTH-1:0] wire_d64_9;
	wire [WIDTH-1:0] wire_d64_10;
	wire [WIDTH-1:0] wire_d64_11;
	wire [WIDTH-1:0] wire_d64_12;
	wire [WIDTH-1:0] wire_d64_13;
	wire [WIDTH-1:0] wire_d64_14;
	wire [WIDTH-1:0] wire_d64_15;
	wire [WIDTH-1:0] wire_d64_16;
	wire [WIDTH-1:0] wire_d64_17;
	wire [WIDTH-1:0] wire_d64_18;
	wire [WIDTH-1:0] wire_d64_19;
	wire [WIDTH-1:0] wire_d64_20;
	wire [WIDTH-1:0] wire_d64_21;
	wire [WIDTH-1:0] wire_d64_22;
	wire [WIDTH-1:0] wire_d64_23;
	wire [WIDTH-1:0] wire_d64_24;
	wire [WIDTH-1:0] wire_d64_25;
	wire [WIDTH-1:0] wire_d64_26;
	wire [WIDTH-1:0] wire_d64_27;
	wire [WIDTH-1:0] wire_d64_28;
	wire [WIDTH-1:0] wire_d64_29;
	wire [WIDTH-1:0] wire_d64_30;
	wire [WIDTH-1:0] wire_d64_31;
	wire [WIDTH-1:0] wire_d64_32;
	wire [WIDTH-1:0] wire_d64_33;
	wire [WIDTH-1:0] wire_d64_34;
	wire [WIDTH-1:0] wire_d64_35;
	wire [WIDTH-1:0] wire_d64_36;
	wire [WIDTH-1:0] wire_d64_37;
	wire [WIDTH-1:0] wire_d64_38;
	wire [WIDTH-1:0] wire_d64_39;
	wire [WIDTH-1:0] wire_d64_40;
	wire [WIDTH-1:0] wire_d64_41;
	wire [WIDTH-1:0] wire_d64_42;
	wire [WIDTH-1:0] wire_d64_43;
	wire [WIDTH-1:0] wire_d64_44;
	wire [WIDTH-1:0] wire_d64_45;
	wire [WIDTH-1:0] wire_d64_46;
	wire [WIDTH-1:0] wire_d64_47;
	wire [WIDTH-1:0] wire_d64_48;
	wire [WIDTH-1:0] wire_d64_49;
	wire [WIDTH-1:0] wire_d64_50;
	wire [WIDTH-1:0] wire_d64_51;
	wire [WIDTH-1:0] wire_d64_52;
	wire [WIDTH-1:0] wire_d64_53;
	wire [WIDTH-1:0] wire_d64_54;
	wire [WIDTH-1:0] wire_d64_55;
	wire [WIDTH-1:0] wire_d64_56;
	wire [WIDTH-1:0] wire_d64_57;
	wire [WIDTH-1:0] wire_d64_58;
	wire [WIDTH-1:0] wire_d64_59;
	wire [WIDTH-1:0] wire_d64_60;
	wire [WIDTH-1:0] wire_d64_61;
	wire [WIDTH-1:0] wire_d64_62;
	wire [WIDTH-1:0] wire_d64_63;
	wire [WIDTH-1:0] wire_d64_64;
	wire [WIDTH-1:0] wire_d64_65;
	wire [WIDTH-1:0] wire_d64_66;
	wire [WIDTH-1:0] wire_d64_67;
	wire [WIDTH-1:0] wire_d64_68;
	wire [WIDTH-1:0] wire_d64_69;
	wire [WIDTH-1:0] wire_d64_70;
	wire [WIDTH-1:0] wire_d64_71;
	wire [WIDTH-1:0] wire_d64_72;
	wire [WIDTH-1:0] wire_d64_73;
	wire [WIDTH-1:0] wire_d64_74;
	wire [WIDTH-1:0] wire_d64_75;
	wire [WIDTH-1:0] wire_d64_76;
	wire [WIDTH-1:0] wire_d64_77;
	wire [WIDTH-1:0] wire_d64_78;
	wire [WIDTH-1:0] wire_d64_79;
	wire [WIDTH-1:0] wire_d64_80;
	wire [WIDTH-1:0] wire_d64_81;
	wire [WIDTH-1:0] wire_d64_82;
	wire [WIDTH-1:0] wire_d64_83;
	wire [WIDTH-1:0] wire_d64_84;
	wire [WIDTH-1:0] wire_d64_85;
	wire [WIDTH-1:0] wire_d64_86;
	wire [WIDTH-1:0] wire_d64_87;
	wire [WIDTH-1:0] wire_d64_88;
	wire [WIDTH-1:0] wire_d64_89;
	wire [WIDTH-1:0] wire_d64_90;
	wire [WIDTH-1:0] wire_d64_91;
	wire [WIDTH-1:0] wire_d64_92;
	wire [WIDTH-1:0] wire_d64_93;
	wire [WIDTH-1:0] wire_d64_94;
	wire [WIDTH-1:0] wire_d64_95;
	wire [WIDTH-1:0] wire_d64_96;
	wire [WIDTH-1:0] wire_d64_97;
	wire [WIDTH-1:0] wire_d64_98;
	wire [WIDTH-1:0] wire_d65_0;
	wire [WIDTH-1:0] wire_d65_1;
	wire [WIDTH-1:0] wire_d65_2;
	wire [WIDTH-1:0] wire_d65_3;
	wire [WIDTH-1:0] wire_d65_4;
	wire [WIDTH-1:0] wire_d65_5;
	wire [WIDTH-1:0] wire_d65_6;
	wire [WIDTH-1:0] wire_d65_7;
	wire [WIDTH-1:0] wire_d65_8;
	wire [WIDTH-1:0] wire_d65_9;
	wire [WIDTH-1:0] wire_d65_10;
	wire [WIDTH-1:0] wire_d65_11;
	wire [WIDTH-1:0] wire_d65_12;
	wire [WIDTH-1:0] wire_d65_13;
	wire [WIDTH-1:0] wire_d65_14;
	wire [WIDTH-1:0] wire_d65_15;
	wire [WIDTH-1:0] wire_d65_16;
	wire [WIDTH-1:0] wire_d65_17;
	wire [WIDTH-1:0] wire_d65_18;
	wire [WIDTH-1:0] wire_d65_19;
	wire [WIDTH-1:0] wire_d65_20;
	wire [WIDTH-1:0] wire_d65_21;
	wire [WIDTH-1:0] wire_d65_22;
	wire [WIDTH-1:0] wire_d65_23;
	wire [WIDTH-1:0] wire_d65_24;
	wire [WIDTH-1:0] wire_d65_25;
	wire [WIDTH-1:0] wire_d65_26;
	wire [WIDTH-1:0] wire_d65_27;
	wire [WIDTH-1:0] wire_d65_28;
	wire [WIDTH-1:0] wire_d65_29;
	wire [WIDTH-1:0] wire_d65_30;
	wire [WIDTH-1:0] wire_d65_31;
	wire [WIDTH-1:0] wire_d65_32;
	wire [WIDTH-1:0] wire_d65_33;
	wire [WIDTH-1:0] wire_d65_34;
	wire [WIDTH-1:0] wire_d65_35;
	wire [WIDTH-1:0] wire_d65_36;
	wire [WIDTH-1:0] wire_d65_37;
	wire [WIDTH-1:0] wire_d65_38;
	wire [WIDTH-1:0] wire_d65_39;
	wire [WIDTH-1:0] wire_d65_40;
	wire [WIDTH-1:0] wire_d65_41;
	wire [WIDTH-1:0] wire_d65_42;
	wire [WIDTH-1:0] wire_d65_43;
	wire [WIDTH-1:0] wire_d65_44;
	wire [WIDTH-1:0] wire_d65_45;
	wire [WIDTH-1:0] wire_d65_46;
	wire [WIDTH-1:0] wire_d65_47;
	wire [WIDTH-1:0] wire_d65_48;
	wire [WIDTH-1:0] wire_d65_49;
	wire [WIDTH-1:0] wire_d65_50;
	wire [WIDTH-1:0] wire_d65_51;
	wire [WIDTH-1:0] wire_d65_52;
	wire [WIDTH-1:0] wire_d65_53;
	wire [WIDTH-1:0] wire_d65_54;
	wire [WIDTH-1:0] wire_d65_55;
	wire [WIDTH-1:0] wire_d65_56;
	wire [WIDTH-1:0] wire_d65_57;
	wire [WIDTH-1:0] wire_d65_58;
	wire [WIDTH-1:0] wire_d65_59;
	wire [WIDTH-1:0] wire_d65_60;
	wire [WIDTH-1:0] wire_d65_61;
	wire [WIDTH-1:0] wire_d65_62;
	wire [WIDTH-1:0] wire_d65_63;
	wire [WIDTH-1:0] wire_d65_64;
	wire [WIDTH-1:0] wire_d65_65;
	wire [WIDTH-1:0] wire_d65_66;
	wire [WIDTH-1:0] wire_d65_67;
	wire [WIDTH-1:0] wire_d65_68;
	wire [WIDTH-1:0] wire_d65_69;
	wire [WIDTH-1:0] wire_d65_70;
	wire [WIDTH-1:0] wire_d65_71;
	wire [WIDTH-1:0] wire_d65_72;
	wire [WIDTH-1:0] wire_d65_73;
	wire [WIDTH-1:0] wire_d65_74;
	wire [WIDTH-1:0] wire_d65_75;
	wire [WIDTH-1:0] wire_d65_76;
	wire [WIDTH-1:0] wire_d65_77;
	wire [WIDTH-1:0] wire_d65_78;
	wire [WIDTH-1:0] wire_d65_79;
	wire [WIDTH-1:0] wire_d65_80;
	wire [WIDTH-1:0] wire_d65_81;
	wire [WIDTH-1:0] wire_d65_82;
	wire [WIDTH-1:0] wire_d65_83;
	wire [WIDTH-1:0] wire_d65_84;
	wire [WIDTH-1:0] wire_d65_85;
	wire [WIDTH-1:0] wire_d65_86;
	wire [WIDTH-1:0] wire_d65_87;
	wire [WIDTH-1:0] wire_d65_88;
	wire [WIDTH-1:0] wire_d65_89;
	wire [WIDTH-1:0] wire_d65_90;
	wire [WIDTH-1:0] wire_d65_91;
	wire [WIDTH-1:0] wire_d65_92;
	wire [WIDTH-1:0] wire_d65_93;
	wire [WIDTH-1:0] wire_d65_94;
	wire [WIDTH-1:0] wire_d65_95;
	wire [WIDTH-1:0] wire_d65_96;
	wire [WIDTH-1:0] wire_d65_97;
	wire [WIDTH-1:0] wire_d65_98;
	wire [WIDTH-1:0] wire_d66_0;
	wire [WIDTH-1:0] wire_d66_1;
	wire [WIDTH-1:0] wire_d66_2;
	wire [WIDTH-1:0] wire_d66_3;
	wire [WIDTH-1:0] wire_d66_4;
	wire [WIDTH-1:0] wire_d66_5;
	wire [WIDTH-1:0] wire_d66_6;
	wire [WIDTH-1:0] wire_d66_7;
	wire [WIDTH-1:0] wire_d66_8;
	wire [WIDTH-1:0] wire_d66_9;
	wire [WIDTH-1:0] wire_d66_10;
	wire [WIDTH-1:0] wire_d66_11;
	wire [WIDTH-1:0] wire_d66_12;
	wire [WIDTH-1:0] wire_d66_13;
	wire [WIDTH-1:0] wire_d66_14;
	wire [WIDTH-1:0] wire_d66_15;
	wire [WIDTH-1:0] wire_d66_16;
	wire [WIDTH-1:0] wire_d66_17;
	wire [WIDTH-1:0] wire_d66_18;
	wire [WIDTH-1:0] wire_d66_19;
	wire [WIDTH-1:0] wire_d66_20;
	wire [WIDTH-1:0] wire_d66_21;
	wire [WIDTH-1:0] wire_d66_22;
	wire [WIDTH-1:0] wire_d66_23;
	wire [WIDTH-1:0] wire_d66_24;
	wire [WIDTH-1:0] wire_d66_25;
	wire [WIDTH-1:0] wire_d66_26;
	wire [WIDTH-1:0] wire_d66_27;
	wire [WIDTH-1:0] wire_d66_28;
	wire [WIDTH-1:0] wire_d66_29;
	wire [WIDTH-1:0] wire_d66_30;
	wire [WIDTH-1:0] wire_d66_31;
	wire [WIDTH-1:0] wire_d66_32;
	wire [WIDTH-1:0] wire_d66_33;
	wire [WIDTH-1:0] wire_d66_34;
	wire [WIDTH-1:0] wire_d66_35;
	wire [WIDTH-1:0] wire_d66_36;
	wire [WIDTH-1:0] wire_d66_37;
	wire [WIDTH-1:0] wire_d66_38;
	wire [WIDTH-1:0] wire_d66_39;
	wire [WIDTH-1:0] wire_d66_40;
	wire [WIDTH-1:0] wire_d66_41;
	wire [WIDTH-1:0] wire_d66_42;
	wire [WIDTH-1:0] wire_d66_43;
	wire [WIDTH-1:0] wire_d66_44;
	wire [WIDTH-1:0] wire_d66_45;
	wire [WIDTH-1:0] wire_d66_46;
	wire [WIDTH-1:0] wire_d66_47;
	wire [WIDTH-1:0] wire_d66_48;
	wire [WIDTH-1:0] wire_d66_49;
	wire [WIDTH-1:0] wire_d66_50;
	wire [WIDTH-1:0] wire_d66_51;
	wire [WIDTH-1:0] wire_d66_52;
	wire [WIDTH-1:0] wire_d66_53;
	wire [WIDTH-1:0] wire_d66_54;
	wire [WIDTH-1:0] wire_d66_55;
	wire [WIDTH-1:0] wire_d66_56;
	wire [WIDTH-1:0] wire_d66_57;
	wire [WIDTH-1:0] wire_d66_58;
	wire [WIDTH-1:0] wire_d66_59;
	wire [WIDTH-1:0] wire_d66_60;
	wire [WIDTH-1:0] wire_d66_61;
	wire [WIDTH-1:0] wire_d66_62;
	wire [WIDTH-1:0] wire_d66_63;
	wire [WIDTH-1:0] wire_d66_64;
	wire [WIDTH-1:0] wire_d66_65;
	wire [WIDTH-1:0] wire_d66_66;
	wire [WIDTH-1:0] wire_d66_67;
	wire [WIDTH-1:0] wire_d66_68;
	wire [WIDTH-1:0] wire_d66_69;
	wire [WIDTH-1:0] wire_d66_70;
	wire [WIDTH-1:0] wire_d66_71;
	wire [WIDTH-1:0] wire_d66_72;
	wire [WIDTH-1:0] wire_d66_73;
	wire [WIDTH-1:0] wire_d66_74;
	wire [WIDTH-1:0] wire_d66_75;
	wire [WIDTH-1:0] wire_d66_76;
	wire [WIDTH-1:0] wire_d66_77;
	wire [WIDTH-1:0] wire_d66_78;
	wire [WIDTH-1:0] wire_d66_79;
	wire [WIDTH-1:0] wire_d66_80;
	wire [WIDTH-1:0] wire_d66_81;
	wire [WIDTH-1:0] wire_d66_82;
	wire [WIDTH-1:0] wire_d66_83;
	wire [WIDTH-1:0] wire_d66_84;
	wire [WIDTH-1:0] wire_d66_85;
	wire [WIDTH-1:0] wire_d66_86;
	wire [WIDTH-1:0] wire_d66_87;
	wire [WIDTH-1:0] wire_d66_88;
	wire [WIDTH-1:0] wire_d66_89;
	wire [WIDTH-1:0] wire_d66_90;
	wire [WIDTH-1:0] wire_d66_91;
	wire [WIDTH-1:0] wire_d66_92;
	wire [WIDTH-1:0] wire_d66_93;
	wire [WIDTH-1:0] wire_d66_94;
	wire [WIDTH-1:0] wire_d66_95;
	wire [WIDTH-1:0] wire_d66_96;
	wire [WIDTH-1:0] wire_d66_97;
	wire [WIDTH-1:0] wire_d66_98;
	wire [WIDTH-1:0] wire_d67_0;
	wire [WIDTH-1:0] wire_d67_1;
	wire [WIDTH-1:0] wire_d67_2;
	wire [WIDTH-1:0] wire_d67_3;
	wire [WIDTH-1:0] wire_d67_4;
	wire [WIDTH-1:0] wire_d67_5;
	wire [WIDTH-1:0] wire_d67_6;
	wire [WIDTH-1:0] wire_d67_7;
	wire [WIDTH-1:0] wire_d67_8;
	wire [WIDTH-1:0] wire_d67_9;
	wire [WIDTH-1:0] wire_d67_10;
	wire [WIDTH-1:0] wire_d67_11;
	wire [WIDTH-1:0] wire_d67_12;
	wire [WIDTH-1:0] wire_d67_13;
	wire [WIDTH-1:0] wire_d67_14;
	wire [WIDTH-1:0] wire_d67_15;
	wire [WIDTH-1:0] wire_d67_16;
	wire [WIDTH-1:0] wire_d67_17;
	wire [WIDTH-1:0] wire_d67_18;
	wire [WIDTH-1:0] wire_d67_19;
	wire [WIDTH-1:0] wire_d67_20;
	wire [WIDTH-1:0] wire_d67_21;
	wire [WIDTH-1:0] wire_d67_22;
	wire [WIDTH-1:0] wire_d67_23;
	wire [WIDTH-1:0] wire_d67_24;
	wire [WIDTH-1:0] wire_d67_25;
	wire [WIDTH-1:0] wire_d67_26;
	wire [WIDTH-1:0] wire_d67_27;
	wire [WIDTH-1:0] wire_d67_28;
	wire [WIDTH-1:0] wire_d67_29;
	wire [WIDTH-1:0] wire_d67_30;
	wire [WIDTH-1:0] wire_d67_31;
	wire [WIDTH-1:0] wire_d67_32;
	wire [WIDTH-1:0] wire_d67_33;
	wire [WIDTH-1:0] wire_d67_34;
	wire [WIDTH-1:0] wire_d67_35;
	wire [WIDTH-1:0] wire_d67_36;
	wire [WIDTH-1:0] wire_d67_37;
	wire [WIDTH-1:0] wire_d67_38;
	wire [WIDTH-1:0] wire_d67_39;
	wire [WIDTH-1:0] wire_d67_40;
	wire [WIDTH-1:0] wire_d67_41;
	wire [WIDTH-1:0] wire_d67_42;
	wire [WIDTH-1:0] wire_d67_43;
	wire [WIDTH-1:0] wire_d67_44;
	wire [WIDTH-1:0] wire_d67_45;
	wire [WIDTH-1:0] wire_d67_46;
	wire [WIDTH-1:0] wire_d67_47;
	wire [WIDTH-1:0] wire_d67_48;
	wire [WIDTH-1:0] wire_d67_49;
	wire [WIDTH-1:0] wire_d67_50;
	wire [WIDTH-1:0] wire_d67_51;
	wire [WIDTH-1:0] wire_d67_52;
	wire [WIDTH-1:0] wire_d67_53;
	wire [WIDTH-1:0] wire_d67_54;
	wire [WIDTH-1:0] wire_d67_55;
	wire [WIDTH-1:0] wire_d67_56;
	wire [WIDTH-1:0] wire_d67_57;
	wire [WIDTH-1:0] wire_d67_58;
	wire [WIDTH-1:0] wire_d67_59;
	wire [WIDTH-1:0] wire_d67_60;
	wire [WIDTH-1:0] wire_d67_61;
	wire [WIDTH-1:0] wire_d67_62;
	wire [WIDTH-1:0] wire_d67_63;
	wire [WIDTH-1:0] wire_d67_64;
	wire [WIDTH-1:0] wire_d67_65;
	wire [WIDTH-1:0] wire_d67_66;
	wire [WIDTH-1:0] wire_d67_67;
	wire [WIDTH-1:0] wire_d67_68;
	wire [WIDTH-1:0] wire_d67_69;
	wire [WIDTH-1:0] wire_d67_70;
	wire [WIDTH-1:0] wire_d67_71;
	wire [WIDTH-1:0] wire_d67_72;
	wire [WIDTH-1:0] wire_d67_73;
	wire [WIDTH-1:0] wire_d67_74;
	wire [WIDTH-1:0] wire_d67_75;
	wire [WIDTH-1:0] wire_d67_76;
	wire [WIDTH-1:0] wire_d67_77;
	wire [WIDTH-1:0] wire_d67_78;
	wire [WIDTH-1:0] wire_d67_79;
	wire [WIDTH-1:0] wire_d67_80;
	wire [WIDTH-1:0] wire_d67_81;
	wire [WIDTH-1:0] wire_d67_82;
	wire [WIDTH-1:0] wire_d67_83;
	wire [WIDTH-1:0] wire_d67_84;
	wire [WIDTH-1:0] wire_d67_85;
	wire [WIDTH-1:0] wire_d67_86;
	wire [WIDTH-1:0] wire_d67_87;
	wire [WIDTH-1:0] wire_d67_88;
	wire [WIDTH-1:0] wire_d67_89;
	wire [WIDTH-1:0] wire_d67_90;
	wire [WIDTH-1:0] wire_d67_91;
	wire [WIDTH-1:0] wire_d67_92;
	wire [WIDTH-1:0] wire_d67_93;
	wire [WIDTH-1:0] wire_d67_94;
	wire [WIDTH-1:0] wire_d67_95;
	wire [WIDTH-1:0] wire_d67_96;
	wire [WIDTH-1:0] wire_d67_97;
	wire [WIDTH-1:0] wire_d67_98;
	wire [WIDTH-1:0] wire_d68_0;
	wire [WIDTH-1:0] wire_d68_1;
	wire [WIDTH-1:0] wire_d68_2;
	wire [WIDTH-1:0] wire_d68_3;
	wire [WIDTH-1:0] wire_d68_4;
	wire [WIDTH-1:0] wire_d68_5;
	wire [WIDTH-1:0] wire_d68_6;
	wire [WIDTH-1:0] wire_d68_7;
	wire [WIDTH-1:0] wire_d68_8;
	wire [WIDTH-1:0] wire_d68_9;
	wire [WIDTH-1:0] wire_d68_10;
	wire [WIDTH-1:0] wire_d68_11;
	wire [WIDTH-1:0] wire_d68_12;
	wire [WIDTH-1:0] wire_d68_13;
	wire [WIDTH-1:0] wire_d68_14;
	wire [WIDTH-1:0] wire_d68_15;
	wire [WIDTH-1:0] wire_d68_16;
	wire [WIDTH-1:0] wire_d68_17;
	wire [WIDTH-1:0] wire_d68_18;
	wire [WIDTH-1:0] wire_d68_19;
	wire [WIDTH-1:0] wire_d68_20;
	wire [WIDTH-1:0] wire_d68_21;
	wire [WIDTH-1:0] wire_d68_22;
	wire [WIDTH-1:0] wire_d68_23;
	wire [WIDTH-1:0] wire_d68_24;
	wire [WIDTH-1:0] wire_d68_25;
	wire [WIDTH-1:0] wire_d68_26;
	wire [WIDTH-1:0] wire_d68_27;
	wire [WIDTH-1:0] wire_d68_28;
	wire [WIDTH-1:0] wire_d68_29;
	wire [WIDTH-1:0] wire_d68_30;
	wire [WIDTH-1:0] wire_d68_31;
	wire [WIDTH-1:0] wire_d68_32;
	wire [WIDTH-1:0] wire_d68_33;
	wire [WIDTH-1:0] wire_d68_34;
	wire [WIDTH-1:0] wire_d68_35;
	wire [WIDTH-1:0] wire_d68_36;
	wire [WIDTH-1:0] wire_d68_37;
	wire [WIDTH-1:0] wire_d68_38;
	wire [WIDTH-1:0] wire_d68_39;
	wire [WIDTH-1:0] wire_d68_40;
	wire [WIDTH-1:0] wire_d68_41;
	wire [WIDTH-1:0] wire_d68_42;
	wire [WIDTH-1:0] wire_d68_43;
	wire [WIDTH-1:0] wire_d68_44;
	wire [WIDTH-1:0] wire_d68_45;
	wire [WIDTH-1:0] wire_d68_46;
	wire [WIDTH-1:0] wire_d68_47;
	wire [WIDTH-1:0] wire_d68_48;
	wire [WIDTH-1:0] wire_d68_49;
	wire [WIDTH-1:0] wire_d68_50;
	wire [WIDTH-1:0] wire_d68_51;
	wire [WIDTH-1:0] wire_d68_52;
	wire [WIDTH-1:0] wire_d68_53;
	wire [WIDTH-1:0] wire_d68_54;
	wire [WIDTH-1:0] wire_d68_55;
	wire [WIDTH-1:0] wire_d68_56;
	wire [WIDTH-1:0] wire_d68_57;
	wire [WIDTH-1:0] wire_d68_58;
	wire [WIDTH-1:0] wire_d68_59;
	wire [WIDTH-1:0] wire_d68_60;
	wire [WIDTH-1:0] wire_d68_61;
	wire [WIDTH-1:0] wire_d68_62;
	wire [WIDTH-1:0] wire_d68_63;
	wire [WIDTH-1:0] wire_d68_64;
	wire [WIDTH-1:0] wire_d68_65;
	wire [WIDTH-1:0] wire_d68_66;
	wire [WIDTH-1:0] wire_d68_67;
	wire [WIDTH-1:0] wire_d68_68;
	wire [WIDTH-1:0] wire_d68_69;
	wire [WIDTH-1:0] wire_d68_70;
	wire [WIDTH-1:0] wire_d68_71;
	wire [WIDTH-1:0] wire_d68_72;
	wire [WIDTH-1:0] wire_d68_73;
	wire [WIDTH-1:0] wire_d68_74;
	wire [WIDTH-1:0] wire_d68_75;
	wire [WIDTH-1:0] wire_d68_76;
	wire [WIDTH-1:0] wire_d68_77;
	wire [WIDTH-1:0] wire_d68_78;
	wire [WIDTH-1:0] wire_d68_79;
	wire [WIDTH-1:0] wire_d68_80;
	wire [WIDTH-1:0] wire_d68_81;
	wire [WIDTH-1:0] wire_d68_82;
	wire [WIDTH-1:0] wire_d68_83;
	wire [WIDTH-1:0] wire_d68_84;
	wire [WIDTH-1:0] wire_d68_85;
	wire [WIDTH-1:0] wire_d68_86;
	wire [WIDTH-1:0] wire_d68_87;
	wire [WIDTH-1:0] wire_d68_88;
	wire [WIDTH-1:0] wire_d68_89;
	wire [WIDTH-1:0] wire_d68_90;
	wire [WIDTH-1:0] wire_d68_91;
	wire [WIDTH-1:0] wire_d68_92;
	wire [WIDTH-1:0] wire_d68_93;
	wire [WIDTH-1:0] wire_d68_94;
	wire [WIDTH-1:0] wire_d68_95;
	wire [WIDTH-1:0] wire_d68_96;
	wire [WIDTH-1:0] wire_d68_97;
	wire [WIDTH-1:0] wire_d68_98;
	wire [WIDTH-1:0] wire_d69_0;
	wire [WIDTH-1:0] wire_d69_1;
	wire [WIDTH-1:0] wire_d69_2;
	wire [WIDTH-1:0] wire_d69_3;
	wire [WIDTH-1:0] wire_d69_4;
	wire [WIDTH-1:0] wire_d69_5;
	wire [WIDTH-1:0] wire_d69_6;
	wire [WIDTH-1:0] wire_d69_7;
	wire [WIDTH-1:0] wire_d69_8;
	wire [WIDTH-1:0] wire_d69_9;
	wire [WIDTH-1:0] wire_d69_10;
	wire [WIDTH-1:0] wire_d69_11;
	wire [WIDTH-1:0] wire_d69_12;
	wire [WIDTH-1:0] wire_d69_13;
	wire [WIDTH-1:0] wire_d69_14;
	wire [WIDTH-1:0] wire_d69_15;
	wire [WIDTH-1:0] wire_d69_16;
	wire [WIDTH-1:0] wire_d69_17;
	wire [WIDTH-1:0] wire_d69_18;
	wire [WIDTH-1:0] wire_d69_19;
	wire [WIDTH-1:0] wire_d69_20;
	wire [WIDTH-1:0] wire_d69_21;
	wire [WIDTH-1:0] wire_d69_22;
	wire [WIDTH-1:0] wire_d69_23;
	wire [WIDTH-1:0] wire_d69_24;
	wire [WIDTH-1:0] wire_d69_25;
	wire [WIDTH-1:0] wire_d69_26;
	wire [WIDTH-1:0] wire_d69_27;
	wire [WIDTH-1:0] wire_d69_28;
	wire [WIDTH-1:0] wire_d69_29;
	wire [WIDTH-1:0] wire_d69_30;
	wire [WIDTH-1:0] wire_d69_31;
	wire [WIDTH-1:0] wire_d69_32;
	wire [WIDTH-1:0] wire_d69_33;
	wire [WIDTH-1:0] wire_d69_34;
	wire [WIDTH-1:0] wire_d69_35;
	wire [WIDTH-1:0] wire_d69_36;
	wire [WIDTH-1:0] wire_d69_37;
	wire [WIDTH-1:0] wire_d69_38;
	wire [WIDTH-1:0] wire_d69_39;
	wire [WIDTH-1:0] wire_d69_40;
	wire [WIDTH-1:0] wire_d69_41;
	wire [WIDTH-1:0] wire_d69_42;
	wire [WIDTH-1:0] wire_d69_43;
	wire [WIDTH-1:0] wire_d69_44;
	wire [WIDTH-1:0] wire_d69_45;
	wire [WIDTH-1:0] wire_d69_46;
	wire [WIDTH-1:0] wire_d69_47;
	wire [WIDTH-1:0] wire_d69_48;
	wire [WIDTH-1:0] wire_d69_49;
	wire [WIDTH-1:0] wire_d69_50;
	wire [WIDTH-1:0] wire_d69_51;
	wire [WIDTH-1:0] wire_d69_52;
	wire [WIDTH-1:0] wire_d69_53;
	wire [WIDTH-1:0] wire_d69_54;
	wire [WIDTH-1:0] wire_d69_55;
	wire [WIDTH-1:0] wire_d69_56;
	wire [WIDTH-1:0] wire_d69_57;
	wire [WIDTH-1:0] wire_d69_58;
	wire [WIDTH-1:0] wire_d69_59;
	wire [WIDTH-1:0] wire_d69_60;
	wire [WIDTH-1:0] wire_d69_61;
	wire [WIDTH-1:0] wire_d69_62;
	wire [WIDTH-1:0] wire_d69_63;
	wire [WIDTH-1:0] wire_d69_64;
	wire [WIDTH-1:0] wire_d69_65;
	wire [WIDTH-1:0] wire_d69_66;
	wire [WIDTH-1:0] wire_d69_67;
	wire [WIDTH-1:0] wire_d69_68;
	wire [WIDTH-1:0] wire_d69_69;
	wire [WIDTH-1:0] wire_d69_70;
	wire [WIDTH-1:0] wire_d69_71;
	wire [WIDTH-1:0] wire_d69_72;
	wire [WIDTH-1:0] wire_d69_73;
	wire [WIDTH-1:0] wire_d69_74;
	wire [WIDTH-1:0] wire_d69_75;
	wire [WIDTH-1:0] wire_d69_76;
	wire [WIDTH-1:0] wire_d69_77;
	wire [WIDTH-1:0] wire_d69_78;
	wire [WIDTH-1:0] wire_d69_79;
	wire [WIDTH-1:0] wire_d69_80;
	wire [WIDTH-1:0] wire_d69_81;
	wire [WIDTH-1:0] wire_d69_82;
	wire [WIDTH-1:0] wire_d69_83;
	wire [WIDTH-1:0] wire_d69_84;
	wire [WIDTH-1:0] wire_d69_85;
	wire [WIDTH-1:0] wire_d69_86;
	wire [WIDTH-1:0] wire_d69_87;
	wire [WIDTH-1:0] wire_d69_88;
	wire [WIDTH-1:0] wire_d69_89;
	wire [WIDTH-1:0] wire_d69_90;
	wire [WIDTH-1:0] wire_d69_91;
	wire [WIDTH-1:0] wire_d69_92;
	wire [WIDTH-1:0] wire_d69_93;
	wire [WIDTH-1:0] wire_d69_94;
	wire [WIDTH-1:0] wire_d69_95;
	wire [WIDTH-1:0] wire_d69_96;
	wire [WIDTH-1:0] wire_d69_97;
	wire [WIDTH-1:0] wire_d69_98;
	wire [WIDTH-1:0] wire_d70_0;
	wire [WIDTH-1:0] wire_d70_1;
	wire [WIDTH-1:0] wire_d70_2;
	wire [WIDTH-1:0] wire_d70_3;
	wire [WIDTH-1:0] wire_d70_4;
	wire [WIDTH-1:0] wire_d70_5;
	wire [WIDTH-1:0] wire_d70_6;
	wire [WIDTH-1:0] wire_d70_7;
	wire [WIDTH-1:0] wire_d70_8;
	wire [WIDTH-1:0] wire_d70_9;
	wire [WIDTH-1:0] wire_d70_10;
	wire [WIDTH-1:0] wire_d70_11;
	wire [WIDTH-1:0] wire_d70_12;
	wire [WIDTH-1:0] wire_d70_13;
	wire [WIDTH-1:0] wire_d70_14;
	wire [WIDTH-1:0] wire_d70_15;
	wire [WIDTH-1:0] wire_d70_16;
	wire [WIDTH-1:0] wire_d70_17;
	wire [WIDTH-1:0] wire_d70_18;
	wire [WIDTH-1:0] wire_d70_19;
	wire [WIDTH-1:0] wire_d70_20;
	wire [WIDTH-1:0] wire_d70_21;
	wire [WIDTH-1:0] wire_d70_22;
	wire [WIDTH-1:0] wire_d70_23;
	wire [WIDTH-1:0] wire_d70_24;
	wire [WIDTH-1:0] wire_d70_25;
	wire [WIDTH-1:0] wire_d70_26;
	wire [WIDTH-1:0] wire_d70_27;
	wire [WIDTH-1:0] wire_d70_28;
	wire [WIDTH-1:0] wire_d70_29;
	wire [WIDTH-1:0] wire_d70_30;
	wire [WIDTH-1:0] wire_d70_31;
	wire [WIDTH-1:0] wire_d70_32;
	wire [WIDTH-1:0] wire_d70_33;
	wire [WIDTH-1:0] wire_d70_34;
	wire [WIDTH-1:0] wire_d70_35;
	wire [WIDTH-1:0] wire_d70_36;
	wire [WIDTH-1:0] wire_d70_37;
	wire [WIDTH-1:0] wire_d70_38;
	wire [WIDTH-1:0] wire_d70_39;
	wire [WIDTH-1:0] wire_d70_40;
	wire [WIDTH-1:0] wire_d70_41;
	wire [WIDTH-1:0] wire_d70_42;
	wire [WIDTH-1:0] wire_d70_43;
	wire [WIDTH-1:0] wire_d70_44;
	wire [WIDTH-1:0] wire_d70_45;
	wire [WIDTH-1:0] wire_d70_46;
	wire [WIDTH-1:0] wire_d70_47;
	wire [WIDTH-1:0] wire_d70_48;
	wire [WIDTH-1:0] wire_d70_49;
	wire [WIDTH-1:0] wire_d70_50;
	wire [WIDTH-1:0] wire_d70_51;
	wire [WIDTH-1:0] wire_d70_52;
	wire [WIDTH-1:0] wire_d70_53;
	wire [WIDTH-1:0] wire_d70_54;
	wire [WIDTH-1:0] wire_d70_55;
	wire [WIDTH-1:0] wire_d70_56;
	wire [WIDTH-1:0] wire_d70_57;
	wire [WIDTH-1:0] wire_d70_58;
	wire [WIDTH-1:0] wire_d70_59;
	wire [WIDTH-1:0] wire_d70_60;
	wire [WIDTH-1:0] wire_d70_61;
	wire [WIDTH-1:0] wire_d70_62;
	wire [WIDTH-1:0] wire_d70_63;
	wire [WIDTH-1:0] wire_d70_64;
	wire [WIDTH-1:0] wire_d70_65;
	wire [WIDTH-1:0] wire_d70_66;
	wire [WIDTH-1:0] wire_d70_67;
	wire [WIDTH-1:0] wire_d70_68;
	wire [WIDTH-1:0] wire_d70_69;
	wire [WIDTH-1:0] wire_d70_70;
	wire [WIDTH-1:0] wire_d70_71;
	wire [WIDTH-1:0] wire_d70_72;
	wire [WIDTH-1:0] wire_d70_73;
	wire [WIDTH-1:0] wire_d70_74;
	wire [WIDTH-1:0] wire_d70_75;
	wire [WIDTH-1:0] wire_d70_76;
	wire [WIDTH-1:0] wire_d70_77;
	wire [WIDTH-1:0] wire_d70_78;
	wire [WIDTH-1:0] wire_d70_79;
	wire [WIDTH-1:0] wire_d70_80;
	wire [WIDTH-1:0] wire_d70_81;
	wire [WIDTH-1:0] wire_d70_82;
	wire [WIDTH-1:0] wire_d70_83;
	wire [WIDTH-1:0] wire_d70_84;
	wire [WIDTH-1:0] wire_d70_85;
	wire [WIDTH-1:0] wire_d70_86;
	wire [WIDTH-1:0] wire_d70_87;
	wire [WIDTH-1:0] wire_d70_88;
	wire [WIDTH-1:0] wire_d70_89;
	wire [WIDTH-1:0] wire_d70_90;
	wire [WIDTH-1:0] wire_d70_91;
	wire [WIDTH-1:0] wire_d70_92;
	wire [WIDTH-1:0] wire_d70_93;
	wire [WIDTH-1:0] wire_d70_94;
	wire [WIDTH-1:0] wire_d70_95;
	wire [WIDTH-1:0] wire_d70_96;
	wire [WIDTH-1:0] wire_d70_97;
	wire [WIDTH-1:0] wire_d70_98;
	wire [WIDTH-1:0] wire_d71_0;
	wire [WIDTH-1:0] wire_d71_1;
	wire [WIDTH-1:0] wire_d71_2;
	wire [WIDTH-1:0] wire_d71_3;
	wire [WIDTH-1:0] wire_d71_4;
	wire [WIDTH-1:0] wire_d71_5;
	wire [WIDTH-1:0] wire_d71_6;
	wire [WIDTH-1:0] wire_d71_7;
	wire [WIDTH-1:0] wire_d71_8;
	wire [WIDTH-1:0] wire_d71_9;
	wire [WIDTH-1:0] wire_d71_10;
	wire [WIDTH-1:0] wire_d71_11;
	wire [WIDTH-1:0] wire_d71_12;
	wire [WIDTH-1:0] wire_d71_13;
	wire [WIDTH-1:0] wire_d71_14;
	wire [WIDTH-1:0] wire_d71_15;
	wire [WIDTH-1:0] wire_d71_16;
	wire [WIDTH-1:0] wire_d71_17;
	wire [WIDTH-1:0] wire_d71_18;
	wire [WIDTH-1:0] wire_d71_19;
	wire [WIDTH-1:0] wire_d71_20;
	wire [WIDTH-1:0] wire_d71_21;
	wire [WIDTH-1:0] wire_d71_22;
	wire [WIDTH-1:0] wire_d71_23;
	wire [WIDTH-1:0] wire_d71_24;
	wire [WIDTH-1:0] wire_d71_25;
	wire [WIDTH-1:0] wire_d71_26;
	wire [WIDTH-1:0] wire_d71_27;
	wire [WIDTH-1:0] wire_d71_28;
	wire [WIDTH-1:0] wire_d71_29;
	wire [WIDTH-1:0] wire_d71_30;
	wire [WIDTH-1:0] wire_d71_31;
	wire [WIDTH-1:0] wire_d71_32;
	wire [WIDTH-1:0] wire_d71_33;
	wire [WIDTH-1:0] wire_d71_34;
	wire [WIDTH-1:0] wire_d71_35;
	wire [WIDTH-1:0] wire_d71_36;
	wire [WIDTH-1:0] wire_d71_37;
	wire [WIDTH-1:0] wire_d71_38;
	wire [WIDTH-1:0] wire_d71_39;
	wire [WIDTH-1:0] wire_d71_40;
	wire [WIDTH-1:0] wire_d71_41;
	wire [WIDTH-1:0] wire_d71_42;
	wire [WIDTH-1:0] wire_d71_43;
	wire [WIDTH-1:0] wire_d71_44;
	wire [WIDTH-1:0] wire_d71_45;
	wire [WIDTH-1:0] wire_d71_46;
	wire [WIDTH-1:0] wire_d71_47;
	wire [WIDTH-1:0] wire_d71_48;
	wire [WIDTH-1:0] wire_d71_49;
	wire [WIDTH-1:0] wire_d71_50;
	wire [WIDTH-1:0] wire_d71_51;
	wire [WIDTH-1:0] wire_d71_52;
	wire [WIDTH-1:0] wire_d71_53;
	wire [WIDTH-1:0] wire_d71_54;
	wire [WIDTH-1:0] wire_d71_55;
	wire [WIDTH-1:0] wire_d71_56;
	wire [WIDTH-1:0] wire_d71_57;
	wire [WIDTH-1:0] wire_d71_58;
	wire [WIDTH-1:0] wire_d71_59;
	wire [WIDTH-1:0] wire_d71_60;
	wire [WIDTH-1:0] wire_d71_61;
	wire [WIDTH-1:0] wire_d71_62;
	wire [WIDTH-1:0] wire_d71_63;
	wire [WIDTH-1:0] wire_d71_64;
	wire [WIDTH-1:0] wire_d71_65;
	wire [WIDTH-1:0] wire_d71_66;
	wire [WIDTH-1:0] wire_d71_67;
	wire [WIDTH-1:0] wire_d71_68;
	wire [WIDTH-1:0] wire_d71_69;
	wire [WIDTH-1:0] wire_d71_70;
	wire [WIDTH-1:0] wire_d71_71;
	wire [WIDTH-1:0] wire_d71_72;
	wire [WIDTH-1:0] wire_d71_73;
	wire [WIDTH-1:0] wire_d71_74;
	wire [WIDTH-1:0] wire_d71_75;
	wire [WIDTH-1:0] wire_d71_76;
	wire [WIDTH-1:0] wire_d71_77;
	wire [WIDTH-1:0] wire_d71_78;
	wire [WIDTH-1:0] wire_d71_79;
	wire [WIDTH-1:0] wire_d71_80;
	wire [WIDTH-1:0] wire_d71_81;
	wire [WIDTH-1:0] wire_d71_82;
	wire [WIDTH-1:0] wire_d71_83;
	wire [WIDTH-1:0] wire_d71_84;
	wire [WIDTH-1:0] wire_d71_85;
	wire [WIDTH-1:0] wire_d71_86;
	wire [WIDTH-1:0] wire_d71_87;
	wire [WIDTH-1:0] wire_d71_88;
	wire [WIDTH-1:0] wire_d71_89;
	wire [WIDTH-1:0] wire_d71_90;
	wire [WIDTH-1:0] wire_d71_91;
	wire [WIDTH-1:0] wire_d71_92;
	wire [WIDTH-1:0] wire_d71_93;
	wire [WIDTH-1:0] wire_d71_94;
	wire [WIDTH-1:0] wire_d71_95;
	wire [WIDTH-1:0] wire_d71_96;
	wire [WIDTH-1:0] wire_d71_97;
	wire [WIDTH-1:0] wire_d71_98;
	wire [WIDTH-1:0] wire_d72_0;
	wire [WIDTH-1:0] wire_d72_1;
	wire [WIDTH-1:0] wire_d72_2;
	wire [WIDTH-1:0] wire_d72_3;
	wire [WIDTH-1:0] wire_d72_4;
	wire [WIDTH-1:0] wire_d72_5;
	wire [WIDTH-1:0] wire_d72_6;
	wire [WIDTH-1:0] wire_d72_7;
	wire [WIDTH-1:0] wire_d72_8;
	wire [WIDTH-1:0] wire_d72_9;
	wire [WIDTH-1:0] wire_d72_10;
	wire [WIDTH-1:0] wire_d72_11;
	wire [WIDTH-1:0] wire_d72_12;
	wire [WIDTH-1:0] wire_d72_13;
	wire [WIDTH-1:0] wire_d72_14;
	wire [WIDTH-1:0] wire_d72_15;
	wire [WIDTH-1:0] wire_d72_16;
	wire [WIDTH-1:0] wire_d72_17;
	wire [WIDTH-1:0] wire_d72_18;
	wire [WIDTH-1:0] wire_d72_19;
	wire [WIDTH-1:0] wire_d72_20;
	wire [WIDTH-1:0] wire_d72_21;
	wire [WIDTH-1:0] wire_d72_22;
	wire [WIDTH-1:0] wire_d72_23;
	wire [WIDTH-1:0] wire_d72_24;
	wire [WIDTH-1:0] wire_d72_25;
	wire [WIDTH-1:0] wire_d72_26;
	wire [WIDTH-1:0] wire_d72_27;
	wire [WIDTH-1:0] wire_d72_28;
	wire [WIDTH-1:0] wire_d72_29;
	wire [WIDTH-1:0] wire_d72_30;
	wire [WIDTH-1:0] wire_d72_31;
	wire [WIDTH-1:0] wire_d72_32;
	wire [WIDTH-1:0] wire_d72_33;
	wire [WIDTH-1:0] wire_d72_34;
	wire [WIDTH-1:0] wire_d72_35;
	wire [WIDTH-1:0] wire_d72_36;
	wire [WIDTH-1:0] wire_d72_37;
	wire [WIDTH-1:0] wire_d72_38;
	wire [WIDTH-1:0] wire_d72_39;
	wire [WIDTH-1:0] wire_d72_40;
	wire [WIDTH-1:0] wire_d72_41;
	wire [WIDTH-1:0] wire_d72_42;
	wire [WIDTH-1:0] wire_d72_43;
	wire [WIDTH-1:0] wire_d72_44;
	wire [WIDTH-1:0] wire_d72_45;
	wire [WIDTH-1:0] wire_d72_46;
	wire [WIDTH-1:0] wire_d72_47;
	wire [WIDTH-1:0] wire_d72_48;
	wire [WIDTH-1:0] wire_d72_49;
	wire [WIDTH-1:0] wire_d72_50;
	wire [WIDTH-1:0] wire_d72_51;
	wire [WIDTH-1:0] wire_d72_52;
	wire [WIDTH-1:0] wire_d72_53;
	wire [WIDTH-1:0] wire_d72_54;
	wire [WIDTH-1:0] wire_d72_55;
	wire [WIDTH-1:0] wire_d72_56;
	wire [WIDTH-1:0] wire_d72_57;
	wire [WIDTH-1:0] wire_d72_58;
	wire [WIDTH-1:0] wire_d72_59;
	wire [WIDTH-1:0] wire_d72_60;
	wire [WIDTH-1:0] wire_d72_61;
	wire [WIDTH-1:0] wire_d72_62;
	wire [WIDTH-1:0] wire_d72_63;
	wire [WIDTH-1:0] wire_d72_64;
	wire [WIDTH-1:0] wire_d72_65;
	wire [WIDTH-1:0] wire_d72_66;
	wire [WIDTH-1:0] wire_d72_67;
	wire [WIDTH-1:0] wire_d72_68;
	wire [WIDTH-1:0] wire_d72_69;
	wire [WIDTH-1:0] wire_d72_70;
	wire [WIDTH-1:0] wire_d72_71;
	wire [WIDTH-1:0] wire_d72_72;
	wire [WIDTH-1:0] wire_d72_73;
	wire [WIDTH-1:0] wire_d72_74;
	wire [WIDTH-1:0] wire_d72_75;
	wire [WIDTH-1:0] wire_d72_76;
	wire [WIDTH-1:0] wire_d72_77;
	wire [WIDTH-1:0] wire_d72_78;
	wire [WIDTH-1:0] wire_d72_79;
	wire [WIDTH-1:0] wire_d72_80;
	wire [WIDTH-1:0] wire_d72_81;
	wire [WIDTH-1:0] wire_d72_82;
	wire [WIDTH-1:0] wire_d72_83;
	wire [WIDTH-1:0] wire_d72_84;
	wire [WIDTH-1:0] wire_d72_85;
	wire [WIDTH-1:0] wire_d72_86;
	wire [WIDTH-1:0] wire_d72_87;
	wire [WIDTH-1:0] wire_d72_88;
	wire [WIDTH-1:0] wire_d72_89;
	wire [WIDTH-1:0] wire_d72_90;
	wire [WIDTH-1:0] wire_d72_91;
	wire [WIDTH-1:0] wire_d72_92;
	wire [WIDTH-1:0] wire_d72_93;
	wire [WIDTH-1:0] wire_d72_94;
	wire [WIDTH-1:0] wire_d72_95;
	wire [WIDTH-1:0] wire_d72_96;
	wire [WIDTH-1:0] wire_d72_97;
	wire [WIDTH-1:0] wire_d72_98;
	wire [WIDTH-1:0] wire_d73_0;
	wire [WIDTH-1:0] wire_d73_1;
	wire [WIDTH-1:0] wire_d73_2;
	wire [WIDTH-1:0] wire_d73_3;
	wire [WIDTH-1:0] wire_d73_4;
	wire [WIDTH-1:0] wire_d73_5;
	wire [WIDTH-1:0] wire_d73_6;
	wire [WIDTH-1:0] wire_d73_7;
	wire [WIDTH-1:0] wire_d73_8;
	wire [WIDTH-1:0] wire_d73_9;
	wire [WIDTH-1:0] wire_d73_10;
	wire [WIDTH-1:0] wire_d73_11;
	wire [WIDTH-1:0] wire_d73_12;
	wire [WIDTH-1:0] wire_d73_13;
	wire [WIDTH-1:0] wire_d73_14;
	wire [WIDTH-1:0] wire_d73_15;
	wire [WIDTH-1:0] wire_d73_16;
	wire [WIDTH-1:0] wire_d73_17;
	wire [WIDTH-1:0] wire_d73_18;
	wire [WIDTH-1:0] wire_d73_19;
	wire [WIDTH-1:0] wire_d73_20;
	wire [WIDTH-1:0] wire_d73_21;
	wire [WIDTH-1:0] wire_d73_22;
	wire [WIDTH-1:0] wire_d73_23;
	wire [WIDTH-1:0] wire_d73_24;
	wire [WIDTH-1:0] wire_d73_25;
	wire [WIDTH-1:0] wire_d73_26;
	wire [WIDTH-1:0] wire_d73_27;
	wire [WIDTH-1:0] wire_d73_28;
	wire [WIDTH-1:0] wire_d73_29;
	wire [WIDTH-1:0] wire_d73_30;
	wire [WIDTH-1:0] wire_d73_31;
	wire [WIDTH-1:0] wire_d73_32;
	wire [WIDTH-1:0] wire_d73_33;
	wire [WIDTH-1:0] wire_d73_34;
	wire [WIDTH-1:0] wire_d73_35;
	wire [WIDTH-1:0] wire_d73_36;
	wire [WIDTH-1:0] wire_d73_37;
	wire [WIDTH-1:0] wire_d73_38;
	wire [WIDTH-1:0] wire_d73_39;
	wire [WIDTH-1:0] wire_d73_40;
	wire [WIDTH-1:0] wire_d73_41;
	wire [WIDTH-1:0] wire_d73_42;
	wire [WIDTH-1:0] wire_d73_43;
	wire [WIDTH-1:0] wire_d73_44;
	wire [WIDTH-1:0] wire_d73_45;
	wire [WIDTH-1:0] wire_d73_46;
	wire [WIDTH-1:0] wire_d73_47;
	wire [WIDTH-1:0] wire_d73_48;
	wire [WIDTH-1:0] wire_d73_49;
	wire [WIDTH-1:0] wire_d73_50;
	wire [WIDTH-1:0] wire_d73_51;
	wire [WIDTH-1:0] wire_d73_52;
	wire [WIDTH-1:0] wire_d73_53;
	wire [WIDTH-1:0] wire_d73_54;
	wire [WIDTH-1:0] wire_d73_55;
	wire [WIDTH-1:0] wire_d73_56;
	wire [WIDTH-1:0] wire_d73_57;
	wire [WIDTH-1:0] wire_d73_58;
	wire [WIDTH-1:0] wire_d73_59;
	wire [WIDTH-1:0] wire_d73_60;
	wire [WIDTH-1:0] wire_d73_61;
	wire [WIDTH-1:0] wire_d73_62;
	wire [WIDTH-1:0] wire_d73_63;
	wire [WIDTH-1:0] wire_d73_64;
	wire [WIDTH-1:0] wire_d73_65;
	wire [WIDTH-1:0] wire_d73_66;
	wire [WIDTH-1:0] wire_d73_67;
	wire [WIDTH-1:0] wire_d73_68;
	wire [WIDTH-1:0] wire_d73_69;
	wire [WIDTH-1:0] wire_d73_70;
	wire [WIDTH-1:0] wire_d73_71;
	wire [WIDTH-1:0] wire_d73_72;
	wire [WIDTH-1:0] wire_d73_73;
	wire [WIDTH-1:0] wire_d73_74;
	wire [WIDTH-1:0] wire_d73_75;
	wire [WIDTH-1:0] wire_d73_76;
	wire [WIDTH-1:0] wire_d73_77;
	wire [WIDTH-1:0] wire_d73_78;
	wire [WIDTH-1:0] wire_d73_79;
	wire [WIDTH-1:0] wire_d73_80;
	wire [WIDTH-1:0] wire_d73_81;
	wire [WIDTH-1:0] wire_d73_82;
	wire [WIDTH-1:0] wire_d73_83;
	wire [WIDTH-1:0] wire_d73_84;
	wire [WIDTH-1:0] wire_d73_85;
	wire [WIDTH-1:0] wire_d73_86;
	wire [WIDTH-1:0] wire_d73_87;
	wire [WIDTH-1:0] wire_d73_88;
	wire [WIDTH-1:0] wire_d73_89;
	wire [WIDTH-1:0] wire_d73_90;
	wire [WIDTH-1:0] wire_d73_91;
	wire [WIDTH-1:0] wire_d73_92;
	wire [WIDTH-1:0] wire_d73_93;
	wire [WIDTH-1:0] wire_d73_94;
	wire [WIDTH-1:0] wire_d73_95;
	wire [WIDTH-1:0] wire_d73_96;
	wire [WIDTH-1:0] wire_d73_97;
	wire [WIDTH-1:0] wire_d73_98;
	wire [WIDTH-1:0] wire_d74_0;
	wire [WIDTH-1:0] wire_d74_1;
	wire [WIDTH-1:0] wire_d74_2;
	wire [WIDTH-1:0] wire_d74_3;
	wire [WIDTH-1:0] wire_d74_4;
	wire [WIDTH-1:0] wire_d74_5;
	wire [WIDTH-1:0] wire_d74_6;
	wire [WIDTH-1:0] wire_d74_7;
	wire [WIDTH-1:0] wire_d74_8;
	wire [WIDTH-1:0] wire_d74_9;
	wire [WIDTH-1:0] wire_d74_10;
	wire [WIDTH-1:0] wire_d74_11;
	wire [WIDTH-1:0] wire_d74_12;
	wire [WIDTH-1:0] wire_d74_13;
	wire [WIDTH-1:0] wire_d74_14;
	wire [WIDTH-1:0] wire_d74_15;
	wire [WIDTH-1:0] wire_d74_16;
	wire [WIDTH-1:0] wire_d74_17;
	wire [WIDTH-1:0] wire_d74_18;
	wire [WIDTH-1:0] wire_d74_19;
	wire [WIDTH-1:0] wire_d74_20;
	wire [WIDTH-1:0] wire_d74_21;
	wire [WIDTH-1:0] wire_d74_22;
	wire [WIDTH-1:0] wire_d74_23;
	wire [WIDTH-1:0] wire_d74_24;
	wire [WIDTH-1:0] wire_d74_25;
	wire [WIDTH-1:0] wire_d74_26;
	wire [WIDTH-1:0] wire_d74_27;
	wire [WIDTH-1:0] wire_d74_28;
	wire [WIDTH-1:0] wire_d74_29;
	wire [WIDTH-1:0] wire_d74_30;
	wire [WIDTH-1:0] wire_d74_31;
	wire [WIDTH-1:0] wire_d74_32;
	wire [WIDTH-1:0] wire_d74_33;
	wire [WIDTH-1:0] wire_d74_34;
	wire [WIDTH-1:0] wire_d74_35;
	wire [WIDTH-1:0] wire_d74_36;
	wire [WIDTH-1:0] wire_d74_37;
	wire [WIDTH-1:0] wire_d74_38;
	wire [WIDTH-1:0] wire_d74_39;
	wire [WIDTH-1:0] wire_d74_40;
	wire [WIDTH-1:0] wire_d74_41;
	wire [WIDTH-1:0] wire_d74_42;
	wire [WIDTH-1:0] wire_d74_43;
	wire [WIDTH-1:0] wire_d74_44;
	wire [WIDTH-1:0] wire_d74_45;
	wire [WIDTH-1:0] wire_d74_46;
	wire [WIDTH-1:0] wire_d74_47;
	wire [WIDTH-1:0] wire_d74_48;
	wire [WIDTH-1:0] wire_d74_49;
	wire [WIDTH-1:0] wire_d74_50;
	wire [WIDTH-1:0] wire_d74_51;
	wire [WIDTH-1:0] wire_d74_52;
	wire [WIDTH-1:0] wire_d74_53;
	wire [WIDTH-1:0] wire_d74_54;
	wire [WIDTH-1:0] wire_d74_55;
	wire [WIDTH-1:0] wire_d74_56;
	wire [WIDTH-1:0] wire_d74_57;
	wire [WIDTH-1:0] wire_d74_58;
	wire [WIDTH-1:0] wire_d74_59;
	wire [WIDTH-1:0] wire_d74_60;
	wire [WIDTH-1:0] wire_d74_61;
	wire [WIDTH-1:0] wire_d74_62;
	wire [WIDTH-1:0] wire_d74_63;
	wire [WIDTH-1:0] wire_d74_64;
	wire [WIDTH-1:0] wire_d74_65;
	wire [WIDTH-1:0] wire_d74_66;
	wire [WIDTH-1:0] wire_d74_67;
	wire [WIDTH-1:0] wire_d74_68;
	wire [WIDTH-1:0] wire_d74_69;
	wire [WIDTH-1:0] wire_d74_70;
	wire [WIDTH-1:0] wire_d74_71;
	wire [WIDTH-1:0] wire_d74_72;
	wire [WIDTH-1:0] wire_d74_73;
	wire [WIDTH-1:0] wire_d74_74;
	wire [WIDTH-1:0] wire_d74_75;
	wire [WIDTH-1:0] wire_d74_76;
	wire [WIDTH-1:0] wire_d74_77;
	wire [WIDTH-1:0] wire_d74_78;
	wire [WIDTH-1:0] wire_d74_79;
	wire [WIDTH-1:0] wire_d74_80;
	wire [WIDTH-1:0] wire_d74_81;
	wire [WIDTH-1:0] wire_d74_82;
	wire [WIDTH-1:0] wire_d74_83;
	wire [WIDTH-1:0] wire_d74_84;
	wire [WIDTH-1:0] wire_d74_85;
	wire [WIDTH-1:0] wire_d74_86;
	wire [WIDTH-1:0] wire_d74_87;
	wire [WIDTH-1:0] wire_d74_88;
	wire [WIDTH-1:0] wire_d74_89;
	wire [WIDTH-1:0] wire_d74_90;
	wire [WIDTH-1:0] wire_d74_91;
	wire [WIDTH-1:0] wire_d74_92;
	wire [WIDTH-1:0] wire_d74_93;
	wire [WIDTH-1:0] wire_d74_94;
	wire [WIDTH-1:0] wire_d74_95;
	wire [WIDTH-1:0] wire_d74_96;
	wire [WIDTH-1:0] wire_d74_97;
	wire [WIDTH-1:0] wire_d74_98;
	wire [WIDTH-1:0] wire_d75_0;
	wire [WIDTH-1:0] wire_d75_1;
	wire [WIDTH-1:0] wire_d75_2;
	wire [WIDTH-1:0] wire_d75_3;
	wire [WIDTH-1:0] wire_d75_4;
	wire [WIDTH-1:0] wire_d75_5;
	wire [WIDTH-1:0] wire_d75_6;
	wire [WIDTH-1:0] wire_d75_7;
	wire [WIDTH-1:0] wire_d75_8;
	wire [WIDTH-1:0] wire_d75_9;
	wire [WIDTH-1:0] wire_d75_10;
	wire [WIDTH-1:0] wire_d75_11;
	wire [WIDTH-1:0] wire_d75_12;
	wire [WIDTH-1:0] wire_d75_13;
	wire [WIDTH-1:0] wire_d75_14;
	wire [WIDTH-1:0] wire_d75_15;
	wire [WIDTH-1:0] wire_d75_16;
	wire [WIDTH-1:0] wire_d75_17;
	wire [WIDTH-1:0] wire_d75_18;
	wire [WIDTH-1:0] wire_d75_19;
	wire [WIDTH-1:0] wire_d75_20;
	wire [WIDTH-1:0] wire_d75_21;
	wire [WIDTH-1:0] wire_d75_22;
	wire [WIDTH-1:0] wire_d75_23;
	wire [WIDTH-1:0] wire_d75_24;
	wire [WIDTH-1:0] wire_d75_25;
	wire [WIDTH-1:0] wire_d75_26;
	wire [WIDTH-1:0] wire_d75_27;
	wire [WIDTH-1:0] wire_d75_28;
	wire [WIDTH-1:0] wire_d75_29;
	wire [WIDTH-1:0] wire_d75_30;
	wire [WIDTH-1:0] wire_d75_31;
	wire [WIDTH-1:0] wire_d75_32;
	wire [WIDTH-1:0] wire_d75_33;
	wire [WIDTH-1:0] wire_d75_34;
	wire [WIDTH-1:0] wire_d75_35;
	wire [WIDTH-1:0] wire_d75_36;
	wire [WIDTH-1:0] wire_d75_37;
	wire [WIDTH-1:0] wire_d75_38;
	wire [WIDTH-1:0] wire_d75_39;
	wire [WIDTH-1:0] wire_d75_40;
	wire [WIDTH-1:0] wire_d75_41;
	wire [WIDTH-1:0] wire_d75_42;
	wire [WIDTH-1:0] wire_d75_43;
	wire [WIDTH-1:0] wire_d75_44;
	wire [WIDTH-1:0] wire_d75_45;
	wire [WIDTH-1:0] wire_d75_46;
	wire [WIDTH-1:0] wire_d75_47;
	wire [WIDTH-1:0] wire_d75_48;
	wire [WIDTH-1:0] wire_d75_49;
	wire [WIDTH-1:0] wire_d75_50;
	wire [WIDTH-1:0] wire_d75_51;
	wire [WIDTH-1:0] wire_d75_52;
	wire [WIDTH-1:0] wire_d75_53;
	wire [WIDTH-1:0] wire_d75_54;
	wire [WIDTH-1:0] wire_d75_55;
	wire [WIDTH-1:0] wire_d75_56;
	wire [WIDTH-1:0] wire_d75_57;
	wire [WIDTH-1:0] wire_d75_58;
	wire [WIDTH-1:0] wire_d75_59;
	wire [WIDTH-1:0] wire_d75_60;
	wire [WIDTH-1:0] wire_d75_61;
	wire [WIDTH-1:0] wire_d75_62;
	wire [WIDTH-1:0] wire_d75_63;
	wire [WIDTH-1:0] wire_d75_64;
	wire [WIDTH-1:0] wire_d75_65;
	wire [WIDTH-1:0] wire_d75_66;
	wire [WIDTH-1:0] wire_d75_67;
	wire [WIDTH-1:0] wire_d75_68;
	wire [WIDTH-1:0] wire_d75_69;
	wire [WIDTH-1:0] wire_d75_70;
	wire [WIDTH-1:0] wire_d75_71;
	wire [WIDTH-1:0] wire_d75_72;
	wire [WIDTH-1:0] wire_d75_73;
	wire [WIDTH-1:0] wire_d75_74;
	wire [WIDTH-1:0] wire_d75_75;
	wire [WIDTH-1:0] wire_d75_76;
	wire [WIDTH-1:0] wire_d75_77;
	wire [WIDTH-1:0] wire_d75_78;
	wire [WIDTH-1:0] wire_d75_79;
	wire [WIDTH-1:0] wire_d75_80;
	wire [WIDTH-1:0] wire_d75_81;
	wire [WIDTH-1:0] wire_d75_82;
	wire [WIDTH-1:0] wire_d75_83;
	wire [WIDTH-1:0] wire_d75_84;
	wire [WIDTH-1:0] wire_d75_85;
	wire [WIDTH-1:0] wire_d75_86;
	wire [WIDTH-1:0] wire_d75_87;
	wire [WIDTH-1:0] wire_d75_88;
	wire [WIDTH-1:0] wire_d75_89;
	wire [WIDTH-1:0] wire_d75_90;
	wire [WIDTH-1:0] wire_d75_91;
	wire [WIDTH-1:0] wire_d75_92;
	wire [WIDTH-1:0] wire_d75_93;
	wire [WIDTH-1:0] wire_d75_94;
	wire [WIDTH-1:0] wire_d75_95;
	wire [WIDTH-1:0] wire_d75_96;
	wire [WIDTH-1:0] wire_d75_97;
	wire [WIDTH-1:0] wire_d75_98;
	wire [WIDTH-1:0] wire_d76_0;
	wire [WIDTH-1:0] wire_d76_1;
	wire [WIDTH-1:0] wire_d76_2;
	wire [WIDTH-1:0] wire_d76_3;
	wire [WIDTH-1:0] wire_d76_4;
	wire [WIDTH-1:0] wire_d76_5;
	wire [WIDTH-1:0] wire_d76_6;
	wire [WIDTH-1:0] wire_d76_7;
	wire [WIDTH-1:0] wire_d76_8;
	wire [WIDTH-1:0] wire_d76_9;
	wire [WIDTH-1:0] wire_d76_10;
	wire [WIDTH-1:0] wire_d76_11;
	wire [WIDTH-1:0] wire_d76_12;
	wire [WIDTH-1:0] wire_d76_13;
	wire [WIDTH-1:0] wire_d76_14;
	wire [WIDTH-1:0] wire_d76_15;
	wire [WIDTH-1:0] wire_d76_16;
	wire [WIDTH-1:0] wire_d76_17;
	wire [WIDTH-1:0] wire_d76_18;
	wire [WIDTH-1:0] wire_d76_19;
	wire [WIDTH-1:0] wire_d76_20;
	wire [WIDTH-1:0] wire_d76_21;
	wire [WIDTH-1:0] wire_d76_22;
	wire [WIDTH-1:0] wire_d76_23;
	wire [WIDTH-1:0] wire_d76_24;
	wire [WIDTH-1:0] wire_d76_25;
	wire [WIDTH-1:0] wire_d76_26;
	wire [WIDTH-1:0] wire_d76_27;
	wire [WIDTH-1:0] wire_d76_28;
	wire [WIDTH-1:0] wire_d76_29;
	wire [WIDTH-1:0] wire_d76_30;
	wire [WIDTH-1:0] wire_d76_31;
	wire [WIDTH-1:0] wire_d76_32;
	wire [WIDTH-1:0] wire_d76_33;
	wire [WIDTH-1:0] wire_d76_34;
	wire [WIDTH-1:0] wire_d76_35;
	wire [WIDTH-1:0] wire_d76_36;
	wire [WIDTH-1:0] wire_d76_37;
	wire [WIDTH-1:0] wire_d76_38;
	wire [WIDTH-1:0] wire_d76_39;
	wire [WIDTH-1:0] wire_d76_40;
	wire [WIDTH-1:0] wire_d76_41;
	wire [WIDTH-1:0] wire_d76_42;
	wire [WIDTH-1:0] wire_d76_43;
	wire [WIDTH-1:0] wire_d76_44;
	wire [WIDTH-1:0] wire_d76_45;
	wire [WIDTH-1:0] wire_d76_46;
	wire [WIDTH-1:0] wire_d76_47;
	wire [WIDTH-1:0] wire_d76_48;
	wire [WIDTH-1:0] wire_d76_49;
	wire [WIDTH-1:0] wire_d76_50;
	wire [WIDTH-1:0] wire_d76_51;
	wire [WIDTH-1:0] wire_d76_52;
	wire [WIDTH-1:0] wire_d76_53;
	wire [WIDTH-1:0] wire_d76_54;
	wire [WIDTH-1:0] wire_d76_55;
	wire [WIDTH-1:0] wire_d76_56;
	wire [WIDTH-1:0] wire_d76_57;
	wire [WIDTH-1:0] wire_d76_58;
	wire [WIDTH-1:0] wire_d76_59;
	wire [WIDTH-1:0] wire_d76_60;
	wire [WIDTH-1:0] wire_d76_61;
	wire [WIDTH-1:0] wire_d76_62;
	wire [WIDTH-1:0] wire_d76_63;
	wire [WIDTH-1:0] wire_d76_64;
	wire [WIDTH-1:0] wire_d76_65;
	wire [WIDTH-1:0] wire_d76_66;
	wire [WIDTH-1:0] wire_d76_67;
	wire [WIDTH-1:0] wire_d76_68;
	wire [WIDTH-1:0] wire_d76_69;
	wire [WIDTH-1:0] wire_d76_70;
	wire [WIDTH-1:0] wire_d76_71;
	wire [WIDTH-1:0] wire_d76_72;
	wire [WIDTH-1:0] wire_d76_73;
	wire [WIDTH-1:0] wire_d76_74;
	wire [WIDTH-1:0] wire_d76_75;
	wire [WIDTH-1:0] wire_d76_76;
	wire [WIDTH-1:0] wire_d76_77;
	wire [WIDTH-1:0] wire_d76_78;
	wire [WIDTH-1:0] wire_d76_79;
	wire [WIDTH-1:0] wire_d76_80;
	wire [WIDTH-1:0] wire_d76_81;
	wire [WIDTH-1:0] wire_d76_82;
	wire [WIDTH-1:0] wire_d76_83;
	wire [WIDTH-1:0] wire_d76_84;
	wire [WIDTH-1:0] wire_d76_85;
	wire [WIDTH-1:0] wire_d76_86;
	wire [WIDTH-1:0] wire_d76_87;
	wire [WIDTH-1:0] wire_d76_88;
	wire [WIDTH-1:0] wire_d76_89;
	wire [WIDTH-1:0] wire_d76_90;
	wire [WIDTH-1:0] wire_d76_91;
	wire [WIDTH-1:0] wire_d76_92;
	wire [WIDTH-1:0] wire_d76_93;
	wire [WIDTH-1:0] wire_d76_94;
	wire [WIDTH-1:0] wire_d76_95;
	wire [WIDTH-1:0] wire_d76_96;
	wire [WIDTH-1:0] wire_d76_97;
	wire [WIDTH-1:0] wire_d76_98;
	wire [WIDTH-1:0] wire_d77_0;
	wire [WIDTH-1:0] wire_d77_1;
	wire [WIDTH-1:0] wire_d77_2;
	wire [WIDTH-1:0] wire_d77_3;
	wire [WIDTH-1:0] wire_d77_4;
	wire [WIDTH-1:0] wire_d77_5;
	wire [WIDTH-1:0] wire_d77_6;
	wire [WIDTH-1:0] wire_d77_7;
	wire [WIDTH-1:0] wire_d77_8;
	wire [WIDTH-1:0] wire_d77_9;
	wire [WIDTH-1:0] wire_d77_10;
	wire [WIDTH-1:0] wire_d77_11;
	wire [WIDTH-1:0] wire_d77_12;
	wire [WIDTH-1:0] wire_d77_13;
	wire [WIDTH-1:0] wire_d77_14;
	wire [WIDTH-1:0] wire_d77_15;
	wire [WIDTH-1:0] wire_d77_16;
	wire [WIDTH-1:0] wire_d77_17;
	wire [WIDTH-1:0] wire_d77_18;
	wire [WIDTH-1:0] wire_d77_19;
	wire [WIDTH-1:0] wire_d77_20;
	wire [WIDTH-1:0] wire_d77_21;
	wire [WIDTH-1:0] wire_d77_22;
	wire [WIDTH-1:0] wire_d77_23;
	wire [WIDTH-1:0] wire_d77_24;
	wire [WIDTH-1:0] wire_d77_25;
	wire [WIDTH-1:0] wire_d77_26;
	wire [WIDTH-1:0] wire_d77_27;
	wire [WIDTH-1:0] wire_d77_28;
	wire [WIDTH-1:0] wire_d77_29;
	wire [WIDTH-1:0] wire_d77_30;
	wire [WIDTH-1:0] wire_d77_31;
	wire [WIDTH-1:0] wire_d77_32;
	wire [WIDTH-1:0] wire_d77_33;
	wire [WIDTH-1:0] wire_d77_34;
	wire [WIDTH-1:0] wire_d77_35;
	wire [WIDTH-1:0] wire_d77_36;
	wire [WIDTH-1:0] wire_d77_37;
	wire [WIDTH-1:0] wire_d77_38;
	wire [WIDTH-1:0] wire_d77_39;
	wire [WIDTH-1:0] wire_d77_40;
	wire [WIDTH-1:0] wire_d77_41;
	wire [WIDTH-1:0] wire_d77_42;
	wire [WIDTH-1:0] wire_d77_43;
	wire [WIDTH-1:0] wire_d77_44;
	wire [WIDTH-1:0] wire_d77_45;
	wire [WIDTH-1:0] wire_d77_46;
	wire [WIDTH-1:0] wire_d77_47;
	wire [WIDTH-1:0] wire_d77_48;
	wire [WIDTH-1:0] wire_d77_49;
	wire [WIDTH-1:0] wire_d77_50;
	wire [WIDTH-1:0] wire_d77_51;
	wire [WIDTH-1:0] wire_d77_52;
	wire [WIDTH-1:0] wire_d77_53;
	wire [WIDTH-1:0] wire_d77_54;
	wire [WIDTH-1:0] wire_d77_55;
	wire [WIDTH-1:0] wire_d77_56;
	wire [WIDTH-1:0] wire_d77_57;
	wire [WIDTH-1:0] wire_d77_58;
	wire [WIDTH-1:0] wire_d77_59;
	wire [WIDTH-1:0] wire_d77_60;
	wire [WIDTH-1:0] wire_d77_61;
	wire [WIDTH-1:0] wire_d77_62;
	wire [WIDTH-1:0] wire_d77_63;
	wire [WIDTH-1:0] wire_d77_64;
	wire [WIDTH-1:0] wire_d77_65;
	wire [WIDTH-1:0] wire_d77_66;
	wire [WIDTH-1:0] wire_d77_67;
	wire [WIDTH-1:0] wire_d77_68;
	wire [WIDTH-1:0] wire_d77_69;
	wire [WIDTH-1:0] wire_d77_70;
	wire [WIDTH-1:0] wire_d77_71;
	wire [WIDTH-1:0] wire_d77_72;
	wire [WIDTH-1:0] wire_d77_73;
	wire [WIDTH-1:0] wire_d77_74;
	wire [WIDTH-1:0] wire_d77_75;
	wire [WIDTH-1:0] wire_d77_76;
	wire [WIDTH-1:0] wire_d77_77;
	wire [WIDTH-1:0] wire_d77_78;
	wire [WIDTH-1:0] wire_d77_79;
	wire [WIDTH-1:0] wire_d77_80;
	wire [WIDTH-1:0] wire_d77_81;
	wire [WIDTH-1:0] wire_d77_82;
	wire [WIDTH-1:0] wire_d77_83;
	wire [WIDTH-1:0] wire_d77_84;
	wire [WIDTH-1:0] wire_d77_85;
	wire [WIDTH-1:0] wire_d77_86;
	wire [WIDTH-1:0] wire_d77_87;
	wire [WIDTH-1:0] wire_d77_88;
	wire [WIDTH-1:0] wire_d77_89;
	wire [WIDTH-1:0] wire_d77_90;
	wire [WIDTH-1:0] wire_d77_91;
	wire [WIDTH-1:0] wire_d77_92;
	wire [WIDTH-1:0] wire_d77_93;
	wire [WIDTH-1:0] wire_d77_94;
	wire [WIDTH-1:0] wire_d77_95;
	wire [WIDTH-1:0] wire_d77_96;
	wire [WIDTH-1:0] wire_d77_97;
	wire [WIDTH-1:0] wire_d77_98;
	wire [WIDTH-1:0] wire_d78_0;
	wire [WIDTH-1:0] wire_d78_1;
	wire [WIDTH-1:0] wire_d78_2;
	wire [WIDTH-1:0] wire_d78_3;
	wire [WIDTH-1:0] wire_d78_4;
	wire [WIDTH-1:0] wire_d78_5;
	wire [WIDTH-1:0] wire_d78_6;
	wire [WIDTH-1:0] wire_d78_7;
	wire [WIDTH-1:0] wire_d78_8;
	wire [WIDTH-1:0] wire_d78_9;
	wire [WIDTH-1:0] wire_d78_10;
	wire [WIDTH-1:0] wire_d78_11;
	wire [WIDTH-1:0] wire_d78_12;
	wire [WIDTH-1:0] wire_d78_13;
	wire [WIDTH-1:0] wire_d78_14;
	wire [WIDTH-1:0] wire_d78_15;
	wire [WIDTH-1:0] wire_d78_16;
	wire [WIDTH-1:0] wire_d78_17;
	wire [WIDTH-1:0] wire_d78_18;
	wire [WIDTH-1:0] wire_d78_19;
	wire [WIDTH-1:0] wire_d78_20;
	wire [WIDTH-1:0] wire_d78_21;
	wire [WIDTH-1:0] wire_d78_22;
	wire [WIDTH-1:0] wire_d78_23;
	wire [WIDTH-1:0] wire_d78_24;
	wire [WIDTH-1:0] wire_d78_25;
	wire [WIDTH-1:0] wire_d78_26;
	wire [WIDTH-1:0] wire_d78_27;
	wire [WIDTH-1:0] wire_d78_28;
	wire [WIDTH-1:0] wire_d78_29;
	wire [WIDTH-1:0] wire_d78_30;
	wire [WIDTH-1:0] wire_d78_31;
	wire [WIDTH-1:0] wire_d78_32;
	wire [WIDTH-1:0] wire_d78_33;
	wire [WIDTH-1:0] wire_d78_34;
	wire [WIDTH-1:0] wire_d78_35;
	wire [WIDTH-1:0] wire_d78_36;
	wire [WIDTH-1:0] wire_d78_37;
	wire [WIDTH-1:0] wire_d78_38;
	wire [WIDTH-1:0] wire_d78_39;
	wire [WIDTH-1:0] wire_d78_40;
	wire [WIDTH-1:0] wire_d78_41;
	wire [WIDTH-1:0] wire_d78_42;
	wire [WIDTH-1:0] wire_d78_43;
	wire [WIDTH-1:0] wire_d78_44;
	wire [WIDTH-1:0] wire_d78_45;
	wire [WIDTH-1:0] wire_d78_46;
	wire [WIDTH-1:0] wire_d78_47;
	wire [WIDTH-1:0] wire_d78_48;
	wire [WIDTH-1:0] wire_d78_49;
	wire [WIDTH-1:0] wire_d78_50;
	wire [WIDTH-1:0] wire_d78_51;
	wire [WIDTH-1:0] wire_d78_52;
	wire [WIDTH-1:0] wire_d78_53;
	wire [WIDTH-1:0] wire_d78_54;
	wire [WIDTH-1:0] wire_d78_55;
	wire [WIDTH-1:0] wire_d78_56;
	wire [WIDTH-1:0] wire_d78_57;
	wire [WIDTH-1:0] wire_d78_58;
	wire [WIDTH-1:0] wire_d78_59;
	wire [WIDTH-1:0] wire_d78_60;
	wire [WIDTH-1:0] wire_d78_61;
	wire [WIDTH-1:0] wire_d78_62;
	wire [WIDTH-1:0] wire_d78_63;
	wire [WIDTH-1:0] wire_d78_64;
	wire [WIDTH-1:0] wire_d78_65;
	wire [WIDTH-1:0] wire_d78_66;
	wire [WIDTH-1:0] wire_d78_67;
	wire [WIDTH-1:0] wire_d78_68;
	wire [WIDTH-1:0] wire_d78_69;
	wire [WIDTH-1:0] wire_d78_70;
	wire [WIDTH-1:0] wire_d78_71;
	wire [WIDTH-1:0] wire_d78_72;
	wire [WIDTH-1:0] wire_d78_73;
	wire [WIDTH-1:0] wire_d78_74;
	wire [WIDTH-1:0] wire_d78_75;
	wire [WIDTH-1:0] wire_d78_76;
	wire [WIDTH-1:0] wire_d78_77;
	wire [WIDTH-1:0] wire_d78_78;
	wire [WIDTH-1:0] wire_d78_79;
	wire [WIDTH-1:0] wire_d78_80;
	wire [WIDTH-1:0] wire_d78_81;
	wire [WIDTH-1:0] wire_d78_82;
	wire [WIDTH-1:0] wire_d78_83;
	wire [WIDTH-1:0] wire_d78_84;
	wire [WIDTH-1:0] wire_d78_85;
	wire [WIDTH-1:0] wire_d78_86;
	wire [WIDTH-1:0] wire_d78_87;
	wire [WIDTH-1:0] wire_d78_88;
	wire [WIDTH-1:0] wire_d78_89;
	wire [WIDTH-1:0] wire_d78_90;
	wire [WIDTH-1:0] wire_d78_91;
	wire [WIDTH-1:0] wire_d78_92;
	wire [WIDTH-1:0] wire_d78_93;
	wire [WIDTH-1:0] wire_d78_94;
	wire [WIDTH-1:0] wire_d78_95;
	wire [WIDTH-1:0] wire_d78_96;
	wire [WIDTH-1:0] wire_d78_97;
	wire [WIDTH-1:0] wire_d78_98;
	wire [WIDTH-1:0] wire_d79_0;
	wire [WIDTH-1:0] wire_d79_1;
	wire [WIDTH-1:0] wire_d79_2;
	wire [WIDTH-1:0] wire_d79_3;
	wire [WIDTH-1:0] wire_d79_4;
	wire [WIDTH-1:0] wire_d79_5;
	wire [WIDTH-1:0] wire_d79_6;
	wire [WIDTH-1:0] wire_d79_7;
	wire [WIDTH-1:0] wire_d79_8;
	wire [WIDTH-1:0] wire_d79_9;
	wire [WIDTH-1:0] wire_d79_10;
	wire [WIDTH-1:0] wire_d79_11;
	wire [WIDTH-1:0] wire_d79_12;
	wire [WIDTH-1:0] wire_d79_13;
	wire [WIDTH-1:0] wire_d79_14;
	wire [WIDTH-1:0] wire_d79_15;
	wire [WIDTH-1:0] wire_d79_16;
	wire [WIDTH-1:0] wire_d79_17;
	wire [WIDTH-1:0] wire_d79_18;
	wire [WIDTH-1:0] wire_d79_19;
	wire [WIDTH-1:0] wire_d79_20;
	wire [WIDTH-1:0] wire_d79_21;
	wire [WIDTH-1:0] wire_d79_22;
	wire [WIDTH-1:0] wire_d79_23;
	wire [WIDTH-1:0] wire_d79_24;
	wire [WIDTH-1:0] wire_d79_25;
	wire [WIDTH-1:0] wire_d79_26;
	wire [WIDTH-1:0] wire_d79_27;
	wire [WIDTH-1:0] wire_d79_28;
	wire [WIDTH-1:0] wire_d79_29;
	wire [WIDTH-1:0] wire_d79_30;
	wire [WIDTH-1:0] wire_d79_31;
	wire [WIDTH-1:0] wire_d79_32;
	wire [WIDTH-1:0] wire_d79_33;
	wire [WIDTH-1:0] wire_d79_34;
	wire [WIDTH-1:0] wire_d79_35;
	wire [WIDTH-1:0] wire_d79_36;
	wire [WIDTH-1:0] wire_d79_37;
	wire [WIDTH-1:0] wire_d79_38;
	wire [WIDTH-1:0] wire_d79_39;
	wire [WIDTH-1:0] wire_d79_40;
	wire [WIDTH-1:0] wire_d79_41;
	wire [WIDTH-1:0] wire_d79_42;
	wire [WIDTH-1:0] wire_d79_43;
	wire [WIDTH-1:0] wire_d79_44;
	wire [WIDTH-1:0] wire_d79_45;
	wire [WIDTH-1:0] wire_d79_46;
	wire [WIDTH-1:0] wire_d79_47;
	wire [WIDTH-1:0] wire_d79_48;
	wire [WIDTH-1:0] wire_d79_49;
	wire [WIDTH-1:0] wire_d79_50;
	wire [WIDTH-1:0] wire_d79_51;
	wire [WIDTH-1:0] wire_d79_52;
	wire [WIDTH-1:0] wire_d79_53;
	wire [WIDTH-1:0] wire_d79_54;
	wire [WIDTH-1:0] wire_d79_55;
	wire [WIDTH-1:0] wire_d79_56;
	wire [WIDTH-1:0] wire_d79_57;
	wire [WIDTH-1:0] wire_d79_58;
	wire [WIDTH-1:0] wire_d79_59;
	wire [WIDTH-1:0] wire_d79_60;
	wire [WIDTH-1:0] wire_d79_61;
	wire [WIDTH-1:0] wire_d79_62;
	wire [WIDTH-1:0] wire_d79_63;
	wire [WIDTH-1:0] wire_d79_64;
	wire [WIDTH-1:0] wire_d79_65;
	wire [WIDTH-1:0] wire_d79_66;
	wire [WIDTH-1:0] wire_d79_67;
	wire [WIDTH-1:0] wire_d79_68;
	wire [WIDTH-1:0] wire_d79_69;
	wire [WIDTH-1:0] wire_d79_70;
	wire [WIDTH-1:0] wire_d79_71;
	wire [WIDTH-1:0] wire_d79_72;
	wire [WIDTH-1:0] wire_d79_73;
	wire [WIDTH-1:0] wire_d79_74;
	wire [WIDTH-1:0] wire_d79_75;
	wire [WIDTH-1:0] wire_d79_76;
	wire [WIDTH-1:0] wire_d79_77;
	wire [WIDTH-1:0] wire_d79_78;
	wire [WIDTH-1:0] wire_d79_79;
	wire [WIDTH-1:0] wire_d79_80;
	wire [WIDTH-1:0] wire_d79_81;
	wire [WIDTH-1:0] wire_d79_82;
	wire [WIDTH-1:0] wire_d79_83;
	wire [WIDTH-1:0] wire_d79_84;
	wire [WIDTH-1:0] wire_d79_85;
	wire [WIDTH-1:0] wire_d79_86;
	wire [WIDTH-1:0] wire_d79_87;
	wire [WIDTH-1:0] wire_d79_88;
	wire [WIDTH-1:0] wire_d79_89;
	wire [WIDTH-1:0] wire_d79_90;
	wire [WIDTH-1:0] wire_d79_91;
	wire [WIDTH-1:0] wire_d79_92;
	wire [WIDTH-1:0] wire_d79_93;
	wire [WIDTH-1:0] wire_d79_94;
	wire [WIDTH-1:0] wire_d79_95;
	wire [WIDTH-1:0] wire_d79_96;
	wire [WIDTH-1:0] wire_d79_97;
	wire [WIDTH-1:0] wire_d79_98;
	wire [WIDTH-1:0] wire_d80_0;
	wire [WIDTH-1:0] wire_d80_1;
	wire [WIDTH-1:0] wire_d80_2;
	wire [WIDTH-1:0] wire_d80_3;
	wire [WIDTH-1:0] wire_d80_4;
	wire [WIDTH-1:0] wire_d80_5;
	wire [WIDTH-1:0] wire_d80_6;
	wire [WIDTH-1:0] wire_d80_7;
	wire [WIDTH-1:0] wire_d80_8;
	wire [WIDTH-1:0] wire_d80_9;
	wire [WIDTH-1:0] wire_d80_10;
	wire [WIDTH-1:0] wire_d80_11;
	wire [WIDTH-1:0] wire_d80_12;
	wire [WIDTH-1:0] wire_d80_13;
	wire [WIDTH-1:0] wire_d80_14;
	wire [WIDTH-1:0] wire_d80_15;
	wire [WIDTH-1:0] wire_d80_16;
	wire [WIDTH-1:0] wire_d80_17;
	wire [WIDTH-1:0] wire_d80_18;
	wire [WIDTH-1:0] wire_d80_19;
	wire [WIDTH-1:0] wire_d80_20;
	wire [WIDTH-1:0] wire_d80_21;
	wire [WIDTH-1:0] wire_d80_22;
	wire [WIDTH-1:0] wire_d80_23;
	wire [WIDTH-1:0] wire_d80_24;
	wire [WIDTH-1:0] wire_d80_25;
	wire [WIDTH-1:0] wire_d80_26;
	wire [WIDTH-1:0] wire_d80_27;
	wire [WIDTH-1:0] wire_d80_28;
	wire [WIDTH-1:0] wire_d80_29;
	wire [WIDTH-1:0] wire_d80_30;
	wire [WIDTH-1:0] wire_d80_31;
	wire [WIDTH-1:0] wire_d80_32;
	wire [WIDTH-1:0] wire_d80_33;
	wire [WIDTH-1:0] wire_d80_34;
	wire [WIDTH-1:0] wire_d80_35;
	wire [WIDTH-1:0] wire_d80_36;
	wire [WIDTH-1:0] wire_d80_37;
	wire [WIDTH-1:0] wire_d80_38;
	wire [WIDTH-1:0] wire_d80_39;
	wire [WIDTH-1:0] wire_d80_40;
	wire [WIDTH-1:0] wire_d80_41;
	wire [WIDTH-1:0] wire_d80_42;
	wire [WIDTH-1:0] wire_d80_43;
	wire [WIDTH-1:0] wire_d80_44;
	wire [WIDTH-1:0] wire_d80_45;
	wire [WIDTH-1:0] wire_d80_46;
	wire [WIDTH-1:0] wire_d80_47;
	wire [WIDTH-1:0] wire_d80_48;
	wire [WIDTH-1:0] wire_d80_49;
	wire [WIDTH-1:0] wire_d80_50;
	wire [WIDTH-1:0] wire_d80_51;
	wire [WIDTH-1:0] wire_d80_52;
	wire [WIDTH-1:0] wire_d80_53;
	wire [WIDTH-1:0] wire_d80_54;
	wire [WIDTH-1:0] wire_d80_55;
	wire [WIDTH-1:0] wire_d80_56;
	wire [WIDTH-1:0] wire_d80_57;
	wire [WIDTH-1:0] wire_d80_58;
	wire [WIDTH-1:0] wire_d80_59;
	wire [WIDTH-1:0] wire_d80_60;
	wire [WIDTH-1:0] wire_d80_61;
	wire [WIDTH-1:0] wire_d80_62;
	wire [WIDTH-1:0] wire_d80_63;
	wire [WIDTH-1:0] wire_d80_64;
	wire [WIDTH-1:0] wire_d80_65;
	wire [WIDTH-1:0] wire_d80_66;
	wire [WIDTH-1:0] wire_d80_67;
	wire [WIDTH-1:0] wire_d80_68;
	wire [WIDTH-1:0] wire_d80_69;
	wire [WIDTH-1:0] wire_d80_70;
	wire [WIDTH-1:0] wire_d80_71;
	wire [WIDTH-1:0] wire_d80_72;
	wire [WIDTH-1:0] wire_d80_73;
	wire [WIDTH-1:0] wire_d80_74;
	wire [WIDTH-1:0] wire_d80_75;
	wire [WIDTH-1:0] wire_d80_76;
	wire [WIDTH-1:0] wire_d80_77;
	wire [WIDTH-1:0] wire_d80_78;
	wire [WIDTH-1:0] wire_d80_79;
	wire [WIDTH-1:0] wire_d80_80;
	wire [WIDTH-1:0] wire_d80_81;
	wire [WIDTH-1:0] wire_d80_82;
	wire [WIDTH-1:0] wire_d80_83;
	wire [WIDTH-1:0] wire_d80_84;
	wire [WIDTH-1:0] wire_d80_85;
	wire [WIDTH-1:0] wire_d80_86;
	wire [WIDTH-1:0] wire_d80_87;
	wire [WIDTH-1:0] wire_d80_88;
	wire [WIDTH-1:0] wire_d80_89;
	wire [WIDTH-1:0] wire_d80_90;
	wire [WIDTH-1:0] wire_d80_91;
	wire [WIDTH-1:0] wire_d80_92;
	wire [WIDTH-1:0] wire_d80_93;
	wire [WIDTH-1:0] wire_d80_94;
	wire [WIDTH-1:0] wire_d80_95;
	wire [WIDTH-1:0] wire_d80_96;
	wire [WIDTH-1:0] wire_d80_97;
	wire [WIDTH-1:0] wire_d80_98;
	wire [WIDTH-1:0] wire_d81_0;
	wire [WIDTH-1:0] wire_d81_1;
	wire [WIDTH-1:0] wire_d81_2;
	wire [WIDTH-1:0] wire_d81_3;
	wire [WIDTH-1:0] wire_d81_4;
	wire [WIDTH-1:0] wire_d81_5;
	wire [WIDTH-1:0] wire_d81_6;
	wire [WIDTH-1:0] wire_d81_7;
	wire [WIDTH-1:0] wire_d81_8;
	wire [WIDTH-1:0] wire_d81_9;
	wire [WIDTH-1:0] wire_d81_10;
	wire [WIDTH-1:0] wire_d81_11;
	wire [WIDTH-1:0] wire_d81_12;
	wire [WIDTH-1:0] wire_d81_13;
	wire [WIDTH-1:0] wire_d81_14;
	wire [WIDTH-1:0] wire_d81_15;
	wire [WIDTH-1:0] wire_d81_16;
	wire [WIDTH-1:0] wire_d81_17;
	wire [WIDTH-1:0] wire_d81_18;
	wire [WIDTH-1:0] wire_d81_19;
	wire [WIDTH-1:0] wire_d81_20;
	wire [WIDTH-1:0] wire_d81_21;
	wire [WIDTH-1:0] wire_d81_22;
	wire [WIDTH-1:0] wire_d81_23;
	wire [WIDTH-1:0] wire_d81_24;
	wire [WIDTH-1:0] wire_d81_25;
	wire [WIDTH-1:0] wire_d81_26;
	wire [WIDTH-1:0] wire_d81_27;
	wire [WIDTH-1:0] wire_d81_28;
	wire [WIDTH-1:0] wire_d81_29;
	wire [WIDTH-1:0] wire_d81_30;
	wire [WIDTH-1:0] wire_d81_31;
	wire [WIDTH-1:0] wire_d81_32;
	wire [WIDTH-1:0] wire_d81_33;
	wire [WIDTH-1:0] wire_d81_34;
	wire [WIDTH-1:0] wire_d81_35;
	wire [WIDTH-1:0] wire_d81_36;
	wire [WIDTH-1:0] wire_d81_37;
	wire [WIDTH-1:0] wire_d81_38;
	wire [WIDTH-1:0] wire_d81_39;
	wire [WIDTH-1:0] wire_d81_40;
	wire [WIDTH-1:0] wire_d81_41;
	wire [WIDTH-1:0] wire_d81_42;
	wire [WIDTH-1:0] wire_d81_43;
	wire [WIDTH-1:0] wire_d81_44;
	wire [WIDTH-1:0] wire_d81_45;
	wire [WIDTH-1:0] wire_d81_46;
	wire [WIDTH-1:0] wire_d81_47;
	wire [WIDTH-1:0] wire_d81_48;
	wire [WIDTH-1:0] wire_d81_49;
	wire [WIDTH-1:0] wire_d81_50;
	wire [WIDTH-1:0] wire_d81_51;
	wire [WIDTH-1:0] wire_d81_52;
	wire [WIDTH-1:0] wire_d81_53;
	wire [WIDTH-1:0] wire_d81_54;
	wire [WIDTH-1:0] wire_d81_55;
	wire [WIDTH-1:0] wire_d81_56;
	wire [WIDTH-1:0] wire_d81_57;
	wire [WIDTH-1:0] wire_d81_58;
	wire [WIDTH-1:0] wire_d81_59;
	wire [WIDTH-1:0] wire_d81_60;
	wire [WIDTH-1:0] wire_d81_61;
	wire [WIDTH-1:0] wire_d81_62;
	wire [WIDTH-1:0] wire_d81_63;
	wire [WIDTH-1:0] wire_d81_64;
	wire [WIDTH-1:0] wire_d81_65;
	wire [WIDTH-1:0] wire_d81_66;
	wire [WIDTH-1:0] wire_d81_67;
	wire [WIDTH-1:0] wire_d81_68;
	wire [WIDTH-1:0] wire_d81_69;
	wire [WIDTH-1:0] wire_d81_70;
	wire [WIDTH-1:0] wire_d81_71;
	wire [WIDTH-1:0] wire_d81_72;
	wire [WIDTH-1:0] wire_d81_73;
	wire [WIDTH-1:0] wire_d81_74;
	wire [WIDTH-1:0] wire_d81_75;
	wire [WIDTH-1:0] wire_d81_76;
	wire [WIDTH-1:0] wire_d81_77;
	wire [WIDTH-1:0] wire_d81_78;
	wire [WIDTH-1:0] wire_d81_79;
	wire [WIDTH-1:0] wire_d81_80;
	wire [WIDTH-1:0] wire_d81_81;
	wire [WIDTH-1:0] wire_d81_82;
	wire [WIDTH-1:0] wire_d81_83;
	wire [WIDTH-1:0] wire_d81_84;
	wire [WIDTH-1:0] wire_d81_85;
	wire [WIDTH-1:0] wire_d81_86;
	wire [WIDTH-1:0] wire_d81_87;
	wire [WIDTH-1:0] wire_d81_88;
	wire [WIDTH-1:0] wire_d81_89;
	wire [WIDTH-1:0] wire_d81_90;
	wire [WIDTH-1:0] wire_d81_91;
	wire [WIDTH-1:0] wire_d81_92;
	wire [WIDTH-1:0] wire_d81_93;
	wire [WIDTH-1:0] wire_d81_94;
	wire [WIDTH-1:0] wire_d81_95;
	wire [WIDTH-1:0] wire_d81_96;
	wire [WIDTH-1:0] wire_d81_97;
	wire [WIDTH-1:0] wire_d81_98;
	wire [WIDTH-1:0] wire_d82_0;
	wire [WIDTH-1:0] wire_d82_1;
	wire [WIDTH-1:0] wire_d82_2;
	wire [WIDTH-1:0] wire_d82_3;
	wire [WIDTH-1:0] wire_d82_4;
	wire [WIDTH-1:0] wire_d82_5;
	wire [WIDTH-1:0] wire_d82_6;
	wire [WIDTH-1:0] wire_d82_7;
	wire [WIDTH-1:0] wire_d82_8;
	wire [WIDTH-1:0] wire_d82_9;
	wire [WIDTH-1:0] wire_d82_10;
	wire [WIDTH-1:0] wire_d82_11;
	wire [WIDTH-1:0] wire_d82_12;
	wire [WIDTH-1:0] wire_d82_13;
	wire [WIDTH-1:0] wire_d82_14;
	wire [WIDTH-1:0] wire_d82_15;
	wire [WIDTH-1:0] wire_d82_16;
	wire [WIDTH-1:0] wire_d82_17;
	wire [WIDTH-1:0] wire_d82_18;
	wire [WIDTH-1:0] wire_d82_19;
	wire [WIDTH-1:0] wire_d82_20;
	wire [WIDTH-1:0] wire_d82_21;
	wire [WIDTH-1:0] wire_d82_22;
	wire [WIDTH-1:0] wire_d82_23;
	wire [WIDTH-1:0] wire_d82_24;
	wire [WIDTH-1:0] wire_d82_25;
	wire [WIDTH-1:0] wire_d82_26;
	wire [WIDTH-1:0] wire_d82_27;
	wire [WIDTH-1:0] wire_d82_28;
	wire [WIDTH-1:0] wire_d82_29;
	wire [WIDTH-1:0] wire_d82_30;
	wire [WIDTH-1:0] wire_d82_31;
	wire [WIDTH-1:0] wire_d82_32;
	wire [WIDTH-1:0] wire_d82_33;
	wire [WIDTH-1:0] wire_d82_34;
	wire [WIDTH-1:0] wire_d82_35;
	wire [WIDTH-1:0] wire_d82_36;
	wire [WIDTH-1:0] wire_d82_37;
	wire [WIDTH-1:0] wire_d82_38;
	wire [WIDTH-1:0] wire_d82_39;
	wire [WIDTH-1:0] wire_d82_40;
	wire [WIDTH-1:0] wire_d82_41;
	wire [WIDTH-1:0] wire_d82_42;
	wire [WIDTH-1:0] wire_d82_43;
	wire [WIDTH-1:0] wire_d82_44;
	wire [WIDTH-1:0] wire_d82_45;
	wire [WIDTH-1:0] wire_d82_46;
	wire [WIDTH-1:0] wire_d82_47;
	wire [WIDTH-1:0] wire_d82_48;
	wire [WIDTH-1:0] wire_d82_49;
	wire [WIDTH-1:0] wire_d82_50;
	wire [WIDTH-1:0] wire_d82_51;
	wire [WIDTH-1:0] wire_d82_52;
	wire [WIDTH-1:0] wire_d82_53;
	wire [WIDTH-1:0] wire_d82_54;
	wire [WIDTH-1:0] wire_d82_55;
	wire [WIDTH-1:0] wire_d82_56;
	wire [WIDTH-1:0] wire_d82_57;
	wire [WIDTH-1:0] wire_d82_58;
	wire [WIDTH-1:0] wire_d82_59;
	wire [WIDTH-1:0] wire_d82_60;
	wire [WIDTH-1:0] wire_d82_61;
	wire [WIDTH-1:0] wire_d82_62;
	wire [WIDTH-1:0] wire_d82_63;
	wire [WIDTH-1:0] wire_d82_64;
	wire [WIDTH-1:0] wire_d82_65;
	wire [WIDTH-1:0] wire_d82_66;
	wire [WIDTH-1:0] wire_d82_67;
	wire [WIDTH-1:0] wire_d82_68;
	wire [WIDTH-1:0] wire_d82_69;
	wire [WIDTH-1:0] wire_d82_70;
	wire [WIDTH-1:0] wire_d82_71;
	wire [WIDTH-1:0] wire_d82_72;
	wire [WIDTH-1:0] wire_d82_73;
	wire [WIDTH-1:0] wire_d82_74;
	wire [WIDTH-1:0] wire_d82_75;
	wire [WIDTH-1:0] wire_d82_76;
	wire [WIDTH-1:0] wire_d82_77;
	wire [WIDTH-1:0] wire_d82_78;
	wire [WIDTH-1:0] wire_d82_79;
	wire [WIDTH-1:0] wire_d82_80;
	wire [WIDTH-1:0] wire_d82_81;
	wire [WIDTH-1:0] wire_d82_82;
	wire [WIDTH-1:0] wire_d82_83;
	wire [WIDTH-1:0] wire_d82_84;
	wire [WIDTH-1:0] wire_d82_85;
	wire [WIDTH-1:0] wire_d82_86;
	wire [WIDTH-1:0] wire_d82_87;
	wire [WIDTH-1:0] wire_d82_88;
	wire [WIDTH-1:0] wire_d82_89;
	wire [WIDTH-1:0] wire_d82_90;
	wire [WIDTH-1:0] wire_d82_91;
	wire [WIDTH-1:0] wire_d82_92;
	wire [WIDTH-1:0] wire_d82_93;
	wire [WIDTH-1:0] wire_d82_94;
	wire [WIDTH-1:0] wire_d82_95;
	wire [WIDTH-1:0] wire_d82_96;
	wire [WIDTH-1:0] wire_d82_97;
	wire [WIDTH-1:0] wire_d82_98;
	wire [WIDTH-1:0] wire_d83_0;
	wire [WIDTH-1:0] wire_d83_1;
	wire [WIDTH-1:0] wire_d83_2;
	wire [WIDTH-1:0] wire_d83_3;
	wire [WIDTH-1:0] wire_d83_4;
	wire [WIDTH-1:0] wire_d83_5;
	wire [WIDTH-1:0] wire_d83_6;
	wire [WIDTH-1:0] wire_d83_7;
	wire [WIDTH-1:0] wire_d83_8;
	wire [WIDTH-1:0] wire_d83_9;
	wire [WIDTH-1:0] wire_d83_10;
	wire [WIDTH-1:0] wire_d83_11;
	wire [WIDTH-1:0] wire_d83_12;
	wire [WIDTH-1:0] wire_d83_13;
	wire [WIDTH-1:0] wire_d83_14;
	wire [WIDTH-1:0] wire_d83_15;
	wire [WIDTH-1:0] wire_d83_16;
	wire [WIDTH-1:0] wire_d83_17;
	wire [WIDTH-1:0] wire_d83_18;
	wire [WIDTH-1:0] wire_d83_19;
	wire [WIDTH-1:0] wire_d83_20;
	wire [WIDTH-1:0] wire_d83_21;
	wire [WIDTH-1:0] wire_d83_22;
	wire [WIDTH-1:0] wire_d83_23;
	wire [WIDTH-1:0] wire_d83_24;
	wire [WIDTH-1:0] wire_d83_25;
	wire [WIDTH-1:0] wire_d83_26;
	wire [WIDTH-1:0] wire_d83_27;
	wire [WIDTH-1:0] wire_d83_28;
	wire [WIDTH-1:0] wire_d83_29;
	wire [WIDTH-1:0] wire_d83_30;
	wire [WIDTH-1:0] wire_d83_31;
	wire [WIDTH-1:0] wire_d83_32;
	wire [WIDTH-1:0] wire_d83_33;
	wire [WIDTH-1:0] wire_d83_34;
	wire [WIDTH-1:0] wire_d83_35;
	wire [WIDTH-1:0] wire_d83_36;
	wire [WIDTH-1:0] wire_d83_37;
	wire [WIDTH-1:0] wire_d83_38;
	wire [WIDTH-1:0] wire_d83_39;
	wire [WIDTH-1:0] wire_d83_40;
	wire [WIDTH-1:0] wire_d83_41;
	wire [WIDTH-1:0] wire_d83_42;
	wire [WIDTH-1:0] wire_d83_43;
	wire [WIDTH-1:0] wire_d83_44;
	wire [WIDTH-1:0] wire_d83_45;
	wire [WIDTH-1:0] wire_d83_46;
	wire [WIDTH-1:0] wire_d83_47;
	wire [WIDTH-1:0] wire_d83_48;
	wire [WIDTH-1:0] wire_d83_49;
	wire [WIDTH-1:0] wire_d83_50;
	wire [WIDTH-1:0] wire_d83_51;
	wire [WIDTH-1:0] wire_d83_52;
	wire [WIDTH-1:0] wire_d83_53;
	wire [WIDTH-1:0] wire_d83_54;
	wire [WIDTH-1:0] wire_d83_55;
	wire [WIDTH-1:0] wire_d83_56;
	wire [WIDTH-1:0] wire_d83_57;
	wire [WIDTH-1:0] wire_d83_58;
	wire [WIDTH-1:0] wire_d83_59;
	wire [WIDTH-1:0] wire_d83_60;
	wire [WIDTH-1:0] wire_d83_61;
	wire [WIDTH-1:0] wire_d83_62;
	wire [WIDTH-1:0] wire_d83_63;
	wire [WIDTH-1:0] wire_d83_64;
	wire [WIDTH-1:0] wire_d83_65;
	wire [WIDTH-1:0] wire_d83_66;
	wire [WIDTH-1:0] wire_d83_67;
	wire [WIDTH-1:0] wire_d83_68;
	wire [WIDTH-1:0] wire_d83_69;
	wire [WIDTH-1:0] wire_d83_70;
	wire [WIDTH-1:0] wire_d83_71;
	wire [WIDTH-1:0] wire_d83_72;
	wire [WIDTH-1:0] wire_d83_73;
	wire [WIDTH-1:0] wire_d83_74;
	wire [WIDTH-1:0] wire_d83_75;
	wire [WIDTH-1:0] wire_d83_76;
	wire [WIDTH-1:0] wire_d83_77;
	wire [WIDTH-1:0] wire_d83_78;
	wire [WIDTH-1:0] wire_d83_79;
	wire [WIDTH-1:0] wire_d83_80;
	wire [WIDTH-1:0] wire_d83_81;
	wire [WIDTH-1:0] wire_d83_82;
	wire [WIDTH-1:0] wire_d83_83;
	wire [WIDTH-1:0] wire_d83_84;
	wire [WIDTH-1:0] wire_d83_85;
	wire [WIDTH-1:0] wire_d83_86;
	wire [WIDTH-1:0] wire_d83_87;
	wire [WIDTH-1:0] wire_d83_88;
	wire [WIDTH-1:0] wire_d83_89;
	wire [WIDTH-1:0] wire_d83_90;
	wire [WIDTH-1:0] wire_d83_91;
	wire [WIDTH-1:0] wire_d83_92;
	wire [WIDTH-1:0] wire_d83_93;
	wire [WIDTH-1:0] wire_d83_94;
	wire [WIDTH-1:0] wire_d83_95;
	wire [WIDTH-1:0] wire_d83_96;
	wire [WIDTH-1:0] wire_d83_97;
	wire [WIDTH-1:0] wire_d83_98;
	wire [WIDTH-1:0] wire_d84_0;
	wire [WIDTH-1:0] wire_d84_1;
	wire [WIDTH-1:0] wire_d84_2;
	wire [WIDTH-1:0] wire_d84_3;
	wire [WIDTH-1:0] wire_d84_4;
	wire [WIDTH-1:0] wire_d84_5;
	wire [WIDTH-1:0] wire_d84_6;
	wire [WIDTH-1:0] wire_d84_7;
	wire [WIDTH-1:0] wire_d84_8;
	wire [WIDTH-1:0] wire_d84_9;
	wire [WIDTH-1:0] wire_d84_10;
	wire [WIDTH-1:0] wire_d84_11;
	wire [WIDTH-1:0] wire_d84_12;
	wire [WIDTH-1:0] wire_d84_13;
	wire [WIDTH-1:0] wire_d84_14;
	wire [WIDTH-1:0] wire_d84_15;
	wire [WIDTH-1:0] wire_d84_16;
	wire [WIDTH-1:0] wire_d84_17;
	wire [WIDTH-1:0] wire_d84_18;
	wire [WIDTH-1:0] wire_d84_19;
	wire [WIDTH-1:0] wire_d84_20;
	wire [WIDTH-1:0] wire_d84_21;
	wire [WIDTH-1:0] wire_d84_22;
	wire [WIDTH-1:0] wire_d84_23;
	wire [WIDTH-1:0] wire_d84_24;
	wire [WIDTH-1:0] wire_d84_25;
	wire [WIDTH-1:0] wire_d84_26;
	wire [WIDTH-1:0] wire_d84_27;
	wire [WIDTH-1:0] wire_d84_28;
	wire [WIDTH-1:0] wire_d84_29;
	wire [WIDTH-1:0] wire_d84_30;
	wire [WIDTH-1:0] wire_d84_31;
	wire [WIDTH-1:0] wire_d84_32;
	wire [WIDTH-1:0] wire_d84_33;
	wire [WIDTH-1:0] wire_d84_34;
	wire [WIDTH-1:0] wire_d84_35;
	wire [WIDTH-1:0] wire_d84_36;
	wire [WIDTH-1:0] wire_d84_37;
	wire [WIDTH-1:0] wire_d84_38;
	wire [WIDTH-1:0] wire_d84_39;
	wire [WIDTH-1:0] wire_d84_40;
	wire [WIDTH-1:0] wire_d84_41;
	wire [WIDTH-1:0] wire_d84_42;
	wire [WIDTH-1:0] wire_d84_43;
	wire [WIDTH-1:0] wire_d84_44;
	wire [WIDTH-1:0] wire_d84_45;
	wire [WIDTH-1:0] wire_d84_46;
	wire [WIDTH-1:0] wire_d84_47;
	wire [WIDTH-1:0] wire_d84_48;
	wire [WIDTH-1:0] wire_d84_49;
	wire [WIDTH-1:0] wire_d84_50;
	wire [WIDTH-1:0] wire_d84_51;
	wire [WIDTH-1:0] wire_d84_52;
	wire [WIDTH-1:0] wire_d84_53;
	wire [WIDTH-1:0] wire_d84_54;
	wire [WIDTH-1:0] wire_d84_55;
	wire [WIDTH-1:0] wire_d84_56;
	wire [WIDTH-1:0] wire_d84_57;
	wire [WIDTH-1:0] wire_d84_58;
	wire [WIDTH-1:0] wire_d84_59;
	wire [WIDTH-1:0] wire_d84_60;
	wire [WIDTH-1:0] wire_d84_61;
	wire [WIDTH-1:0] wire_d84_62;
	wire [WIDTH-1:0] wire_d84_63;
	wire [WIDTH-1:0] wire_d84_64;
	wire [WIDTH-1:0] wire_d84_65;
	wire [WIDTH-1:0] wire_d84_66;
	wire [WIDTH-1:0] wire_d84_67;
	wire [WIDTH-1:0] wire_d84_68;
	wire [WIDTH-1:0] wire_d84_69;
	wire [WIDTH-1:0] wire_d84_70;
	wire [WIDTH-1:0] wire_d84_71;
	wire [WIDTH-1:0] wire_d84_72;
	wire [WIDTH-1:0] wire_d84_73;
	wire [WIDTH-1:0] wire_d84_74;
	wire [WIDTH-1:0] wire_d84_75;
	wire [WIDTH-1:0] wire_d84_76;
	wire [WIDTH-1:0] wire_d84_77;
	wire [WIDTH-1:0] wire_d84_78;
	wire [WIDTH-1:0] wire_d84_79;
	wire [WIDTH-1:0] wire_d84_80;
	wire [WIDTH-1:0] wire_d84_81;
	wire [WIDTH-1:0] wire_d84_82;
	wire [WIDTH-1:0] wire_d84_83;
	wire [WIDTH-1:0] wire_d84_84;
	wire [WIDTH-1:0] wire_d84_85;
	wire [WIDTH-1:0] wire_d84_86;
	wire [WIDTH-1:0] wire_d84_87;
	wire [WIDTH-1:0] wire_d84_88;
	wire [WIDTH-1:0] wire_d84_89;
	wire [WIDTH-1:0] wire_d84_90;
	wire [WIDTH-1:0] wire_d84_91;
	wire [WIDTH-1:0] wire_d84_92;
	wire [WIDTH-1:0] wire_d84_93;
	wire [WIDTH-1:0] wire_d84_94;
	wire [WIDTH-1:0] wire_d84_95;
	wire [WIDTH-1:0] wire_d84_96;
	wire [WIDTH-1:0] wire_d84_97;
	wire [WIDTH-1:0] wire_d84_98;
	wire [WIDTH-1:0] wire_d85_0;
	wire [WIDTH-1:0] wire_d85_1;
	wire [WIDTH-1:0] wire_d85_2;
	wire [WIDTH-1:0] wire_d85_3;
	wire [WIDTH-1:0] wire_d85_4;
	wire [WIDTH-1:0] wire_d85_5;
	wire [WIDTH-1:0] wire_d85_6;
	wire [WIDTH-1:0] wire_d85_7;
	wire [WIDTH-1:0] wire_d85_8;
	wire [WIDTH-1:0] wire_d85_9;
	wire [WIDTH-1:0] wire_d85_10;
	wire [WIDTH-1:0] wire_d85_11;
	wire [WIDTH-1:0] wire_d85_12;
	wire [WIDTH-1:0] wire_d85_13;
	wire [WIDTH-1:0] wire_d85_14;
	wire [WIDTH-1:0] wire_d85_15;
	wire [WIDTH-1:0] wire_d85_16;
	wire [WIDTH-1:0] wire_d85_17;
	wire [WIDTH-1:0] wire_d85_18;
	wire [WIDTH-1:0] wire_d85_19;
	wire [WIDTH-1:0] wire_d85_20;
	wire [WIDTH-1:0] wire_d85_21;
	wire [WIDTH-1:0] wire_d85_22;
	wire [WIDTH-1:0] wire_d85_23;
	wire [WIDTH-1:0] wire_d85_24;
	wire [WIDTH-1:0] wire_d85_25;
	wire [WIDTH-1:0] wire_d85_26;
	wire [WIDTH-1:0] wire_d85_27;
	wire [WIDTH-1:0] wire_d85_28;
	wire [WIDTH-1:0] wire_d85_29;
	wire [WIDTH-1:0] wire_d85_30;
	wire [WIDTH-1:0] wire_d85_31;
	wire [WIDTH-1:0] wire_d85_32;
	wire [WIDTH-1:0] wire_d85_33;
	wire [WIDTH-1:0] wire_d85_34;
	wire [WIDTH-1:0] wire_d85_35;
	wire [WIDTH-1:0] wire_d85_36;
	wire [WIDTH-1:0] wire_d85_37;
	wire [WIDTH-1:0] wire_d85_38;
	wire [WIDTH-1:0] wire_d85_39;
	wire [WIDTH-1:0] wire_d85_40;
	wire [WIDTH-1:0] wire_d85_41;
	wire [WIDTH-1:0] wire_d85_42;
	wire [WIDTH-1:0] wire_d85_43;
	wire [WIDTH-1:0] wire_d85_44;
	wire [WIDTH-1:0] wire_d85_45;
	wire [WIDTH-1:0] wire_d85_46;
	wire [WIDTH-1:0] wire_d85_47;
	wire [WIDTH-1:0] wire_d85_48;
	wire [WIDTH-1:0] wire_d85_49;
	wire [WIDTH-1:0] wire_d85_50;
	wire [WIDTH-1:0] wire_d85_51;
	wire [WIDTH-1:0] wire_d85_52;
	wire [WIDTH-1:0] wire_d85_53;
	wire [WIDTH-1:0] wire_d85_54;
	wire [WIDTH-1:0] wire_d85_55;
	wire [WIDTH-1:0] wire_d85_56;
	wire [WIDTH-1:0] wire_d85_57;
	wire [WIDTH-1:0] wire_d85_58;
	wire [WIDTH-1:0] wire_d85_59;
	wire [WIDTH-1:0] wire_d85_60;
	wire [WIDTH-1:0] wire_d85_61;
	wire [WIDTH-1:0] wire_d85_62;
	wire [WIDTH-1:0] wire_d85_63;
	wire [WIDTH-1:0] wire_d85_64;
	wire [WIDTH-1:0] wire_d85_65;
	wire [WIDTH-1:0] wire_d85_66;
	wire [WIDTH-1:0] wire_d85_67;
	wire [WIDTH-1:0] wire_d85_68;
	wire [WIDTH-1:0] wire_d85_69;
	wire [WIDTH-1:0] wire_d85_70;
	wire [WIDTH-1:0] wire_d85_71;
	wire [WIDTH-1:0] wire_d85_72;
	wire [WIDTH-1:0] wire_d85_73;
	wire [WIDTH-1:0] wire_d85_74;
	wire [WIDTH-1:0] wire_d85_75;
	wire [WIDTH-1:0] wire_d85_76;
	wire [WIDTH-1:0] wire_d85_77;
	wire [WIDTH-1:0] wire_d85_78;
	wire [WIDTH-1:0] wire_d85_79;
	wire [WIDTH-1:0] wire_d85_80;
	wire [WIDTH-1:0] wire_d85_81;
	wire [WIDTH-1:0] wire_d85_82;
	wire [WIDTH-1:0] wire_d85_83;
	wire [WIDTH-1:0] wire_d85_84;
	wire [WIDTH-1:0] wire_d85_85;
	wire [WIDTH-1:0] wire_d85_86;
	wire [WIDTH-1:0] wire_d85_87;
	wire [WIDTH-1:0] wire_d85_88;
	wire [WIDTH-1:0] wire_d85_89;
	wire [WIDTH-1:0] wire_d85_90;
	wire [WIDTH-1:0] wire_d85_91;
	wire [WIDTH-1:0] wire_d85_92;
	wire [WIDTH-1:0] wire_d85_93;
	wire [WIDTH-1:0] wire_d85_94;
	wire [WIDTH-1:0] wire_d85_95;
	wire [WIDTH-1:0] wire_d85_96;
	wire [WIDTH-1:0] wire_d85_97;
	wire [WIDTH-1:0] wire_d85_98;
	wire [WIDTH-1:0] wire_d86_0;
	wire [WIDTH-1:0] wire_d86_1;
	wire [WIDTH-1:0] wire_d86_2;
	wire [WIDTH-1:0] wire_d86_3;
	wire [WIDTH-1:0] wire_d86_4;
	wire [WIDTH-1:0] wire_d86_5;
	wire [WIDTH-1:0] wire_d86_6;
	wire [WIDTH-1:0] wire_d86_7;
	wire [WIDTH-1:0] wire_d86_8;
	wire [WIDTH-1:0] wire_d86_9;
	wire [WIDTH-1:0] wire_d86_10;
	wire [WIDTH-1:0] wire_d86_11;
	wire [WIDTH-1:0] wire_d86_12;
	wire [WIDTH-1:0] wire_d86_13;
	wire [WIDTH-1:0] wire_d86_14;
	wire [WIDTH-1:0] wire_d86_15;
	wire [WIDTH-1:0] wire_d86_16;
	wire [WIDTH-1:0] wire_d86_17;
	wire [WIDTH-1:0] wire_d86_18;
	wire [WIDTH-1:0] wire_d86_19;
	wire [WIDTH-1:0] wire_d86_20;
	wire [WIDTH-1:0] wire_d86_21;
	wire [WIDTH-1:0] wire_d86_22;
	wire [WIDTH-1:0] wire_d86_23;
	wire [WIDTH-1:0] wire_d86_24;
	wire [WIDTH-1:0] wire_d86_25;
	wire [WIDTH-1:0] wire_d86_26;
	wire [WIDTH-1:0] wire_d86_27;
	wire [WIDTH-1:0] wire_d86_28;
	wire [WIDTH-1:0] wire_d86_29;
	wire [WIDTH-1:0] wire_d86_30;
	wire [WIDTH-1:0] wire_d86_31;
	wire [WIDTH-1:0] wire_d86_32;
	wire [WIDTH-1:0] wire_d86_33;
	wire [WIDTH-1:0] wire_d86_34;
	wire [WIDTH-1:0] wire_d86_35;
	wire [WIDTH-1:0] wire_d86_36;
	wire [WIDTH-1:0] wire_d86_37;
	wire [WIDTH-1:0] wire_d86_38;
	wire [WIDTH-1:0] wire_d86_39;
	wire [WIDTH-1:0] wire_d86_40;
	wire [WIDTH-1:0] wire_d86_41;
	wire [WIDTH-1:0] wire_d86_42;
	wire [WIDTH-1:0] wire_d86_43;
	wire [WIDTH-1:0] wire_d86_44;
	wire [WIDTH-1:0] wire_d86_45;
	wire [WIDTH-1:0] wire_d86_46;
	wire [WIDTH-1:0] wire_d86_47;
	wire [WIDTH-1:0] wire_d86_48;
	wire [WIDTH-1:0] wire_d86_49;
	wire [WIDTH-1:0] wire_d86_50;
	wire [WIDTH-1:0] wire_d86_51;
	wire [WIDTH-1:0] wire_d86_52;
	wire [WIDTH-1:0] wire_d86_53;
	wire [WIDTH-1:0] wire_d86_54;
	wire [WIDTH-1:0] wire_d86_55;
	wire [WIDTH-1:0] wire_d86_56;
	wire [WIDTH-1:0] wire_d86_57;
	wire [WIDTH-1:0] wire_d86_58;
	wire [WIDTH-1:0] wire_d86_59;
	wire [WIDTH-1:0] wire_d86_60;
	wire [WIDTH-1:0] wire_d86_61;
	wire [WIDTH-1:0] wire_d86_62;
	wire [WIDTH-1:0] wire_d86_63;
	wire [WIDTH-1:0] wire_d86_64;
	wire [WIDTH-1:0] wire_d86_65;
	wire [WIDTH-1:0] wire_d86_66;
	wire [WIDTH-1:0] wire_d86_67;
	wire [WIDTH-1:0] wire_d86_68;
	wire [WIDTH-1:0] wire_d86_69;
	wire [WIDTH-1:0] wire_d86_70;
	wire [WIDTH-1:0] wire_d86_71;
	wire [WIDTH-1:0] wire_d86_72;
	wire [WIDTH-1:0] wire_d86_73;
	wire [WIDTH-1:0] wire_d86_74;
	wire [WIDTH-1:0] wire_d86_75;
	wire [WIDTH-1:0] wire_d86_76;
	wire [WIDTH-1:0] wire_d86_77;
	wire [WIDTH-1:0] wire_d86_78;
	wire [WIDTH-1:0] wire_d86_79;
	wire [WIDTH-1:0] wire_d86_80;
	wire [WIDTH-1:0] wire_d86_81;
	wire [WIDTH-1:0] wire_d86_82;
	wire [WIDTH-1:0] wire_d86_83;
	wire [WIDTH-1:0] wire_d86_84;
	wire [WIDTH-1:0] wire_d86_85;
	wire [WIDTH-1:0] wire_d86_86;
	wire [WIDTH-1:0] wire_d86_87;
	wire [WIDTH-1:0] wire_d86_88;
	wire [WIDTH-1:0] wire_d86_89;
	wire [WIDTH-1:0] wire_d86_90;
	wire [WIDTH-1:0] wire_d86_91;
	wire [WIDTH-1:0] wire_d86_92;
	wire [WIDTH-1:0] wire_d86_93;
	wire [WIDTH-1:0] wire_d86_94;
	wire [WIDTH-1:0] wire_d86_95;
	wire [WIDTH-1:0] wire_d86_96;
	wire [WIDTH-1:0] wire_d86_97;
	wire [WIDTH-1:0] wire_d86_98;
	wire [WIDTH-1:0] wire_d87_0;
	wire [WIDTH-1:0] wire_d87_1;
	wire [WIDTH-1:0] wire_d87_2;
	wire [WIDTH-1:0] wire_d87_3;
	wire [WIDTH-1:0] wire_d87_4;
	wire [WIDTH-1:0] wire_d87_5;
	wire [WIDTH-1:0] wire_d87_6;
	wire [WIDTH-1:0] wire_d87_7;
	wire [WIDTH-1:0] wire_d87_8;
	wire [WIDTH-1:0] wire_d87_9;
	wire [WIDTH-1:0] wire_d87_10;
	wire [WIDTH-1:0] wire_d87_11;
	wire [WIDTH-1:0] wire_d87_12;
	wire [WIDTH-1:0] wire_d87_13;
	wire [WIDTH-1:0] wire_d87_14;
	wire [WIDTH-1:0] wire_d87_15;
	wire [WIDTH-1:0] wire_d87_16;
	wire [WIDTH-1:0] wire_d87_17;
	wire [WIDTH-1:0] wire_d87_18;
	wire [WIDTH-1:0] wire_d87_19;
	wire [WIDTH-1:0] wire_d87_20;
	wire [WIDTH-1:0] wire_d87_21;
	wire [WIDTH-1:0] wire_d87_22;
	wire [WIDTH-1:0] wire_d87_23;
	wire [WIDTH-1:0] wire_d87_24;
	wire [WIDTH-1:0] wire_d87_25;
	wire [WIDTH-1:0] wire_d87_26;
	wire [WIDTH-1:0] wire_d87_27;
	wire [WIDTH-1:0] wire_d87_28;
	wire [WIDTH-1:0] wire_d87_29;
	wire [WIDTH-1:0] wire_d87_30;
	wire [WIDTH-1:0] wire_d87_31;
	wire [WIDTH-1:0] wire_d87_32;
	wire [WIDTH-1:0] wire_d87_33;
	wire [WIDTH-1:0] wire_d87_34;
	wire [WIDTH-1:0] wire_d87_35;
	wire [WIDTH-1:0] wire_d87_36;
	wire [WIDTH-1:0] wire_d87_37;
	wire [WIDTH-1:0] wire_d87_38;
	wire [WIDTH-1:0] wire_d87_39;
	wire [WIDTH-1:0] wire_d87_40;
	wire [WIDTH-1:0] wire_d87_41;
	wire [WIDTH-1:0] wire_d87_42;
	wire [WIDTH-1:0] wire_d87_43;
	wire [WIDTH-1:0] wire_d87_44;
	wire [WIDTH-1:0] wire_d87_45;
	wire [WIDTH-1:0] wire_d87_46;
	wire [WIDTH-1:0] wire_d87_47;
	wire [WIDTH-1:0] wire_d87_48;
	wire [WIDTH-1:0] wire_d87_49;
	wire [WIDTH-1:0] wire_d87_50;
	wire [WIDTH-1:0] wire_d87_51;
	wire [WIDTH-1:0] wire_d87_52;
	wire [WIDTH-1:0] wire_d87_53;
	wire [WIDTH-1:0] wire_d87_54;
	wire [WIDTH-1:0] wire_d87_55;
	wire [WIDTH-1:0] wire_d87_56;
	wire [WIDTH-1:0] wire_d87_57;
	wire [WIDTH-1:0] wire_d87_58;
	wire [WIDTH-1:0] wire_d87_59;
	wire [WIDTH-1:0] wire_d87_60;
	wire [WIDTH-1:0] wire_d87_61;
	wire [WIDTH-1:0] wire_d87_62;
	wire [WIDTH-1:0] wire_d87_63;
	wire [WIDTH-1:0] wire_d87_64;
	wire [WIDTH-1:0] wire_d87_65;
	wire [WIDTH-1:0] wire_d87_66;
	wire [WIDTH-1:0] wire_d87_67;
	wire [WIDTH-1:0] wire_d87_68;
	wire [WIDTH-1:0] wire_d87_69;
	wire [WIDTH-1:0] wire_d87_70;
	wire [WIDTH-1:0] wire_d87_71;
	wire [WIDTH-1:0] wire_d87_72;
	wire [WIDTH-1:0] wire_d87_73;
	wire [WIDTH-1:0] wire_d87_74;
	wire [WIDTH-1:0] wire_d87_75;
	wire [WIDTH-1:0] wire_d87_76;
	wire [WIDTH-1:0] wire_d87_77;
	wire [WIDTH-1:0] wire_d87_78;
	wire [WIDTH-1:0] wire_d87_79;
	wire [WIDTH-1:0] wire_d87_80;
	wire [WIDTH-1:0] wire_d87_81;
	wire [WIDTH-1:0] wire_d87_82;
	wire [WIDTH-1:0] wire_d87_83;
	wire [WIDTH-1:0] wire_d87_84;
	wire [WIDTH-1:0] wire_d87_85;
	wire [WIDTH-1:0] wire_d87_86;
	wire [WIDTH-1:0] wire_d87_87;
	wire [WIDTH-1:0] wire_d87_88;
	wire [WIDTH-1:0] wire_d87_89;
	wire [WIDTH-1:0] wire_d87_90;
	wire [WIDTH-1:0] wire_d87_91;
	wire [WIDTH-1:0] wire_d87_92;
	wire [WIDTH-1:0] wire_d87_93;
	wire [WIDTH-1:0] wire_d87_94;
	wire [WIDTH-1:0] wire_d87_95;
	wire [WIDTH-1:0] wire_d87_96;
	wire [WIDTH-1:0] wire_d87_97;
	wire [WIDTH-1:0] wire_d87_98;
	wire [WIDTH-1:0] wire_d88_0;
	wire [WIDTH-1:0] wire_d88_1;
	wire [WIDTH-1:0] wire_d88_2;
	wire [WIDTH-1:0] wire_d88_3;
	wire [WIDTH-1:0] wire_d88_4;
	wire [WIDTH-1:0] wire_d88_5;
	wire [WIDTH-1:0] wire_d88_6;
	wire [WIDTH-1:0] wire_d88_7;
	wire [WIDTH-1:0] wire_d88_8;
	wire [WIDTH-1:0] wire_d88_9;
	wire [WIDTH-1:0] wire_d88_10;
	wire [WIDTH-1:0] wire_d88_11;
	wire [WIDTH-1:0] wire_d88_12;
	wire [WIDTH-1:0] wire_d88_13;
	wire [WIDTH-1:0] wire_d88_14;
	wire [WIDTH-1:0] wire_d88_15;
	wire [WIDTH-1:0] wire_d88_16;
	wire [WIDTH-1:0] wire_d88_17;
	wire [WIDTH-1:0] wire_d88_18;
	wire [WIDTH-1:0] wire_d88_19;
	wire [WIDTH-1:0] wire_d88_20;
	wire [WIDTH-1:0] wire_d88_21;
	wire [WIDTH-1:0] wire_d88_22;
	wire [WIDTH-1:0] wire_d88_23;
	wire [WIDTH-1:0] wire_d88_24;
	wire [WIDTH-1:0] wire_d88_25;
	wire [WIDTH-1:0] wire_d88_26;
	wire [WIDTH-1:0] wire_d88_27;
	wire [WIDTH-1:0] wire_d88_28;
	wire [WIDTH-1:0] wire_d88_29;
	wire [WIDTH-1:0] wire_d88_30;
	wire [WIDTH-1:0] wire_d88_31;
	wire [WIDTH-1:0] wire_d88_32;
	wire [WIDTH-1:0] wire_d88_33;
	wire [WIDTH-1:0] wire_d88_34;
	wire [WIDTH-1:0] wire_d88_35;
	wire [WIDTH-1:0] wire_d88_36;
	wire [WIDTH-1:0] wire_d88_37;
	wire [WIDTH-1:0] wire_d88_38;
	wire [WIDTH-1:0] wire_d88_39;
	wire [WIDTH-1:0] wire_d88_40;
	wire [WIDTH-1:0] wire_d88_41;
	wire [WIDTH-1:0] wire_d88_42;
	wire [WIDTH-1:0] wire_d88_43;
	wire [WIDTH-1:0] wire_d88_44;
	wire [WIDTH-1:0] wire_d88_45;
	wire [WIDTH-1:0] wire_d88_46;
	wire [WIDTH-1:0] wire_d88_47;
	wire [WIDTH-1:0] wire_d88_48;
	wire [WIDTH-1:0] wire_d88_49;
	wire [WIDTH-1:0] wire_d88_50;
	wire [WIDTH-1:0] wire_d88_51;
	wire [WIDTH-1:0] wire_d88_52;
	wire [WIDTH-1:0] wire_d88_53;
	wire [WIDTH-1:0] wire_d88_54;
	wire [WIDTH-1:0] wire_d88_55;
	wire [WIDTH-1:0] wire_d88_56;
	wire [WIDTH-1:0] wire_d88_57;
	wire [WIDTH-1:0] wire_d88_58;
	wire [WIDTH-1:0] wire_d88_59;
	wire [WIDTH-1:0] wire_d88_60;
	wire [WIDTH-1:0] wire_d88_61;
	wire [WIDTH-1:0] wire_d88_62;
	wire [WIDTH-1:0] wire_d88_63;
	wire [WIDTH-1:0] wire_d88_64;
	wire [WIDTH-1:0] wire_d88_65;
	wire [WIDTH-1:0] wire_d88_66;
	wire [WIDTH-1:0] wire_d88_67;
	wire [WIDTH-1:0] wire_d88_68;
	wire [WIDTH-1:0] wire_d88_69;
	wire [WIDTH-1:0] wire_d88_70;
	wire [WIDTH-1:0] wire_d88_71;
	wire [WIDTH-1:0] wire_d88_72;
	wire [WIDTH-1:0] wire_d88_73;
	wire [WIDTH-1:0] wire_d88_74;
	wire [WIDTH-1:0] wire_d88_75;
	wire [WIDTH-1:0] wire_d88_76;
	wire [WIDTH-1:0] wire_d88_77;
	wire [WIDTH-1:0] wire_d88_78;
	wire [WIDTH-1:0] wire_d88_79;
	wire [WIDTH-1:0] wire_d88_80;
	wire [WIDTH-1:0] wire_d88_81;
	wire [WIDTH-1:0] wire_d88_82;
	wire [WIDTH-1:0] wire_d88_83;
	wire [WIDTH-1:0] wire_d88_84;
	wire [WIDTH-1:0] wire_d88_85;
	wire [WIDTH-1:0] wire_d88_86;
	wire [WIDTH-1:0] wire_d88_87;
	wire [WIDTH-1:0] wire_d88_88;
	wire [WIDTH-1:0] wire_d88_89;
	wire [WIDTH-1:0] wire_d88_90;
	wire [WIDTH-1:0] wire_d88_91;
	wire [WIDTH-1:0] wire_d88_92;
	wire [WIDTH-1:0] wire_d88_93;
	wire [WIDTH-1:0] wire_d88_94;
	wire [WIDTH-1:0] wire_d88_95;
	wire [WIDTH-1:0] wire_d88_96;
	wire [WIDTH-1:0] wire_d88_97;
	wire [WIDTH-1:0] wire_d88_98;
	wire [WIDTH-1:0] wire_d89_0;
	wire [WIDTH-1:0] wire_d89_1;
	wire [WIDTH-1:0] wire_d89_2;
	wire [WIDTH-1:0] wire_d89_3;
	wire [WIDTH-1:0] wire_d89_4;
	wire [WIDTH-1:0] wire_d89_5;
	wire [WIDTH-1:0] wire_d89_6;
	wire [WIDTH-1:0] wire_d89_7;
	wire [WIDTH-1:0] wire_d89_8;
	wire [WIDTH-1:0] wire_d89_9;
	wire [WIDTH-1:0] wire_d89_10;
	wire [WIDTH-1:0] wire_d89_11;
	wire [WIDTH-1:0] wire_d89_12;
	wire [WIDTH-1:0] wire_d89_13;
	wire [WIDTH-1:0] wire_d89_14;
	wire [WIDTH-1:0] wire_d89_15;
	wire [WIDTH-1:0] wire_d89_16;
	wire [WIDTH-1:0] wire_d89_17;
	wire [WIDTH-1:0] wire_d89_18;
	wire [WIDTH-1:0] wire_d89_19;
	wire [WIDTH-1:0] wire_d89_20;
	wire [WIDTH-1:0] wire_d89_21;
	wire [WIDTH-1:0] wire_d89_22;
	wire [WIDTH-1:0] wire_d89_23;
	wire [WIDTH-1:0] wire_d89_24;
	wire [WIDTH-1:0] wire_d89_25;
	wire [WIDTH-1:0] wire_d89_26;
	wire [WIDTH-1:0] wire_d89_27;
	wire [WIDTH-1:0] wire_d89_28;
	wire [WIDTH-1:0] wire_d89_29;
	wire [WIDTH-1:0] wire_d89_30;
	wire [WIDTH-1:0] wire_d89_31;
	wire [WIDTH-1:0] wire_d89_32;
	wire [WIDTH-1:0] wire_d89_33;
	wire [WIDTH-1:0] wire_d89_34;
	wire [WIDTH-1:0] wire_d89_35;
	wire [WIDTH-1:0] wire_d89_36;
	wire [WIDTH-1:0] wire_d89_37;
	wire [WIDTH-1:0] wire_d89_38;
	wire [WIDTH-1:0] wire_d89_39;
	wire [WIDTH-1:0] wire_d89_40;
	wire [WIDTH-1:0] wire_d89_41;
	wire [WIDTH-1:0] wire_d89_42;
	wire [WIDTH-1:0] wire_d89_43;
	wire [WIDTH-1:0] wire_d89_44;
	wire [WIDTH-1:0] wire_d89_45;
	wire [WIDTH-1:0] wire_d89_46;
	wire [WIDTH-1:0] wire_d89_47;
	wire [WIDTH-1:0] wire_d89_48;
	wire [WIDTH-1:0] wire_d89_49;
	wire [WIDTH-1:0] wire_d89_50;
	wire [WIDTH-1:0] wire_d89_51;
	wire [WIDTH-1:0] wire_d89_52;
	wire [WIDTH-1:0] wire_d89_53;
	wire [WIDTH-1:0] wire_d89_54;
	wire [WIDTH-1:0] wire_d89_55;
	wire [WIDTH-1:0] wire_d89_56;
	wire [WIDTH-1:0] wire_d89_57;
	wire [WIDTH-1:0] wire_d89_58;
	wire [WIDTH-1:0] wire_d89_59;
	wire [WIDTH-1:0] wire_d89_60;
	wire [WIDTH-1:0] wire_d89_61;
	wire [WIDTH-1:0] wire_d89_62;
	wire [WIDTH-1:0] wire_d89_63;
	wire [WIDTH-1:0] wire_d89_64;
	wire [WIDTH-1:0] wire_d89_65;
	wire [WIDTH-1:0] wire_d89_66;
	wire [WIDTH-1:0] wire_d89_67;
	wire [WIDTH-1:0] wire_d89_68;
	wire [WIDTH-1:0] wire_d89_69;
	wire [WIDTH-1:0] wire_d89_70;
	wire [WIDTH-1:0] wire_d89_71;
	wire [WIDTH-1:0] wire_d89_72;
	wire [WIDTH-1:0] wire_d89_73;
	wire [WIDTH-1:0] wire_d89_74;
	wire [WIDTH-1:0] wire_d89_75;
	wire [WIDTH-1:0] wire_d89_76;
	wire [WIDTH-1:0] wire_d89_77;
	wire [WIDTH-1:0] wire_d89_78;
	wire [WIDTH-1:0] wire_d89_79;
	wire [WIDTH-1:0] wire_d89_80;
	wire [WIDTH-1:0] wire_d89_81;
	wire [WIDTH-1:0] wire_d89_82;
	wire [WIDTH-1:0] wire_d89_83;
	wire [WIDTH-1:0] wire_d89_84;
	wire [WIDTH-1:0] wire_d89_85;
	wire [WIDTH-1:0] wire_d89_86;
	wire [WIDTH-1:0] wire_d89_87;
	wire [WIDTH-1:0] wire_d89_88;
	wire [WIDTH-1:0] wire_d89_89;
	wire [WIDTH-1:0] wire_d89_90;
	wire [WIDTH-1:0] wire_d89_91;
	wire [WIDTH-1:0] wire_d89_92;
	wire [WIDTH-1:0] wire_d89_93;
	wire [WIDTH-1:0] wire_d89_94;
	wire [WIDTH-1:0] wire_d89_95;
	wire [WIDTH-1:0] wire_d89_96;
	wire [WIDTH-1:0] wire_d89_97;
	wire [WIDTH-1:0] wire_d89_98;

	large_mux #(.WIDTH(WIDTH)) large_mux_instance100(.data_in(d_in0),.data_out(wire_d0_0),.clk(clk),.rst(rst));            //channel 1
	invertion #(.WIDTH(WIDTH)) invertion_instance101(.data_in(wire_d0_0),.data_out(wire_d0_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance102(.data_in(wire_d0_1),.data_out(wire_d0_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance103(.data_in(wire_d0_2),.data_out(wire_d0_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance104(.data_in(wire_d0_3),.data_out(wire_d0_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance105(.data_in(wire_d0_4),.data_out(wire_d0_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance106(.data_in(wire_d0_5),.data_out(wire_d0_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance107(.data_in(wire_d0_6),.data_out(wire_d0_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance108(.data_in(wire_d0_7),.data_out(wire_d0_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance109(.data_in(wire_d0_8),.data_out(wire_d0_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1010(.data_in(wire_d0_9),.data_out(wire_d0_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1011(.data_in(wire_d0_10),.data_out(wire_d0_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1012(.data_in(wire_d0_11),.data_out(wire_d0_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1013(.data_in(wire_d0_12),.data_out(wire_d0_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1014(.data_in(wire_d0_13),.data_out(wire_d0_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1015(.data_in(wire_d0_14),.data_out(wire_d0_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1016(.data_in(wire_d0_15),.data_out(wire_d0_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1017(.data_in(wire_d0_16),.data_out(wire_d0_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1018(.data_in(wire_d0_17),.data_out(wire_d0_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1019(.data_in(wire_d0_18),.data_out(wire_d0_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1020(.data_in(wire_d0_19),.data_out(wire_d0_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1021(.data_in(wire_d0_20),.data_out(wire_d0_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1022(.data_in(wire_d0_21),.data_out(wire_d0_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1023(.data_in(wire_d0_22),.data_out(wire_d0_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1024(.data_in(wire_d0_23),.data_out(wire_d0_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1025(.data_in(wire_d0_24),.data_out(wire_d0_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1026(.data_in(wire_d0_25),.data_out(wire_d0_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1027(.data_in(wire_d0_26),.data_out(wire_d0_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1028(.data_in(wire_d0_27),.data_out(wire_d0_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1029(.data_in(wire_d0_28),.data_out(wire_d0_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1030(.data_in(wire_d0_29),.data_out(wire_d0_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1031(.data_in(wire_d0_30),.data_out(wire_d0_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1032(.data_in(wire_d0_31),.data_out(wire_d0_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1033(.data_in(wire_d0_32),.data_out(wire_d0_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1034(.data_in(wire_d0_33),.data_out(wire_d0_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1035(.data_in(wire_d0_34),.data_out(wire_d0_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1036(.data_in(wire_d0_35),.data_out(wire_d0_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1037(.data_in(wire_d0_36),.data_out(wire_d0_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1038(.data_in(wire_d0_37),.data_out(wire_d0_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1039(.data_in(wire_d0_38),.data_out(wire_d0_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1040(.data_in(wire_d0_39),.data_out(wire_d0_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1041(.data_in(wire_d0_40),.data_out(wire_d0_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1042(.data_in(wire_d0_41),.data_out(wire_d0_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1043(.data_in(wire_d0_42),.data_out(wire_d0_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1044(.data_in(wire_d0_43),.data_out(wire_d0_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1045(.data_in(wire_d0_44),.data_out(wire_d0_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1046(.data_in(wire_d0_45),.data_out(wire_d0_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1047(.data_in(wire_d0_46),.data_out(wire_d0_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1048(.data_in(wire_d0_47),.data_out(wire_d0_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1049(.data_in(wire_d0_48),.data_out(wire_d0_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1050(.data_in(wire_d0_49),.data_out(wire_d0_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1051(.data_in(wire_d0_50),.data_out(wire_d0_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1052(.data_in(wire_d0_51),.data_out(wire_d0_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1053(.data_in(wire_d0_52),.data_out(wire_d0_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1054(.data_in(wire_d0_53),.data_out(wire_d0_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1055(.data_in(wire_d0_54),.data_out(wire_d0_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1056(.data_in(wire_d0_55),.data_out(wire_d0_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1057(.data_in(wire_d0_56),.data_out(wire_d0_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1058(.data_in(wire_d0_57),.data_out(wire_d0_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1059(.data_in(wire_d0_58),.data_out(wire_d0_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1060(.data_in(wire_d0_59),.data_out(wire_d0_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1061(.data_in(wire_d0_60),.data_out(wire_d0_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1062(.data_in(wire_d0_61),.data_out(wire_d0_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1063(.data_in(wire_d0_62),.data_out(wire_d0_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1064(.data_in(wire_d0_63),.data_out(wire_d0_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1065(.data_in(wire_d0_64),.data_out(wire_d0_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1066(.data_in(wire_d0_65),.data_out(wire_d0_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1067(.data_in(wire_d0_66),.data_out(wire_d0_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1068(.data_in(wire_d0_67),.data_out(wire_d0_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1069(.data_in(wire_d0_68),.data_out(wire_d0_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1070(.data_in(wire_d0_69),.data_out(wire_d0_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1071(.data_in(wire_d0_70),.data_out(wire_d0_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1072(.data_in(wire_d0_71),.data_out(wire_d0_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1073(.data_in(wire_d0_72),.data_out(wire_d0_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1074(.data_in(wire_d0_73),.data_out(wire_d0_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1075(.data_in(wire_d0_74),.data_out(wire_d0_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1076(.data_in(wire_d0_75),.data_out(wire_d0_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1077(.data_in(wire_d0_76),.data_out(wire_d0_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1078(.data_in(wire_d0_77),.data_out(wire_d0_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1079(.data_in(wire_d0_78),.data_out(wire_d0_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1080(.data_in(wire_d0_79),.data_out(wire_d0_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1081(.data_in(wire_d0_80),.data_out(wire_d0_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1082(.data_in(wire_d0_81),.data_out(wire_d0_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1083(.data_in(wire_d0_82),.data_out(wire_d0_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1084(.data_in(wire_d0_83),.data_out(wire_d0_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1085(.data_in(wire_d0_84),.data_out(wire_d0_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1086(.data_in(wire_d0_85),.data_out(wire_d0_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1087(.data_in(wire_d0_86),.data_out(wire_d0_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1088(.data_in(wire_d0_87),.data_out(wire_d0_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1089(.data_in(wire_d0_88),.data_out(wire_d0_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1090(.data_in(wire_d0_89),.data_out(wire_d0_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1091(.data_in(wire_d0_90),.data_out(wire_d0_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1092(.data_in(wire_d0_91),.data_out(wire_d0_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1093(.data_in(wire_d0_92),.data_out(wire_d0_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1094(.data_in(wire_d0_93),.data_out(wire_d0_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1095(.data_in(wire_d0_94),.data_out(wire_d0_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1096(.data_in(wire_d0_95),.data_out(wire_d0_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1097(.data_in(wire_d0_96),.data_out(wire_d0_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1098(.data_in(wire_d0_97),.data_out(wire_d0_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1099(.data_in(wire_d0_98),.data_out(d_out0),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance210(.data_in(d_in1),.data_out(wire_d1_0),.clk(clk),.rst(rst));            //channel 2
	encoder #(.WIDTH(WIDTH)) encoder_instance211(.data_in(wire_d1_0),.data_out(wire_d1_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212(.data_in(wire_d1_1),.data_out(wire_d1_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance213(.data_in(wire_d1_2),.data_out(wire_d1_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance214(.data_in(wire_d1_3),.data_out(wire_d1_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance215(.data_in(wire_d1_4),.data_out(wire_d1_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance216(.data_in(wire_d1_5),.data_out(wire_d1_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance217(.data_in(wire_d1_6),.data_out(wire_d1_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance218(.data_in(wire_d1_7),.data_out(wire_d1_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance219(.data_in(wire_d1_8),.data_out(wire_d1_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2110(.data_in(wire_d1_9),.data_out(wire_d1_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2111(.data_in(wire_d1_10),.data_out(wire_d1_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2112(.data_in(wire_d1_11),.data_out(wire_d1_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2113(.data_in(wire_d1_12),.data_out(wire_d1_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2114(.data_in(wire_d1_13),.data_out(wire_d1_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2115(.data_in(wire_d1_14),.data_out(wire_d1_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2116(.data_in(wire_d1_15),.data_out(wire_d1_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2117(.data_in(wire_d1_16),.data_out(wire_d1_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2118(.data_in(wire_d1_17),.data_out(wire_d1_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2119(.data_in(wire_d1_18),.data_out(wire_d1_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2120(.data_in(wire_d1_19),.data_out(wire_d1_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2121(.data_in(wire_d1_20),.data_out(wire_d1_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2122(.data_in(wire_d1_21),.data_out(wire_d1_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2123(.data_in(wire_d1_22),.data_out(wire_d1_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2124(.data_in(wire_d1_23),.data_out(wire_d1_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2125(.data_in(wire_d1_24),.data_out(wire_d1_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2126(.data_in(wire_d1_25),.data_out(wire_d1_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2127(.data_in(wire_d1_26),.data_out(wire_d1_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2128(.data_in(wire_d1_27),.data_out(wire_d1_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2129(.data_in(wire_d1_28),.data_out(wire_d1_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2130(.data_in(wire_d1_29),.data_out(wire_d1_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2131(.data_in(wire_d1_30),.data_out(wire_d1_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2132(.data_in(wire_d1_31),.data_out(wire_d1_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2133(.data_in(wire_d1_32),.data_out(wire_d1_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2134(.data_in(wire_d1_33),.data_out(wire_d1_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2135(.data_in(wire_d1_34),.data_out(wire_d1_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2136(.data_in(wire_d1_35),.data_out(wire_d1_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2137(.data_in(wire_d1_36),.data_out(wire_d1_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2138(.data_in(wire_d1_37),.data_out(wire_d1_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2139(.data_in(wire_d1_38),.data_out(wire_d1_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2140(.data_in(wire_d1_39),.data_out(wire_d1_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2141(.data_in(wire_d1_40),.data_out(wire_d1_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2142(.data_in(wire_d1_41),.data_out(wire_d1_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2143(.data_in(wire_d1_42),.data_out(wire_d1_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2144(.data_in(wire_d1_43),.data_out(wire_d1_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2145(.data_in(wire_d1_44),.data_out(wire_d1_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2146(.data_in(wire_d1_45),.data_out(wire_d1_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2147(.data_in(wire_d1_46),.data_out(wire_d1_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2148(.data_in(wire_d1_47),.data_out(wire_d1_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2149(.data_in(wire_d1_48),.data_out(wire_d1_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2150(.data_in(wire_d1_49),.data_out(wire_d1_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2151(.data_in(wire_d1_50),.data_out(wire_d1_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2152(.data_in(wire_d1_51),.data_out(wire_d1_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2153(.data_in(wire_d1_52),.data_out(wire_d1_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2154(.data_in(wire_d1_53),.data_out(wire_d1_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2155(.data_in(wire_d1_54),.data_out(wire_d1_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2156(.data_in(wire_d1_55),.data_out(wire_d1_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2157(.data_in(wire_d1_56),.data_out(wire_d1_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2158(.data_in(wire_d1_57),.data_out(wire_d1_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2159(.data_in(wire_d1_58),.data_out(wire_d1_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2160(.data_in(wire_d1_59),.data_out(wire_d1_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2161(.data_in(wire_d1_60),.data_out(wire_d1_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2162(.data_in(wire_d1_61),.data_out(wire_d1_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2163(.data_in(wire_d1_62),.data_out(wire_d1_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2164(.data_in(wire_d1_63),.data_out(wire_d1_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2165(.data_in(wire_d1_64),.data_out(wire_d1_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2166(.data_in(wire_d1_65),.data_out(wire_d1_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2167(.data_in(wire_d1_66),.data_out(wire_d1_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2168(.data_in(wire_d1_67),.data_out(wire_d1_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2169(.data_in(wire_d1_68),.data_out(wire_d1_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2170(.data_in(wire_d1_69),.data_out(wire_d1_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2171(.data_in(wire_d1_70),.data_out(wire_d1_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2172(.data_in(wire_d1_71),.data_out(wire_d1_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2173(.data_in(wire_d1_72),.data_out(wire_d1_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2174(.data_in(wire_d1_73),.data_out(wire_d1_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2175(.data_in(wire_d1_74),.data_out(wire_d1_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2176(.data_in(wire_d1_75),.data_out(wire_d1_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2177(.data_in(wire_d1_76),.data_out(wire_d1_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2178(.data_in(wire_d1_77),.data_out(wire_d1_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2179(.data_in(wire_d1_78),.data_out(wire_d1_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2180(.data_in(wire_d1_79),.data_out(wire_d1_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2181(.data_in(wire_d1_80),.data_out(wire_d1_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2182(.data_in(wire_d1_81),.data_out(wire_d1_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2183(.data_in(wire_d1_82),.data_out(wire_d1_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2184(.data_in(wire_d1_83),.data_out(wire_d1_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2185(.data_in(wire_d1_84),.data_out(wire_d1_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2186(.data_in(wire_d1_85),.data_out(wire_d1_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2187(.data_in(wire_d1_86),.data_out(wire_d1_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2188(.data_in(wire_d1_87),.data_out(wire_d1_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2189(.data_in(wire_d1_88),.data_out(wire_d1_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2190(.data_in(wire_d1_89),.data_out(wire_d1_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2191(.data_in(wire_d1_90),.data_out(wire_d1_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2192(.data_in(wire_d1_91),.data_out(wire_d1_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2193(.data_in(wire_d1_92),.data_out(wire_d1_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2194(.data_in(wire_d1_93),.data_out(wire_d1_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2195(.data_in(wire_d1_94),.data_out(wire_d1_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2196(.data_in(wire_d1_95),.data_out(wire_d1_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2197(.data_in(wire_d1_96),.data_out(wire_d1_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2198(.data_in(wire_d1_97),.data_out(wire_d1_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2199(.data_in(wire_d1_98),.data_out(d_out1),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance320(.data_in(d_in2),.data_out(wire_d2_0),.clk(clk),.rst(rst));            //channel 3
	encoder #(.WIDTH(WIDTH)) encoder_instance321(.data_in(wire_d2_0),.data_out(wire_d2_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance322(.data_in(wire_d2_1),.data_out(wire_d2_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323(.data_in(wire_d2_2),.data_out(wire_d2_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance324(.data_in(wire_d2_3),.data_out(wire_d2_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance325(.data_in(wire_d2_4),.data_out(wire_d2_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance326(.data_in(wire_d2_5),.data_out(wire_d2_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance327(.data_in(wire_d2_6),.data_out(wire_d2_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance328(.data_in(wire_d2_7),.data_out(wire_d2_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance329(.data_in(wire_d2_8),.data_out(wire_d2_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3210(.data_in(wire_d2_9),.data_out(wire_d2_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3211(.data_in(wire_d2_10),.data_out(wire_d2_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3212(.data_in(wire_d2_11),.data_out(wire_d2_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3213(.data_in(wire_d2_12),.data_out(wire_d2_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3214(.data_in(wire_d2_13),.data_out(wire_d2_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3215(.data_in(wire_d2_14),.data_out(wire_d2_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3216(.data_in(wire_d2_15),.data_out(wire_d2_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3217(.data_in(wire_d2_16),.data_out(wire_d2_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3218(.data_in(wire_d2_17),.data_out(wire_d2_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3219(.data_in(wire_d2_18),.data_out(wire_d2_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3220(.data_in(wire_d2_19),.data_out(wire_d2_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3221(.data_in(wire_d2_20),.data_out(wire_d2_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3222(.data_in(wire_d2_21),.data_out(wire_d2_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3223(.data_in(wire_d2_22),.data_out(wire_d2_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3224(.data_in(wire_d2_23),.data_out(wire_d2_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3225(.data_in(wire_d2_24),.data_out(wire_d2_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3226(.data_in(wire_d2_25),.data_out(wire_d2_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3227(.data_in(wire_d2_26),.data_out(wire_d2_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3228(.data_in(wire_d2_27),.data_out(wire_d2_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3229(.data_in(wire_d2_28),.data_out(wire_d2_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3230(.data_in(wire_d2_29),.data_out(wire_d2_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3231(.data_in(wire_d2_30),.data_out(wire_d2_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3232(.data_in(wire_d2_31),.data_out(wire_d2_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3233(.data_in(wire_d2_32),.data_out(wire_d2_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3234(.data_in(wire_d2_33),.data_out(wire_d2_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3235(.data_in(wire_d2_34),.data_out(wire_d2_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3236(.data_in(wire_d2_35),.data_out(wire_d2_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3237(.data_in(wire_d2_36),.data_out(wire_d2_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3238(.data_in(wire_d2_37),.data_out(wire_d2_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3239(.data_in(wire_d2_38),.data_out(wire_d2_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3240(.data_in(wire_d2_39),.data_out(wire_d2_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3241(.data_in(wire_d2_40),.data_out(wire_d2_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3242(.data_in(wire_d2_41),.data_out(wire_d2_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3243(.data_in(wire_d2_42),.data_out(wire_d2_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3244(.data_in(wire_d2_43),.data_out(wire_d2_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3245(.data_in(wire_d2_44),.data_out(wire_d2_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3246(.data_in(wire_d2_45),.data_out(wire_d2_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3247(.data_in(wire_d2_46),.data_out(wire_d2_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3248(.data_in(wire_d2_47),.data_out(wire_d2_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3249(.data_in(wire_d2_48),.data_out(wire_d2_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3250(.data_in(wire_d2_49),.data_out(wire_d2_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3251(.data_in(wire_d2_50),.data_out(wire_d2_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3252(.data_in(wire_d2_51),.data_out(wire_d2_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3253(.data_in(wire_d2_52),.data_out(wire_d2_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3254(.data_in(wire_d2_53),.data_out(wire_d2_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3255(.data_in(wire_d2_54),.data_out(wire_d2_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3256(.data_in(wire_d2_55),.data_out(wire_d2_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3257(.data_in(wire_d2_56),.data_out(wire_d2_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3258(.data_in(wire_d2_57),.data_out(wire_d2_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3259(.data_in(wire_d2_58),.data_out(wire_d2_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3260(.data_in(wire_d2_59),.data_out(wire_d2_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3261(.data_in(wire_d2_60),.data_out(wire_d2_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3262(.data_in(wire_d2_61),.data_out(wire_d2_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3263(.data_in(wire_d2_62),.data_out(wire_d2_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3264(.data_in(wire_d2_63),.data_out(wire_d2_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3265(.data_in(wire_d2_64),.data_out(wire_d2_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3266(.data_in(wire_d2_65),.data_out(wire_d2_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3267(.data_in(wire_d2_66),.data_out(wire_d2_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3268(.data_in(wire_d2_67),.data_out(wire_d2_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3269(.data_in(wire_d2_68),.data_out(wire_d2_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3270(.data_in(wire_d2_69),.data_out(wire_d2_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3271(.data_in(wire_d2_70),.data_out(wire_d2_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3272(.data_in(wire_d2_71),.data_out(wire_d2_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3273(.data_in(wire_d2_72),.data_out(wire_d2_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3274(.data_in(wire_d2_73),.data_out(wire_d2_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3275(.data_in(wire_d2_74),.data_out(wire_d2_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3276(.data_in(wire_d2_75),.data_out(wire_d2_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3277(.data_in(wire_d2_76),.data_out(wire_d2_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3278(.data_in(wire_d2_77),.data_out(wire_d2_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3279(.data_in(wire_d2_78),.data_out(wire_d2_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3280(.data_in(wire_d2_79),.data_out(wire_d2_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3281(.data_in(wire_d2_80),.data_out(wire_d2_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3282(.data_in(wire_d2_81),.data_out(wire_d2_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3283(.data_in(wire_d2_82),.data_out(wire_d2_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3284(.data_in(wire_d2_83),.data_out(wire_d2_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3285(.data_in(wire_d2_84),.data_out(wire_d2_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3286(.data_in(wire_d2_85),.data_out(wire_d2_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3287(.data_in(wire_d2_86),.data_out(wire_d2_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3288(.data_in(wire_d2_87),.data_out(wire_d2_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3289(.data_in(wire_d2_88),.data_out(wire_d2_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3290(.data_in(wire_d2_89),.data_out(wire_d2_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3291(.data_in(wire_d2_90),.data_out(wire_d2_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3292(.data_in(wire_d2_91),.data_out(wire_d2_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3293(.data_in(wire_d2_92),.data_out(wire_d2_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3294(.data_in(wire_d2_93),.data_out(wire_d2_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3295(.data_in(wire_d2_94),.data_out(wire_d2_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3296(.data_in(wire_d2_95),.data_out(wire_d2_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3297(.data_in(wire_d2_96),.data_out(wire_d2_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3298(.data_in(wire_d2_97),.data_out(wire_d2_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3299(.data_in(wire_d2_98),.data_out(d_out2),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance430(.data_in(d_in3),.data_out(wire_d3_0),.clk(clk),.rst(rst));            //channel 4
	encoder #(.WIDTH(WIDTH)) encoder_instance431(.data_in(wire_d3_0),.data_out(wire_d3_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance432(.data_in(wire_d3_1),.data_out(wire_d3_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance433(.data_in(wire_d3_2),.data_out(wire_d3_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434(.data_in(wire_d3_3),.data_out(wire_d3_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance435(.data_in(wire_d3_4),.data_out(wire_d3_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance436(.data_in(wire_d3_5),.data_out(wire_d3_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance437(.data_in(wire_d3_6),.data_out(wire_d3_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance438(.data_in(wire_d3_7),.data_out(wire_d3_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance439(.data_in(wire_d3_8),.data_out(wire_d3_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4310(.data_in(wire_d3_9),.data_out(wire_d3_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4311(.data_in(wire_d3_10),.data_out(wire_d3_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4312(.data_in(wire_d3_11),.data_out(wire_d3_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4313(.data_in(wire_d3_12),.data_out(wire_d3_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4314(.data_in(wire_d3_13),.data_out(wire_d3_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4315(.data_in(wire_d3_14),.data_out(wire_d3_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4316(.data_in(wire_d3_15),.data_out(wire_d3_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4317(.data_in(wire_d3_16),.data_out(wire_d3_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4318(.data_in(wire_d3_17),.data_out(wire_d3_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4319(.data_in(wire_d3_18),.data_out(wire_d3_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4320(.data_in(wire_d3_19),.data_out(wire_d3_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4321(.data_in(wire_d3_20),.data_out(wire_d3_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4322(.data_in(wire_d3_21),.data_out(wire_d3_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4323(.data_in(wire_d3_22),.data_out(wire_d3_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4324(.data_in(wire_d3_23),.data_out(wire_d3_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4325(.data_in(wire_d3_24),.data_out(wire_d3_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4326(.data_in(wire_d3_25),.data_out(wire_d3_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4327(.data_in(wire_d3_26),.data_out(wire_d3_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4328(.data_in(wire_d3_27),.data_out(wire_d3_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4329(.data_in(wire_d3_28),.data_out(wire_d3_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4330(.data_in(wire_d3_29),.data_out(wire_d3_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4331(.data_in(wire_d3_30),.data_out(wire_d3_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4332(.data_in(wire_d3_31),.data_out(wire_d3_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4333(.data_in(wire_d3_32),.data_out(wire_d3_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4334(.data_in(wire_d3_33),.data_out(wire_d3_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4335(.data_in(wire_d3_34),.data_out(wire_d3_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4336(.data_in(wire_d3_35),.data_out(wire_d3_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4337(.data_in(wire_d3_36),.data_out(wire_d3_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4338(.data_in(wire_d3_37),.data_out(wire_d3_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4339(.data_in(wire_d3_38),.data_out(wire_d3_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4340(.data_in(wire_d3_39),.data_out(wire_d3_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4341(.data_in(wire_d3_40),.data_out(wire_d3_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4342(.data_in(wire_d3_41),.data_out(wire_d3_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4343(.data_in(wire_d3_42),.data_out(wire_d3_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4344(.data_in(wire_d3_43),.data_out(wire_d3_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4345(.data_in(wire_d3_44),.data_out(wire_d3_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4346(.data_in(wire_d3_45),.data_out(wire_d3_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4347(.data_in(wire_d3_46),.data_out(wire_d3_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4348(.data_in(wire_d3_47),.data_out(wire_d3_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4349(.data_in(wire_d3_48),.data_out(wire_d3_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4350(.data_in(wire_d3_49),.data_out(wire_d3_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4351(.data_in(wire_d3_50),.data_out(wire_d3_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4352(.data_in(wire_d3_51),.data_out(wire_d3_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4353(.data_in(wire_d3_52),.data_out(wire_d3_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4354(.data_in(wire_d3_53),.data_out(wire_d3_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4355(.data_in(wire_d3_54),.data_out(wire_d3_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4356(.data_in(wire_d3_55),.data_out(wire_d3_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4357(.data_in(wire_d3_56),.data_out(wire_d3_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4358(.data_in(wire_d3_57),.data_out(wire_d3_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4359(.data_in(wire_d3_58),.data_out(wire_d3_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4360(.data_in(wire_d3_59),.data_out(wire_d3_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4361(.data_in(wire_d3_60),.data_out(wire_d3_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4362(.data_in(wire_d3_61),.data_out(wire_d3_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4363(.data_in(wire_d3_62),.data_out(wire_d3_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4364(.data_in(wire_d3_63),.data_out(wire_d3_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4365(.data_in(wire_d3_64),.data_out(wire_d3_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4366(.data_in(wire_d3_65),.data_out(wire_d3_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4367(.data_in(wire_d3_66),.data_out(wire_d3_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4368(.data_in(wire_d3_67),.data_out(wire_d3_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4369(.data_in(wire_d3_68),.data_out(wire_d3_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4370(.data_in(wire_d3_69),.data_out(wire_d3_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4371(.data_in(wire_d3_70),.data_out(wire_d3_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4372(.data_in(wire_d3_71),.data_out(wire_d3_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4373(.data_in(wire_d3_72),.data_out(wire_d3_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4374(.data_in(wire_d3_73),.data_out(wire_d3_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4375(.data_in(wire_d3_74),.data_out(wire_d3_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4376(.data_in(wire_d3_75),.data_out(wire_d3_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4377(.data_in(wire_d3_76),.data_out(wire_d3_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4378(.data_in(wire_d3_77),.data_out(wire_d3_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4379(.data_in(wire_d3_78),.data_out(wire_d3_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4380(.data_in(wire_d3_79),.data_out(wire_d3_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4381(.data_in(wire_d3_80),.data_out(wire_d3_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4382(.data_in(wire_d3_81),.data_out(wire_d3_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4383(.data_in(wire_d3_82),.data_out(wire_d3_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4384(.data_in(wire_d3_83),.data_out(wire_d3_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4385(.data_in(wire_d3_84),.data_out(wire_d3_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4386(.data_in(wire_d3_85),.data_out(wire_d3_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4387(.data_in(wire_d3_86),.data_out(wire_d3_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4388(.data_in(wire_d3_87),.data_out(wire_d3_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4389(.data_in(wire_d3_88),.data_out(wire_d3_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4390(.data_in(wire_d3_89),.data_out(wire_d3_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4391(.data_in(wire_d3_90),.data_out(wire_d3_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4392(.data_in(wire_d3_91),.data_out(wire_d3_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4393(.data_in(wire_d3_92),.data_out(wire_d3_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4394(.data_in(wire_d3_93),.data_out(wire_d3_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4395(.data_in(wire_d3_94),.data_out(wire_d3_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4396(.data_in(wire_d3_95),.data_out(wire_d3_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4397(.data_in(wire_d3_96),.data_out(wire_d3_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4398(.data_in(wire_d3_97),.data_out(wire_d3_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4399(.data_in(wire_d3_98),.data_out(d_out3),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance540(.data_in(d_in4),.data_out(wire_d4_0),.clk(clk),.rst(rst));            //channel 5
	invertion #(.WIDTH(WIDTH)) invertion_instance541(.data_in(wire_d4_0),.data_out(wire_d4_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance542(.data_in(wire_d4_1),.data_out(wire_d4_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance543(.data_in(wire_d4_2),.data_out(wire_d4_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance544(.data_in(wire_d4_3),.data_out(wire_d4_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545(.data_in(wire_d4_4),.data_out(wire_d4_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance546(.data_in(wire_d4_5),.data_out(wire_d4_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance547(.data_in(wire_d4_6),.data_out(wire_d4_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance548(.data_in(wire_d4_7),.data_out(wire_d4_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance549(.data_in(wire_d4_8),.data_out(wire_d4_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5410(.data_in(wire_d4_9),.data_out(wire_d4_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5411(.data_in(wire_d4_10),.data_out(wire_d4_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5412(.data_in(wire_d4_11),.data_out(wire_d4_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5413(.data_in(wire_d4_12),.data_out(wire_d4_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5414(.data_in(wire_d4_13),.data_out(wire_d4_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5415(.data_in(wire_d4_14),.data_out(wire_d4_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5416(.data_in(wire_d4_15),.data_out(wire_d4_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5417(.data_in(wire_d4_16),.data_out(wire_d4_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5418(.data_in(wire_d4_17),.data_out(wire_d4_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5419(.data_in(wire_d4_18),.data_out(wire_d4_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5420(.data_in(wire_d4_19),.data_out(wire_d4_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5421(.data_in(wire_d4_20),.data_out(wire_d4_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5422(.data_in(wire_d4_21),.data_out(wire_d4_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5423(.data_in(wire_d4_22),.data_out(wire_d4_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5424(.data_in(wire_d4_23),.data_out(wire_d4_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5425(.data_in(wire_d4_24),.data_out(wire_d4_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5426(.data_in(wire_d4_25),.data_out(wire_d4_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5427(.data_in(wire_d4_26),.data_out(wire_d4_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5428(.data_in(wire_d4_27),.data_out(wire_d4_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5429(.data_in(wire_d4_28),.data_out(wire_d4_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5430(.data_in(wire_d4_29),.data_out(wire_d4_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5431(.data_in(wire_d4_30),.data_out(wire_d4_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5432(.data_in(wire_d4_31),.data_out(wire_d4_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5433(.data_in(wire_d4_32),.data_out(wire_d4_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5434(.data_in(wire_d4_33),.data_out(wire_d4_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5435(.data_in(wire_d4_34),.data_out(wire_d4_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5436(.data_in(wire_d4_35),.data_out(wire_d4_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5437(.data_in(wire_d4_36),.data_out(wire_d4_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5438(.data_in(wire_d4_37),.data_out(wire_d4_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5439(.data_in(wire_d4_38),.data_out(wire_d4_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5440(.data_in(wire_d4_39),.data_out(wire_d4_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5441(.data_in(wire_d4_40),.data_out(wire_d4_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5442(.data_in(wire_d4_41),.data_out(wire_d4_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5443(.data_in(wire_d4_42),.data_out(wire_d4_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5444(.data_in(wire_d4_43),.data_out(wire_d4_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5445(.data_in(wire_d4_44),.data_out(wire_d4_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5446(.data_in(wire_d4_45),.data_out(wire_d4_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5447(.data_in(wire_d4_46),.data_out(wire_d4_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5448(.data_in(wire_d4_47),.data_out(wire_d4_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5449(.data_in(wire_d4_48),.data_out(wire_d4_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5450(.data_in(wire_d4_49),.data_out(wire_d4_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5451(.data_in(wire_d4_50),.data_out(wire_d4_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5452(.data_in(wire_d4_51),.data_out(wire_d4_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5453(.data_in(wire_d4_52),.data_out(wire_d4_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5454(.data_in(wire_d4_53),.data_out(wire_d4_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5455(.data_in(wire_d4_54),.data_out(wire_d4_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5456(.data_in(wire_d4_55),.data_out(wire_d4_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5457(.data_in(wire_d4_56),.data_out(wire_d4_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5458(.data_in(wire_d4_57),.data_out(wire_d4_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5459(.data_in(wire_d4_58),.data_out(wire_d4_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5460(.data_in(wire_d4_59),.data_out(wire_d4_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5461(.data_in(wire_d4_60),.data_out(wire_d4_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5462(.data_in(wire_d4_61),.data_out(wire_d4_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5463(.data_in(wire_d4_62),.data_out(wire_d4_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5464(.data_in(wire_d4_63),.data_out(wire_d4_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5465(.data_in(wire_d4_64),.data_out(wire_d4_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5466(.data_in(wire_d4_65),.data_out(wire_d4_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5467(.data_in(wire_d4_66),.data_out(wire_d4_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5468(.data_in(wire_d4_67),.data_out(wire_d4_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5469(.data_in(wire_d4_68),.data_out(wire_d4_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5470(.data_in(wire_d4_69),.data_out(wire_d4_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5471(.data_in(wire_d4_70),.data_out(wire_d4_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5472(.data_in(wire_d4_71),.data_out(wire_d4_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5473(.data_in(wire_d4_72),.data_out(wire_d4_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5474(.data_in(wire_d4_73),.data_out(wire_d4_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5475(.data_in(wire_d4_74),.data_out(wire_d4_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5476(.data_in(wire_d4_75),.data_out(wire_d4_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5477(.data_in(wire_d4_76),.data_out(wire_d4_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5478(.data_in(wire_d4_77),.data_out(wire_d4_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5479(.data_in(wire_d4_78),.data_out(wire_d4_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5480(.data_in(wire_d4_79),.data_out(wire_d4_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5481(.data_in(wire_d4_80),.data_out(wire_d4_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5482(.data_in(wire_d4_81),.data_out(wire_d4_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5483(.data_in(wire_d4_82),.data_out(wire_d4_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5484(.data_in(wire_d4_83),.data_out(wire_d4_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5485(.data_in(wire_d4_84),.data_out(wire_d4_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5486(.data_in(wire_d4_85),.data_out(wire_d4_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5487(.data_in(wire_d4_86),.data_out(wire_d4_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5488(.data_in(wire_d4_87),.data_out(wire_d4_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5489(.data_in(wire_d4_88),.data_out(wire_d4_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5490(.data_in(wire_d4_89),.data_out(wire_d4_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5491(.data_in(wire_d4_90),.data_out(wire_d4_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5492(.data_in(wire_d4_91),.data_out(wire_d4_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5493(.data_in(wire_d4_92),.data_out(wire_d4_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5494(.data_in(wire_d4_93),.data_out(wire_d4_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5495(.data_in(wire_d4_94),.data_out(wire_d4_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5496(.data_in(wire_d4_95),.data_out(wire_d4_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5497(.data_in(wire_d4_96),.data_out(wire_d4_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5498(.data_in(wire_d4_97),.data_out(wire_d4_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5499(.data_in(wire_d4_98),.data_out(d_out4),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance650(.data_in(d_in5),.data_out(wire_d5_0),.clk(clk),.rst(rst));            //channel 6
	register #(.WIDTH(WIDTH)) register_instance651(.data_in(wire_d5_0),.data_out(wire_d5_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance652(.data_in(wire_d5_1),.data_out(wire_d5_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance653(.data_in(wire_d5_2),.data_out(wire_d5_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance654(.data_in(wire_d5_3),.data_out(wire_d5_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance655(.data_in(wire_d5_4),.data_out(wire_d5_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656(.data_in(wire_d5_5),.data_out(wire_d5_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance657(.data_in(wire_d5_6),.data_out(wire_d5_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance658(.data_in(wire_d5_7),.data_out(wire_d5_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance659(.data_in(wire_d5_8),.data_out(wire_d5_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6510(.data_in(wire_d5_9),.data_out(wire_d5_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6511(.data_in(wire_d5_10),.data_out(wire_d5_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6512(.data_in(wire_d5_11),.data_out(wire_d5_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6513(.data_in(wire_d5_12),.data_out(wire_d5_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6514(.data_in(wire_d5_13),.data_out(wire_d5_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6515(.data_in(wire_d5_14),.data_out(wire_d5_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6516(.data_in(wire_d5_15),.data_out(wire_d5_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6517(.data_in(wire_d5_16),.data_out(wire_d5_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6518(.data_in(wire_d5_17),.data_out(wire_d5_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6519(.data_in(wire_d5_18),.data_out(wire_d5_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6520(.data_in(wire_d5_19),.data_out(wire_d5_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6521(.data_in(wire_d5_20),.data_out(wire_d5_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6522(.data_in(wire_d5_21),.data_out(wire_d5_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6523(.data_in(wire_d5_22),.data_out(wire_d5_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6524(.data_in(wire_d5_23),.data_out(wire_d5_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6525(.data_in(wire_d5_24),.data_out(wire_d5_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6526(.data_in(wire_d5_25),.data_out(wire_d5_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6527(.data_in(wire_d5_26),.data_out(wire_d5_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6528(.data_in(wire_d5_27),.data_out(wire_d5_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6529(.data_in(wire_d5_28),.data_out(wire_d5_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6530(.data_in(wire_d5_29),.data_out(wire_d5_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6531(.data_in(wire_d5_30),.data_out(wire_d5_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6532(.data_in(wire_d5_31),.data_out(wire_d5_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6533(.data_in(wire_d5_32),.data_out(wire_d5_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6534(.data_in(wire_d5_33),.data_out(wire_d5_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6535(.data_in(wire_d5_34),.data_out(wire_d5_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6536(.data_in(wire_d5_35),.data_out(wire_d5_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6537(.data_in(wire_d5_36),.data_out(wire_d5_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6538(.data_in(wire_d5_37),.data_out(wire_d5_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6539(.data_in(wire_d5_38),.data_out(wire_d5_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6540(.data_in(wire_d5_39),.data_out(wire_d5_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6541(.data_in(wire_d5_40),.data_out(wire_d5_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6542(.data_in(wire_d5_41),.data_out(wire_d5_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6543(.data_in(wire_d5_42),.data_out(wire_d5_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6544(.data_in(wire_d5_43),.data_out(wire_d5_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6545(.data_in(wire_d5_44),.data_out(wire_d5_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6546(.data_in(wire_d5_45),.data_out(wire_d5_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6547(.data_in(wire_d5_46),.data_out(wire_d5_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6548(.data_in(wire_d5_47),.data_out(wire_d5_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6549(.data_in(wire_d5_48),.data_out(wire_d5_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6550(.data_in(wire_d5_49),.data_out(wire_d5_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6551(.data_in(wire_d5_50),.data_out(wire_d5_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6552(.data_in(wire_d5_51),.data_out(wire_d5_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6553(.data_in(wire_d5_52),.data_out(wire_d5_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6554(.data_in(wire_d5_53),.data_out(wire_d5_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6555(.data_in(wire_d5_54),.data_out(wire_d5_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6556(.data_in(wire_d5_55),.data_out(wire_d5_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6557(.data_in(wire_d5_56),.data_out(wire_d5_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6558(.data_in(wire_d5_57),.data_out(wire_d5_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6559(.data_in(wire_d5_58),.data_out(wire_d5_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6560(.data_in(wire_d5_59),.data_out(wire_d5_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6561(.data_in(wire_d5_60),.data_out(wire_d5_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6562(.data_in(wire_d5_61),.data_out(wire_d5_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6563(.data_in(wire_d5_62),.data_out(wire_d5_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6564(.data_in(wire_d5_63),.data_out(wire_d5_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6565(.data_in(wire_d5_64),.data_out(wire_d5_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6566(.data_in(wire_d5_65),.data_out(wire_d5_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6567(.data_in(wire_d5_66),.data_out(wire_d5_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6568(.data_in(wire_d5_67),.data_out(wire_d5_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6569(.data_in(wire_d5_68),.data_out(wire_d5_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6570(.data_in(wire_d5_69),.data_out(wire_d5_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6571(.data_in(wire_d5_70),.data_out(wire_d5_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6572(.data_in(wire_d5_71),.data_out(wire_d5_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6573(.data_in(wire_d5_72),.data_out(wire_d5_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6574(.data_in(wire_d5_73),.data_out(wire_d5_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6575(.data_in(wire_d5_74),.data_out(wire_d5_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6576(.data_in(wire_d5_75),.data_out(wire_d5_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6577(.data_in(wire_d5_76),.data_out(wire_d5_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6578(.data_in(wire_d5_77),.data_out(wire_d5_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6579(.data_in(wire_d5_78),.data_out(wire_d5_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6580(.data_in(wire_d5_79),.data_out(wire_d5_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6581(.data_in(wire_d5_80),.data_out(wire_d5_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6582(.data_in(wire_d5_81),.data_out(wire_d5_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6583(.data_in(wire_d5_82),.data_out(wire_d5_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6584(.data_in(wire_d5_83),.data_out(wire_d5_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6585(.data_in(wire_d5_84),.data_out(wire_d5_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6586(.data_in(wire_d5_85),.data_out(wire_d5_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6587(.data_in(wire_d5_86),.data_out(wire_d5_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6588(.data_in(wire_d5_87),.data_out(wire_d5_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6589(.data_in(wire_d5_88),.data_out(wire_d5_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6590(.data_in(wire_d5_89),.data_out(wire_d5_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6591(.data_in(wire_d5_90),.data_out(wire_d5_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6592(.data_in(wire_d5_91),.data_out(wire_d5_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6593(.data_in(wire_d5_92),.data_out(wire_d5_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6594(.data_in(wire_d5_93),.data_out(wire_d5_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6595(.data_in(wire_d5_94),.data_out(wire_d5_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6596(.data_in(wire_d5_95),.data_out(wire_d5_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6597(.data_in(wire_d5_96),.data_out(wire_d5_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6598(.data_in(wire_d5_97),.data_out(wire_d5_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6599(.data_in(wire_d5_98),.data_out(d_out5),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance760(.data_in(d_in6),.data_out(wire_d6_0),.clk(clk),.rst(rst));            //channel 7
	register #(.WIDTH(WIDTH)) register_instance761(.data_in(wire_d6_0),.data_out(wire_d6_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance762(.data_in(wire_d6_1),.data_out(wire_d6_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance763(.data_in(wire_d6_2),.data_out(wire_d6_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance764(.data_in(wire_d6_3),.data_out(wire_d6_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance765(.data_in(wire_d6_4),.data_out(wire_d6_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance766(.data_in(wire_d6_5),.data_out(wire_d6_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767(.data_in(wire_d6_6),.data_out(wire_d6_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance768(.data_in(wire_d6_7),.data_out(wire_d6_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance769(.data_in(wire_d6_8),.data_out(wire_d6_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7610(.data_in(wire_d6_9),.data_out(wire_d6_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7611(.data_in(wire_d6_10),.data_out(wire_d6_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7612(.data_in(wire_d6_11),.data_out(wire_d6_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7613(.data_in(wire_d6_12),.data_out(wire_d6_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7614(.data_in(wire_d6_13),.data_out(wire_d6_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7615(.data_in(wire_d6_14),.data_out(wire_d6_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7616(.data_in(wire_d6_15),.data_out(wire_d6_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7617(.data_in(wire_d6_16),.data_out(wire_d6_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7618(.data_in(wire_d6_17),.data_out(wire_d6_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7619(.data_in(wire_d6_18),.data_out(wire_d6_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7620(.data_in(wire_d6_19),.data_out(wire_d6_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7621(.data_in(wire_d6_20),.data_out(wire_d6_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7622(.data_in(wire_d6_21),.data_out(wire_d6_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7623(.data_in(wire_d6_22),.data_out(wire_d6_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7624(.data_in(wire_d6_23),.data_out(wire_d6_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7625(.data_in(wire_d6_24),.data_out(wire_d6_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7626(.data_in(wire_d6_25),.data_out(wire_d6_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7627(.data_in(wire_d6_26),.data_out(wire_d6_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7628(.data_in(wire_d6_27),.data_out(wire_d6_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7629(.data_in(wire_d6_28),.data_out(wire_d6_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7630(.data_in(wire_d6_29),.data_out(wire_d6_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7631(.data_in(wire_d6_30),.data_out(wire_d6_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7632(.data_in(wire_d6_31),.data_out(wire_d6_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7633(.data_in(wire_d6_32),.data_out(wire_d6_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7634(.data_in(wire_d6_33),.data_out(wire_d6_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7635(.data_in(wire_d6_34),.data_out(wire_d6_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7636(.data_in(wire_d6_35),.data_out(wire_d6_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7637(.data_in(wire_d6_36),.data_out(wire_d6_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7638(.data_in(wire_d6_37),.data_out(wire_d6_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7639(.data_in(wire_d6_38),.data_out(wire_d6_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7640(.data_in(wire_d6_39),.data_out(wire_d6_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7641(.data_in(wire_d6_40),.data_out(wire_d6_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7642(.data_in(wire_d6_41),.data_out(wire_d6_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7643(.data_in(wire_d6_42),.data_out(wire_d6_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7644(.data_in(wire_d6_43),.data_out(wire_d6_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7645(.data_in(wire_d6_44),.data_out(wire_d6_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7646(.data_in(wire_d6_45),.data_out(wire_d6_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7647(.data_in(wire_d6_46),.data_out(wire_d6_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7648(.data_in(wire_d6_47),.data_out(wire_d6_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7649(.data_in(wire_d6_48),.data_out(wire_d6_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7650(.data_in(wire_d6_49),.data_out(wire_d6_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7651(.data_in(wire_d6_50),.data_out(wire_d6_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7652(.data_in(wire_d6_51),.data_out(wire_d6_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7653(.data_in(wire_d6_52),.data_out(wire_d6_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7654(.data_in(wire_d6_53),.data_out(wire_d6_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7655(.data_in(wire_d6_54),.data_out(wire_d6_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7656(.data_in(wire_d6_55),.data_out(wire_d6_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7657(.data_in(wire_d6_56),.data_out(wire_d6_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7658(.data_in(wire_d6_57),.data_out(wire_d6_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7659(.data_in(wire_d6_58),.data_out(wire_d6_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7660(.data_in(wire_d6_59),.data_out(wire_d6_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7661(.data_in(wire_d6_60),.data_out(wire_d6_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7662(.data_in(wire_d6_61),.data_out(wire_d6_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7663(.data_in(wire_d6_62),.data_out(wire_d6_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7664(.data_in(wire_d6_63),.data_out(wire_d6_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7665(.data_in(wire_d6_64),.data_out(wire_d6_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7666(.data_in(wire_d6_65),.data_out(wire_d6_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7667(.data_in(wire_d6_66),.data_out(wire_d6_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7668(.data_in(wire_d6_67),.data_out(wire_d6_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7669(.data_in(wire_d6_68),.data_out(wire_d6_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7670(.data_in(wire_d6_69),.data_out(wire_d6_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7671(.data_in(wire_d6_70),.data_out(wire_d6_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7672(.data_in(wire_d6_71),.data_out(wire_d6_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7673(.data_in(wire_d6_72),.data_out(wire_d6_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7674(.data_in(wire_d6_73),.data_out(wire_d6_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7675(.data_in(wire_d6_74),.data_out(wire_d6_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7676(.data_in(wire_d6_75),.data_out(wire_d6_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7677(.data_in(wire_d6_76),.data_out(wire_d6_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7678(.data_in(wire_d6_77),.data_out(wire_d6_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7679(.data_in(wire_d6_78),.data_out(wire_d6_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7680(.data_in(wire_d6_79),.data_out(wire_d6_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7681(.data_in(wire_d6_80),.data_out(wire_d6_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7682(.data_in(wire_d6_81),.data_out(wire_d6_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7683(.data_in(wire_d6_82),.data_out(wire_d6_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7684(.data_in(wire_d6_83),.data_out(wire_d6_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7685(.data_in(wire_d6_84),.data_out(wire_d6_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7686(.data_in(wire_d6_85),.data_out(wire_d6_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7687(.data_in(wire_d6_86),.data_out(wire_d6_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7688(.data_in(wire_d6_87),.data_out(wire_d6_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7689(.data_in(wire_d6_88),.data_out(wire_d6_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7690(.data_in(wire_d6_89),.data_out(wire_d6_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7691(.data_in(wire_d6_90),.data_out(wire_d6_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7692(.data_in(wire_d6_91),.data_out(wire_d6_92),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7693(.data_in(wire_d6_92),.data_out(wire_d6_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7694(.data_in(wire_d6_93),.data_out(wire_d6_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7695(.data_in(wire_d6_94),.data_out(wire_d6_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7696(.data_in(wire_d6_95),.data_out(wire_d6_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7697(.data_in(wire_d6_96),.data_out(wire_d6_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7698(.data_in(wire_d6_97),.data_out(wire_d6_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7699(.data_in(wire_d6_98),.data_out(d_out6),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance870(.data_in(d_in7),.data_out(wire_d7_0),.clk(clk),.rst(rst));            //channel 8
	encoder #(.WIDTH(WIDTH)) encoder_instance871(.data_in(wire_d7_0),.data_out(wire_d7_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance872(.data_in(wire_d7_1),.data_out(wire_d7_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance873(.data_in(wire_d7_2),.data_out(wire_d7_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance874(.data_in(wire_d7_3),.data_out(wire_d7_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance875(.data_in(wire_d7_4),.data_out(wire_d7_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance876(.data_in(wire_d7_5),.data_out(wire_d7_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance877(.data_in(wire_d7_6),.data_out(wire_d7_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878(.data_in(wire_d7_7),.data_out(wire_d7_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance879(.data_in(wire_d7_8),.data_out(wire_d7_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8710(.data_in(wire_d7_9),.data_out(wire_d7_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8711(.data_in(wire_d7_10),.data_out(wire_d7_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8712(.data_in(wire_d7_11),.data_out(wire_d7_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8713(.data_in(wire_d7_12),.data_out(wire_d7_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8714(.data_in(wire_d7_13),.data_out(wire_d7_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8715(.data_in(wire_d7_14),.data_out(wire_d7_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8716(.data_in(wire_d7_15),.data_out(wire_d7_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8717(.data_in(wire_d7_16),.data_out(wire_d7_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8718(.data_in(wire_d7_17),.data_out(wire_d7_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8719(.data_in(wire_d7_18),.data_out(wire_d7_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8720(.data_in(wire_d7_19),.data_out(wire_d7_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8721(.data_in(wire_d7_20),.data_out(wire_d7_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8722(.data_in(wire_d7_21),.data_out(wire_d7_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8723(.data_in(wire_d7_22),.data_out(wire_d7_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8724(.data_in(wire_d7_23),.data_out(wire_d7_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8725(.data_in(wire_d7_24),.data_out(wire_d7_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8726(.data_in(wire_d7_25),.data_out(wire_d7_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8727(.data_in(wire_d7_26),.data_out(wire_d7_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8728(.data_in(wire_d7_27),.data_out(wire_d7_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8729(.data_in(wire_d7_28),.data_out(wire_d7_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8730(.data_in(wire_d7_29),.data_out(wire_d7_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8731(.data_in(wire_d7_30),.data_out(wire_d7_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8732(.data_in(wire_d7_31),.data_out(wire_d7_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8733(.data_in(wire_d7_32),.data_out(wire_d7_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8734(.data_in(wire_d7_33),.data_out(wire_d7_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8735(.data_in(wire_d7_34),.data_out(wire_d7_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8736(.data_in(wire_d7_35),.data_out(wire_d7_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8737(.data_in(wire_d7_36),.data_out(wire_d7_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8738(.data_in(wire_d7_37),.data_out(wire_d7_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8739(.data_in(wire_d7_38),.data_out(wire_d7_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8740(.data_in(wire_d7_39),.data_out(wire_d7_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8741(.data_in(wire_d7_40),.data_out(wire_d7_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8742(.data_in(wire_d7_41),.data_out(wire_d7_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8743(.data_in(wire_d7_42),.data_out(wire_d7_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8744(.data_in(wire_d7_43),.data_out(wire_d7_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8745(.data_in(wire_d7_44),.data_out(wire_d7_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8746(.data_in(wire_d7_45),.data_out(wire_d7_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8747(.data_in(wire_d7_46),.data_out(wire_d7_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8748(.data_in(wire_d7_47),.data_out(wire_d7_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8749(.data_in(wire_d7_48),.data_out(wire_d7_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8750(.data_in(wire_d7_49),.data_out(wire_d7_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8751(.data_in(wire_d7_50),.data_out(wire_d7_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8752(.data_in(wire_d7_51),.data_out(wire_d7_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8753(.data_in(wire_d7_52),.data_out(wire_d7_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8754(.data_in(wire_d7_53),.data_out(wire_d7_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8755(.data_in(wire_d7_54),.data_out(wire_d7_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8756(.data_in(wire_d7_55),.data_out(wire_d7_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8757(.data_in(wire_d7_56),.data_out(wire_d7_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8758(.data_in(wire_d7_57),.data_out(wire_d7_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8759(.data_in(wire_d7_58),.data_out(wire_d7_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8760(.data_in(wire_d7_59),.data_out(wire_d7_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8761(.data_in(wire_d7_60),.data_out(wire_d7_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8762(.data_in(wire_d7_61),.data_out(wire_d7_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8763(.data_in(wire_d7_62),.data_out(wire_d7_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8764(.data_in(wire_d7_63),.data_out(wire_d7_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8765(.data_in(wire_d7_64),.data_out(wire_d7_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8766(.data_in(wire_d7_65),.data_out(wire_d7_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8767(.data_in(wire_d7_66),.data_out(wire_d7_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8768(.data_in(wire_d7_67),.data_out(wire_d7_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8769(.data_in(wire_d7_68),.data_out(wire_d7_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8770(.data_in(wire_d7_69),.data_out(wire_d7_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8771(.data_in(wire_d7_70),.data_out(wire_d7_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8772(.data_in(wire_d7_71),.data_out(wire_d7_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8773(.data_in(wire_d7_72),.data_out(wire_d7_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8774(.data_in(wire_d7_73),.data_out(wire_d7_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8775(.data_in(wire_d7_74),.data_out(wire_d7_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8776(.data_in(wire_d7_75),.data_out(wire_d7_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8777(.data_in(wire_d7_76),.data_out(wire_d7_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8778(.data_in(wire_d7_77),.data_out(wire_d7_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8779(.data_in(wire_d7_78),.data_out(wire_d7_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8780(.data_in(wire_d7_79),.data_out(wire_d7_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8781(.data_in(wire_d7_80),.data_out(wire_d7_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8782(.data_in(wire_d7_81),.data_out(wire_d7_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8783(.data_in(wire_d7_82),.data_out(wire_d7_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8784(.data_in(wire_d7_83),.data_out(wire_d7_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8785(.data_in(wire_d7_84),.data_out(wire_d7_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8786(.data_in(wire_d7_85),.data_out(wire_d7_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8787(.data_in(wire_d7_86),.data_out(wire_d7_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8788(.data_in(wire_d7_87),.data_out(wire_d7_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8789(.data_in(wire_d7_88),.data_out(wire_d7_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8790(.data_in(wire_d7_89),.data_out(wire_d7_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8791(.data_in(wire_d7_90),.data_out(wire_d7_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8792(.data_in(wire_d7_91),.data_out(wire_d7_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8793(.data_in(wire_d7_92),.data_out(wire_d7_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8794(.data_in(wire_d7_93),.data_out(wire_d7_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8795(.data_in(wire_d7_94),.data_out(wire_d7_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8796(.data_in(wire_d7_95),.data_out(wire_d7_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8797(.data_in(wire_d7_96),.data_out(wire_d7_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8798(.data_in(wire_d7_97),.data_out(wire_d7_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8799(.data_in(wire_d7_98),.data_out(d_out7),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance980(.data_in(d_in8),.data_out(wire_d8_0),.clk(clk),.rst(rst));            //channel 9
	invertion #(.WIDTH(WIDTH)) invertion_instance981(.data_in(wire_d8_0),.data_out(wire_d8_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance982(.data_in(wire_d8_1),.data_out(wire_d8_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance983(.data_in(wire_d8_2),.data_out(wire_d8_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance984(.data_in(wire_d8_3),.data_out(wire_d8_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance985(.data_in(wire_d8_4),.data_out(wire_d8_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance986(.data_in(wire_d8_5),.data_out(wire_d8_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance987(.data_in(wire_d8_6),.data_out(wire_d8_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance988(.data_in(wire_d8_7),.data_out(wire_d8_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance989(.data_in(wire_d8_8),.data_out(wire_d8_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9810(.data_in(wire_d8_9),.data_out(wire_d8_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9811(.data_in(wire_d8_10),.data_out(wire_d8_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9812(.data_in(wire_d8_11),.data_out(wire_d8_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9813(.data_in(wire_d8_12),.data_out(wire_d8_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9814(.data_in(wire_d8_13),.data_out(wire_d8_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9815(.data_in(wire_d8_14),.data_out(wire_d8_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9816(.data_in(wire_d8_15),.data_out(wire_d8_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9817(.data_in(wire_d8_16),.data_out(wire_d8_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9818(.data_in(wire_d8_17),.data_out(wire_d8_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9819(.data_in(wire_d8_18),.data_out(wire_d8_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9820(.data_in(wire_d8_19),.data_out(wire_d8_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9821(.data_in(wire_d8_20),.data_out(wire_d8_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9822(.data_in(wire_d8_21),.data_out(wire_d8_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9823(.data_in(wire_d8_22),.data_out(wire_d8_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9824(.data_in(wire_d8_23),.data_out(wire_d8_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9825(.data_in(wire_d8_24),.data_out(wire_d8_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9826(.data_in(wire_d8_25),.data_out(wire_d8_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9827(.data_in(wire_d8_26),.data_out(wire_d8_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9828(.data_in(wire_d8_27),.data_out(wire_d8_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9829(.data_in(wire_d8_28),.data_out(wire_d8_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9830(.data_in(wire_d8_29),.data_out(wire_d8_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9831(.data_in(wire_d8_30),.data_out(wire_d8_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9832(.data_in(wire_d8_31),.data_out(wire_d8_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9833(.data_in(wire_d8_32),.data_out(wire_d8_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9834(.data_in(wire_d8_33),.data_out(wire_d8_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9835(.data_in(wire_d8_34),.data_out(wire_d8_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9836(.data_in(wire_d8_35),.data_out(wire_d8_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9837(.data_in(wire_d8_36),.data_out(wire_d8_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9838(.data_in(wire_d8_37),.data_out(wire_d8_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9839(.data_in(wire_d8_38),.data_out(wire_d8_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9840(.data_in(wire_d8_39),.data_out(wire_d8_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9841(.data_in(wire_d8_40),.data_out(wire_d8_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9842(.data_in(wire_d8_41),.data_out(wire_d8_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9843(.data_in(wire_d8_42),.data_out(wire_d8_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9844(.data_in(wire_d8_43),.data_out(wire_d8_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9845(.data_in(wire_d8_44),.data_out(wire_d8_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9846(.data_in(wire_d8_45),.data_out(wire_d8_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9847(.data_in(wire_d8_46),.data_out(wire_d8_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9848(.data_in(wire_d8_47),.data_out(wire_d8_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9849(.data_in(wire_d8_48),.data_out(wire_d8_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9850(.data_in(wire_d8_49),.data_out(wire_d8_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9851(.data_in(wire_d8_50),.data_out(wire_d8_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9852(.data_in(wire_d8_51),.data_out(wire_d8_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9853(.data_in(wire_d8_52),.data_out(wire_d8_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9854(.data_in(wire_d8_53),.data_out(wire_d8_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9855(.data_in(wire_d8_54),.data_out(wire_d8_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9856(.data_in(wire_d8_55),.data_out(wire_d8_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9857(.data_in(wire_d8_56),.data_out(wire_d8_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9858(.data_in(wire_d8_57),.data_out(wire_d8_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9859(.data_in(wire_d8_58),.data_out(wire_d8_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9860(.data_in(wire_d8_59),.data_out(wire_d8_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9861(.data_in(wire_d8_60),.data_out(wire_d8_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9862(.data_in(wire_d8_61),.data_out(wire_d8_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9863(.data_in(wire_d8_62),.data_out(wire_d8_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9864(.data_in(wire_d8_63),.data_out(wire_d8_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9865(.data_in(wire_d8_64),.data_out(wire_d8_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9866(.data_in(wire_d8_65),.data_out(wire_d8_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9867(.data_in(wire_d8_66),.data_out(wire_d8_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9868(.data_in(wire_d8_67),.data_out(wire_d8_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9869(.data_in(wire_d8_68),.data_out(wire_d8_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9870(.data_in(wire_d8_69),.data_out(wire_d8_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9871(.data_in(wire_d8_70),.data_out(wire_d8_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9872(.data_in(wire_d8_71),.data_out(wire_d8_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9873(.data_in(wire_d8_72),.data_out(wire_d8_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9874(.data_in(wire_d8_73),.data_out(wire_d8_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9875(.data_in(wire_d8_74),.data_out(wire_d8_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9876(.data_in(wire_d8_75),.data_out(wire_d8_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9877(.data_in(wire_d8_76),.data_out(wire_d8_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9878(.data_in(wire_d8_77),.data_out(wire_d8_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9879(.data_in(wire_d8_78),.data_out(wire_d8_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9880(.data_in(wire_d8_79),.data_out(wire_d8_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9881(.data_in(wire_d8_80),.data_out(wire_d8_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9882(.data_in(wire_d8_81),.data_out(wire_d8_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9883(.data_in(wire_d8_82),.data_out(wire_d8_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9884(.data_in(wire_d8_83),.data_out(wire_d8_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9885(.data_in(wire_d8_84),.data_out(wire_d8_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9886(.data_in(wire_d8_85),.data_out(wire_d8_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9887(.data_in(wire_d8_86),.data_out(wire_d8_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9888(.data_in(wire_d8_87),.data_out(wire_d8_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9889(.data_in(wire_d8_88),.data_out(wire_d8_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9890(.data_in(wire_d8_89),.data_out(wire_d8_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9891(.data_in(wire_d8_90),.data_out(wire_d8_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9892(.data_in(wire_d8_91),.data_out(wire_d8_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9893(.data_in(wire_d8_92),.data_out(wire_d8_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9894(.data_in(wire_d8_93),.data_out(wire_d8_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9895(.data_in(wire_d8_94),.data_out(wire_d8_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9896(.data_in(wire_d8_95),.data_out(wire_d8_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9897(.data_in(wire_d8_96),.data_out(wire_d8_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9898(.data_in(wire_d8_97),.data_out(wire_d8_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9899(.data_in(wire_d8_98),.data_out(d_out8),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance1090(.data_in(d_in9),.data_out(wire_d9_0),.clk(clk),.rst(rst));            //channel 10
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1091(.data_in(wire_d9_0),.data_out(wire_d9_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1092(.data_in(wire_d9_1),.data_out(wire_d9_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1093(.data_in(wire_d9_2),.data_out(wire_d9_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1094(.data_in(wire_d9_3),.data_out(wire_d9_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1095(.data_in(wire_d9_4),.data_out(wire_d9_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1096(.data_in(wire_d9_5),.data_out(wire_d9_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1097(.data_in(wire_d9_6),.data_out(wire_d9_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1098(.data_in(wire_d9_7),.data_out(wire_d9_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1099(.data_in(wire_d9_8),.data_out(wire_d9_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10910(.data_in(wire_d9_9),.data_out(wire_d9_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10911(.data_in(wire_d9_10),.data_out(wire_d9_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10912(.data_in(wire_d9_11),.data_out(wire_d9_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10913(.data_in(wire_d9_12),.data_out(wire_d9_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10914(.data_in(wire_d9_13),.data_out(wire_d9_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10915(.data_in(wire_d9_14),.data_out(wire_d9_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10916(.data_in(wire_d9_15),.data_out(wire_d9_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10917(.data_in(wire_d9_16),.data_out(wire_d9_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10918(.data_in(wire_d9_17),.data_out(wire_d9_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10919(.data_in(wire_d9_18),.data_out(wire_d9_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10920(.data_in(wire_d9_19),.data_out(wire_d9_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10921(.data_in(wire_d9_20),.data_out(wire_d9_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10922(.data_in(wire_d9_21),.data_out(wire_d9_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10923(.data_in(wire_d9_22),.data_out(wire_d9_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10924(.data_in(wire_d9_23),.data_out(wire_d9_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10925(.data_in(wire_d9_24),.data_out(wire_d9_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10926(.data_in(wire_d9_25),.data_out(wire_d9_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10927(.data_in(wire_d9_26),.data_out(wire_d9_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10928(.data_in(wire_d9_27),.data_out(wire_d9_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10929(.data_in(wire_d9_28),.data_out(wire_d9_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10930(.data_in(wire_d9_29),.data_out(wire_d9_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10931(.data_in(wire_d9_30),.data_out(wire_d9_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10932(.data_in(wire_d9_31),.data_out(wire_d9_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10933(.data_in(wire_d9_32),.data_out(wire_d9_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10934(.data_in(wire_d9_33),.data_out(wire_d9_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10935(.data_in(wire_d9_34),.data_out(wire_d9_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10936(.data_in(wire_d9_35),.data_out(wire_d9_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10937(.data_in(wire_d9_36),.data_out(wire_d9_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10938(.data_in(wire_d9_37),.data_out(wire_d9_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10939(.data_in(wire_d9_38),.data_out(wire_d9_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10940(.data_in(wire_d9_39),.data_out(wire_d9_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10941(.data_in(wire_d9_40),.data_out(wire_d9_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10942(.data_in(wire_d9_41),.data_out(wire_d9_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10943(.data_in(wire_d9_42),.data_out(wire_d9_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10944(.data_in(wire_d9_43),.data_out(wire_d9_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10945(.data_in(wire_d9_44),.data_out(wire_d9_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10946(.data_in(wire_d9_45),.data_out(wire_d9_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10947(.data_in(wire_d9_46),.data_out(wire_d9_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10948(.data_in(wire_d9_47),.data_out(wire_d9_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10949(.data_in(wire_d9_48),.data_out(wire_d9_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10950(.data_in(wire_d9_49),.data_out(wire_d9_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10951(.data_in(wire_d9_50),.data_out(wire_d9_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10952(.data_in(wire_d9_51),.data_out(wire_d9_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10953(.data_in(wire_d9_52),.data_out(wire_d9_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10954(.data_in(wire_d9_53),.data_out(wire_d9_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10955(.data_in(wire_d9_54),.data_out(wire_d9_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10956(.data_in(wire_d9_55),.data_out(wire_d9_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10957(.data_in(wire_d9_56),.data_out(wire_d9_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10958(.data_in(wire_d9_57),.data_out(wire_d9_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10959(.data_in(wire_d9_58),.data_out(wire_d9_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10960(.data_in(wire_d9_59),.data_out(wire_d9_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10961(.data_in(wire_d9_60),.data_out(wire_d9_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10962(.data_in(wire_d9_61),.data_out(wire_d9_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10963(.data_in(wire_d9_62),.data_out(wire_d9_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10964(.data_in(wire_d9_63),.data_out(wire_d9_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10965(.data_in(wire_d9_64),.data_out(wire_d9_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10966(.data_in(wire_d9_65),.data_out(wire_d9_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10967(.data_in(wire_d9_66),.data_out(wire_d9_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10968(.data_in(wire_d9_67),.data_out(wire_d9_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10969(.data_in(wire_d9_68),.data_out(wire_d9_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10970(.data_in(wire_d9_69),.data_out(wire_d9_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10971(.data_in(wire_d9_70),.data_out(wire_d9_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10972(.data_in(wire_d9_71),.data_out(wire_d9_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10973(.data_in(wire_d9_72),.data_out(wire_d9_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10974(.data_in(wire_d9_73),.data_out(wire_d9_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10975(.data_in(wire_d9_74),.data_out(wire_d9_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10976(.data_in(wire_d9_75),.data_out(wire_d9_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10977(.data_in(wire_d9_76),.data_out(wire_d9_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10978(.data_in(wire_d9_77),.data_out(wire_d9_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10979(.data_in(wire_d9_78),.data_out(wire_d9_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10980(.data_in(wire_d9_79),.data_out(wire_d9_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10981(.data_in(wire_d9_80),.data_out(wire_d9_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10982(.data_in(wire_d9_81),.data_out(wire_d9_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10983(.data_in(wire_d9_82),.data_out(wire_d9_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10984(.data_in(wire_d9_83),.data_out(wire_d9_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10985(.data_in(wire_d9_84),.data_out(wire_d9_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10986(.data_in(wire_d9_85),.data_out(wire_d9_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10987(.data_in(wire_d9_86),.data_out(wire_d9_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10988(.data_in(wire_d9_87),.data_out(wire_d9_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10989(.data_in(wire_d9_88),.data_out(wire_d9_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10990(.data_in(wire_d9_89),.data_out(wire_d9_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10991(.data_in(wire_d9_90),.data_out(wire_d9_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10992(.data_in(wire_d9_91),.data_out(wire_d9_92),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10993(.data_in(wire_d9_92),.data_out(wire_d9_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10994(.data_in(wire_d9_93),.data_out(wire_d9_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10995(.data_in(wire_d9_94),.data_out(wire_d9_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10996(.data_in(wire_d9_95),.data_out(wire_d9_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10997(.data_in(wire_d9_96),.data_out(wire_d9_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10998(.data_in(wire_d9_97),.data_out(wire_d9_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10999(.data_in(wire_d9_98),.data_out(d_out9),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance11100(.data_in(d_in10),.data_out(wire_d10_0),.clk(clk),.rst(rst));            //channel 11
	encoder #(.WIDTH(WIDTH)) encoder_instance11101(.data_in(wire_d10_0),.data_out(wire_d10_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance11102(.data_in(wire_d10_1),.data_out(wire_d10_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance11103(.data_in(wire_d10_2),.data_out(wire_d10_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance11104(.data_in(wire_d10_3),.data_out(wire_d10_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance11105(.data_in(wire_d10_4),.data_out(wire_d10_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance11106(.data_in(wire_d10_5),.data_out(wire_d10_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance11107(.data_in(wire_d10_6),.data_out(wire_d10_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance11108(.data_in(wire_d10_7),.data_out(wire_d10_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance11109(.data_in(wire_d10_8),.data_out(wire_d10_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111010(.data_in(wire_d10_9),.data_out(wire_d10_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111011(.data_in(wire_d10_10),.data_out(wire_d10_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111012(.data_in(wire_d10_11),.data_out(wire_d10_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111013(.data_in(wire_d10_12),.data_out(wire_d10_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111014(.data_in(wire_d10_13),.data_out(wire_d10_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111015(.data_in(wire_d10_14),.data_out(wire_d10_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111016(.data_in(wire_d10_15),.data_out(wire_d10_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111017(.data_in(wire_d10_16),.data_out(wire_d10_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111018(.data_in(wire_d10_17),.data_out(wire_d10_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111019(.data_in(wire_d10_18),.data_out(wire_d10_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111020(.data_in(wire_d10_19),.data_out(wire_d10_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111021(.data_in(wire_d10_20),.data_out(wire_d10_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111022(.data_in(wire_d10_21),.data_out(wire_d10_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111023(.data_in(wire_d10_22),.data_out(wire_d10_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111024(.data_in(wire_d10_23),.data_out(wire_d10_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111025(.data_in(wire_d10_24),.data_out(wire_d10_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111026(.data_in(wire_d10_25),.data_out(wire_d10_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111027(.data_in(wire_d10_26),.data_out(wire_d10_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111028(.data_in(wire_d10_27),.data_out(wire_d10_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111029(.data_in(wire_d10_28),.data_out(wire_d10_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111030(.data_in(wire_d10_29),.data_out(wire_d10_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111031(.data_in(wire_d10_30),.data_out(wire_d10_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111032(.data_in(wire_d10_31),.data_out(wire_d10_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111033(.data_in(wire_d10_32),.data_out(wire_d10_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111034(.data_in(wire_d10_33),.data_out(wire_d10_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111035(.data_in(wire_d10_34),.data_out(wire_d10_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111036(.data_in(wire_d10_35),.data_out(wire_d10_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111037(.data_in(wire_d10_36),.data_out(wire_d10_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111038(.data_in(wire_d10_37),.data_out(wire_d10_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111039(.data_in(wire_d10_38),.data_out(wire_d10_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111040(.data_in(wire_d10_39),.data_out(wire_d10_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111041(.data_in(wire_d10_40),.data_out(wire_d10_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111042(.data_in(wire_d10_41),.data_out(wire_d10_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111043(.data_in(wire_d10_42),.data_out(wire_d10_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111044(.data_in(wire_d10_43),.data_out(wire_d10_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111045(.data_in(wire_d10_44),.data_out(wire_d10_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111046(.data_in(wire_d10_45),.data_out(wire_d10_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111047(.data_in(wire_d10_46),.data_out(wire_d10_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111048(.data_in(wire_d10_47),.data_out(wire_d10_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111049(.data_in(wire_d10_48),.data_out(wire_d10_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111050(.data_in(wire_d10_49),.data_out(wire_d10_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111051(.data_in(wire_d10_50),.data_out(wire_d10_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111052(.data_in(wire_d10_51),.data_out(wire_d10_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111053(.data_in(wire_d10_52),.data_out(wire_d10_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111054(.data_in(wire_d10_53),.data_out(wire_d10_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111055(.data_in(wire_d10_54),.data_out(wire_d10_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111056(.data_in(wire_d10_55),.data_out(wire_d10_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111057(.data_in(wire_d10_56),.data_out(wire_d10_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111058(.data_in(wire_d10_57),.data_out(wire_d10_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111059(.data_in(wire_d10_58),.data_out(wire_d10_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111060(.data_in(wire_d10_59),.data_out(wire_d10_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111061(.data_in(wire_d10_60),.data_out(wire_d10_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111062(.data_in(wire_d10_61),.data_out(wire_d10_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111063(.data_in(wire_d10_62),.data_out(wire_d10_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111064(.data_in(wire_d10_63),.data_out(wire_d10_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111065(.data_in(wire_d10_64),.data_out(wire_d10_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111066(.data_in(wire_d10_65),.data_out(wire_d10_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111067(.data_in(wire_d10_66),.data_out(wire_d10_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111068(.data_in(wire_d10_67),.data_out(wire_d10_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111069(.data_in(wire_d10_68),.data_out(wire_d10_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111070(.data_in(wire_d10_69),.data_out(wire_d10_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111071(.data_in(wire_d10_70),.data_out(wire_d10_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111072(.data_in(wire_d10_71),.data_out(wire_d10_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111073(.data_in(wire_d10_72),.data_out(wire_d10_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111074(.data_in(wire_d10_73),.data_out(wire_d10_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111075(.data_in(wire_d10_74),.data_out(wire_d10_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111076(.data_in(wire_d10_75),.data_out(wire_d10_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111077(.data_in(wire_d10_76),.data_out(wire_d10_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111078(.data_in(wire_d10_77),.data_out(wire_d10_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111079(.data_in(wire_d10_78),.data_out(wire_d10_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111080(.data_in(wire_d10_79),.data_out(wire_d10_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111081(.data_in(wire_d10_80),.data_out(wire_d10_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111082(.data_in(wire_d10_81),.data_out(wire_d10_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111083(.data_in(wire_d10_82),.data_out(wire_d10_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111084(.data_in(wire_d10_83),.data_out(wire_d10_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111085(.data_in(wire_d10_84),.data_out(wire_d10_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111086(.data_in(wire_d10_85),.data_out(wire_d10_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111087(.data_in(wire_d10_86),.data_out(wire_d10_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111088(.data_in(wire_d10_87),.data_out(wire_d10_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111089(.data_in(wire_d10_88),.data_out(wire_d10_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111090(.data_in(wire_d10_89),.data_out(wire_d10_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111091(.data_in(wire_d10_90),.data_out(wire_d10_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111092(.data_in(wire_d10_91),.data_out(wire_d10_92),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111093(.data_in(wire_d10_92),.data_out(wire_d10_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111094(.data_in(wire_d10_93),.data_out(wire_d10_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111095(.data_in(wire_d10_94),.data_out(wire_d10_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111096(.data_in(wire_d10_95),.data_out(wire_d10_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111097(.data_in(wire_d10_96),.data_out(wire_d10_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111098(.data_in(wire_d10_97),.data_out(wire_d10_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111099(.data_in(wire_d10_98),.data_out(d_out10),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance12110(.data_in(d_in11),.data_out(wire_d11_0),.clk(clk),.rst(rst));            //channel 12
	invertion #(.WIDTH(WIDTH)) invertion_instance12111(.data_in(wire_d11_0),.data_out(wire_d11_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance12112(.data_in(wire_d11_1),.data_out(wire_d11_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance12113(.data_in(wire_d11_2),.data_out(wire_d11_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance12114(.data_in(wire_d11_3),.data_out(wire_d11_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance12115(.data_in(wire_d11_4),.data_out(wire_d11_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance12116(.data_in(wire_d11_5),.data_out(wire_d11_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance12117(.data_in(wire_d11_6),.data_out(wire_d11_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance12118(.data_in(wire_d11_7),.data_out(wire_d11_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance12119(.data_in(wire_d11_8),.data_out(wire_d11_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121110(.data_in(wire_d11_9),.data_out(wire_d11_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121111(.data_in(wire_d11_10),.data_out(wire_d11_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121112(.data_in(wire_d11_11),.data_out(wire_d11_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121113(.data_in(wire_d11_12),.data_out(wire_d11_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121114(.data_in(wire_d11_13),.data_out(wire_d11_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121115(.data_in(wire_d11_14),.data_out(wire_d11_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121116(.data_in(wire_d11_15),.data_out(wire_d11_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121117(.data_in(wire_d11_16),.data_out(wire_d11_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121118(.data_in(wire_d11_17),.data_out(wire_d11_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121119(.data_in(wire_d11_18),.data_out(wire_d11_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121120(.data_in(wire_d11_19),.data_out(wire_d11_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121121(.data_in(wire_d11_20),.data_out(wire_d11_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121122(.data_in(wire_d11_21),.data_out(wire_d11_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121123(.data_in(wire_d11_22),.data_out(wire_d11_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121124(.data_in(wire_d11_23),.data_out(wire_d11_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121125(.data_in(wire_d11_24),.data_out(wire_d11_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121126(.data_in(wire_d11_25),.data_out(wire_d11_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121127(.data_in(wire_d11_26),.data_out(wire_d11_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121128(.data_in(wire_d11_27),.data_out(wire_d11_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121129(.data_in(wire_d11_28),.data_out(wire_d11_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121130(.data_in(wire_d11_29),.data_out(wire_d11_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121131(.data_in(wire_d11_30),.data_out(wire_d11_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121132(.data_in(wire_d11_31),.data_out(wire_d11_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121133(.data_in(wire_d11_32),.data_out(wire_d11_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121134(.data_in(wire_d11_33),.data_out(wire_d11_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121135(.data_in(wire_d11_34),.data_out(wire_d11_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121136(.data_in(wire_d11_35),.data_out(wire_d11_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121137(.data_in(wire_d11_36),.data_out(wire_d11_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121138(.data_in(wire_d11_37),.data_out(wire_d11_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121139(.data_in(wire_d11_38),.data_out(wire_d11_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121140(.data_in(wire_d11_39),.data_out(wire_d11_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121141(.data_in(wire_d11_40),.data_out(wire_d11_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121142(.data_in(wire_d11_41),.data_out(wire_d11_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121143(.data_in(wire_d11_42),.data_out(wire_d11_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121144(.data_in(wire_d11_43),.data_out(wire_d11_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121145(.data_in(wire_d11_44),.data_out(wire_d11_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121146(.data_in(wire_d11_45),.data_out(wire_d11_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121147(.data_in(wire_d11_46),.data_out(wire_d11_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121148(.data_in(wire_d11_47),.data_out(wire_d11_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121149(.data_in(wire_d11_48),.data_out(wire_d11_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121150(.data_in(wire_d11_49),.data_out(wire_d11_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121151(.data_in(wire_d11_50),.data_out(wire_d11_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121152(.data_in(wire_d11_51),.data_out(wire_d11_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121153(.data_in(wire_d11_52),.data_out(wire_d11_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121154(.data_in(wire_d11_53),.data_out(wire_d11_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121155(.data_in(wire_d11_54),.data_out(wire_d11_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121156(.data_in(wire_d11_55),.data_out(wire_d11_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121157(.data_in(wire_d11_56),.data_out(wire_d11_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121158(.data_in(wire_d11_57),.data_out(wire_d11_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121159(.data_in(wire_d11_58),.data_out(wire_d11_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121160(.data_in(wire_d11_59),.data_out(wire_d11_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121161(.data_in(wire_d11_60),.data_out(wire_d11_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121162(.data_in(wire_d11_61),.data_out(wire_d11_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121163(.data_in(wire_d11_62),.data_out(wire_d11_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121164(.data_in(wire_d11_63),.data_out(wire_d11_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121165(.data_in(wire_d11_64),.data_out(wire_d11_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121166(.data_in(wire_d11_65),.data_out(wire_d11_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121167(.data_in(wire_d11_66),.data_out(wire_d11_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121168(.data_in(wire_d11_67),.data_out(wire_d11_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121169(.data_in(wire_d11_68),.data_out(wire_d11_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121170(.data_in(wire_d11_69),.data_out(wire_d11_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121171(.data_in(wire_d11_70),.data_out(wire_d11_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121172(.data_in(wire_d11_71),.data_out(wire_d11_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121173(.data_in(wire_d11_72),.data_out(wire_d11_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121174(.data_in(wire_d11_73),.data_out(wire_d11_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121175(.data_in(wire_d11_74),.data_out(wire_d11_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121176(.data_in(wire_d11_75),.data_out(wire_d11_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121177(.data_in(wire_d11_76),.data_out(wire_d11_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121178(.data_in(wire_d11_77),.data_out(wire_d11_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121179(.data_in(wire_d11_78),.data_out(wire_d11_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121180(.data_in(wire_d11_79),.data_out(wire_d11_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121181(.data_in(wire_d11_80),.data_out(wire_d11_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121182(.data_in(wire_d11_81),.data_out(wire_d11_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121183(.data_in(wire_d11_82),.data_out(wire_d11_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121184(.data_in(wire_d11_83),.data_out(wire_d11_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121185(.data_in(wire_d11_84),.data_out(wire_d11_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121186(.data_in(wire_d11_85),.data_out(wire_d11_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121187(.data_in(wire_d11_86),.data_out(wire_d11_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121188(.data_in(wire_d11_87),.data_out(wire_d11_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121189(.data_in(wire_d11_88),.data_out(wire_d11_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121190(.data_in(wire_d11_89),.data_out(wire_d11_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121191(.data_in(wire_d11_90),.data_out(wire_d11_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121192(.data_in(wire_d11_91),.data_out(wire_d11_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121193(.data_in(wire_d11_92),.data_out(wire_d11_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121194(.data_in(wire_d11_93),.data_out(wire_d11_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121195(.data_in(wire_d11_94),.data_out(wire_d11_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121196(.data_in(wire_d11_95),.data_out(wire_d11_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121197(.data_in(wire_d11_96),.data_out(wire_d11_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121198(.data_in(wire_d11_97),.data_out(wire_d11_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121199(.data_in(wire_d11_98),.data_out(d_out11),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance13120(.data_in(d_in12),.data_out(wire_d12_0),.clk(clk),.rst(rst));            //channel 13
	encoder #(.WIDTH(WIDTH)) encoder_instance13121(.data_in(wire_d12_0),.data_out(wire_d12_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance13122(.data_in(wire_d12_1),.data_out(wire_d12_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance13123(.data_in(wire_d12_2),.data_out(wire_d12_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance13124(.data_in(wire_d12_3),.data_out(wire_d12_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance13125(.data_in(wire_d12_4),.data_out(wire_d12_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance13126(.data_in(wire_d12_5),.data_out(wire_d12_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance13127(.data_in(wire_d12_6),.data_out(wire_d12_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance13128(.data_in(wire_d12_7),.data_out(wire_d12_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance13129(.data_in(wire_d12_8),.data_out(wire_d12_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131210(.data_in(wire_d12_9),.data_out(wire_d12_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131211(.data_in(wire_d12_10),.data_out(wire_d12_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131212(.data_in(wire_d12_11),.data_out(wire_d12_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131213(.data_in(wire_d12_12),.data_out(wire_d12_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131214(.data_in(wire_d12_13),.data_out(wire_d12_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131215(.data_in(wire_d12_14),.data_out(wire_d12_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131216(.data_in(wire_d12_15),.data_out(wire_d12_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131217(.data_in(wire_d12_16),.data_out(wire_d12_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131218(.data_in(wire_d12_17),.data_out(wire_d12_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131219(.data_in(wire_d12_18),.data_out(wire_d12_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131220(.data_in(wire_d12_19),.data_out(wire_d12_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131221(.data_in(wire_d12_20),.data_out(wire_d12_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131222(.data_in(wire_d12_21),.data_out(wire_d12_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131223(.data_in(wire_d12_22),.data_out(wire_d12_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131224(.data_in(wire_d12_23),.data_out(wire_d12_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131225(.data_in(wire_d12_24),.data_out(wire_d12_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131226(.data_in(wire_d12_25),.data_out(wire_d12_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131227(.data_in(wire_d12_26),.data_out(wire_d12_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131228(.data_in(wire_d12_27),.data_out(wire_d12_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131229(.data_in(wire_d12_28),.data_out(wire_d12_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131230(.data_in(wire_d12_29),.data_out(wire_d12_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131231(.data_in(wire_d12_30),.data_out(wire_d12_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131232(.data_in(wire_d12_31),.data_out(wire_d12_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131233(.data_in(wire_d12_32),.data_out(wire_d12_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131234(.data_in(wire_d12_33),.data_out(wire_d12_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131235(.data_in(wire_d12_34),.data_out(wire_d12_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131236(.data_in(wire_d12_35),.data_out(wire_d12_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131237(.data_in(wire_d12_36),.data_out(wire_d12_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131238(.data_in(wire_d12_37),.data_out(wire_d12_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131239(.data_in(wire_d12_38),.data_out(wire_d12_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131240(.data_in(wire_d12_39),.data_out(wire_d12_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131241(.data_in(wire_d12_40),.data_out(wire_d12_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131242(.data_in(wire_d12_41),.data_out(wire_d12_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131243(.data_in(wire_d12_42),.data_out(wire_d12_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131244(.data_in(wire_d12_43),.data_out(wire_d12_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131245(.data_in(wire_d12_44),.data_out(wire_d12_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131246(.data_in(wire_d12_45),.data_out(wire_d12_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131247(.data_in(wire_d12_46),.data_out(wire_d12_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131248(.data_in(wire_d12_47),.data_out(wire_d12_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131249(.data_in(wire_d12_48),.data_out(wire_d12_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131250(.data_in(wire_d12_49),.data_out(wire_d12_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131251(.data_in(wire_d12_50),.data_out(wire_d12_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131252(.data_in(wire_d12_51),.data_out(wire_d12_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131253(.data_in(wire_d12_52),.data_out(wire_d12_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131254(.data_in(wire_d12_53),.data_out(wire_d12_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131255(.data_in(wire_d12_54),.data_out(wire_d12_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131256(.data_in(wire_d12_55),.data_out(wire_d12_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131257(.data_in(wire_d12_56),.data_out(wire_d12_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131258(.data_in(wire_d12_57),.data_out(wire_d12_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131259(.data_in(wire_d12_58),.data_out(wire_d12_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131260(.data_in(wire_d12_59),.data_out(wire_d12_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131261(.data_in(wire_d12_60),.data_out(wire_d12_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131262(.data_in(wire_d12_61),.data_out(wire_d12_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131263(.data_in(wire_d12_62),.data_out(wire_d12_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131264(.data_in(wire_d12_63),.data_out(wire_d12_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131265(.data_in(wire_d12_64),.data_out(wire_d12_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131266(.data_in(wire_d12_65),.data_out(wire_d12_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131267(.data_in(wire_d12_66),.data_out(wire_d12_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131268(.data_in(wire_d12_67),.data_out(wire_d12_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131269(.data_in(wire_d12_68),.data_out(wire_d12_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131270(.data_in(wire_d12_69),.data_out(wire_d12_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131271(.data_in(wire_d12_70),.data_out(wire_d12_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131272(.data_in(wire_d12_71),.data_out(wire_d12_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131273(.data_in(wire_d12_72),.data_out(wire_d12_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131274(.data_in(wire_d12_73),.data_out(wire_d12_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131275(.data_in(wire_d12_74),.data_out(wire_d12_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131276(.data_in(wire_d12_75),.data_out(wire_d12_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131277(.data_in(wire_d12_76),.data_out(wire_d12_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131278(.data_in(wire_d12_77),.data_out(wire_d12_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131279(.data_in(wire_d12_78),.data_out(wire_d12_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131280(.data_in(wire_d12_79),.data_out(wire_d12_80),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131281(.data_in(wire_d12_80),.data_out(wire_d12_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131282(.data_in(wire_d12_81),.data_out(wire_d12_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131283(.data_in(wire_d12_82),.data_out(wire_d12_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131284(.data_in(wire_d12_83),.data_out(wire_d12_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131285(.data_in(wire_d12_84),.data_out(wire_d12_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131286(.data_in(wire_d12_85),.data_out(wire_d12_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131287(.data_in(wire_d12_86),.data_out(wire_d12_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131288(.data_in(wire_d12_87),.data_out(wire_d12_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131289(.data_in(wire_d12_88),.data_out(wire_d12_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131290(.data_in(wire_d12_89),.data_out(wire_d12_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131291(.data_in(wire_d12_90),.data_out(wire_d12_91),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131292(.data_in(wire_d12_91),.data_out(wire_d12_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131293(.data_in(wire_d12_92),.data_out(wire_d12_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131294(.data_in(wire_d12_93),.data_out(wire_d12_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131295(.data_in(wire_d12_94),.data_out(wire_d12_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131296(.data_in(wire_d12_95),.data_out(wire_d12_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131297(.data_in(wire_d12_96),.data_out(wire_d12_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131298(.data_in(wire_d12_97),.data_out(wire_d12_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131299(.data_in(wire_d12_98),.data_out(d_out12),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance14130(.data_in(d_in13),.data_out(wire_d13_0),.clk(clk),.rst(rst));            //channel 14
	encoder #(.WIDTH(WIDTH)) encoder_instance14131(.data_in(wire_d13_0),.data_out(wire_d13_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance14132(.data_in(wire_d13_1),.data_out(wire_d13_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance14133(.data_in(wire_d13_2),.data_out(wire_d13_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance14134(.data_in(wire_d13_3),.data_out(wire_d13_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance14135(.data_in(wire_d13_4),.data_out(wire_d13_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance14136(.data_in(wire_d13_5),.data_out(wire_d13_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance14137(.data_in(wire_d13_6),.data_out(wire_d13_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance14138(.data_in(wire_d13_7),.data_out(wire_d13_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance14139(.data_in(wire_d13_8),.data_out(wire_d13_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141310(.data_in(wire_d13_9),.data_out(wire_d13_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141311(.data_in(wire_d13_10),.data_out(wire_d13_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141312(.data_in(wire_d13_11),.data_out(wire_d13_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141313(.data_in(wire_d13_12),.data_out(wire_d13_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141314(.data_in(wire_d13_13),.data_out(wire_d13_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141315(.data_in(wire_d13_14),.data_out(wire_d13_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141316(.data_in(wire_d13_15),.data_out(wire_d13_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141317(.data_in(wire_d13_16),.data_out(wire_d13_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141318(.data_in(wire_d13_17),.data_out(wire_d13_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141319(.data_in(wire_d13_18),.data_out(wire_d13_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141320(.data_in(wire_d13_19),.data_out(wire_d13_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141321(.data_in(wire_d13_20),.data_out(wire_d13_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141322(.data_in(wire_d13_21),.data_out(wire_d13_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141323(.data_in(wire_d13_22),.data_out(wire_d13_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141324(.data_in(wire_d13_23),.data_out(wire_d13_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141325(.data_in(wire_d13_24),.data_out(wire_d13_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141326(.data_in(wire_d13_25),.data_out(wire_d13_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141327(.data_in(wire_d13_26),.data_out(wire_d13_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141328(.data_in(wire_d13_27),.data_out(wire_d13_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141329(.data_in(wire_d13_28),.data_out(wire_d13_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141330(.data_in(wire_d13_29),.data_out(wire_d13_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141331(.data_in(wire_d13_30),.data_out(wire_d13_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141332(.data_in(wire_d13_31),.data_out(wire_d13_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141333(.data_in(wire_d13_32),.data_out(wire_d13_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141334(.data_in(wire_d13_33),.data_out(wire_d13_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141335(.data_in(wire_d13_34),.data_out(wire_d13_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141336(.data_in(wire_d13_35),.data_out(wire_d13_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141337(.data_in(wire_d13_36),.data_out(wire_d13_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141338(.data_in(wire_d13_37),.data_out(wire_d13_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141339(.data_in(wire_d13_38),.data_out(wire_d13_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141340(.data_in(wire_d13_39),.data_out(wire_d13_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141341(.data_in(wire_d13_40),.data_out(wire_d13_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141342(.data_in(wire_d13_41),.data_out(wire_d13_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141343(.data_in(wire_d13_42),.data_out(wire_d13_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141344(.data_in(wire_d13_43),.data_out(wire_d13_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141345(.data_in(wire_d13_44),.data_out(wire_d13_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141346(.data_in(wire_d13_45),.data_out(wire_d13_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141347(.data_in(wire_d13_46),.data_out(wire_d13_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141348(.data_in(wire_d13_47),.data_out(wire_d13_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141349(.data_in(wire_d13_48),.data_out(wire_d13_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141350(.data_in(wire_d13_49),.data_out(wire_d13_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141351(.data_in(wire_d13_50),.data_out(wire_d13_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141352(.data_in(wire_d13_51),.data_out(wire_d13_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141353(.data_in(wire_d13_52),.data_out(wire_d13_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141354(.data_in(wire_d13_53),.data_out(wire_d13_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141355(.data_in(wire_d13_54),.data_out(wire_d13_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141356(.data_in(wire_d13_55),.data_out(wire_d13_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141357(.data_in(wire_d13_56),.data_out(wire_d13_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141358(.data_in(wire_d13_57),.data_out(wire_d13_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141359(.data_in(wire_d13_58),.data_out(wire_d13_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141360(.data_in(wire_d13_59),.data_out(wire_d13_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141361(.data_in(wire_d13_60),.data_out(wire_d13_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141362(.data_in(wire_d13_61),.data_out(wire_d13_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141363(.data_in(wire_d13_62),.data_out(wire_d13_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141364(.data_in(wire_d13_63),.data_out(wire_d13_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141365(.data_in(wire_d13_64),.data_out(wire_d13_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141366(.data_in(wire_d13_65),.data_out(wire_d13_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141367(.data_in(wire_d13_66),.data_out(wire_d13_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141368(.data_in(wire_d13_67),.data_out(wire_d13_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141369(.data_in(wire_d13_68),.data_out(wire_d13_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141370(.data_in(wire_d13_69),.data_out(wire_d13_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141371(.data_in(wire_d13_70),.data_out(wire_d13_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141372(.data_in(wire_d13_71),.data_out(wire_d13_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141373(.data_in(wire_d13_72),.data_out(wire_d13_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141374(.data_in(wire_d13_73),.data_out(wire_d13_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141375(.data_in(wire_d13_74),.data_out(wire_d13_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141376(.data_in(wire_d13_75),.data_out(wire_d13_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141377(.data_in(wire_d13_76),.data_out(wire_d13_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141378(.data_in(wire_d13_77),.data_out(wire_d13_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141379(.data_in(wire_d13_78),.data_out(wire_d13_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141380(.data_in(wire_d13_79),.data_out(wire_d13_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141381(.data_in(wire_d13_80),.data_out(wire_d13_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141382(.data_in(wire_d13_81),.data_out(wire_d13_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141383(.data_in(wire_d13_82),.data_out(wire_d13_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141384(.data_in(wire_d13_83),.data_out(wire_d13_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141385(.data_in(wire_d13_84),.data_out(wire_d13_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141386(.data_in(wire_d13_85),.data_out(wire_d13_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141387(.data_in(wire_d13_86),.data_out(wire_d13_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141388(.data_in(wire_d13_87),.data_out(wire_d13_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141389(.data_in(wire_d13_88),.data_out(wire_d13_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141390(.data_in(wire_d13_89),.data_out(wire_d13_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141391(.data_in(wire_d13_90),.data_out(wire_d13_91),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141392(.data_in(wire_d13_91),.data_out(wire_d13_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141393(.data_in(wire_d13_92),.data_out(wire_d13_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141394(.data_in(wire_d13_93),.data_out(wire_d13_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141395(.data_in(wire_d13_94),.data_out(wire_d13_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141396(.data_in(wire_d13_95),.data_out(wire_d13_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141397(.data_in(wire_d13_96),.data_out(wire_d13_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141398(.data_in(wire_d13_97),.data_out(wire_d13_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141399(.data_in(wire_d13_98),.data_out(d_out13),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance15140(.data_in(d_in14),.data_out(wire_d14_0),.clk(clk),.rst(rst));            //channel 15
	encoder #(.WIDTH(WIDTH)) encoder_instance15141(.data_in(wire_d14_0),.data_out(wire_d14_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance15142(.data_in(wire_d14_1),.data_out(wire_d14_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance15143(.data_in(wire_d14_2),.data_out(wire_d14_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance15144(.data_in(wire_d14_3),.data_out(wire_d14_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance15145(.data_in(wire_d14_4),.data_out(wire_d14_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance15146(.data_in(wire_d14_5),.data_out(wire_d14_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance15147(.data_in(wire_d14_6),.data_out(wire_d14_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance15148(.data_in(wire_d14_7),.data_out(wire_d14_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance15149(.data_in(wire_d14_8),.data_out(wire_d14_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151410(.data_in(wire_d14_9),.data_out(wire_d14_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151411(.data_in(wire_d14_10),.data_out(wire_d14_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151412(.data_in(wire_d14_11),.data_out(wire_d14_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151413(.data_in(wire_d14_12),.data_out(wire_d14_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151414(.data_in(wire_d14_13),.data_out(wire_d14_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151415(.data_in(wire_d14_14),.data_out(wire_d14_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151416(.data_in(wire_d14_15),.data_out(wire_d14_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151417(.data_in(wire_d14_16),.data_out(wire_d14_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151418(.data_in(wire_d14_17),.data_out(wire_d14_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151419(.data_in(wire_d14_18),.data_out(wire_d14_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151420(.data_in(wire_d14_19),.data_out(wire_d14_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151421(.data_in(wire_d14_20),.data_out(wire_d14_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151422(.data_in(wire_d14_21),.data_out(wire_d14_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151423(.data_in(wire_d14_22),.data_out(wire_d14_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151424(.data_in(wire_d14_23),.data_out(wire_d14_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151425(.data_in(wire_d14_24),.data_out(wire_d14_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151426(.data_in(wire_d14_25),.data_out(wire_d14_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151427(.data_in(wire_d14_26),.data_out(wire_d14_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151428(.data_in(wire_d14_27),.data_out(wire_d14_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151429(.data_in(wire_d14_28),.data_out(wire_d14_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151430(.data_in(wire_d14_29),.data_out(wire_d14_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151431(.data_in(wire_d14_30),.data_out(wire_d14_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151432(.data_in(wire_d14_31),.data_out(wire_d14_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151433(.data_in(wire_d14_32),.data_out(wire_d14_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151434(.data_in(wire_d14_33),.data_out(wire_d14_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151435(.data_in(wire_d14_34),.data_out(wire_d14_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151436(.data_in(wire_d14_35),.data_out(wire_d14_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151437(.data_in(wire_d14_36),.data_out(wire_d14_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151438(.data_in(wire_d14_37),.data_out(wire_d14_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151439(.data_in(wire_d14_38),.data_out(wire_d14_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151440(.data_in(wire_d14_39),.data_out(wire_d14_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151441(.data_in(wire_d14_40),.data_out(wire_d14_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151442(.data_in(wire_d14_41),.data_out(wire_d14_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151443(.data_in(wire_d14_42),.data_out(wire_d14_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151444(.data_in(wire_d14_43),.data_out(wire_d14_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151445(.data_in(wire_d14_44),.data_out(wire_d14_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151446(.data_in(wire_d14_45),.data_out(wire_d14_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151447(.data_in(wire_d14_46),.data_out(wire_d14_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151448(.data_in(wire_d14_47),.data_out(wire_d14_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151449(.data_in(wire_d14_48),.data_out(wire_d14_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151450(.data_in(wire_d14_49),.data_out(wire_d14_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151451(.data_in(wire_d14_50),.data_out(wire_d14_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151452(.data_in(wire_d14_51),.data_out(wire_d14_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151453(.data_in(wire_d14_52),.data_out(wire_d14_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151454(.data_in(wire_d14_53),.data_out(wire_d14_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151455(.data_in(wire_d14_54),.data_out(wire_d14_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151456(.data_in(wire_d14_55),.data_out(wire_d14_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151457(.data_in(wire_d14_56),.data_out(wire_d14_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151458(.data_in(wire_d14_57),.data_out(wire_d14_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151459(.data_in(wire_d14_58),.data_out(wire_d14_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151460(.data_in(wire_d14_59),.data_out(wire_d14_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151461(.data_in(wire_d14_60),.data_out(wire_d14_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151462(.data_in(wire_d14_61),.data_out(wire_d14_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151463(.data_in(wire_d14_62),.data_out(wire_d14_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151464(.data_in(wire_d14_63),.data_out(wire_d14_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151465(.data_in(wire_d14_64),.data_out(wire_d14_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151466(.data_in(wire_d14_65),.data_out(wire_d14_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151467(.data_in(wire_d14_66),.data_out(wire_d14_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151468(.data_in(wire_d14_67),.data_out(wire_d14_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151469(.data_in(wire_d14_68),.data_out(wire_d14_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151470(.data_in(wire_d14_69),.data_out(wire_d14_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151471(.data_in(wire_d14_70),.data_out(wire_d14_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151472(.data_in(wire_d14_71),.data_out(wire_d14_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151473(.data_in(wire_d14_72),.data_out(wire_d14_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151474(.data_in(wire_d14_73),.data_out(wire_d14_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151475(.data_in(wire_d14_74),.data_out(wire_d14_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151476(.data_in(wire_d14_75),.data_out(wire_d14_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151477(.data_in(wire_d14_76),.data_out(wire_d14_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151478(.data_in(wire_d14_77),.data_out(wire_d14_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151479(.data_in(wire_d14_78),.data_out(wire_d14_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151480(.data_in(wire_d14_79),.data_out(wire_d14_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151481(.data_in(wire_d14_80),.data_out(wire_d14_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151482(.data_in(wire_d14_81),.data_out(wire_d14_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151483(.data_in(wire_d14_82),.data_out(wire_d14_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151484(.data_in(wire_d14_83),.data_out(wire_d14_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151485(.data_in(wire_d14_84),.data_out(wire_d14_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151486(.data_in(wire_d14_85),.data_out(wire_d14_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151487(.data_in(wire_d14_86),.data_out(wire_d14_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151488(.data_in(wire_d14_87),.data_out(wire_d14_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151489(.data_in(wire_d14_88),.data_out(wire_d14_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151490(.data_in(wire_d14_89),.data_out(wire_d14_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151491(.data_in(wire_d14_90),.data_out(wire_d14_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151492(.data_in(wire_d14_91),.data_out(wire_d14_92),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151493(.data_in(wire_d14_92),.data_out(wire_d14_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151494(.data_in(wire_d14_93),.data_out(wire_d14_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151495(.data_in(wire_d14_94),.data_out(wire_d14_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151496(.data_in(wire_d14_95),.data_out(wire_d14_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151497(.data_in(wire_d14_96),.data_out(wire_d14_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151498(.data_in(wire_d14_97),.data_out(wire_d14_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151499(.data_in(wire_d14_98),.data_out(d_out14),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance16150(.data_in(d_in15),.data_out(wire_d15_0),.clk(clk),.rst(rst));            //channel 16
	register #(.WIDTH(WIDTH)) register_instance16151(.data_in(wire_d15_0),.data_out(wire_d15_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance16152(.data_in(wire_d15_1),.data_out(wire_d15_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance16153(.data_in(wire_d15_2),.data_out(wire_d15_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance16154(.data_in(wire_d15_3),.data_out(wire_d15_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance16155(.data_in(wire_d15_4),.data_out(wire_d15_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance16156(.data_in(wire_d15_5),.data_out(wire_d15_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance16157(.data_in(wire_d15_6),.data_out(wire_d15_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance16158(.data_in(wire_d15_7),.data_out(wire_d15_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance16159(.data_in(wire_d15_8),.data_out(wire_d15_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161510(.data_in(wire_d15_9),.data_out(wire_d15_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161511(.data_in(wire_d15_10),.data_out(wire_d15_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161512(.data_in(wire_d15_11),.data_out(wire_d15_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161513(.data_in(wire_d15_12),.data_out(wire_d15_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161514(.data_in(wire_d15_13),.data_out(wire_d15_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161515(.data_in(wire_d15_14),.data_out(wire_d15_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161516(.data_in(wire_d15_15),.data_out(wire_d15_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161517(.data_in(wire_d15_16),.data_out(wire_d15_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161518(.data_in(wire_d15_17),.data_out(wire_d15_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161519(.data_in(wire_d15_18),.data_out(wire_d15_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161520(.data_in(wire_d15_19),.data_out(wire_d15_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161521(.data_in(wire_d15_20),.data_out(wire_d15_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161522(.data_in(wire_d15_21),.data_out(wire_d15_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161523(.data_in(wire_d15_22),.data_out(wire_d15_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161524(.data_in(wire_d15_23),.data_out(wire_d15_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161525(.data_in(wire_d15_24),.data_out(wire_d15_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161526(.data_in(wire_d15_25),.data_out(wire_d15_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161527(.data_in(wire_d15_26),.data_out(wire_d15_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161528(.data_in(wire_d15_27),.data_out(wire_d15_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161529(.data_in(wire_d15_28),.data_out(wire_d15_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161530(.data_in(wire_d15_29),.data_out(wire_d15_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161531(.data_in(wire_d15_30),.data_out(wire_d15_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161532(.data_in(wire_d15_31),.data_out(wire_d15_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161533(.data_in(wire_d15_32),.data_out(wire_d15_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161534(.data_in(wire_d15_33),.data_out(wire_d15_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161535(.data_in(wire_d15_34),.data_out(wire_d15_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161536(.data_in(wire_d15_35),.data_out(wire_d15_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161537(.data_in(wire_d15_36),.data_out(wire_d15_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161538(.data_in(wire_d15_37),.data_out(wire_d15_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161539(.data_in(wire_d15_38),.data_out(wire_d15_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161540(.data_in(wire_d15_39),.data_out(wire_d15_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161541(.data_in(wire_d15_40),.data_out(wire_d15_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161542(.data_in(wire_d15_41),.data_out(wire_d15_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161543(.data_in(wire_d15_42),.data_out(wire_d15_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161544(.data_in(wire_d15_43),.data_out(wire_d15_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161545(.data_in(wire_d15_44),.data_out(wire_d15_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161546(.data_in(wire_d15_45),.data_out(wire_d15_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161547(.data_in(wire_d15_46),.data_out(wire_d15_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161548(.data_in(wire_d15_47),.data_out(wire_d15_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161549(.data_in(wire_d15_48),.data_out(wire_d15_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161550(.data_in(wire_d15_49),.data_out(wire_d15_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161551(.data_in(wire_d15_50),.data_out(wire_d15_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161552(.data_in(wire_d15_51),.data_out(wire_d15_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161553(.data_in(wire_d15_52),.data_out(wire_d15_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161554(.data_in(wire_d15_53),.data_out(wire_d15_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161555(.data_in(wire_d15_54),.data_out(wire_d15_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161556(.data_in(wire_d15_55),.data_out(wire_d15_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161557(.data_in(wire_d15_56),.data_out(wire_d15_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161558(.data_in(wire_d15_57),.data_out(wire_d15_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161559(.data_in(wire_d15_58),.data_out(wire_d15_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161560(.data_in(wire_d15_59),.data_out(wire_d15_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161561(.data_in(wire_d15_60),.data_out(wire_d15_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161562(.data_in(wire_d15_61),.data_out(wire_d15_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161563(.data_in(wire_d15_62),.data_out(wire_d15_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161564(.data_in(wire_d15_63),.data_out(wire_d15_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161565(.data_in(wire_d15_64),.data_out(wire_d15_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161566(.data_in(wire_d15_65),.data_out(wire_d15_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161567(.data_in(wire_d15_66),.data_out(wire_d15_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161568(.data_in(wire_d15_67),.data_out(wire_d15_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161569(.data_in(wire_d15_68),.data_out(wire_d15_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161570(.data_in(wire_d15_69),.data_out(wire_d15_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161571(.data_in(wire_d15_70),.data_out(wire_d15_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161572(.data_in(wire_d15_71),.data_out(wire_d15_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161573(.data_in(wire_d15_72),.data_out(wire_d15_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161574(.data_in(wire_d15_73),.data_out(wire_d15_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161575(.data_in(wire_d15_74),.data_out(wire_d15_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161576(.data_in(wire_d15_75),.data_out(wire_d15_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161577(.data_in(wire_d15_76),.data_out(wire_d15_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161578(.data_in(wire_d15_77),.data_out(wire_d15_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161579(.data_in(wire_d15_78),.data_out(wire_d15_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161580(.data_in(wire_d15_79),.data_out(wire_d15_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161581(.data_in(wire_d15_80),.data_out(wire_d15_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161582(.data_in(wire_d15_81),.data_out(wire_d15_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161583(.data_in(wire_d15_82),.data_out(wire_d15_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161584(.data_in(wire_d15_83),.data_out(wire_d15_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161585(.data_in(wire_d15_84),.data_out(wire_d15_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161586(.data_in(wire_d15_85),.data_out(wire_d15_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161587(.data_in(wire_d15_86),.data_out(wire_d15_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161588(.data_in(wire_d15_87),.data_out(wire_d15_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161589(.data_in(wire_d15_88),.data_out(wire_d15_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161590(.data_in(wire_d15_89),.data_out(wire_d15_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161591(.data_in(wire_d15_90),.data_out(wire_d15_91),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161592(.data_in(wire_d15_91),.data_out(wire_d15_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161593(.data_in(wire_d15_92),.data_out(wire_d15_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161594(.data_in(wire_d15_93),.data_out(wire_d15_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161595(.data_in(wire_d15_94),.data_out(wire_d15_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161596(.data_in(wire_d15_95),.data_out(wire_d15_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161597(.data_in(wire_d15_96),.data_out(wire_d15_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161598(.data_in(wire_d15_97),.data_out(wire_d15_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161599(.data_in(wire_d15_98),.data_out(d_out15),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance17160(.data_in(d_in16),.data_out(wire_d16_0),.clk(clk),.rst(rst));            //channel 17
	encoder #(.WIDTH(WIDTH)) encoder_instance17161(.data_in(wire_d16_0),.data_out(wire_d16_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance17162(.data_in(wire_d16_1),.data_out(wire_d16_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance17163(.data_in(wire_d16_2),.data_out(wire_d16_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance17164(.data_in(wire_d16_3),.data_out(wire_d16_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance17165(.data_in(wire_d16_4),.data_out(wire_d16_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance17166(.data_in(wire_d16_5),.data_out(wire_d16_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance17167(.data_in(wire_d16_6),.data_out(wire_d16_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance17168(.data_in(wire_d16_7),.data_out(wire_d16_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance17169(.data_in(wire_d16_8),.data_out(wire_d16_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171610(.data_in(wire_d16_9),.data_out(wire_d16_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171611(.data_in(wire_d16_10),.data_out(wire_d16_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171612(.data_in(wire_d16_11),.data_out(wire_d16_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171613(.data_in(wire_d16_12),.data_out(wire_d16_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171614(.data_in(wire_d16_13),.data_out(wire_d16_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171615(.data_in(wire_d16_14),.data_out(wire_d16_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171616(.data_in(wire_d16_15),.data_out(wire_d16_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171617(.data_in(wire_d16_16),.data_out(wire_d16_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171618(.data_in(wire_d16_17),.data_out(wire_d16_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171619(.data_in(wire_d16_18),.data_out(wire_d16_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171620(.data_in(wire_d16_19),.data_out(wire_d16_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171621(.data_in(wire_d16_20),.data_out(wire_d16_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171622(.data_in(wire_d16_21),.data_out(wire_d16_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171623(.data_in(wire_d16_22),.data_out(wire_d16_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171624(.data_in(wire_d16_23),.data_out(wire_d16_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171625(.data_in(wire_d16_24),.data_out(wire_d16_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171626(.data_in(wire_d16_25),.data_out(wire_d16_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171627(.data_in(wire_d16_26),.data_out(wire_d16_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171628(.data_in(wire_d16_27),.data_out(wire_d16_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171629(.data_in(wire_d16_28),.data_out(wire_d16_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171630(.data_in(wire_d16_29),.data_out(wire_d16_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171631(.data_in(wire_d16_30),.data_out(wire_d16_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171632(.data_in(wire_d16_31),.data_out(wire_d16_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171633(.data_in(wire_d16_32),.data_out(wire_d16_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171634(.data_in(wire_d16_33),.data_out(wire_d16_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171635(.data_in(wire_d16_34),.data_out(wire_d16_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171636(.data_in(wire_d16_35),.data_out(wire_d16_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171637(.data_in(wire_d16_36),.data_out(wire_d16_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171638(.data_in(wire_d16_37),.data_out(wire_d16_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171639(.data_in(wire_d16_38),.data_out(wire_d16_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171640(.data_in(wire_d16_39),.data_out(wire_d16_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171641(.data_in(wire_d16_40),.data_out(wire_d16_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171642(.data_in(wire_d16_41),.data_out(wire_d16_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171643(.data_in(wire_d16_42),.data_out(wire_d16_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171644(.data_in(wire_d16_43),.data_out(wire_d16_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171645(.data_in(wire_d16_44),.data_out(wire_d16_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171646(.data_in(wire_d16_45),.data_out(wire_d16_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171647(.data_in(wire_d16_46),.data_out(wire_d16_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171648(.data_in(wire_d16_47),.data_out(wire_d16_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171649(.data_in(wire_d16_48),.data_out(wire_d16_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171650(.data_in(wire_d16_49),.data_out(wire_d16_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171651(.data_in(wire_d16_50),.data_out(wire_d16_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171652(.data_in(wire_d16_51),.data_out(wire_d16_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171653(.data_in(wire_d16_52),.data_out(wire_d16_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171654(.data_in(wire_d16_53),.data_out(wire_d16_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171655(.data_in(wire_d16_54),.data_out(wire_d16_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171656(.data_in(wire_d16_55),.data_out(wire_d16_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171657(.data_in(wire_d16_56),.data_out(wire_d16_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171658(.data_in(wire_d16_57),.data_out(wire_d16_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171659(.data_in(wire_d16_58),.data_out(wire_d16_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171660(.data_in(wire_d16_59),.data_out(wire_d16_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171661(.data_in(wire_d16_60),.data_out(wire_d16_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171662(.data_in(wire_d16_61),.data_out(wire_d16_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171663(.data_in(wire_d16_62),.data_out(wire_d16_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171664(.data_in(wire_d16_63),.data_out(wire_d16_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171665(.data_in(wire_d16_64),.data_out(wire_d16_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171666(.data_in(wire_d16_65),.data_out(wire_d16_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171667(.data_in(wire_d16_66),.data_out(wire_d16_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171668(.data_in(wire_d16_67),.data_out(wire_d16_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171669(.data_in(wire_d16_68),.data_out(wire_d16_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171670(.data_in(wire_d16_69),.data_out(wire_d16_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171671(.data_in(wire_d16_70),.data_out(wire_d16_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171672(.data_in(wire_d16_71),.data_out(wire_d16_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171673(.data_in(wire_d16_72),.data_out(wire_d16_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171674(.data_in(wire_d16_73),.data_out(wire_d16_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171675(.data_in(wire_d16_74),.data_out(wire_d16_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171676(.data_in(wire_d16_75),.data_out(wire_d16_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171677(.data_in(wire_d16_76),.data_out(wire_d16_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171678(.data_in(wire_d16_77),.data_out(wire_d16_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171679(.data_in(wire_d16_78),.data_out(wire_d16_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171680(.data_in(wire_d16_79),.data_out(wire_d16_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171681(.data_in(wire_d16_80),.data_out(wire_d16_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171682(.data_in(wire_d16_81),.data_out(wire_d16_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171683(.data_in(wire_d16_82),.data_out(wire_d16_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171684(.data_in(wire_d16_83),.data_out(wire_d16_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171685(.data_in(wire_d16_84),.data_out(wire_d16_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171686(.data_in(wire_d16_85),.data_out(wire_d16_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171687(.data_in(wire_d16_86),.data_out(wire_d16_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171688(.data_in(wire_d16_87),.data_out(wire_d16_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171689(.data_in(wire_d16_88),.data_out(wire_d16_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171690(.data_in(wire_d16_89),.data_out(wire_d16_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171691(.data_in(wire_d16_90),.data_out(wire_d16_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171692(.data_in(wire_d16_91),.data_out(wire_d16_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171693(.data_in(wire_d16_92),.data_out(wire_d16_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171694(.data_in(wire_d16_93),.data_out(wire_d16_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171695(.data_in(wire_d16_94),.data_out(wire_d16_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171696(.data_in(wire_d16_95),.data_out(wire_d16_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171697(.data_in(wire_d16_96),.data_out(wire_d16_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171698(.data_in(wire_d16_97),.data_out(wire_d16_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171699(.data_in(wire_d16_98),.data_out(d_out16),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance18170(.data_in(d_in17),.data_out(wire_d17_0),.clk(clk),.rst(rst));            //channel 18
	large_mux #(.WIDTH(WIDTH)) large_mux_instance18171(.data_in(wire_d17_0),.data_out(wire_d17_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance18172(.data_in(wire_d17_1),.data_out(wire_d17_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance18173(.data_in(wire_d17_2),.data_out(wire_d17_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance18174(.data_in(wire_d17_3),.data_out(wire_d17_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance18175(.data_in(wire_d17_4),.data_out(wire_d17_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance18176(.data_in(wire_d17_5),.data_out(wire_d17_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance18177(.data_in(wire_d17_6),.data_out(wire_d17_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance18178(.data_in(wire_d17_7),.data_out(wire_d17_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance18179(.data_in(wire_d17_8),.data_out(wire_d17_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181710(.data_in(wire_d17_9),.data_out(wire_d17_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181711(.data_in(wire_d17_10),.data_out(wire_d17_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181712(.data_in(wire_d17_11),.data_out(wire_d17_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181713(.data_in(wire_d17_12),.data_out(wire_d17_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181714(.data_in(wire_d17_13),.data_out(wire_d17_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181715(.data_in(wire_d17_14),.data_out(wire_d17_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181716(.data_in(wire_d17_15),.data_out(wire_d17_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181717(.data_in(wire_d17_16),.data_out(wire_d17_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181718(.data_in(wire_d17_17),.data_out(wire_d17_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181719(.data_in(wire_d17_18),.data_out(wire_d17_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181720(.data_in(wire_d17_19),.data_out(wire_d17_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181721(.data_in(wire_d17_20),.data_out(wire_d17_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181722(.data_in(wire_d17_21),.data_out(wire_d17_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181723(.data_in(wire_d17_22),.data_out(wire_d17_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181724(.data_in(wire_d17_23),.data_out(wire_d17_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181725(.data_in(wire_d17_24),.data_out(wire_d17_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181726(.data_in(wire_d17_25),.data_out(wire_d17_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181727(.data_in(wire_d17_26),.data_out(wire_d17_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181728(.data_in(wire_d17_27),.data_out(wire_d17_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181729(.data_in(wire_d17_28),.data_out(wire_d17_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181730(.data_in(wire_d17_29),.data_out(wire_d17_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181731(.data_in(wire_d17_30),.data_out(wire_d17_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181732(.data_in(wire_d17_31),.data_out(wire_d17_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181733(.data_in(wire_d17_32),.data_out(wire_d17_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181734(.data_in(wire_d17_33),.data_out(wire_d17_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181735(.data_in(wire_d17_34),.data_out(wire_d17_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181736(.data_in(wire_d17_35),.data_out(wire_d17_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181737(.data_in(wire_d17_36),.data_out(wire_d17_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181738(.data_in(wire_d17_37),.data_out(wire_d17_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181739(.data_in(wire_d17_38),.data_out(wire_d17_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181740(.data_in(wire_d17_39),.data_out(wire_d17_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181741(.data_in(wire_d17_40),.data_out(wire_d17_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181742(.data_in(wire_d17_41),.data_out(wire_d17_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181743(.data_in(wire_d17_42),.data_out(wire_d17_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181744(.data_in(wire_d17_43),.data_out(wire_d17_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181745(.data_in(wire_d17_44),.data_out(wire_d17_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181746(.data_in(wire_d17_45),.data_out(wire_d17_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181747(.data_in(wire_d17_46),.data_out(wire_d17_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181748(.data_in(wire_d17_47),.data_out(wire_d17_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181749(.data_in(wire_d17_48),.data_out(wire_d17_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181750(.data_in(wire_d17_49),.data_out(wire_d17_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181751(.data_in(wire_d17_50),.data_out(wire_d17_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181752(.data_in(wire_d17_51),.data_out(wire_d17_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181753(.data_in(wire_d17_52),.data_out(wire_d17_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181754(.data_in(wire_d17_53),.data_out(wire_d17_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181755(.data_in(wire_d17_54),.data_out(wire_d17_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181756(.data_in(wire_d17_55),.data_out(wire_d17_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181757(.data_in(wire_d17_56),.data_out(wire_d17_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181758(.data_in(wire_d17_57),.data_out(wire_d17_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181759(.data_in(wire_d17_58),.data_out(wire_d17_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181760(.data_in(wire_d17_59),.data_out(wire_d17_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181761(.data_in(wire_d17_60),.data_out(wire_d17_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181762(.data_in(wire_d17_61),.data_out(wire_d17_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181763(.data_in(wire_d17_62),.data_out(wire_d17_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181764(.data_in(wire_d17_63),.data_out(wire_d17_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181765(.data_in(wire_d17_64),.data_out(wire_d17_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181766(.data_in(wire_d17_65),.data_out(wire_d17_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181767(.data_in(wire_d17_66),.data_out(wire_d17_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181768(.data_in(wire_d17_67),.data_out(wire_d17_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181769(.data_in(wire_d17_68),.data_out(wire_d17_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181770(.data_in(wire_d17_69),.data_out(wire_d17_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181771(.data_in(wire_d17_70),.data_out(wire_d17_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181772(.data_in(wire_d17_71),.data_out(wire_d17_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181773(.data_in(wire_d17_72),.data_out(wire_d17_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181774(.data_in(wire_d17_73),.data_out(wire_d17_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181775(.data_in(wire_d17_74),.data_out(wire_d17_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181776(.data_in(wire_d17_75),.data_out(wire_d17_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181777(.data_in(wire_d17_76),.data_out(wire_d17_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181778(.data_in(wire_d17_77),.data_out(wire_d17_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181779(.data_in(wire_d17_78),.data_out(wire_d17_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181780(.data_in(wire_d17_79),.data_out(wire_d17_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181781(.data_in(wire_d17_80),.data_out(wire_d17_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181782(.data_in(wire_d17_81),.data_out(wire_d17_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181783(.data_in(wire_d17_82),.data_out(wire_d17_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181784(.data_in(wire_d17_83),.data_out(wire_d17_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181785(.data_in(wire_d17_84),.data_out(wire_d17_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181786(.data_in(wire_d17_85),.data_out(wire_d17_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181787(.data_in(wire_d17_86),.data_out(wire_d17_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181788(.data_in(wire_d17_87),.data_out(wire_d17_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181789(.data_in(wire_d17_88),.data_out(wire_d17_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181790(.data_in(wire_d17_89),.data_out(wire_d17_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181791(.data_in(wire_d17_90),.data_out(wire_d17_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181792(.data_in(wire_d17_91),.data_out(wire_d17_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181793(.data_in(wire_d17_92),.data_out(wire_d17_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181794(.data_in(wire_d17_93),.data_out(wire_d17_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181795(.data_in(wire_d17_94),.data_out(wire_d17_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181796(.data_in(wire_d17_95),.data_out(wire_d17_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181797(.data_in(wire_d17_96),.data_out(wire_d17_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181798(.data_in(wire_d17_97),.data_out(wire_d17_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181799(.data_in(wire_d17_98),.data_out(d_out17),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance19180(.data_in(d_in18),.data_out(wire_d18_0),.clk(clk),.rst(rst));            //channel 19
	encoder #(.WIDTH(WIDTH)) encoder_instance19181(.data_in(wire_d18_0),.data_out(wire_d18_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance19182(.data_in(wire_d18_1),.data_out(wire_d18_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance19183(.data_in(wire_d18_2),.data_out(wire_d18_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance19184(.data_in(wire_d18_3),.data_out(wire_d18_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance19185(.data_in(wire_d18_4),.data_out(wire_d18_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance19186(.data_in(wire_d18_5),.data_out(wire_d18_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance19187(.data_in(wire_d18_6),.data_out(wire_d18_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance19188(.data_in(wire_d18_7),.data_out(wire_d18_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance19189(.data_in(wire_d18_8),.data_out(wire_d18_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191810(.data_in(wire_d18_9),.data_out(wire_d18_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191811(.data_in(wire_d18_10),.data_out(wire_d18_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191812(.data_in(wire_d18_11),.data_out(wire_d18_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191813(.data_in(wire_d18_12),.data_out(wire_d18_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191814(.data_in(wire_d18_13),.data_out(wire_d18_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191815(.data_in(wire_d18_14),.data_out(wire_d18_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191816(.data_in(wire_d18_15),.data_out(wire_d18_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191817(.data_in(wire_d18_16),.data_out(wire_d18_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191818(.data_in(wire_d18_17),.data_out(wire_d18_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191819(.data_in(wire_d18_18),.data_out(wire_d18_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191820(.data_in(wire_d18_19),.data_out(wire_d18_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191821(.data_in(wire_d18_20),.data_out(wire_d18_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191822(.data_in(wire_d18_21),.data_out(wire_d18_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191823(.data_in(wire_d18_22),.data_out(wire_d18_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191824(.data_in(wire_d18_23),.data_out(wire_d18_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191825(.data_in(wire_d18_24),.data_out(wire_d18_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191826(.data_in(wire_d18_25),.data_out(wire_d18_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191827(.data_in(wire_d18_26),.data_out(wire_d18_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191828(.data_in(wire_d18_27),.data_out(wire_d18_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191829(.data_in(wire_d18_28),.data_out(wire_d18_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191830(.data_in(wire_d18_29),.data_out(wire_d18_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191831(.data_in(wire_d18_30),.data_out(wire_d18_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191832(.data_in(wire_d18_31),.data_out(wire_d18_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191833(.data_in(wire_d18_32),.data_out(wire_d18_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191834(.data_in(wire_d18_33),.data_out(wire_d18_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191835(.data_in(wire_d18_34),.data_out(wire_d18_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191836(.data_in(wire_d18_35),.data_out(wire_d18_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191837(.data_in(wire_d18_36),.data_out(wire_d18_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191838(.data_in(wire_d18_37),.data_out(wire_d18_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191839(.data_in(wire_d18_38),.data_out(wire_d18_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191840(.data_in(wire_d18_39),.data_out(wire_d18_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191841(.data_in(wire_d18_40),.data_out(wire_d18_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191842(.data_in(wire_d18_41),.data_out(wire_d18_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191843(.data_in(wire_d18_42),.data_out(wire_d18_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191844(.data_in(wire_d18_43),.data_out(wire_d18_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191845(.data_in(wire_d18_44),.data_out(wire_d18_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191846(.data_in(wire_d18_45),.data_out(wire_d18_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191847(.data_in(wire_d18_46),.data_out(wire_d18_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191848(.data_in(wire_d18_47),.data_out(wire_d18_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191849(.data_in(wire_d18_48),.data_out(wire_d18_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191850(.data_in(wire_d18_49),.data_out(wire_d18_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191851(.data_in(wire_d18_50),.data_out(wire_d18_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191852(.data_in(wire_d18_51),.data_out(wire_d18_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191853(.data_in(wire_d18_52),.data_out(wire_d18_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191854(.data_in(wire_d18_53),.data_out(wire_d18_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191855(.data_in(wire_d18_54),.data_out(wire_d18_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191856(.data_in(wire_d18_55),.data_out(wire_d18_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191857(.data_in(wire_d18_56),.data_out(wire_d18_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191858(.data_in(wire_d18_57),.data_out(wire_d18_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191859(.data_in(wire_d18_58),.data_out(wire_d18_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191860(.data_in(wire_d18_59),.data_out(wire_d18_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191861(.data_in(wire_d18_60),.data_out(wire_d18_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191862(.data_in(wire_d18_61),.data_out(wire_d18_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191863(.data_in(wire_d18_62),.data_out(wire_d18_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191864(.data_in(wire_d18_63),.data_out(wire_d18_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191865(.data_in(wire_d18_64),.data_out(wire_d18_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191866(.data_in(wire_d18_65),.data_out(wire_d18_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191867(.data_in(wire_d18_66),.data_out(wire_d18_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191868(.data_in(wire_d18_67),.data_out(wire_d18_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191869(.data_in(wire_d18_68),.data_out(wire_d18_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191870(.data_in(wire_d18_69),.data_out(wire_d18_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191871(.data_in(wire_d18_70),.data_out(wire_d18_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191872(.data_in(wire_d18_71),.data_out(wire_d18_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191873(.data_in(wire_d18_72),.data_out(wire_d18_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191874(.data_in(wire_d18_73),.data_out(wire_d18_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191875(.data_in(wire_d18_74),.data_out(wire_d18_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191876(.data_in(wire_d18_75),.data_out(wire_d18_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191877(.data_in(wire_d18_76),.data_out(wire_d18_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191878(.data_in(wire_d18_77),.data_out(wire_d18_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191879(.data_in(wire_d18_78),.data_out(wire_d18_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191880(.data_in(wire_d18_79),.data_out(wire_d18_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191881(.data_in(wire_d18_80),.data_out(wire_d18_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191882(.data_in(wire_d18_81),.data_out(wire_d18_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191883(.data_in(wire_d18_82),.data_out(wire_d18_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191884(.data_in(wire_d18_83),.data_out(wire_d18_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191885(.data_in(wire_d18_84),.data_out(wire_d18_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191886(.data_in(wire_d18_85),.data_out(wire_d18_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191887(.data_in(wire_d18_86),.data_out(wire_d18_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191888(.data_in(wire_d18_87),.data_out(wire_d18_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191889(.data_in(wire_d18_88),.data_out(wire_d18_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191890(.data_in(wire_d18_89),.data_out(wire_d18_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191891(.data_in(wire_d18_90),.data_out(wire_d18_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191892(.data_in(wire_d18_91),.data_out(wire_d18_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191893(.data_in(wire_d18_92),.data_out(wire_d18_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191894(.data_in(wire_d18_93),.data_out(wire_d18_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191895(.data_in(wire_d18_94),.data_out(wire_d18_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191896(.data_in(wire_d18_95),.data_out(wire_d18_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191897(.data_in(wire_d18_96),.data_out(wire_d18_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191898(.data_in(wire_d18_97),.data_out(wire_d18_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191899(.data_in(wire_d18_98),.data_out(d_out18),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance20190(.data_in(d_in19),.data_out(wire_d19_0),.clk(clk),.rst(rst));            //channel 20
	encoder #(.WIDTH(WIDTH)) encoder_instance20191(.data_in(wire_d19_0),.data_out(wire_d19_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance20192(.data_in(wire_d19_1),.data_out(wire_d19_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance20193(.data_in(wire_d19_2),.data_out(wire_d19_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance20194(.data_in(wire_d19_3),.data_out(wire_d19_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance20195(.data_in(wire_d19_4),.data_out(wire_d19_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance20196(.data_in(wire_d19_5),.data_out(wire_d19_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance20197(.data_in(wire_d19_6),.data_out(wire_d19_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance20198(.data_in(wire_d19_7),.data_out(wire_d19_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance20199(.data_in(wire_d19_8),.data_out(wire_d19_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201910(.data_in(wire_d19_9),.data_out(wire_d19_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201911(.data_in(wire_d19_10),.data_out(wire_d19_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201912(.data_in(wire_d19_11),.data_out(wire_d19_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201913(.data_in(wire_d19_12),.data_out(wire_d19_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201914(.data_in(wire_d19_13),.data_out(wire_d19_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201915(.data_in(wire_d19_14),.data_out(wire_d19_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201916(.data_in(wire_d19_15),.data_out(wire_d19_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201917(.data_in(wire_d19_16),.data_out(wire_d19_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201918(.data_in(wire_d19_17),.data_out(wire_d19_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201919(.data_in(wire_d19_18),.data_out(wire_d19_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201920(.data_in(wire_d19_19),.data_out(wire_d19_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201921(.data_in(wire_d19_20),.data_out(wire_d19_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201922(.data_in(wire_d19_21),.data_out(wire_d19_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201923(.data_in(wire_d19_22),.data_out(wire_d19_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201924(.data_in(wire_d19_23),.data_out(wire_d19_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201925(.data_in(wire_d19_24),.data_out(wire_d19_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201926(.data_in(wire_d19_25),.data_out(wire_d19_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201927(.data_in(wire_d19_26),.data_out(wire_d19_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201928(.data_in(wire_d19_27),.data_out(wire_d19_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201929(.data_in(wire_d19_28),.data_out(wire_d19_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201930(.data_in(wire_d19_29),.data_out(wire_d19_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201931(.data_in(wire_d19_30),.data_out(wire_d19_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201932(.data_in(wire_d19_31),.data_out(wire_d19_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201933(.data_in(wire_d19_32),.data_out(wire_d19_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201934(.data_in(wire_d19_33),.data_out(wire_d19_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201935(.data_in(wire_d19_34),.data_out(wire_d19_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201936(.data_in(wire_d19_35),.data_out(wire_d19_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201937(.data_in(wire_d19_36),.data_out(wire_d19_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201938(.data_in(wire_d19_37),.data_out(wire_d19_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201939(.data_in(wire_d19_38),.data_out(wire_d19_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201940(.data_in(wire_d19_39),.data_out(wire_d19_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201941(.data_in(wire_d19_40),.data_out(wire_d19_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201942(.data_in(wire_d19_41),.data_out(wire_d19_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201943(.data_in(wire_d19_42),.data_out(wire_d19_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201944(.data_in(wire_d19_43),.data_out(wire_d19_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201945(.data_in(wire_d19_44),.data_out(wire_d19_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201946(.data_in(wire_d19_45),.data_out(wire_d19_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201947(.data_in(wire_d19_46),.data_out(wire_d19_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201948(.data_in(wire_d19_47),.data_out(wire_d19_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201949(.data_in(wire_d19_48),.data_out(wire_d19_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201950(.data_in(wire_d19_49),.data_out(wire_d19_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201951(.data_in(wire_d19_50),.data_out(wire_d19_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201952(.data_in(wire_d19_51),.data_out(wire_d19_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201953(.data_in(wire_d19_52),.data_out(wire_d19_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201954(.data_in(wire_d19_53),.data_out(wire_d19_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201955(.data_in(wire_d19_54),.data_out(wire_d19_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201956(.data_in(wire_d19_55),.data_out(wire_d19_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201957(.data_in(wire_d19_56),.data_out(wire_d19_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201958(.data_in(wire_d19_57),.data_out(wire_d19_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201959(.data_in(wire_d19_58),.data_out(wire_d19_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201960(.data_in(wire_d19_59),.data_out(wire_d19_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201961(.data_in(wire_d19_60),.data_out(wire_d19_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201962(.data_in(wire_d19_61),.data_out(wire_d19_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201963(.data_in(wire_d19_62),.data_out(wire_d19_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201964(.data_in(wire_d19_63),.data_out(wire_d19_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201965(.data_in(wire_d19_64),.data_out(wire_d19_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201966(.data_in(wire_d19_65),.data_out(wire_d19_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201967(.data_in(wire_d19_66),.data_out(wire_d19_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201968(.data_in(wire_d19_67),.data_out(wire_d19_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201969(.data_in(wire_d19_68),.data_out(wire_d19_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201970(.data_in(wire_d19_69),.data_out(wire_d19_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201971(.data_in(wire_d19_70),.data_out(wire_d19_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201972(.data_in(wire_d19_71),.data_out(wire_d19_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201973(.data_in(wire_d19_72),.data_out(wire_d19_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201974(.data_in(wire_d19_73),.data_out(wire_d19_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201975(.data_in(wire_d19_74),.data_out(wire_d19_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201976(.data_in(wire_d19_75),.data_out(wire_d19_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201977(.data_in(wire_d19_76),.data_out(wire_d19_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201978(.data_in(wire_d19_77),.data_out(wire_d19_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201979(.data_in(wire_d19_78),.data_out(wire_d19_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201980(.data_in(wire_d19_79),.data_out(wire_d19_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201981(.data_in(wire_d19_80),.data_out(wire_d19_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201982(.data_in(wire_d19_81),.data_out(wire_d19_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201983(.data_in(wire_d19_82),.data_out(wire_d19_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201984(.data_in(wire_d19_83),.data_out(wire_d19_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201985(.data_in(wire_d19_84),.data_out(wire_d19_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201986(.data_in(wire_d19_85),.data_out(wire_d19_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201987(.data_in(wire_d19_86),.data_out(wire_d19_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201988(.data_in(wire_d19_87),.data_out(wire_d19_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201989(.data_in(wire_d19_88),.data_out(wire_d19_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201990(.data_in(wire_d19_89),.data_out(wire_d19_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201991(.data_in(wire_d19_90),.data_out(wire_d19_91),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201992(.data_in(wire_d19_91),.data_out(wire_d19_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201993(.data_in(wire_d19_92),.data_out(wire_d19_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201994(.data_in(wire_d19_93),.data_out(wire_d19_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201995(.data_in(wire_d19_94),.data_out(wire_d19_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201996(.data_in(wire_d19_95),.data_out(wire_d19_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201997(.data_in(wire_d19_96),.data_out(wire_d19_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201998(.data_in(wire_d19_97),.data_out(wire_d19_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201999(.data_in(wire_d19_98),.data_out(d_out19),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance21200(.data_in(d_in20),.data_out(wire_d20_0),.clk(clk),.rst(rst));            //channel 21
	large_mux #(.WIDTH(WIDTH)) large_mux_instance21201(.data_in(wire_d20_0),.data_out(wire_d20_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance21202(.data_in(wire_d20_1),.data_out(wire_d20_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance21203(.data_in(wire_d20_2),.data_out(wire_d20_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21204(.data_in(wire_d20_3),.data_out(wire_d20_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance21205(.data_in(wire_d20_4),.data_out(wire_d20_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance21206(.data_in(wire_d20_5),.data_out(wire_d20_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance21207(.data_in(wire_d20_6),.data_out(wire_d20_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance21208(.data_in(wire_d20_7),.data_out(wire_d20_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance21209(.data_in(wire_d20_8),.data_out(wire_d20_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212010(.data_in(wire_d20_9),.data_out(wire_d20_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212011(.data_in(wire_d20_10),.data_out(wire_d20_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212012(.data_in(wire_d20_11),.data_out(wire_d20_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212013(.data_in(wire_d20_12),.data_out(wire_d20_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212014(.data_in(wire_d20_13),.data_out(wire_d20_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212015(.data_in(wire_d20_14),.data_out(wire_d20_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212016(.data_in(wire_d20_15),.data_out(wire_d20_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212017(.data_in(wire_d20_16),.data_out(wire_d20_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212018(.data_in(wire_d20_17),.data_out(wire_d20_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212019(.data_in(wire_d20_18),.data_out(wire_d20_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212020(.data_in(wire_d20_19),.data_out(wire_d20_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212021(.data_in(wire_d20_20),.data_out(wire_d20_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212022(.data_in(wire_d20_21),.data_out(wire_d20_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212023(.data_in(wire_d20_22),.data_out(wire_d20_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212024(.data_in(wire_d20_23),.data_out(wire_d20_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212025(.data_in(wire_d20_24),.data_out(wire_d20_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212026(.data_in(wire_d20_25),.data_out(wire_d20_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212027(.data_in(wire_d20_26),.data_out(wire_d20_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212028(.data_in(wire_d20_27),.data_out(wire_d20_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212029(.data_in(wire_d20_28),.data_out(wire_d20_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212030(.data_in(wire_d20_29),.data_out(wire_d20_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212031(.data_in(wire_d20_30),.data_out(wire_d20_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212032(.data_in(wire_d20_31),.data_out(wire_d20_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212033(.data_in(wire_d20_32),.data_out(wire_d20_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212034(.data_in(wire_d20_33),.data_out(wire_d20_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212035(.data_in(wire_d20_34),.data_out(wire_d20_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212036(.data_in(wire_d20_35),.data_out(wire_d20_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212037(.data_in(wire_d20_36),.data_out(wire_d20_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212038(.data_in(wire_d20_37),.data_out(wire_d20_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212039(.data_in(wire_d20_38),.data_out(wire_d20_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212040(.data_in(wire_d20_39),.data_out(wire_d20_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212041(.data_in(wire_d20_40),.data_out(wire_d20_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212042(.data_in(wire_d20_41),.data_out(wire_d20_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212043(.data_in(wire_d20_42),.data_out(wire_d20_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212044(.data_in(wire_d20_43),.data_out(wire_d20_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212045(.data_in(wire_d20_44),.data_out(wire_d20_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212046(.data_in(wire_d20_45),.data_out(wire_d20_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212047(.data_in(wire_d20_46),.data_out(wire_d20_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212048(.data_in(wire_d20_47),.data_out(wire_d20_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212049(.data_in(wire_d20_48),.data_out(wire_d20_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212050(.data_in(wire_d20_49),.data_out(wire_d20_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212051(.data_in(wire_d20_50),.data_out(wire_d20_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212052(.data_in(wire_d20_51),.data_out(wire_d20_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212053(.data_in(wire_d20_52),.data_out(wire_d20_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212054(.data_in(wire_d20_53),.data_out(wire_d20_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212055(.data_in(wire_d20_54),.data_out(wire_d20_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212056(.data_in(wire_d20_55),.data_out(wire_d20_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212057(.data_in(wire_d20_56),.data_out(wire_d20_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212058(.data_in(wire_d20_57),.data_out(wire_d20_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212059(.data_in(wire_d20_58),.data_out(wire_d20_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212060(.data_in(wire_d20_59),.data_out(wire_d20_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212061(.data_in(wire_d20_60),.data_out(wire_d20_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212062(.data_in(wire_d20_61),.data_out(wire_d20_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212063(.data_in(wire_d20_62),.data_out(wire_d20_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212064(.data_in(wire_d20_63),.data_out(wire_d20_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212065(.data_in(wire_d20_64),.data_out(wire_d20_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212066(.data_in(wire_d20_65),.data_out(wire_d20_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212067(.data_in(wire_d20_66),.data_out(wire_d20_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212068(.data_in(wire_d20_67),.data_out(wire_d20_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212069(.data_in(wire_d20_68),.data_out(wire_d20_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212070(.data_in(wire_d20_69),.data_out(wire_d20_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212071(.data_in(wire_d20_70),.data_out(wire_d20_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212072(.data_in(wire_d20_71),.data_out(wire_d20_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212073(.data_in(wire_d20_72),.data_out(wire_d20_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212074(.data_in(wire_d20_73),.data_out(wire_d20_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212075(.data_in(wire_d20_74),.data_out(wire_d20_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212076(.data_in(wire_d20_75),.data_out(wire_d20_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212077(.data_in(wire_d20_76),.data_out(wire_d20_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212078(.data_in(wire_d20_77),.data_out(wire_d20_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212079(.data_in(wire_d20_78),.data_out(wire_d20_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212080(.data_in(wire_d20_79),.data_out(wire_d20_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212081(.data_in(wire_d20_80),.data_out(wire_d20_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212082(.data_in(wire_d20_81),.data_out(wire_d20_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212083(.data_in(wire_d20_82),.data_out(wire_d20_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212084(.data_in(wire_d20_83),.data_out(wire_d20_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212085(.data_in(wire_d20_84),.data_out(wire_d20_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212086(.data_in(wire_d20_85),.data_out(wire_d20_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212087(.data_in(wire_d20_86),.data_out(wire_d20_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212088(.data_in(wire_d20_87),.data_out(wire_d20_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212089(.data_in(wire_d20_88),.data_out(wire_d20_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212090(.data_in(wire_d20_89),.data_out(wire_d20_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212091(.data_in(wire_d20_90),.data_out(wire_d20_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212092(.data_in(wire_d20_91),.data_out(wire_d20_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212093(.data_in(wire_d20_92),.data_out(wire_d20_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212094(.data_in(wire_d20_93),.data_out(wire_d20_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212095(.data_in(wire_d20_94),.data_out(wire_d20_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212096(.data_in(wire_d20_95),.data_out(wire_d20_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212097(.data_in(wire_d20_96),.data_out(wire_d20_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212098(.data_in(wire_d20_97),.data_out(wire_d20_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212099(.data_in(wire_d20_98),.data_out(d_out20),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance22210(.data_in(d_in21),.data_out(wire_d21_0),.clk(clk),.rst(rst));            //channel 22
	invertion #(.WIDTH(WIDTH)) invertion_instance22211(.data_in(wire_d21_0),.data_out(wire_d21_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance22212(.data_in(wire_d21_1),.data_out(wire_d21_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance22213(.data_in(wire_d21_2),.data_out(wire_d21_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance22214(.data_in(wire_d21_3),.data_out(wire_d21_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance22215(.data_in(wire_d21_4),.data_out(wire_d21_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance22216(.data_in(wire_d21_5),.data_out(wire_d21_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance22217(.data_in(wire_d21_6),.data_out(wire_d21_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance22218(.data_in(wire_d21_7),.data_out(wire_d21_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance22219(.data_in(wire_d21_8),.data_out(wire_d21_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222110(.data_in(wire_d21_9),.data_out(wire_d21_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222111(.data_in(wire_d21_10),.data_out(wire_d21_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222112(.data_in(wire_d21_11),.data_out(wire_d21_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222113(.data_in(wire_d21_12),.data_out(wire_d21_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222114(.data_in(wire_d21_13),.data_out(wire_d21_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222115(.data_in(wire_d21_14),.data_out(wire_d21_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222116(.data_in(wire_d21_15),.data_out(wire_d21_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222117(.data_in(wire_d21_16),.data_out(wire_d21_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222118(.data_in(wire_d21_17),.data_out(wire_d21_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222119(.data_in(wire_d21_18),.data_out(wire_d21_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222120(.data_in(wire_d21_19),.data_out(wire_d21_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222121(.data_in(wire_d21_20),.data_out(wire_d21_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222122(.data_in(wire_d21_21),.data_out(wire_d21_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222123(.data_in(wire_d21_22),.data_out(wire_d21_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222124(.data_in(wire_d21_23),.data_out(wire_d21_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222125(.data_in(wire_d21_24),.data_out(wire_d21_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222126(.data_in(wire_d21_25),.data_out(wire_d21_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222127(.data_in(wire_d21_26),.data_out(wire_d21_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222128(.data_in(wire_d21_27),.data_out(wire_d21_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222129(.data_in(wire_d21_28),.data_out(wire_d21_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222130(.data_in(wire_d21_29),.data_out(wire_d21_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222131(.data_in(wire_d21_30),.data_out(wire_d21_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222132(.data_in(wire_d21_31),.data_out(wire_d21_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222133(.data_in(wire_d21_32),.data_out(wire_d21_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222134(.data_in(wire_d21_33),.data_out(wire_d21_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222135(.data_in(wire_d21_34),.data_out(wire_d21_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222136(.data_in(wire_d21_35),.data_out(wire_d21_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222137(.data_in(wire_d21_36),.data_out(wire_d21_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222138(.data_in(wire_d21_37),.data_out(wire_d21_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222139(.data_in(wire_d21_38),.data_out(wire_d21_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222140(.data_in(wire_d21_39),.data_out(wire_d21_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222141(.data_in(wire_d21_40),.data_out(wire_d21_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222142(.data_in(wire_d21_41),.data_out(wire_d21_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222143(.data_in(wire_d21_42),.data_out(wire_d21_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222144(.data_in(wire_d21_43),.data_out(wire_d21_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222145(.data_in(wire_d21_44),.data_out(wire_d21_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222146(.data_in(wire_d21_45),.data_out(wire_d21_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222147(.data_in(wire_d21_46),.data_out(wire_d21_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222148(.data_in(wire_d21_47),.data_out(wire_d21_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222149(.data_in(wire_d21_48),.data_out(wire_d21_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222150(.data_in(wire_d21_49),.data_out(wire_d21_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222151(.data_in(wire_d21_50),.data_out(wire_d21_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222152(.data_in(wire_d21_51),.data_out(wire_d21_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222153(.data_in(wire_d21_52),.data_out(wire_d21_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222154(.data_in(wire_d21_53),.data_out(wire_d21_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222155(.data_in(wire_d21_54),.data_out(wire_d21_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222156(.data_in(wire_d21_55),.data_out(wire_d21_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222157(.data_in(wire_d21_56),.data_out(wire_d21_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222158(.data_in(wire_d21_57),.data_out(wire_d21_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222159(.data_in(wire_d21_58),.data_out(wire_d21_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222160(.data_in(wire_d21_59),.data_out(wire_d21_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222161(.data_in(wire_d21_60),.data_out(wire_d21_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222162(.data_in(wire_d21_61),.data_out(wire_d21_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222163(.data_in(wire_d21_62),.data_out(wire_d21_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222164(.data_in(wire_d21_63),.data_out(wire_d21_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222165(.data_in(wire_d21_64),.data_out(wire_d21_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222166(.data_in(wire_d21_65),.data_out(wire_d21_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222167(.data_in(wire_d21_66),.data_out(wire_d21_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222168(.data_in(wire_d21_67),.data_out(wire_d21_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222169(.data_in(wire_d21_68),.data_out(wire_d21_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222170(.data_in(wire_d21_69),.data_out(wire_d21_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222171(.data_in(wire_d21_70),.data_out(wire_d21_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222172(.data_in(wire_d21_71),.data_out(wire_d21_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222173(.data_in(wire_d21_72),.data_out(wire_d21_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222174(.data_in(wire_d21_73),.data_out(wire_d21_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222175(.data_in(wire_d21_74),.data_out(wire_d21_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222176(.data_in(wire_d21_75),.data_out(wire_d21_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222177(.data_in(wire_d21_76),.data_out(wire_d21_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222178(.data_in(wire_d21_77),.data_out(wire_d21_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222179(.data_in(wire_d21_78),.data_out(wire_d21_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222180(.data_in(wire_d21_79),.data_out(wire_d21_80),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222181(.data_in(wire_d21_80),.data_out(wire_d21_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222182(.data_in(wire_d21_81),.data_out(wire_d21_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222183(.data_in(wire_d21_82),.data_out(wire_d21_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222184(.data_in(wire_d21_83),.data_out(wire_d21_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222185(.data_in(wire_d21_84),.data_out(wire_d21_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222186(.data_in(wire_d21_85),.data_out(wire_d21_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222187(.data_in(wire_d21_86),.data_out(wire_d21_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222188(.data_in(wire_d21_87),.data_out(wire_d21_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222189(.data_in(wire_d21_88),.data_out(wire_d21_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222190(.data_in(wire_d21_89),.data_out(wire_d21_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222191(.data_in(wire_d21_90),.data_out(wire_d21_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222192(.data_in(wire_d21_91),.data_out(wire_d21_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222193(.data_in(wire_d21_92),.data_out(wire_d21_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222194(.data_in(wire_d21_93),.data_out(wire_d21_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222195(.data_in(wire_d21_94),.data_out(wire_d21_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222196(.data_in(wire_d21_95),.data_out(wire_d21_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222197(.data_in(wire_d21_96),.data_out(wire_d21_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222198(.data_in(wire_d21_97),.data_out(wire_d21_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222199(.data_in(wire_d21_98),.data_out(d_out21),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance23220(.data_in(d_in22),.data_out(wire_d22_0),.clk(clk),.rst(rst));            //channel 23
	register #(.WIDTH(WIDTH)) register_instance23221(.data_in(wire_d22_0),.data_out(wire_d22_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance23222(.data_in(wire_d22_1),.data_out(wire_d22_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance23223(.data_in(wire_d22_2),.data_out(wire_d22_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance23224(.data_in(wire_d22_3),.data_out(wire_d22_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance23225(.data_in(wire_d22_4),.data_out(wire_d22_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance23226(.data_in(wire_d22_5),.data_out(wire_d22_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance23227(.data_in(wire_d22_6),.data_out(wire_d22_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance23228(.data_in(wire_d22_7),.data_out(wire_d22_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance23229(.data_in(wire_d22_8),.data_out(wire_d22_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232210(.data_in(wire_d22_9),.data_out(wire_d22_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232211(.data_in(wire_d22_10),.data_out(wire_d22_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232212(.data_in(wire_d22_11),.data_out(wire_d22_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232213(.data_in(wire_d22_12),.data_out(wire_d22_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232214(.data_in(wire_d22_13),.data_out(wire_d22_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232215(.data_in(wire_d22_14),.data_out(wire_d22_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232216(.data_in(wire_d22_15),.data_out(wire_d22_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232217(.data_in(wire_d22_16),.data_out(wire_d22_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232218(.data_in(wire_d22_17),.data_out(wire_d22_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232219(.data_in(wire_d22_18),.data_out(wire_d22_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232220(.data_in(wire_d22_19),.data_out(wire_d22_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232221(.data_in(wire_d22_20),.data_out(wire_d22_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232222(.data_in(wire_d22_21),.data_out(wire_d22_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232223(.data_in(wire_d22_22),.data_out(wire_d22_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232224(.data_in(wire_d22_23),.data_out(wire_d22_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232225(.data_in(wire_d22_24),.data_out(wire_d22_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232226(.data_in(wire_d22_25),.data_out(wire_d22_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232227(.data_in(wire_d22_26),.data_out(wire_d22_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232228(.data_in(wire_d22_27),.data_out(wire_d22_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232229(.data_in(wire_d22_28),.data_out(wire_d22_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232230(.data_in(wire_d22_29),.data_out(wire_d22_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232231(.data_in(wire_d22_30),.data_out(wire_d22_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232232(.data_in(wire_d22_31),.data_out(wire_d22_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232233(.data_in(wire_d22_32),.data_out(wire_d22_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232234(.data_in(wire_d22_33),.data_out(wire_d22_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232235(.data_in(wire_d22_34),.data_out(wire_d22_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232236(.data_in(wire_d22_35),.data_out(wire_d22_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232237(.data_in(wire_d22_36),.data_out(wire_d22_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232238(.data_in(wire_d22_37),.data_out(wire_d22_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232239(.data_in(wire_d22_38),.data_out(wire_d22_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232240(.data_in(wire_d22_39),.data_out(wire_d22_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232241(.data_in(wire_d22_40),.data_out(wire_d22_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232242(.data_in(wire_d22_41),.data_out(wire_d22_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232243(.data_in(wire_d22_42),.data_out(wire_d22_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232244(.data_in(wire_d22_43),.data_out(wire_d22_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232245(.data_in(wire_d22_44),.data_out(wire_d22_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232246(.data_in(wire_d22_45),.data_out(wire_d22_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232247(.data_in(wire_d22_46),.data_out(wire_d22_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232248(.data_in(wire_d22_47),.data_out(wire_d22_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232249(.data_in(wire_d22_48),.data_out(wire_d22_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232250(.data_in(wire_d22_49),.data_out(wire_d22_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232251(.data_in(wire_d22_50),.data_out(wire_d22_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232252(.data_in(wire_d22_51),.data_out(wire_d22_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232253(.data_in(wire_d22_52),.data_out(wire_d22_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232254(.data_in(wire_d22_53),.data_out(wire_d22_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232255(.data_in(wire_d22_54),.data_out(wire_d22_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232256(.data_in(wire_d22_55),.data_out(wire_d22_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232257(.data_in(wire_d22_56),.data_out(wire_d22_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232258(.data_in(wire_d22_57),.data_out(wire_d22_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232259(.data_in(wire_d22_58),.data_out(wire_d22_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232260(.data_in(wire_d22_59),.data_out(wire_d22_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232261(.data_in(wire_d22_60),.data_out(wire_d22_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232262(.data_in(wire_d22_61),.data_out(wire_d22_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232263(.data_in(wire_d22_62),.data_out(wire_d22_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232264(.data_in(wire_d22_63),.data_out(wire_d22_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232265(.data_in(wire_d22_64),.data_out(wire_d22_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232266(.data_in(wire_d22_65),.data_out(wire_d22_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232267(.data_in(wire_d22_66),.data_out(wire_d22_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232268(.data_in(wire_d22_67),.data_out(wire_d22_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232269(.data_in(wire_d22_68),.data_out(wire_d22_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232270(.data_in(wire_d22_69),.data_out(wire_d22_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232271(.data_in(wire_d22_70),.data_out(wire_d22_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232272(.data_in(wire_d22_71),.data_out(wire_d22_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232273(.data_in(wire_d22_72),.data_out(wire_d22_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232274(.data_in(wire_d22_73),.data_out(wire_d22_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232275(.data_in(wire_d22_74),.data_out(wire_d22_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232276(.data_in(wire_d22_75),.data_out(wire_d22_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232277(.data_in(wire_d22_76),.data_out(wire_d22_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232278(.data_in(wire_d22_77),.data_out(wire_d22_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232279(.data_in(wire_d22_78),.data_out(wire_d22_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232280(.data_in(wire_d22_79),.data_out(wire_d22_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232281(.data_in(wire_d22_80),.data_out(wire_d22_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232282(.data_in(wire_d22_81),.data_out(wire_d22_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232283(.data_in(wire_d22_82),.data_out(wire_d22_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232284(.data_in(wire_d22_83),.data_out(wire_d22_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232285(.data_in(wire_d22_84),.data_out(wire_d22_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232286(.data_in(wire_d22_85),.data_out(wire_d22_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232287(.data_in(wire_d22_86),.data_out(wire_d22_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232288(.data_in(wire_d22_87),.data_out(wire_d22_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232289(.data_in(wire_d22_88),.data_out(wire_d22_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232290(.data_in(wire_d22_89),.data_out(wire_d22_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232291(.data_in(wire_d22_90),.data_out(wire_d22_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232292(.data_in(wire_d22_91),.data_out(wire_d22_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232293(.data_in(wire_d22_92),.data_out(wire_d22_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232294(.data_in(wire_d22_93),.data_out(wire_d22_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232295(.data_in(wire_d22_94),.data_out(wire_d22_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232296(.data_in(wire_d22_95),.data_out(wire_d22_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232297(.data_in(wire_d22_96),.data_out(wire_d22_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232298(.data_in(wire_d22_97),.data_out(wire_d22_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232299(.data_in(wire_d22_98),.data_out(d_out22),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance24230(.data_in(d_in23),.data_out(wire_d23_0),.clk(clk),.rst(rst));            //channel 24
	large_mux #(.WIDTH(WIDTH)) large_mux_instance24231(.data_in(wire_d23_0),.data_out(wire_d23_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance24232(.data_in(wire_d23_1),.data_out(wire_d23_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance24233(.data_in(wire_d23_2),.data_out(wire_d23_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance24234(.data_in(wire_d23_3),.data_out(wire_d23_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance24235(.data_in(wire_d23_4),.data_out(wire_d23_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance24236(.data_in(wire_d23_5),.data_out(wire_d23_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance24237(.data_in(wire_d23_6),.data_out(wire_d23_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance24238(.data_in(wire_d23_7),.data_out(wire_d23_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance24239(.data_in(wire_d23_8),.data_out(wire_d23_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242310(.data_in(wire_d23_9),.data_out(wire_d23_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242311(.data_in(wire_d23_10),.data_out(wire_d23_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242312(.data_in(wire_d23_11),.data_out(wire_d23_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242313(.data_in(wire_d23_12),.data_out(wire_d23_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242314(.data_in(wire_d23_13),.data_out(wire_d23_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242315(.data_in(wire_d23_14),.data_out(wire_d23_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242316(.data_in(wire_d23_15),.data_out(wire_d23_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242317(.data_in(wire_d23_16),.data_out(wire_d23_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242318(.data_in(wire_d23_17),.data_out(wire_d23_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242319(.data_in(wire_d23_18),.data_out(wire_d23_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242320(.data_in(wire_d23_19),.data_out(wire_d23_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242321(.data_in(wire_d23_20),.data_out(wire_d23_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242322(.data_in(wire_d23_21),.data_out(wire_d23_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242323(.data_in(wire_d23_22),.data_out(wire_d23_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242324(.data_in(wire_d23_23),.data_out(wire_d23_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242325(.data_in(wire_d23_24),.data_out(wire_d23_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242326(.data_in(wire_d23_25),.data_out(wire_d23_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242327(.data_in(wire_d23_26),.data_out(wire_d23_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242328(.data_in(wire_d23_27),.data_out(wire_d23_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242329(.data_in(wire_d23_28),.data_out(wire_d23_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242330(.data_in(wire_d23_29),.data_out(wire_d23_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242331(.data_in(wire_d23_30),.data_out(wire_d23_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242332(.data_in(wire_d23_31),.data_out(wire_d23_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242333(.data_in(wire_d23_32),.data_out(wire_d23_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242334(.data_in(wire_d23_33),.data_out(wire_d23_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242335(.data_in(wire_d23_34),.data_out(wire_d23_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242336(.data_in(wire_d23_35),.data_out(wire_d23_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242337(.data_in(wire_d23_36),.data_out(wire_d23_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242338(.data_in(wire_d23_37),.data_out(wire_d23_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242339(.data_in(wire_d23_38),.data_out(wire_d23_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242340(.data_in(wire_d23_39),.data_out(wire_d23_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242341(.data_in(wire_d23_40),.data_out(wire_d23_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242342(.data_in(wire_d23_41),.data_out(wire_d23_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242343(.data_in(wire_d23_42),.data_out(wire_d23_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242344(.data_in(wire_d23_43),.data_out(wire_d23_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242345(.data_in(wire_d23_44),.data_out(wire_d23_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242346(.data_in(wire_d23_45),.data_out(wire_d23_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242347(.data_in(wire_d23_46),.data_out(wire_d23_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242348(.data_in(wire_d23_47),.data_out(wire_d23_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242349(.data_in(wire_d23_48),.data_out(wire_d23_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242350(.data_in(wire_d23_49),.data_out(wire_d23_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242351(.data_in(wire_d23_50),.data_out(wire_d23_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242352(.data_in(wire_d23_51),.data_out(wire_d23_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242353(.data_in(wire_d23_52),.data_out(wire_d23_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242354(.data_in(wire_d23_53),.data_out(wire_d23_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242355(.data_in(wire_d23_54),.data_out(wire_d23_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242356(.data_in(wire_d23_55),.data_out(wire_d23_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242357(.data_in(wire_d23_56),.data_out(wire_d23_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242358(.data_in(wire_d23_57),.data_out(wire_d23_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242359(.data_in(wire_d23_58),.data_out(wire_d23_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242360(.data_in(wire_d23_59),.data_out(wire_d23_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242361(.data_in(wire_d23_60),.data_out(wire_d23_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242362(.data_in(wire_d23_61),.data_out(wire_d23_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242363(.data_in(wire_d23_62),.data_out(wire_d23_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242364(.data_in(wire_d23_63),.data_out(wire_d23_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242365(.data_in(wire_d23_64),.data_out(wire_d23_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242366(.data_in(wire_d23_65),.data_out(wire_d23_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242367(.data_in(wire_d23_66),.data_out(wire_d23_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242368(.data_in(wire_d23_67),.data_out(wire_d23_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242369(.data_in(wire_d23_68),.data_out(wire_d23_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242370(.data_in(wire_d23_69),.data_out(wire_d23_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242371(.data_in(wire_d23_70),.data_out(wire_d23_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242372(.data_in(wire_d23_71),.data_out(wire_d23_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242373(.data_in(wire_d23_72),.data_out(wire_d23_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242374(.data_in(wire_d23_73),.data_out(wire_d23_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242375(.data_in(wire_d23_74),.data_out(wire_d23_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242376(.data_in(wire_d23_75),.data_out(wire_d23_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242377(.data_in(wire_d23_76),.data_out(wire_d23_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242378(.data_in(wire_d23_77),.data_out(wire_d23_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242379(.data_in(wire_d23_78),.data_out(wire_d23_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242380(.data_in(wire_d23_79),.data_out(wire_d23_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242381(.data_in(wire_d23_80),.data_out(wire_d23_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242382(.data_in(wire_d23_81),.data_out(wire_d23_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242383(.data_in(wire_d23_82),.data_out(wire_d23_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242384(.data_in(wire_d23_83),.data_out(wire_d23_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242385(.data_in(wire_d23_84),.data_out(wire_d23_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242386(.data_in(wire_d23_85),.data_out(wire_d23_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242387(.data_in(wire_d23_86),.data_out(wire_d23_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242388(.data_in(wire_d23_87),.data_out(wire_d23_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242389(.data_in(wire_d23_88),.data_out(wire_d23_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242390(.data_in(wire_d23_89),.data_out(wire_d23_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242391(.data_in(wire_d23_90),.data_out(wire_d23_91),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242392(.data_in(wire_d23_91),.data_out(wire_d23_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242393(.data_in(wire_d23_92),.data_out(wire_d23_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242394(.data_in(wire_d23_93),.data_out(wire_d23_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242395(.data_in(wire_d23_94),.data_out(wire_d23_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242396(.data_in(wire_d23_95),.data_out(wire_d23_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242397(.data_in(wire_d23_96),.data_out(wire_d23_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242398(.data_in(wire_d23_97),.data_out(wire_d23_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242399(.data_in(wire_d23_98),.data_out(d_out23),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance25240(.data_in(d_in24),.data_out(wire_d24_0),.clk(clk),.rst(rst));            //channel 25
	large_mux #(.WIDTH(WIDTH)) large_mux_instance25241(.data_in(wire_d24_0),.data_out(wire_d24_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance25242(.data_in(wire_d24_1),.data_out(wire_d24_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance25243(.data_in(wire_d24_2),.data_out(wire_d24_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance25244(.data_in(wire_d24_3),.data_out(wire_d24_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance25245(.data_in(wire_d24_4),.data_out(wire_d24_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance25246(.data_in(wire_d24_5),.data_out(wire_d24_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance25247(.data_in(wire_d24_6),.data_out(wire_d24_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance25248(.data_in(wire_d24_7),.data_out(wire_d24_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance25249(.data_in(wire_d24_8),.data_out(wire_d24_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252410(.data_in(wire_d24_9),.data_out(wire_d24_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252411(.data_in(wire_d24_10),.data_out(wire_d24_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252412(.data_in(wire_d24_11),.data_out(wire_d24_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252413(.data_in(wire_d24_12),.data_out(wire_d24_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252414(.data_in(wire_d24_13),.data_out(wire_d24_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252415(.data_in(wire_d24_14),.data_out(wire_d24_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252416(.data_in(wire_d24_15),.data_out(wire_d24_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252417(.data_in(wire_d24_16),.data_out(wire_d24_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252418(.data_in(wire_d24_17),.data_out(wire_d24_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252419(.data_in(wire_d24_18),.data_out(wire_d24_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252420(.data_in(wire_d24_19),.data_out(wire_d24_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252421(.data_in(wire_d24_20),.data_out(wire_d24_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252422(.data_in(wire_d24_21),.data_out(wire_d24_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252423(.data_in(wire_d24_22),.data_out(wire_d24_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252424(.data_in(wire_d24_23),.data_out(wire_d24_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252425(.data_in(wire_d24_24),.data_out(wire_d24_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252426(.data_in(wire_d24_25),.data_out(wire_d24_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252427(.data_in(wire_d24_26),.data_out(wire_d24_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252428(.data_in(wire_d24_27),.data_out(wire_d24_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252429(.data_in(wire_d24_28),.data_out(wire_d24_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252430(.data_in(wire_d24_29),.data_out(wire_d24_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252431(.data_in(wire_d24_30),.data_out(wire_d24_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252432(.data_in(wire_d24_31),.data_out(wire_d24_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252433(.data_in(wire_d24_32),.data_out(wire_d24_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252434(.data_in(wire_d24_33),.data_out(wire_d24_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252435(.data_in(wire_d24_34),.data_out(wire_d24_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252436(.data_in(wire_d24_35),.data_out(wire_d24_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252437(.data_in(wire_d24_36),.data_out(wire_d24_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252438(.data_in(wire_d24_37),.data_out(wire_d24_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252439(.data_in(wire_d24_38),.data_out(wire_d24_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252440(.data_in(wire_d24_39),.data_out(wire_d24_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252441(.data_in(wire_d24_40),.data_out(wire_d24_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252442(.data_in(wire_d24_41),.data_out(wire_d24_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252443(.data_in(wire_d24_42),.data_out(wire_d24_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252444(.data_in(wire_d24_43),.data_out(wire_d24_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252445(.data_in(wire_d24_44),.data_out(wire_d24_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252446(.data_in(wire_d24_45),.data_out(wire_d24_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252447(.data_in(wire_d24_46),.data_out(wire_d24_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252448(.data_in(wire_d24_47),.data_out(wire_d24_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252449(.data_in(wire_d24_48),.data_out(wire_d24_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252450(.data_in(wire_d24_49),.data_out(wire_d24_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252451(.data_in(wire_d24_50),.data_out(wire_d24_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252452(.data_in(wire_d24_51),.data_out(wire_d24_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252453(.data_in(wire_d24_52),.data_out(wire_d24_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252454(.data_in(wire_d24_53),.data_out(wire_d24_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252455(.data_in(wire_d24_54),.data_out(wire_d24_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252456(.data_in(wire_d24_55),.data_out(wire_d24_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252457(.data_in(wire_d24_56),.data_out(wire_d24_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252458(.data_in(wire_d24_57),.data_out(wire_d24_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252459(.data_in(wire_d24_58),.data_out(wire_d24_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252460(.data_in(wire_d24_59),.data_out(wire_d24_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252461(.data_in(wire_d24_60),.data_out(wire_d24_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252462(.data_in(wire_d24_61),.data_out(wire_d24_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252463(.data_in(wire_d24_62),.data_out(wire_d24_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252464(.data_in(wire_d24_63),.data_out(wire_d24_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252465(.data_in(wire_d24_64),.data_out(wire_d24_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252466(.data_in(wire_d24_65),.data_out(wire_d24_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252467(.data_in(wire_d24_66),.data_out(wire_d24_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252468(.data_in(wire_d24_67),.data_out(wire_d24_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252469(.data_in(wire_d24_68),.data_out(wire_d24_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252470(.data_in(wire_d24_69),.data_out(wire_d24_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252471(.data_in(wire_d24_70),.data_out(wire_d24_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252472(.data_in(wire_d24_71),.data_out(wire_d24_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252473(.data_in(wire_d24_72),.data_out(wire_d24_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252474(.data_in(wire_d24_73),.data_out(wire_d24_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252475(.data_in(wire_d24_74),.data_out(wire_d24_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252476(.data_in(wire_d24_75),.data_out(wire_d24_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252477(.data_in(wire_d24_76),.data_out(wire_d24_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252478(.data_in(wire_d24_77),.data_out(wire_d24_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252479(.data_in(wire_d24_78),.data_out(wire_d24_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252480(.data_in(wire_d24_79),.data_out(wire_d24_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252481(.data_in(wire_d24_80),.data_out(wire_d24_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252482(.data_in(wire_d24_81),.data_out(wire_d24_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252483(.data_in(wire_d24_82),.data_out(wire_d24_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252484(.data_in(wire_d24_83),.data_out(wire_d24_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252485(.data_in(wire_d24_84),.data_out(wire_d24_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252486(.data_in(wire_d24_85),.data_out(wire_d24_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252487(.data_in(wire_d24_86),.data_out(wire_d24_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252488(.data_in(wire_d24_87),.data_out(wire_d24_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252489(.data_in(wire_d24_88),.data_out(wire_d24_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252490(.data_in(wire_d24_89),.data_out(wire_d24_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252491(.data_in(wire_d24_90),.data_out(wire_d24_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252492(.data_in(wire_d24_91),.data_out(wire_d24_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252493(.data_in(wire_d24_92),.data_out(wire_d24_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252494(.data_in(wire_d24_93),.data_out(wire_d24_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252495(.data_in(wire_d24_94),.data_out(wire_d24_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252496(.data_in(wire_d24_95),.data_out(wire_d24_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252497(.data_in(wire_d24_96),.data_out(wire_d24_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252498(.data_in(wire_d24_97),.data_out(wire_d24_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252499(.data_in(wire_d24_98),.data_out(d_out24),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance26250(.data_in(d_in25),.data_out(wire_d25_0),.clk(clk),.rst(rst));            //channel 26
	large_mux #(.WIDTH(WIDTH)) large_mux_instance26251(.data_in(wire_d25_0),.data_out(wire_d25_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance26252(.data_in(wire_d25_1),.data_out(wire_d25_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance26253(.data_in(wire_d25_2),.data_out(wire_d25_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance26254(.data_in(wire_d25_3),.data_out(wire_d25_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance26255(.data_in(wire_d25_4),.data_out(wire_d25_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance26256(.data_in(wire_d25_5),.data_out(wire_d25_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance26257(.data_in(wire_d25_6),.data_out(wire_d25_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance26258(.data_in(wire_d25_7),.data_out(wire_d25_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance26259(.data_in(wire_d25_8),.data_out(wire_d25_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262510(.data_in(wire_d25_9),.data_out(wire_d25_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262511(.data_in(wire_d25_10),.data_out(wire_d25_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262512(.data_in(wire_d25_11),.data_out(wire_d25_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262513(.data_in(wire_d25_12),.data_out(wire_d25_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262514(.data_in(wire_d25_13),.data_out(wire_d25_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262515(.data_in(wire_d25_14),.data_out(wire_d25_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262516(.data_in(wire_d25_15),.data_out(wire_d25_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262517(.data_in(wire_d25_16),.data_out(wire_d25_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262518(.data_in(wire_d25_17),.data_out(wire_d25_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262519(.data_in(wire_d25_18),.data_out(wire_d25_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262520(.data_in(wire_d25_19),.data_out(wire_d25_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262521(.data_in(wire_d25_20),.data_out(wire_d25_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262522(.data_in(wire_d25_21),.data_out(wire_d25_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262523(.data_in(wire_d25_22),.data_out(wire_d25_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262524(.data_in(wire_d25_23),.data_out(wire_d25_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262525(.data_in(wire_d25_24),.data_out(wire_d25_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262526(.data_in(wire_d25_25),.data_out(wire_d25_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262527(.data_in(wire_d25_26),.data_out(wire_d25_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262528(.data_in(wire_d25_27),.data_out(wire_d25_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262529(.data_in(wire_d25_28),.data_out(wire_d25_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262530(.data_in(wire_d25_29),.data_out(wire_d25_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262531(.data_in(wire_d25_30),.data_out(wire_d25_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262532(.data_in(wire_d25_31),.data_out(wire_d25_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262533(.data_in(wire_d25_32),.data_out(wire_d25_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262534(.data_in(wire_d25_33),.data_out(wire_d25_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262535(.data_in(wire_d25_34),.data_out(wire_d25_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262536(.data_in(wire_d25_35),.data_out(wire_d25_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262537(.data_in(wire_d25_36),.data_out(wire_d25_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262538(.data_in(wire_d25_37),.data_out(wire_d25_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262539(.data_in(wire_d25_38),.data_out(wire_d25_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262540(.data_in(wire_d25_39),.data_out(wire_d25_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262541(.data_in(wire_d25_40),.data_out(wire_d25_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262542(.data_in(wire_d25_41),.data_out(wire_d25_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262543(.data_in(wire_d25_42),.data_out(wire_d25_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262544(.data_in(wire_d25_43),.data_out(wire_d25_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262545(.data_in(wire_d25_44),.data_out(wire_d25_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262546(.data_in(wire_d25_45),.data_out(wire_d25_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262547(.data_in(wire_d25_46),.data_out(wire_d25_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262548(.data_in(wire_d25_47),.data_out(wire_d25_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262549(.data_in(wire_d25_48),.data_out(wire_d25_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262550(.data_in(wire_d25_49),.data_out(wire_d25_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262551(.data_in(wire_d25_50),.data_out(wire_d25_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262552(.data_in(wire_d25_51),.data_out(wire_d25_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262553(.data_in(wire_d25_52),.data_out(wire_d25_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262554(.data_in(wire_d25_53),.data_out(wire_d25_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262555(.data_in(wire_d25_54),.data_out(wire_d25_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262556(.data_in(wire_d25_55),.data_out(wire_d25_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262557(.data_in(wire_d25_56),.data_out(wire_d25_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262558(.data_in(wire_d25_57),.data_out(wire_d25_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262559(.data_in(wire_d25_58),.data_out(wire_d25_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262560(.data_in(wire_d25_59),.data_out(wire_d25_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262561(.data_in(wire_d25_60),.data_out(wire_d25_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262562(.data_in(wire_d25_61),.data_out(wire_d25_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262563(.data_in(wire_d25_62),.data_out(wire_d25_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262564(.data_in(wire_d25_63),.data_out(wire_d25_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262565(.data_in(wire_d25_64),.data_out(wire_d25_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262566(.data_in(wire_d25_65),.data_out(wire_d25_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262567(.data_in(wire_d25_66),.data_out(wire_d25_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262568(.data_in(wire_d25_67),.data_out(wire_d25_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262569(.data_in(wire_d25_68),.data_out(wire_d25_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262570(.data_in(wire_d25_69),.data_out(wire_d25_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262571(.data_in(wire_d25_70),.data_out(wire_d25_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262572(.data_in(wire_d25_71),.data_out(wire_d25_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262573(.data_in(wire_d25_72),.data_out(wire_d25_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262574(.data_in(wire_d25_73),.data_out(wire_d25_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262575(.data_in(wire_d25_74),.data_out(wire_d25_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262576(.data_in(wire_d25_75),.data_out(wire_d25_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262577(.data_in(wire_d25_76),.data_out(wire_d25_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262578(.data_in(wire_d25_77),.data_out(wire_d25_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262579(.data_in(wire_d25_78),.data_out(wire_d25_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262580(.data_in(wire_d25_79),.data_out(wire_d25_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262581(.data_in(wire_d25_80),.data_out(wire_d25_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262582(.data_in(wire_d25_81),.data_out(wire_d25_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262583(.data_in(wire_d25_82),.data_out(wire_d25_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262584(.data_in(wire_d25_83),.data_out(wire_d25_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262585(.data_in(wire_d25_84),.data_out(wire_d25_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262586(.data_in(wire_d25_85),.data_out(wire_d25_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262587(.data_in(wire_d25_86),.data_out(wire_d25_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262588(.data_in(wire_d25_87),.data_out(wire_d25_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262589(.data_in(wire_d25_88),.data_out(wire_d25_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262590(.data_in(wire_d25_89),.data_out(wire_d25_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262591(.data_in(wire_d25_90),.data_out(wire_d25_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262592(.data_in(wire_d25_91),.data_out(wire_d25_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262593(.data_in(wire_d25_92),.data_out(wire_d25_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262594(.data_in(wire_d25_93),.data_out(wire_d25_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262595(.data_in(wire_d25_94),.data_out(wire_d25_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262596(.data_in(wire_d25_95),.data_out(wire_d25_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262597(.data_in(wire_d25_96),.data_out(wire_d25_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262598(.data_in(wire_d25_97),.data_out(wire_d25_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262599(.data_in(wire_d25_98),.data_out(d_out25),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance27260(.data_in(d_in26),.data_out(wire_d26_0),.clk(clk),.rst(rst));            //channel 27
	invertion #(.WIDTH(WIDTH)) invertion_instance27261(.data_in(wire_d26_0),.data_out(wire_d26_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance27262(.data_in(wire_d26_1),.data_out(wire_d26_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance27263(.data_in(wire_d26_2),.data_out(wire_d26_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance27264(.data_in(wire_d26_3),.data_out(wire_d26_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance27265(.data_in(wire_d26_4),.data_out(wire_d26_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance27266(.data_in(wire_d26_5),.data_out(wire_d26_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance27267(.data_in(wire_d26_6),.data_out(wire_d26_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance27268(.data_in(wire_d26_7),.data_out(wire_d26_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance27269(.data_in(wire_d26_8),.data_out(wire_d26_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272610(.data_in(wire_d26_9),.data_out(wire_d26_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272611(.data_in(wire_d26_10),.data_out(wire_d26_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272612(.data_in(wire_d26_11),.data_out(wire_d26_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272613(.data_in(wire_d26_12),.data_out(wire_d26_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272614(.data_in(wire_d26_13),.data_out(wire_d26_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272615(.data_in(wire_d26_14),.data_out(wire_d26_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272616(.data_in(wire_d26_15),.data_out(wire_d26_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272617(.data_in(wire_d26_16),.data_out(wire_d26_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272618(.data_in(wire_d26_17),.data_out(wire_d26_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272619(.data_in(wire_d26_18),.data_out(wire_d26_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272620(.data_in(wire_d26_19),.data_out(wire_d26_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272621(.data_in(wire_d26_20),.data_out(wire_d26_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272622(.data_in(wire_d26_21),.data_out(wire_d26_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272623(.data_in(wire_d26_22),.data_out(wire_d26_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272624(.data_in(wire_d26_23),.data_out(wire_d26_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272625(.data_in(wire_d26_24),.data_out(wire_d26_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272626(.data_in(wire_d26_25),.data_out(wire_d26_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272627(.data_in(wire_d26_26),.data_out(wire_d26_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272628(.data_in(wire_d26_27),.data_out(wire_d26_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272629(.data_in(wire_d26_28),.data_out(wire_d26_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272630(.data_in(wire_d26_29),.data_out(wire_d26_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272631(.data_in(wire_d26_30),.data_out(wire_d26_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272632(.data_in(wire_d26_31),.data_out(wire_d26_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272633(.data_in(wire_d26_32),.data_out(wire_d26_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272634(.data_in(wire_d26_33),.data_out(wire_d26_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272635(.data_in(wire_d26_34),.data_out(wire_d26_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272636(.data_in(wire_d26_35),.data_out(wire_d26_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272637(.data_in(wire_d26_36),.data_out(wire_d26_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272638(.data_in(wire_d26_37),.data_out(wire_d26_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272639(.data_in(wire_d26_38),.data_out(wire_d26_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272640(.data_in(wire_d26_39),.data_out(wire_d26_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272641(.data_in(wire_d26_40),.data_out(wire_d26_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272642(.data_in(wire_d26_41),.data_out(wire_d26_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272643(.data_in(wire_d26_42),.data_out(wire_d26_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272644(.data_in(wire_d26_43),.data_out(wire_d26_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272645(.data_in(wire_d26_44),.data_out(wire_d26_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272646(.data_in(wire_d26_45),.data_out(wire_d26_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272647(.data_in(wire_d26_46),.data_out(wire_d26_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272648(.data_in(wire_d26_47),.data_out(wire_d26_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272649(.data_in(wire_d26_48),.data_out(wire_d26_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272650(.data_in(wire_d26_49),.data_out(wire_d26_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272651(.data_in(wire_d26_50),.data_out(wire_d26_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272652(.data_in(wire_d26_51),.data_out(wire_d26_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272653(.data_in(wire_d26_52),.data_out(wire_d26_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272654(.data_in(wire_d26_53),.data_out(wire_d26_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272655(.data_in(wire_d26_54),.data_out(wire_d26_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272656(.data_in(wire_d26_55),.data_out(wire_d26_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272657(.data_in(wire_d26_56),.data_out(wire_d26_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272658(.data_in(wire_d26_57),.data_out(wire_d26_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272659(.data_in(wire_d26_58),.data_out(wire_d26_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272660(.data_in(wire_d26_59),.data_out(wire_d26_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272661(.data_in(wire_d26_60),.data_out(wire_d26_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272662(.data_in(wire_d26_61),.data_out(wire_d26_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272663(.data_in(wire_d26_62),.data_out(wire_d26_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272664(.data_in(wire_d26_63),.data_out(wire_d26_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272665(.data_in(wire_d26_64),.data_out(wire_d26_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272666(.data_in(wire_d26_65),.data_out(wire_d26_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272667(.data_in(wire_d26_66),.data_out(wire_d26_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272668(.data_in(wire_d26_67),.data_out(wire_d26_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272669(.data_in(wire_d26_68),.data_out(wire_d26_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272670(.data_in(wire_d26_69),.data_out(wire_d26_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272671(.data_in(wire_d26_70),.data_out(wire_d26_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272672(.data_in(wire_d26_71),.data_out(wire_d26_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272673(.data_in(wire_d26_72),.data_out(wire_d26_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272674(.data_in(wire_d26_73),.data_out(wire_d26_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272675(.data_in(wire_d26_74),.data_out(wire_d26_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272676(.data_in(wire_d26_75),.data_out(wire_d26_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272677(.data_in(wire_d26_76),.data_out(wire_d26_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272678(.data_in(wire_d26_77),.data_out(wire_d26_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272679(.data_in(wire_d26_78),.data_out(wire_d26_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272680(.data_in(wire_d26_79),.data_out(wire_d26_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272681(.data_in(wire_d26_80),.data_out(wire_d26_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272682(.data_in(wire_d26_81),.data_out(wire_d26_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272683(.data_in(wire_d26_82),.data_out(wire_d26_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272684(.data_in(wire_d26_83),.data_out(wire_d26_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272685(.data_in(wire_d26_84),.data_out(wire_d26_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272686(.data_in(wire_d26_85),.data_out(wire_d26_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272687(.data_in(wire_d26_86),.data_out(wire_d26_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272688(.data_in(wire_d26_87),.data_out(wire_d26_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272689(.data_in(wire_d26_88),.data_out(wire_d26_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272690(.data_in(wire_d26_89),.data_out(wire_d26_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272691(.data_in(wire_d26_90),.data_out(wire_d26_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272692(.data_in(wire_d26_91),.data_out(wire_d26_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272693(.data_in(wire_d26_92),.data_out(wire_d26_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272694(.data_in(wire_d26_93),.data_out(wire_d26_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272695(.data_in(wire_d26_94),.data_out(wire_d26_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272696(.data_in(wire_d26_95),.data_out(wire_d26_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272697(.data_in(wire_d26_96),.data_out(wire_d26_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272698(.data_in(wire_d26_97),.data_out(wire_d26_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272699(.data_in(wire_d26_98),.data_out(d_out26),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance28270(.data_in(d_in27),.data_out(wire_d27_0),.clk(clk),.rst(rst));            //channel 28
	register #(.WIDTH(WIDTH)) register_instance28271(.data_in(wire_d27_0),.data_out(wire_d27_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance28272(.data_in(wire_d27_1),.data_out(wire_d27_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance28273(.data_in(wire_d27_2),.data_out(wire_d27_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance28274(.data_in(wire_d27_3),.data_out(wire_d27_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance28275(.data_in(wire_d27_4),.data_out(wire_d27_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance28276(.data_in(wire_d27_5),.data_out(wire_d27_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance28277(.data_in(wire_d27_6),.data_out(wire_d27_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance28278(.data_in(wire_d27_7),.data_out(wire_d27_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance28279(.data_in(wire_d27_8),.data_out(wire_d27_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282710(.data_in(wire_d27_9),.data_out(wire_d27_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282711(.data_in(wire_d27_10),.data_out(wire_d27_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282712(.data_in(wire_d27_11),.data_out(wire_d27_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282713(.data_in(wire_d27_12),.data_out(wire_d27_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282714(.data_in(wire_d27_13),.data_out(wire_d27_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282715(.data_in(wire_d27_14),.data_out(wire_d27_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282716(.data_in(wire_d27_15),.data_out(wire_d27_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282717(.data_in(wire_d27_16),.data_out(wire_d27_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282718(.data_in(wire_d27_17),.data_out(wire_d27_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282719(.data_in(wire_d27_18),.data_out(wire_d27_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282720(.data_in(wire_d27_19),.data_out(wire_d27_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282721(.data_in(wire_d27_20),.data_out(wire_d27_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282722(.data_in(wire_d27_21),.data_out(wire_d27_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282723(.data_in(wire_d27_22),.data_out(wire_d27_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282724(.data_in(wire_d27_23),.data_out(wire_d27_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282725(.data_in(wire_d27_24),.data_out(wire_d27_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282726(.data_in(wire_d27_25),.data_out(wire_d27_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282727(.data_in(wire_d27_26),.data_out(wire_d27_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282728(.data_in(wire_d27_27),.data_out(wire_d27_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282729(.data_in(wire_d27_28),.data_out(wire_d27_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282730(.data_in(wire_d27_29),.data_out(wire_d27_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282731(.data_in(wire_d27_30),.data_out(wire_d27_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282732(.data_in(wire_d27_31),.data_out(wire_d27_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282733(.data_in(wire_d27_32),.data_out(wire_d27_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282734(.data_in(wire_d27_33),.data_out(wire_d27_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282735(.data_in(wire_d27_34),.data_out(wire_d27_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282736(.data_in(wire_d27_35),.data_out(wire_d27_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282737(.data_in(wire_d27_36),.data_out(wire_d27_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282738(.data_in(wire_d27_37),.data_out(wire_d27_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282739(.data_in(wire_d27_38),.data_out(wire_d27_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282740(.data_in(wire_d27_39),.data_out(wire_d27_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282741(.data_in(wire_d27_40),.data_out(wire_d27_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282742(.data_in(wire_d27_41),.data_out(wire_d27_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282743(.data_in(wire_d27_42),.data_out(wire_d27_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282744(.data_in(wire_d27_43),.data_out(wire_d27_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282745(.data_in(wire_d27_44),.data_out(wire_d27_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282746(.data_in(wire_d27_45),.data_out(wire_d27_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282747(.data_in(wire_d27_46),.data_out(wire_d27_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282748(.data_in(wire_d27_47),.data_out(wire_d27_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282749(.data_in(wire_d27_48),.data_out(wire_d27_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282750(.data_in(wire_d27_49),.data_out(wire_d27_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282751(.data_in(wire_d27_50),.data_out(wire_d27_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282752(.data_in(wire_d27_51),.data_out(wire_d27_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282753(.data_in(wire_d27_52),.data_out(wire_d27_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282754(.data_in(wire_d27_53),.data_out(wire_d27_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282755(.data_in(wire_d27_54),.data_out(wire_d27_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282756(.data_in(wire_d27_55),.data_out(wire_d27_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282757(.data_in(wire_d27_56),.data_out(wire_d27_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282758(.data_in(wire_d27_57),.data_out(wire_d27_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282759(.data_in(wire_d27_58),.data_out(wire_d27_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282760(.data_in(wire_d27_59),.data_out(wire_d27_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282761(.data_in(wire_d27_60),.data_out(wire_d27_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282762(.data_in(wire_d27_61),.data_out(wire_d27_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282763(.data_in(wire_d27_62),.data_out(wire_d27_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282764(.data_in(wire_d27_63),.data_out(wire_d27_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282765(.data_in(wire_d27_64),.data_out(wire_d27_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282766(.data_in(wire_d27_65),.data_out(wire_d27_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282767(.data_in(wire_d27_66),.data_out(wire_d27_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282768(.data_in(wire_d27_67),.data_out(wire_d27_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282769(.data_in(wire_d27_68),.data_out(wire_d27_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282770(.data_in(wire_d27_69),.data_out(wire_d27_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282771(.data_in(wire_d27_70),.data_out(wire_d27_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282772(.data_in(wire_d27_71),.data_out(wire_d27_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282773(.data_in(wire_d27_72),.data_out(wire_d27_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282774(.data_in(wire_d27_73),.data_out(wire_d27_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282775(.data_in(wire_d27_74),.data_out(wire_d27_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282776(.data_in(wire_d27_75),.data_out(wire_d27_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282777(.data_in(wire_d27_76),.data_out(wire_d27_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282778(.data_in(wire_d27_77),.data_out(wire_d27_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282779(.data_in(wire_d27_78),.data_out(wire_d27_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282780(.data_in(wire_d27_79),.data_out(wire_d27_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282781(.data_in(wire_d27_80),.data_out(wire_d27_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282782(.data_in(wire_d27_81),.data_out(wire_d27_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282783(.data_in(wire_d27_82),.data_out(wire_d27_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282784(.data_in(wire_d27_83),.data_out(wire_d27_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282785(.data_in(wire_d27_84),.data_out(wire_d27_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282786(.data_in(wire_d27_85),.data_out(wire_d27_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282787(.data_in(wire_d27_86),.data_out(wire_d27_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282788(.data_in(wire_d27_87),.data_out(wire_d27_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282789(.data_in(wire_d27_88),.data_out(wire_d27_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282790(.data_in(wire_d27_89),.data_out(wire_d27_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282791(.data_in(wire_d27_90),.data_out(wire_d27_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282792(.data_in(wire_d27_91),.data_out(wire_d27_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282793(.data_in(wire_d27_92),.data_out(wire_d27_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282794(.data_in(wire_d27_93),.data_out(wire_d27_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282795(.data_in(wire_d27_94),.data_out(wire_d27_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282796(.data_in(wire_d27_95),.data_out(wire_d27_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282797(.data_in(wire_d27_96),.data_out(wire_d27_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282798(.data_in(wire_d27_97),.data_out(wire_d27_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282799(.data_in(wire_d27_98),.data_out(d_out27),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance29280(.data_in(d_in28),.data_out(wire_d28_0),.clk(clk),.rst(rst));            //channel 29
	invertion #(.WIDTH(WIDTH)) invertion_instance29281(.data_in(wire_d28_0),.data_out(wire_d28_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance29282(.data_in(wire_d28_1),.data_out(wire_d28_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance29283(.data_in(wire_d28_2),.data_out(wire_d28_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance29284(.data_in(wire_d28_3),.data_out(wire_d28_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance29285(.data_in(wire_d28_4),.data_out(wire_d28_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance29286(.data_in(wire_d28_5),.data_out(wire_d28_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance29287(.data_in(wire_d28_6),.data_out(wire_d28_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance29288(.data_in(wire_d28_7),.data_out(wire_d28_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance29289(.data_in(wire_d28_8),.data_out(wire_d28_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292810(.data_in(wire_d28_9),.data_out(wire_d28_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292811(.data_in(wire_d28_10),.data_out(wire_d28_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292812(.data_in(wire_d28_11),.data_out(wire_d28_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292813(.data_in(wire_d28_12),.data_out(wire_d28_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292814(.data_in(wire_d28_13),.data_out(wire_d28_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292815(.data_in(wire_d28_14),.data_out(wire_d28_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292816(.data_in(wire_d28_15),.data_out(wire_d28_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292817(.data_in(wire_d28_16),.data_out(wire_d28_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292818(.data_in(wire_d28_17),.data_out(wire_d28_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292819(.data_in(wire_d28_18),.data_out(wire_d28_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292820(.data_in(wire_d28_19),.data_out(wire_d28_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292821(.data_in(wire_d28_20),.data_out(wire_d28_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292822(.data_in(wire_d28_21),.data_out(wire_d28_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292823(.data_in(wire_d28_22),.data_out(wire_d28_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292824(.data_in(wire_d28_23),.data_out(wire_d28_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292825(.data_in(wire_d28_24),.data_out(wire_d28_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292826(.data_in(wire_d28_25),.data_out(wire_d28_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292827(.data_in(wire_d28_26),.data_out(wire_d28_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292828(.data_in(wire_d28_27),.data_out(wire_d28_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292829(.data_in(wire_d28_28),.data_out(wire_d28_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292830(.data_in(wire_d28_29),.data_out(wire_d28_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292831(.data_in(wire_d28_30),.data_out(wire_d28_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292832(.data_in(wire_d28_31),.data_out(wire_d28_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292833(.data_in(wire_d28_32),.data_out(wire_d28_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292834(.data_in(wire_d28_33),.data_out(wire_d28_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292835(.data_in(wire_d28_34),.data_out(wire_d28_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292836(.data_in(wire_d28_35),.data_out(wire_d28_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292837(.data_in(wire_d28_36),.data_out(wire_d28_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292838(.data_in(wire_d28_37),.data_out(wire_d28_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292839(.data_in(wire_d28_38),.data_out(wire_d28_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292840(.data_in(wire_d28_39),.data_out(wire_d28_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292841(.data_in(wire_d28_40),.data_out(wire_d28_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292842(.data_in(wire_d28_41),.data_out(wire_d28_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292843(.data_in(wire_d28_42),.data_out(wire_d28_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292844(.data_in(wire_d28_43),.data_out(wire_d28_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292845(.data_in(wire_d28_44),.data_out(wire_d28_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292846(.data_in(wire_d28_45),.data_out(wire_d28_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292847(.data_in(wire_d28_46),.data_out(wire_d28_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292848(.data_in(wire_d28_47),.data_out(wire_d28_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292849(.data_in(wire_d28_48),.data_out(wire_d28_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292850(.data_in(wire_d28_49),.data_out(wire_d28_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292851(.data_in(wire_d28_50),.data_out(wire_d28_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292852(.data_in(wire_d28_51),.data_out(wire_d28_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292853(.data_in(wire_d28_52),.data_out(wire_d28_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292854(.data_in(wire_d28_53),.data_out(wire_d28_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292855(.data_in(wire_d28_54),.data_out(wire_d28_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292856(.data_in(wire_d28_55),.data_out(wire_d28_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292857(.data_in(wire_d28_56),.data_out(wire_d28_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292858(.data_in(wire_d28_57),.data_out(wire_d28_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292859(.data_in(wire_d28_58),.data_out(wire_d28_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292860(.data_in(wire_d28_59),.data_out(wire_d28_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292861(.data_in(wire_d28_60),.data_out(wire_d28_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292862(.data_in(wire_d28_61),.data_out(wire_d28_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292863(.data_in(wire_d28_62),.data_out(wire_d28_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292864(.data_in(wire_d28_63),.data_out(wire_d28_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292865(.data_in(wire_d28_64),.data_out(wire_d28_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292866(.data_in(wire_d28_65),.data_out(wire_d28_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292867(.data_in(wire_d28_66),.data_out(wire_d28_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292868(.data_in(wire_d28_67),.data_out(wire_d28_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292869(.data_in(wire_d28_68),.data_out(wire_d28_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292870(.data_in(wire_d28_69),.data_out(wire_d28_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292871(.data_in(wire_d28_70),.data_out(wire_d28_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292872(.data_in(wire_d28_71),.data_out(wire_d28_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292873(.data_in(wire_d28_72),.data_out(wire_d28_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292874(.data_in(wire_d28_73),.data_out(wire_d28_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292875(.data_in(wire_d28_74),.data_out(wire_d28_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292876(.data_in(wire_d28_75),.data_out(wire_d28_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292877(.data_in(wire_d28_76),.data_out(wire_d28_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292878(.data_in(wire_d28_77),.data_out(wire_d28_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292879(.data_in(wire_d28_78),.data_out(wire_d28_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292880(.data_in(wire_d28_79),.data_out(wire_d28_80),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292881(.data_in(wire_d28_80),.data_out(wire_d28_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292882(.data_in(wire_d28_81),.data_out(wire_d28_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292883(.data_in(wire_d28_82),.data_out(wire_d28_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292884(.data_in(wire_d28_83),.data_out(wire_d28_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292885(.data_in(wire_d28_84),.data_out(wire_d28_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292886(.data_in(wire_d28_85),.data_out(wire_d28_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292887(.data_in(wire_d28_86),.data_out(wire_d28_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292888(.data_in(wire_d28_87),.data_out(wire_d28_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292889(.data_in(wire_d28_88),.data_out(wire_d28_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292890(.data_in(wire_d28_89),.data_out(wire_d28_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292891(.data_in(wire_d28_90),.data_out(wire_d28_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292892(.data_in(wire_d28_91),.data_out(wire_d28_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292893(.data_in(wire_d28_92),.data_out(wire_d28_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292894(.data_in(wire_d28_93),.data_out(wire_d28_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292895(.data_in(wire_d28_94),.data_out(wire_d28_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292896(.data_in(wire_d28_95),.data_out(wire_d28_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292897(.data_in(wire_d28_96),.data_out(wire_d28_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292898(.data_in(wire_d28_97),.data_out(wire_d28_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292899(.data_in(wire_d28_98),.data_out(d_out28),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance30290(.data_in(d_in29),.data_out(wire_d29_0),.clk(clk),.rst(rst));            //channel 30
	register #(.WIDTH(WIDTH)) register_instance30291(.data_in(wire_d29_0),.data_out(wire_d29_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance30292(.data_in(wire_d29_1),.data_out(wire_d29_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance30293(.data_in(wire_d29_2),.data_out(wire_d29_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance30294(.data_in(wire_d29_3),.data_out(wire_d29_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance30295(.data_in(wire_d29_4),.data_out(wire_d29_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance30296(.data_in(wire_d29_5),.data_out(wire_d29_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance30297(.data_in(wire_d29_6),.data_out(wire_d29_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance30298(.data_in(wire_d29_7),.data_out(wire_d29_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance30299(.data_in(wire_d29_8),.data_out(wire_d29_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302910(.data_in(wire_d29_9),.data_out(wire_d29_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302911(.data_in(wire_d29_10),.data_out(wire_d29_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302912(.data_in(wire_d29_11),.data_out(wire_d29_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302913(.data_in(wire_d29_12),.data_out(wire_d29_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302914(.data_in(wire_d29_13),.data_out(wire_d29_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302915(.data_in(wire_d29_14),.data_out(wire_d29_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302916(.data_in(wire_d29_15),.data_out(wire_d29_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302917(.data_in(wire_d29_16),.data_out(wire_d29_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302918(.data_in(wire_d29_17),.data_out(wire_d29_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302919(.data_in(wire_d29_18),.data_out(wire_d29_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302920(.data_in(wire_d29_19),.data_out(wire_d29_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302921(.data_in(wire_d29_20),.data_out(wire_d29_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302922(.data_in(wire_d29_21),.data_out(wire_d29_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302923(.data_in(wire_d29_22),.data_out(wire_d29_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302924(.data_in(wire_d29_23),.data_out(wire_d29_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302925(.data_in(wire_d29_24),.data_out(wire_d29_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302926(.data_in(wire_d29_25),.data_out(wire_d29_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302927(.data_in(wire_d29_26),.data_out(wire_d29_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302928(.data_in(wire_d29_27),.data_out(wire_d29_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302929(.data_in(wire_d29_28),.data_out(wire_d29_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302930(.data_in(wire_d29_29),.data_out(wire_d29_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302931(.data_in(wire_d29_30),.data_out(wire_d29_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302932(.data_in(wire_d29_31),.data_out(wire_d29_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302933(.data_in(wire_d29_32),.data_out(wire_d29_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302934(.data_in(wire_d29_33),.data_out(wire_d29_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302935(.data_in(wire_d29_34),.data_out(wire_d29_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302936(.data_in(wire_d29_35),.data_out(wire_d29_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302937(.data_in(wire_d29_36),.data_out(wire_d29_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302938(.data_in(wire_d29_37),.data_out(wire_d29_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302939(.data_in(wire_d29_38),.data_out(wire_d29_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302940(.data_in(wire_d29_39),.data_out(wire_d29_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302941(.data_in(wire_d29_40),.data_out(wire_d29_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302942(.data_in(wire_d29_41),.data_out(wire_d29_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302943(.data_in(wire_d29_42),.data_out(wire_d29_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302944(.data_in(wire_d29_43),.data_out(wire_d29_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302945(.data_in(wire_d29_44),.data_out(wire_d29_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302946(.data_in(wire_d29_45),.data_out(wire_d29_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302947(.data_in(wire_d29_46),.data_out(wire_d29_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302948(.data_in(wire_d29_47),.data_out(wire_d29_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302949(.data_in(wire_d29_48),.data_out(wire_d29_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302950(.data_in(wire_d29_49),.data_out(wire_d29_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302951(.data_in(wire_d29_50),.data_out(wire_d29_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302952(.data_in(wire_d29_51),.data_out(wire_d29_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302953(.data_in(wire_d29_52),.data_out(wire_d29_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302954(.data_in(wire_d29_53),.data_out(wire_d29_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302955(.data_in(wire_d29_54),.data_out(wire_d29_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302956(.data_in(wire_d29_55),.data_out(wire_d29_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302957(.data_in(wire_d29_56),.data_out(wire_d29_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302958(.data_in(wire_d29_57),.data_out(wire_d29_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302959(.data_in(wire_d29_58),.data_out(wire_d29_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302960(.data_in(wire_d29_59),.data_out(wire_d29_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302961(.data_in(wire_d29_60),.data_out(wire_d29_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302962(.data_in(wire_d29_61),.data_out(wire_d29_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302963(.data_in(wire_d29_62),.data_out(wire_d29_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302964(.data_in(wire_d29_63),.data_out(wire_d29_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302965(.data_in(wire_d29_64),.data_out(wire_d29_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302966(.data_in(wire_d29_65),.data_out(wire_d29_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302967(.data_in(wire_d29_66),.data_out(wire_d29_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302968(.data_in(wire_d29_67),.data_out(wire_d29_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302969(.data_in(wire_d29_68),.data_out(wire_d29_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302970(.data_in(wire_d29_69),.data_out(wire_d29_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302971(.data_in(wire_d29_70),.data_out(wire_d29_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302972(.data_in(wire_d29_71),.data_out(wire_d29_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302973(.data_in(wire_d29_72),.data_out(wire_d29_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302974(.data_in(wire_d29_73),.data_out(wire_d29_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302975(.data_in(wire_d29_74),.data_out(wire_d29_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302976(.data_in(wire_d29_75),.data_out(wire_d29_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302977(.data_in(wire_d29_76),.data_out(wire_d29_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302978(.data_in(wire_d29_77),.data_out(wire_d29_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302979(.data_in(wire_d29_78),.data_out(wire_d29_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302980(.data_in(wire_d29_79),.data_out(wire_d29_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302981(.data_in(wire_d29_80),.data_out(wire_d29_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302982(.data_in(wire_d29_81),.data_out(wire_d29_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302983(.data_in(wire_d29_82),.data_out(wire_d29_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302984(.data_in(wire_d29_83),.data_out(wire_d29_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302985(.data_in(wire_d29_84),.data_out(wire_d29_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302986(.data_in(wire_d29_85),.data_out(wire_d29_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302987(.data_in(wire_d29_86),.data_out(wire_d29_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302988(.data_in(wire_d29_87),.data_out(wire_d29_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302989(.data_in(wire_d29_88),.data_out(wire_d29_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302990(.data_in(wire_d29_89),.data_out(wire_d29_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302991(.data_in(wire_d29_90),.data_out(wire_d29_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302992(.data_in(wire_d29_91),.data_out(wire_d29_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302993(.data_in(wire_d29_92),.data_out(wire_d29_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302994(.data_in(wire_d29_93),.data_out(wire_d29_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302995(.data_in(wire_d29_94),.data_out(wire_d29_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302996(.data_in(wire_d29_95),.data_out(wire_d29_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302997(.data_in(wire_d29_96),.data_out(wire_d29_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302998(.data_in(wire_d29_97),.data_out(wire_d29_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302999(.data_in(wire_d29_98),.data_out(d_out29),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance31300(.data_in(d_in30),.data_out(wire_d30_0),.clk(clk),.rst(rst));            //channel 31
	encoder #(.WIDTH(WIDTH)) encoder_instance31301(.data_in(wire_d30_0),.data_out(wire_d30_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance31302(.data_in(wire_d30_1),.data_out(wire_d30_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance31303(.data_in(wire_d30_2),.data_out(wire_d30_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance31304(.data_in(wire_d30_3),.data_out(wire_d30_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance31305(.data_in(wire_d30_4),.data_out(wire_d30_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance31306(.data_in(wire_d30_5),.data_out(wire_d30_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance31307(.data_in(wire_d30_6),.data_out(wire_d30_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance31308(.data_in(wire_d30_7),.data_out(wire_d30_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance31309(.data_in(wire_d30_8),.data_out(wire_d30_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313010(.data_in(wire_d30_9),.data_out(wire_d30_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313011(.data_in(wire_d30_10),.data_out(wire_d30_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313012(.data_in(wire_d30_11),.data_out(wire_d30_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313013(.data_in(wire_d30_12),.data_out(wire_d30_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313014(.data_in(wire_d30_13),.data_out(wire_d30_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313015(.data_in(wire_d30_14),.data_out(wire_d30_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313016(.data_in(wire_d30_15),.data_out(wire_d30_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313017(.data_in(wire_d30_16),.data_out(wire_d30_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313018(.data_in(wire_d30_17),.data_out(wire_d30_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313019(.data_in(wire_d30_18),.data_out(wire_d30_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313020(.data_in(wire_d30_19),.data_out(wire_d30_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313021(.data_in(wire_d30_20),.data_out(wire_d30_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313022(.data_in(wire_d30_21),.data_out(wire_d30_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313023(.data_in(wire_d30_22),.data_out(wire_d30_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313024(.data_in(wire_d30_23),.data_out(wire_d30_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313025(.data_in(wire_d30_24),.data_out(wire_d30_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313026(.data_in(wire_d30_25),.data_out(wire_d30_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313027(.data_in(wire_d30_26),.data_out(wire_d30_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313028(.data_in(wire_d30_27),.data_out(wire_d30_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313029(.data_in(wire_d30_28),.data_out(wire_d30_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313030(.data_in(wire_d30_29),.data_out(wire_d30_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313031(.data_in(wire_d30_30),.data_out(wire_d30_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313032(.data_in(wire_d30_31),.data_out(wire_d30_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313033(.data_in(wire_d30_32),.data_out(wire_d30_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313034(.data_in(wire_d30_33),.data_out(wire_d30_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313035(.data_in(wire_d30_34),.data_out(wire_d30_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313036(.data_in(wire_d30_35),.data_out(wire_d30_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313037(.data_in(wire_d30_36),.data_out(wire_d30_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313038(.data_in(wire_d30_37),.data_out(wire_d30_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313039(.data_in(wire_d30_38),.data_out(wire_d30_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313040(.data_in(wire_d30_39),.data_out(wire_d30_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313041(.data_in(wire_d30_40),.data_out(wire_d30_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313042(.data_in(wire_d30_41),.data_out(wire_d30_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313043(.data_in(wire_d30_42),.data_out(wire_d30_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313044(.data_in(wire_d30_43),.data_out(wire_d30_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313045(.data_in(wire_d30_44),.data_out(wire_d30_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313046(.data_in(wire_d30_45),.data_out(wire_d30_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313047(.data_in(wire_d30_46),.data_out(wire_d30_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313048(.data_in(wire_d30_47),.data_out(wire_d30_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313049(.data_in(wire_d30_48),.data_out(wire_d30_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313050(.data_in(wire_d30_49),.data_out(wire_d30_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313051(.data_in(wire_d30_50),.data_out(wire_d30_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313052(.data_in(wire_d30_51),.data_out(wire_d30_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313053(.data_in(wire_d30_52),.data_out(wire_d30_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313054(.data_in(wire_d30_53),.data_out(wire_d30_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313055(.data_in(wire_d30_54),.data_out(wire_d30_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313056(.data_in(wire_d30_55),.data_out(wire_d30_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313057(.data_in(wire_d30_56),.data_out(wire_d30_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313058(.data_in(wire_d30_57),.data_out(wire_d30_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313059(.data_in(wire_d30_58),.data_out(wire_d30_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313060(.data_in(wire_d30_59),.data_out(wire_d30_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313061(.data_in(wire_d30_60),.data_out(wire_d30_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313062(.data_in(wire_d30_61),.data_out(wire_d30_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313063(.data_in(wire_d30_62),.data_out(wire_d30_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313064(.data_in(wire_d30_63),.data_out(wire_d30_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313065(.data_in(wire_d30_64),.data_out(wire_d30_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313066(.data_in(wire_d30_65),.data_out(wire_d30_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313067(.data_in(wire_d30_66),.data_out(wire_d30_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313068(.data_in(wire_d30_67),.data_out(wire_d30_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313069(.data_in(wire_d30_68),.data_out(wire_d30_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313070(.data_in(wire_d30_69),.data_out(wire_d30_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313071(.data_in(wire_d30_70),.data_out(wire_d30_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313072(.data_in(wire_d30_71),.data_out(wire_d30_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313073(.data_in(wire_d30_72),.data_out(wire_d30_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313074(.data_in(wire_d30_73),.data_out(wire_d30_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313075(.data_in(wire_d30_74),.data_out(wire_d30_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313076(.data_in(wire_d30_75),.data_out(wire_d30_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313077(.data_in(wire_d30_76),.data_out(wire_d30_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313078(.data_in(wire_d30_77),.data_out(wire_d30_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313079(.data_in(wire_d30_78),.data_out(wire_d30_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313080(.data_in(wire_d30_79),.data_out(wire_d30_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313081(.data_in(wire_d30_80),.data_out(wire_d30_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313082(.data_in(wire_d30_81),.data_out(wire_d30_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313083(.data_in(wire_d30_82),.data_out(wire_d30_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313084(.data_in(wire_d30_83),.data_out(wire_d30_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313085(.data_in(wire_d30_84),.data_out(wire_d30_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313086(.data_in(wire_d30_85),.data_out(wire_d30_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313087(.data_in(wire_d30_86),.data_out(wire_d30_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313088(.data_in(wire_d30_87),.data_out(wire_d30_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313089(.data_in(wire_d30_88),.data_out(wire_d30_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313090(.data_in(wire_d30_89),.data_out(wire_d30_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313091(.data_in(wire_d30_90),.data_out(wire_d30_91),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313092(.data_in(wire_d30_91),.data_out(wire_d30_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313093(.data_in(wire_d30_92),.data_out(wire_d30_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313094(.data_in(wire_d30_93),.data_out(wire_d30_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313095(.data_in(wire_d30_94),.data_out(wire_d30_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313096(.data_in(wire_d30_95),.data_out(wire_d30_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313097(.data_in(wire_d30_96),.data_out(wire_d30_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313098(.data_in(wire_d30_97),.data_out(wire_d30_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313099(.data_in(wire_d30_98),.data_out(d_out30),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance32310(.data_in(d_in31),.data_out(wire_d31_0),.clk(clk),.rst(rst));            //channel 32
	large_mux #(.WIDTH(WIDTH)) large_mux_instance32311(.data_in(wire_d31_0),.data_out(wire_d31_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance32312(.data_in(wire_d31_1),.data_out(wire_d31_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance32313(.data_in(wire_d31_2),.data_out(wire_d31_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance32314(.data_in(wire_d31_3),.data_out(wire_d31_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance32315(.data_in(wire_d31_4),.data_out(wire_d31_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance32316(.data_in(wire_d31_5),.data_out(wire_d31_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance32317(.data_in(wire_d31_6),.data_out(wire_d31_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance32318(.data_in(wire_d31_7),.data_out(wire_d31_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32319(.data_in(wire_d31_8),.data_out(wire_d31_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323110(.data_in(wire_d31_9),.data_out(wire_d31_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323111(.data_in(wire_d31_10),.data_out(wire_d31_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323112(.data_in(wire_d31_11),.data_out(wire_d31_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323113(.data_in(wire_d31_12),.data_out(wire_d31_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323114(.data_in(wire_d31_13),.data_out(wire_d31_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323115(.data_in(wire_d31_14),.data_out(wire_d31_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323116(.data_in(wire_d31_15),.data_out(wire_d31_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323117(.data_in(wire_d31_16),.data_out(wire_d31_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323118(.data_in(wire_d31_17),.data_out(wire_d31_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323119(.data_in(wire_d31_18),.data_out(wire_d31_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323120(.data_in(wire_d31_19),.data_out(wire_d31_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323121(.data_in(wire_d31_20),.data_out(wire_d31_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323122(.data_in(wire_d31_21),.data_out(wire_d31_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323123(.data_in(wire_d31_22),.data_out(wire_d31_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323124(.data_in(wire_d31_23),.data_out(wire_d31_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323125(.data_in(wire_d31_24),.data_out(wire_d31_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323126(.data_in(wire_d31_25),.data_out(wire_d31_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323127(.data_in(wire_d31_26),.data_out(wire_d31_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323128(.data_in(wire_d31_27),.data_out(wire_d31_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323129(.data_in(wire_d31_28),.data_out(wire_d31_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323130(.data_in(wire_d31_29),.data_out(wire_d31_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323131(.data_in(wire_d31_30),.data_out(wire_d31_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323132(.data_in(wire_d31_31),.data_out(wire_d31_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323133(.data_in(wire_d31_32),.data_out(wire_d31_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323134(.data_in(wire_d31_33),.data_out(wire_d31_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323135(.data_in(wire_d31_34),.data_out(wire_d31_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323136(.data_in(wire_d31_35),.data_out(wire_d31_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323137(.data_in(wire_d31_36),.data_out(wire_d31_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323138(.data_in(wire_d31_37),.data_out(wire_d31_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323139(.data_in(wire_d31_38),.data_out(wire_d31_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323140(.data_in(wire_d31_39),.data_out(wire_d31_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323141(.data_in(wire_d31_40),.data_out(wire_d31_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323142(.data_in(wire_d31_41),.data_out(wire_d31_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323143(.data_in(wire_d31_42),.data_out(wire_d31_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323144(.data_in(wire_d31_43),.data_out(wire_d31_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323145(.data_in(wire_d31_44),.data_out(wire_d31_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323146(.data_in(wire_d31_45),.data_out(wire_d31_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323147(.data_in(wire_d31_46),.data_out(wire_d31_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323148(.data_in(wire_d31_47),.data_out(wire_d31_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323149(.data_in(wire_d31_48),.data_out(wire_d31_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323150(.data_in(wire_d31_49),.data_out(wire_d31_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323151(.data_in(wire_d31_50),.data_out(wire_d31_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323152(.data_in(wire_d31_51),.data_out(wire_d31_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323153(.data_in(wire_d31_52),.data_out(wire_d31_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323154(.data_in(wire_d31_53),.data_out(wire_d31_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323155(.data_in(wire_d31_54),.data_out(wire_d31_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323156(.data_in(wire_d31_55),.data_out(wire_d31_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323157(.data_in(wire_d31_56),.data_out(wire_d31_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323158(.data_in(wire_d31_57),.data_out(wire_d31_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323159(.data_in(wire_d31_58),.data_out(wire_d31_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323160(.data_in(wire_d31_59),.data_out(wire_d31_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323161(.data_in(wire_d31_60),.data_out(wire_d31_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323162(.data_in(wire_d31_61),.data_out(wire_d31_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323163(.data_in(wire_d31_62),.data_out(wire_d31_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323164(.data_in(wire_d31_63),.data_out(wire_d31_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323165(.data_in(wire_d31_64),.data_out(wire_d31_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323166(.data_in(wire_d31_65),.data_out(wire_d31_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323167(.data_in(wire_d31_66),.data_out(wire_d31_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323168(.data_in(wire_d31_67),.data_out(wire_d31_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323169(.data_in(wire_d31_68),.data_out(wire_d31_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323170(.data_in(wire_d31_69),.data_out(wire_d31_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323171(.data_in(wire_d31_70),.data_out(wire_d31_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323172(.data_in(wire_d31_71),.data_out(wire_d31_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323173(.data_in(wire_d31_72),.data_out(wire_d31_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323174(.data_in(wire_d31_73),.data_out(wire_d31_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323175(.data_in(wire_d31_74),.data_out(wire_d31_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323176(.data_in(wire_d31_75),.data_out(wire_d31_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323177(.data_in(wire_d31_76),.data_out(wire_d31_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323178(.data_in(wire_d31_77),.data_out(wire_d31_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323179(.data_in(wire_d31_78),.data_out(wire_d31_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323180(.data_in(wire_d31_79),.data_out(wire_d31_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323181(.data_in(wire_d31_80),.data_out(wire_d31_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323182(.data_in(wire_d31_81),.data_out(wire_d31_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323183(.data_in(wire_d31_82),.data_out(wire_d31_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323184(.data_in(wire_d31_83),.data_out(wire_d31_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323185(.data_in(wire_d31_84),.data_out(wire_d31_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323186(.data_in(wire_d31_85),.data_out(wire_d31_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323187(.data_in(wire_d31_86),.data_out(wire_d31_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323188(.data_in(wire_d31_87),.data_out(wire_d31_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323189(.data_in(wire_d31_88),.data_out(wire_d31_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323190(.data_in(wire_d31_89),.data_out(wire_d31_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323191(.data_in(wire_d31_90),.data_out(wire_d31_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323192(.data_in(wire_d31_91),.data_out(wire_d31_92),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323193(.data_in(wire_d31_92),.data_out(wire_d31_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323194(.data_in(wire_d31_93),.data_out(wire_d31_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323195(.data_in(wire_d31_94),.data_out(wire_d31_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323196(.data_in(wire_d31_95),.data_out(wire_d31_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323197(.data_in(wire_d31_96),.data_out(wire_d31_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323198(.data_in(wire_d31_97),.data_out(wire_d31_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323199(.data_in(wire_d31_98),.data_out(d_out31),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance33320(.data_in(d_in32),.data_out(wire_d32_0),.clk(clk),.rst(rst));            //channel 33
	encoder #(.WIDTH(WIDTH)) encoder_instance33321(.data_in(wire_d32_0),.data_out(wire_d32_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance33322(.data_in(wire_d32_1),.data_out(wire_d32_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance33323(.data_in(wire_d32_2),.data_out(wire_d32_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance33324(.data_in(wire_d32_3),.data_out(wire_d32_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance33325(.data_in(wire_d32_4),.data_out(wire_d32_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance33326(.data_in(wire_d32_5),.data_out(wire_d32_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance33327(.data_in(wire_d32_6),.data_out(wire_d32_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance33328(.data_in(wire_d32_7),.data_out(wire_d32_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance33329(.data_in(wire_d32_8),.data_out(wire_d32_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333210(.data_in(wire_d32_9),.data_out(wire_d32_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333211(.data_in(wire_d32_10),.data_out(wire_d32_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333212(.data_in(wire_d32_11),.data_out(wire_d32_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333213(.data_in(wire_d32_12),.data_out(wire_d32_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333214(.data_in(wire_d32_13),.data_out(wire_d32_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333215(.data_in(wire_d32_14),.data_out(wire_d32_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333216(.data_in(wire_d32_15),.data_out(wire_d32_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333217(.data_in(wire_d32_16),.data_out(wire_d32_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333218(.data_in(wire_d32_17),.data_out(wire_d32_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333219(.data_in(wire_d32_18),.data_out(wire_d32_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333220(.data_in(wire_d32_19),.data_out(wire_d32_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333221(.data_in(wire_d32_20),.data_out(wire_d32_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333222(.data_in(wire_d32_21),.data_out(wire_d32_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333223(.data_in(wire_d32_22),.data_out(wire_d32_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333224(.data_in(wire_d32_23),.data_out(wire_d32_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333225(.data_in(wire_d32_24),.data_out(wire_d32_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333226(.data_in(wire_d32_25),.data_out(wire_d32_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333227(.data_in(wire_d32_26),.data_out(wire_d32_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333228(.data_in(wire_d32_27),.data_out(wire_d32_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333229(.data_in(wire_d32_28),.data_out(wire_d32_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333230(.data_in(wire_d32_29),.data_out(wire_d32_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333231(.data_in(wire_d32_30),.data_out(wire_d32_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333232(.data_in(wire_d32_31),.data_out(wire_d32_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333233(.data_in(wire_d32_32),.data_out(wire_d32_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333234(.data_in(wire_d32_33),.data_out(wire_d32_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333235(.data_in(wire_d32_34),.data_out(wire_d32_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333236(.data_in(wire_d32_35),.data_out(wire_d32_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333237(.data_in(wire_d32_36),.data_out(wire_d32_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333238(.data_in(wire_d32_37),.data_out(wire_d32_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333239(.data_in(wire_d32_38),.data_out(wire_d32_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333240(.data_in(wire_d32_39),.data_out(wire_d32_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333241(.data_in(wire_d32_40),.data_out(wire_d32_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333242(.data_in(wire_d32_41),.data_out(wire_d32_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333243(.data_in(wire_d32_42),.data_out(wire_d32_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333244(.data_in(wire_d32_43),.data_out(wire_d32_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333245(.data_in(wire_d32_44),.data_out(wire_d32_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333246(.data_in(wire_d32_45),.data_out(wire_d32_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333247(.data_in(wire_d32_46),.data_out(wire_d32_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333248(.data_in(wire_d32_47),.data_out(wire_d32_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333249(.data_in(wire_d32_48),.data_out(wire_d32_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333250(.data_in(wire_d32_49),.data_out(wire_d32_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333251(.data_in(wire_d32_50),.data_out(wire_d32_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333252(.data_in(wire_d32_51),.data_out(wire_d32_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333253(.data_in(wire_d32_52),.data_out(wire_d32_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333254(.data_in(wire_d32_53),.data_out(wire_d32_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333255(.data_in(wire_d32_54),.data_out(wire_d32_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333256(.data_in(wire_d32_55),.data_out(wire_d32_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333257(.data_in(wire_d32_56),.data_out(wire_d32_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333258(.data_in(wire_d32_57),.data_out(wire_d32_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333259(.data_in(wire_d32_58),.data_out(wire_d32_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333260(.data_in(wire_d32_59),.data_out(wire_d32_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333261(.data_in(wire_d32_60),.data_out(wire_d32_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333262(.data_in(wire_d32_61),.data_out(wire_d32_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333263(.data_in(wire_d32_62),.data_out(wire_d32_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333264(.data_in(wire_d32_63),.data_out(wire_d32_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333265(.data_in(wire_d32_64),.data_out(wire_d32_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333266(.data_in(wire_d32_65),.data_out(wire_d32_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333267(.data_in(wire_d32_66),.data_out(wire_d32_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333268(.data_in(wire_d32_67),.data_out(wire_d32_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333269(.data_in(wire_d32_68),.data_out(wire_d32_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333270(.data_in(wire_d32_69),.data_out(wire_d32_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333271(.data_in(wire_d32_70),.data_out(wire_d32_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333272(.data_in(wire_d32_71),.data_out(wire_d32_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333273(.data_in(wire_d32_72),.data_out(wire_d32_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333274(.data_in(wire_d32_73),.data_out(wire_d32_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333275(.data_in(wire_d32_74),.data_out(wire_d32_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333276(.data_in(wire_d32_75),.data_out(wire_d32_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333277(.data_in(wire_d32_76),.data_out(wire_d32_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333278(.data_in(wire_d32_77),.data_out(wire_d32_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333279(.data_in(wire_d32_78),.data_out(wire_d32_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333280(.data_in(wire_d32_79),.data_out(wire_d32_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333281(.data_in(wire_d32_80),.data_out(wire_d32_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333282(.data_in(wire_d32_81),.data_out(wire_d32_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333283(.data_in(wire_d32_82),.data_out(wire_d32_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333284(.data_in(wire_d32_83),.data_out(wire_d32_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333285(.data_in(wire_d32_84),.data_out(wire_d32_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333286(.data_in(wire_d32_85),.data_out(wire_d32_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333287(.data_in(wire_d32_86),.data_out(wire_d32_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333288(.data_in(wire_d32_87),.data_out(wire_d32_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333289(.data_in(wire_d32_88),.data_out(wire_d32_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333290(.data_in(wire_d32_89),.data_out(wire_d32_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333291(.data_in(wire_d32_90),.data_out(wire_d32_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333292(.data_in(wire_d32_91),.data_out(wire_d32_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333293(.data_in(wire_d32_92),.data_out(wire_d32_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333294(.data_in(wire_d32_93),.data_out(wire_d32_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333295(.data_in(wire_d32_94),.data_out(wire_d32_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333296(.data_in(wire_d32_95),.data_out(wire_d32_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333297(.data_in(wire_d32_96),.data_out(wire_d32_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333298(.data_in(wire_d32_97),.data_out(wire_d32_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333299(.data_in(wire_d32_98),.data_out(d_out32),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance34330(.data_in(d_in33),.data_out(wire_d33_0),.clk(clk),.rst(rst));            //channel 34
	encoder #(.WIDTH(WIDTH)) encoder_instance34331(.data_in(wire_d33_0),.data_out(wire_d33_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance34332(.data_in(wire_d33_1),.data_out(wire_d33_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance34333(.data_in(wire_d33_2),.data_out(wire_d33_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance34334(.data_in(wire_d33_3),.data_out(wire_d33_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance34335(.data_in(wire_d33_4),.data_out(wire_d33_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance34336(.data_in(wire_d33_5),.data_out(wire_d33_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance34337(.data_in(wire_d33_6),.data_out(wire_d33_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance34338(.data_in(wire_d33_7),.data_out(wire_d33_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance34339(.data_in(wire_d33_8),.data_out(wire_d33_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343310(.data_in(wire_d33_9),.data_out(wire_d33_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343311(.data_in(wire_d33_10),.data_out(wire_d33_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343312(.data_in(wire_d33_11),.data_out(wire_d33_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343313(.data_in(wire_d33_12),.data_out(wire_d33_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343314(.data_in(wire_d33_13),.data_out(wire_d33_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343315(.data_in(wire_d33_14),.data_out(wire_d33_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343316(.data_in(wire_d33_15),.data_out(wire_d33_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343317(.data_in(wire_d33_16),.data_out(wire_d33_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343318(.data_in(wire_d33_17),.data_out(wire_d33_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343319(.data_in(wire_d33_18),.data_out(wire_d33_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343320(.data_in(wire_d33_19),.data_out(wire_d33_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343321(.data_in(wire_d33_20),.data_out(wire_d33_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343322(.data_in(wire_d33_21),.data_out(wire_d33_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343323(.data_in(wire_d33_22),.data_out(wire_d33_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343324(.data_in(wire_d33_23),.data_out(wire_d33_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343325(.data_in(wire_d33_24),.data_out(wire_d33_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343326(.data_in(wire_d33_25),.data_out(wire_d33_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343327(.data_in(wire_d33_26),.data_out(wire_d33_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343328(.data_in(wire_d33_27),.data_out(wire_d33_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343329(.data_in(wire_d33_28),.data_out(wire_d33_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343330(.data_in(wire_d33_29),.data_out(wire_d33_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343331(.data_in(wire_d33_30),.data_out(wire_d33_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343332(.data_in(wire_d33_31),.data_out(wire_d33_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343333(.data_in(wire_d33_32),.data_out(wire_d33_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343334(.data_in(wire_d33_33),.data_out(wire_d33_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343335(.data_in(wire_d33_34),.data_out(wire_d33_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343336(.data_in(wire_d33_35),.data_out(wire_d33_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343337(.data_in(wire_d33_36),.data_out(wire_d33_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343338(.data_in(wire_d33_37),.data_out(wire_d33_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343339(.data_in(wire_d33_38),.data_out(wire_d33_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343340(.data_in(wire_d33_39),.data_out(wire_d33_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343341(.data_in(wire_d33_40),.data_out(wire_d33_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343342(.data_in(wire_d33_41),.data_out(wire_d33_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343343(.data_in(wire_d33_42),.data_out(wire_d33_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343344(.data_in(wire_d33_43),.data_out(wire_d33_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343345(.data_in(wire_d33_44),.data_out(wire_d33_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343346(.data_in(wire_d33_45),.data_out(wire_d33_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343347(.data_in(wire_d33_46),.data_out(wire_d33_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343348(.data_in(wire_d33_47),.data_out(wire_d33_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343349(.data_in(wire_d33_48),.data_out(wire_d33_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343350(.data_in(wire_d33_49),.data_out(wire_d33_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343351(.data_in(wire_d33_50),.data_out(wire_d33_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343352(.data_in(wire_d33_51),.data_out(wire_d33_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343353(.data_in(wire_d33_52),.data_out(wire_d33_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343354(.data_in(wire_d33_53),.data_out(wire_d33_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343355(.data_in(wire_d33_54),.data_out(wire_d33_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343356(.data_in(wire_d33_55),.data_out(wire_d33_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343357(.data_in(wire_d33_56),.data_out(wire_d33_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343358(.data_in(wire_d33_57),.data_out(wire_d33_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343359(.data_in(wire_d33_58),.data_out(wire_d33_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343360(.data_in(wire_d33_59),.data_out(wire_d33_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343361(.data_in(wire_d33_60),.data_out(wire_d33_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343362(.data_in(wire_d33_61),.data_out(wire_d33_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343363(.data_in(wire_d33_62),.data_out(wire_d33_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343364(.data_in(wire_d33_63),.data_out(wire_d33_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343365(.data_in(wire_d33_64),.data_out(wire_d33_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343366(.data_in(wire_d33_65),.data_out(wire_d33_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343367(.data_in(wire_d33_66),.data_out(wire_d33_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343368(.data_in(wire_d33_67),.data_out(wire_d33_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343369(.data_in(wire_d33_68),.data_out(wire_d33_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343370(.data_in(wire_d33_69),.data_out(wire_d33_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343371(.data_in(wire_d33_70),.data_out(wire_d33_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343372(.data_in(wire_d33_71),.data_out(wire_d33_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343373(.data_in(wire_d33_72),.data_out(wire_d33_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343374(.data_in(wire_d33_73),.data_out(wire_d33_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343375(.data_in(wire_d33_74),.data_out(wire_d33_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343376(.data_in(wire_d33_75),.data_out(wire_d33_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343377(.data_in(wire_d33_76),.data_out(wire_d33_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343378(.data_in(wire_d33_77),.data_out(wire_d33_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343379(.data_in(wire_d33_78),.data_out(wire_d33_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343380(.data_in(wire_d33_79),.data_out(wire_d33_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343381(.data_in(wire_d33_80),.data_out(wire_d33_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343382(.data_in(wire_d33_81),.data_out(wire_d33_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343383(.data_in(wire_d33_82),.data_out(wire_d33_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343384(.data_in(wire_d33_83),.data_out(wire_d33_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343385(.data_in(wire_d33_84),.data_out(wire_d33_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343386(.data_in(wire_d33_85),.data_out(wire_d33_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343387(.data_in(wire_d33_86),.data_out(wire_d33_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343388(.data_in(wire_d33_87),.data_out(wire_d33_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343389(.data_in(wire_d33_88),.data_out(wire_d33_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343390(.data_in(wire_d33_89),.data_out(wire_d33_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343391(.data_in(wire_d33_90),.data_out(wire_d33_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343392(.data_in(wire_d33_91),.data_out(wire_d33_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343393(.data_in(wire_d33_92),.data_out(wire_d33_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343394(.data_in(wire_d33_93),.data_out(wire_d33_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343395(.data_in(wire_d33_94),.data_out(wire_d33_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343396(.data_in(wire_d33_95),.data_out(wire_d33_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343397(.data_in(wire_d33_96),.data_out(wire_d33_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343398(.data_in(wire_d33_97),.data_out(wire_d33_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343399(.data_in(wire_d33_98),.data_out(d_out33),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance35340(.data_in(d_in34),.data_out(wire_d34_0),.clk(clk),.rst(rst));            //channel 35
	large_mux #(.WIDTH(WIDTH)) large_mux_instance35341(.data_in(wire_d34_0),.data_out(wire_d34_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance35342(.data_in(wire_d34_1),.data_out(wire_d34_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance35343(.data_in(wire_d34_2),.data_out(wire_d34_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance35344(.data_in(wire_d34_3),.data_out(wire_d34_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance35345(.data_in(wire_d34_4),.data_out(wire_d34_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance35346(.data_in(wire_d34_5),.data_out(wire_d34_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance35347(.data_in(wire_d34_6),.data_out(wire_d34_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance35348(.data_in(wire_d34_7),.data_out(wire_d34_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance35349(.data_in(wire_d34_8),.data_out(wire_d34_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353410(.data_in(wire_d34_9),.data_out(wire_d34_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353411(.data_in(wire_d34_10),.data_out(wire_d34_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353412(.data_in(wire_d34_11),.data_out(wire_d34_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353413(.data_in(wire_d34_12),.data_out(wire_d34_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353414(.data_in(wire_d34_13),.data_out(wire_d34_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353415(.data_in(wire_d34_14),.data_out(wire_d34_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353416(.data_in(wire_d34_15),.data_out(wire_d34_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353417(.data_in(wire_d34_16),.data_out(wire_d34_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353418(.data_in(wire_d34_17),.data_out(wire_d34_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353419(.data_in(wire_d34_18),.data_out(wire_d34_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353420(.data_in(wire_d34_19),.data_out(wire_d34_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353421(.data_in(wire_d34_20),.data_out(wire_d34_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353422(.data_in(wire_d34_21),.data_out(wire_d34_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353423(.data_in(wire_d34_22),.data_out(wire_d34_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353424(.data_in(wire_d34_23),.data_out(wire_d34_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353425(.data_in(wire_d34_24),.data_out(wire_d34_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353426(.data_in(wire_d34_25),.data_out(wire_d34_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353427(.data_in(wire_d34_26),.data_out(wire_d34_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353428(.data_in(wire_d34_27),.data_out(wire_d34_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353429(.data_in(wire_d34_28),.data_out(wire_d34_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353430(.data_in(wire_d34_29),.data_out(wire_d34_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353431(.data_in(wire_d34_30),.data_out(wire_d34_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353432(.data_in(wire_d34_31),.data_out(wire_d34_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353433(.data_in(wire_d34_32),.data_out(wire_d34_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353434(.data_in(wire_d34_33),.data_out(wire_d34_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353435(.data_in(wire_d34_34),.data_out(wire_d34_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353436(.data_in(wire_d34_35),.data_out(wire_d34_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353437(.data_in(wire_d34_36),.data_out(wire_d34_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353438(.data_in(wire_d34_37),.data_out(wire_d34_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353439(.data_in(wire_d34_38),.data_out(wire_d34_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353440(.data_in(wire_d34_39),.data_out(wire_d34_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353441(.data_in(wire_d34_40),.data_out(wire_d34_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353442(.data_in(wire_d34_41),.data_out(wire_d34_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353443(.data_in(wire_d34_42),.data_out(wire_d34_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353444(.data_in(wire_d34_43),.data_out(wire_d34_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353445(.data_in(wire_d34_44),.data_out(wire_d34_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353446(.data_in(wire_d34_45),.data_out(wire_d34_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353447(.data_in(wire_d34_46),.data_out(wire_d34_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353448(.data_in(wire_d34_47),.data_out(wire_d34_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353449(.data_in(wire_d34_48),.data_out(wire_d34_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353450(.data_in(wire_d34_49),.data_out(wire_d34_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353451(.data_in(wire_d34_50),.data_out(wire_d34_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353452(.data_in(wire_d34_51),.data_out(wire_d34_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353453(.data_in(wire_d34_52),.data_out(wire_d34_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353454(.data_in(wire_d34_53),.data_out(wire_d34_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353455(.data_in(wire_d34_54),.data_out(wire_d34_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353456(.data_in(wire_d34_55),.data_out(wire_d34_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353457(.data_in(wire_d34_56),.data_out(wire_d34_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353458(.data_in(wire_d34_57),.data_out(wire_d34_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353459(.data_in(wire_d34_58),.data_out(wire_d34_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353460(.data_in(wire_d34_59),.data_out(wire_d34_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353461(.data_in(wire_d34_60),.data_out(wire_d34_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353462(.data_in(wire_d34_61),.data_out(wire_d34_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353463(.data_in(wire_d34_62),.data_out(wire_d34_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353464(.data_in(wire_d34_63),.data_out(wire_d34_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353465(.data_in(wire_d34_64),.data_out(wire_d34_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353466(.data_in(wire_d34_65),.data_out(wire_d34_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353467(.data_in(wire_d34_66),.data_out(wire_d34_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353468(.data_in(wire_d34_67),.data_out(wire_d34_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353469(.data_in(wire_d34_68),.data_out(wire_d34_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353470(.data_in(wire_d34_69),.data_out(wire_d34_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353471(.data_in(wire_d34_70),.data_out(wire_d34_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353472(.data_in(wire_d34_71),.data_out(wire_d34_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353473(.data_in(wire_d34_72),.data_out(wire_d34_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353474(.data_in(wire_d34_73),.data_out(wire_d34_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353475(.data_in(wire_d34_74),.data_out(wire_d34_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353476(.data_in(wire_d34_75),.data_out(wire_d34_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353477(.data_in(wire_d34_76),.data_out(wire_d34_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353478(.data_in(wire_d34_77),.data_out(wire_d34_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353479(.data_in(wire_d34_78),.data_out(wire_d34_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353480(.data_in(wire_d34_79),.data_out(wire_d34_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353481(.data_in(wire_d34_80),.data_out(wire_d34_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353482(.data_in(wire_d34_81),.data_out(wire_d34_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353483(.data_in(wire_d34_82),.data_out(wire_d34_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353484(.data_in(wire_d34_83),.data_out(wire_d34_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353485(.data_in(wire_d34_84),.data_out(wire_d34_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353486(.data_in(wire_d34_85),.data_out(wire_d34_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353487(.data_in(wire_d34_86),.data_out(wire_d34_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353488(.data_in(wire_d34_87),.data_out(wire_d34_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353489(.data_in(wire_d34_88),.data_out(wire_d34_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353490(.data_in(wire_d34_89),.data_out(wire_d34_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353491(.data_in(wire_d34_90),.data_out(wire_d34_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353492(.data_in(wire_d34_91),.data_out(wire_d34_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353493(.data_in(wire_d34_92),.data_out(wire_d34_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353494(.data_in(wire_d34_93),.data_out(wire_d34_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353495(.data_in(wire_d34_94),.data_out(wire_d34_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353496(.data_in(wire_d34_95),.data_out(wire_d34_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353497(.data_in(wire_d34_96),.data_out(wire_d34_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353498(.data_in(wire_d34_97),.data_out(wire_d34_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353499(.data_in(wire_d34_98),.data_out(d_out34),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance36350(.data_in(d_in35),.data_out(wire_d35_0),.clk(clk),.rst(rst));            //channel 36
	invertion #(.WIDTH(WIDTH)) invertion_instance36351(.data_in(wire_d35_0),.data_out(wire_d35_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance36352(.data_in(wire_d35_1),.data_out(wire_d35_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance36353(.data_in(wire_d35_2),.data_out(wire_d35_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance36354(.data_in(wire_d35_3),.data_out(wire_d35_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance36355(.data_in(wire_d35_4),.data_out(wire_d35_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance36356(.data_in(wire_d35_5),.data_out(wire_d35_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance36357(.data_in(wire_d35_6),.data_out(wire_d35_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance36358(.data_in(wire_d35_7),.data_out(wire_d35_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance36359(.data_in(wire_d35_8),.data_out(wire_d35_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363510(.data_in(wire_d35_9),.data_out(wire_d35_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363511(.data_in(wire_d35_10),.data_out(wire_d35_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363512(.data_in(wire_d35_11),.data_out(wire_d35_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363513(.data_in(wire_d35_12),.data_out(wire_d35_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363514(.data_in(wire_d35_13),.data_out(wire_d35_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363515(.data_in(wire_d35_14),.data_out(wire_d35_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363516(.data_in(wire_d35_15),.data_out(wire_d35_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363517(.data_in(wire_d35_16),.data_out(wire_d35_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363518(.data_in(wire_d35_17),.data_out(wire_d35_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363519(.data_in(wire_d35_18),.data_out(wire_d35_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363520(.data_in(wire_d35_19),.data_out(wire_d35_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363521(.data_in(wire_d35_20),.data_out(wire_d35_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363522(.data_in(wire_d35_21),.data_out(wire_d35_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363523(.data_in(wire_d35_22),.data_out(wire_d35_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363524(.data_in(wire_d35_23),.data_out(wire_d35_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363525(.data_in(wire_d35_24),.data_out(wire_d35_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363526(.data_in(wire_d35_25),.data_out(wire_d35_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363527(.data_in(wire_d35_26),.data_out(wire_d35_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363528(.data_in(wire_d35_27),.data_out(wire_d35_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363529(.data_in(wire_d35_28),.data_out(wire_d35_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363530(.data_in(wire_d35_29),.data_out(wire_d35_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363531(.data_in(wire_d35_30),.data_out(wire_d35_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363532(.data_in(wire_d35_31),.data_out(wire_d35_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363533(.data_in(wire_d35_32),.data_out(wire_d35_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363534(.data_in(wire_d35_33),.data_out(wire_d35_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363535(.data_in(wire_d35_34),.data_out(wire_d35_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363536(.data_in(wire_d35_35),.data_out(wire_d35_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363537(.data_in(wire_d35_36),.data_out(wire_d35_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363538(.data_in(wire_d35_37),.data_out(wire_d35_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363539(.data_in(wire_d35_38),.data_out(wire_d35_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363540(.data_in(wire_d35_39),.data_out(wire_d35_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363541(.data_in(wire_d35_40),.data_out(wire_d35_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363542(.data_in(wire_d35_41),.data_out(wire_d35_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363543(.data_in(wire_d35_42),.data_out(wire_d35_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363544(.data_in(wire_d35_43),.data_out(wire_d35_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363545(.data_in(wire_d35_44),.data_out(wire_d35_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363546(.data_in(wire_d35_45),.data_out(wire_d35_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363547(.data_in(wire_d35_46),.data_out(wire_d35_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363548(.data_in(wire_d35_47),.data_out(wire_d35_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363549(.data_in(wire_d35_48),.data_out(wire_d35_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363550(.data_in(wire_d35_49),.data_out(wire_d35_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363551(.data_in(wire_d35_50),.data_out(wire_d35_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363552(.data_in(wire_d35_51),.data_out(wire_d35_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363553(.data_in(wire_d35_52),.data_out(wire_d35_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363554(.data_in(wire_d35_53),.data_out(wire_d35_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363555(.data_in(wire_d35_54),.data_out(wire_d35_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363556(.data_in(wire_d35_55),.data_out(wire_d35_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363557(.data_in(wire_d35_56),.data_out(wire_d35_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363558(.data_in(wire_d35_57),.data_out(wire_d35_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363559(.data_in(wire_d35_58),.data_out(wire_d35_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363560(.data_in(wire_d35_59),.data_out(wire_d35_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363561(.data_in(wire_d35_60),.data_out(wire_d35_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363562(.data_in(wire_d35_61),.data_out(wire_d35_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363563(.data_in(wire_d35_62),.data_out(wire_d35_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363564(.data_in(wire_d35_63),.data_out(wire_d35_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363565(.data_in(wire_d35_64),.data_out(wire_d35_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363566(.data_in(wire_d35_65),.data_out(wire_d35_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363567(.data_in(wire_d35_66),.data_out(wire_d35_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363568(.data_in(wire_d35_67),.data_out(wire_d35_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363569(.data_in(wire_d35_68),.data_out(wire_d35_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363570(.data_in(wire_d35_69),.data_out(wire_d35_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363571(.data_in(wire_d35_70),.data_out(wire_d35_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363572(.data_in(wire_d35_71),.data_out(wire_d35_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363573(.data_in(wire_d35_72),.data_out(wire_d35_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363574(.data_in(wire_d35_73),.data_out(wire_d35_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363575(.data_in(wire_d35_74),.data_out(wire_d35_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363576(.data_in(wire_d35_75),.data_out(wire_d35_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363577(.data_in(wire_d35_76),.data_out(wire_d35_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363578(.data_in(wire_d35_77),.data_out(wire_d35_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363579(.data_in(wire_d35_78),.data_out(wire_d35_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363580(.data_in(wire_d35_79),.data_out(wire_d35_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363581(.data_in(wire_d35_80),.data_out(wire_d35_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363582(.data_in(wire_d35_81),.data_out(wire_d35_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363583(.data_in(wire_d35_82),.data_out(wire_d35_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363584(.data_in(wire_d35_83),.data_out(wire_d35_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363585(.data_in(wire_d35_84),.data_out(wire_d35_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363586(.data_in(wire_d35_85),.data_out(wire_d35_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363587(.data_in(wire_d35_86),.data_out(wire_d35_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363588(.data_in(wire_d35_87),.data_out(wire_d35_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363589(.data_in(wire_d35_88),.data_out(wire_d35_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363590(.data_in(wire_d35_89),.data_out(wire_d35_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363591(.data_in(wire_d35_90),.data_out(wire_d35_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363592(.data_in(wire_d35_91),.data_out(wire_d35_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363593(.data_in(wire_d35_92),.data_out(wire_d35_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363594(.data_in(wire_d35_93),.data_out(wire_d35_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363595(.data_in(wire_d35_94),.data_out(wire_d35_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363596(.data_in(wire_d35_95),.data_out(wire_d35_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363597(.data_in(wire_d35_96),.data_out(wire_d35_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363598(.data_in(wire_d35_97),.data_out(wire_d35_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363599(.data_in(wire_d35_98),.data_out(d_out35),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance37360(.data_in(d_in36),.data_out(wire_d36_0),.clk(clk),.rst(rst));            //channel 37
	register #(.WIDTH(WIDTH)) register_instance37361(.data_in(wire_d36_0),.data_out(wire_d36_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance37362(.data_in(wire_d36_1),.data_out(wire_d36_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance37363(.data_in(wire_d36_2),.data_out(wire_d36_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance37364(.data_in(wire_d36_3),.data_out(wire_d36_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance37365(.data_in(wire_d36_4),.data_out(wire_d36_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance37366(.data_in(wire_d36_5),.data_out(wire_d36_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance37367(.data_in(wire_d36_6),.data_out(wire_d36_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance37368(.data_in(wire_d36_7),.data_out(wire_d36_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance37369(.data_in(wire_d36_8),.data_out(wire_d36_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373610(.data_in(wire_d36_9),.data_out(wire_d36_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373611(.data_in(wire_d36_10),.data_out(wire_d36_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373612(.data_in(wire_d36_11),.data_out(wire_d36_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373613(.data_in(wire_d36_12),.data_out(wire_d36_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373614(.data_in(wire_d36_13),.data_out(wire_d36_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373615(.data_in(wire_d36_14),.data_out(wire_d36_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373616(.data_in(wire_d36_15),.data_out(wire_d36_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373617(.data_in(wire_d36_16),.data_out(wire_d36_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373618(.data_in(wire_d36_17),.data_out(wire_d36_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373619(.data_in(wire_d36_18),.data_out(wire_d36_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373620(.data_in(wire_d36_19),.data_out(wire_d36_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373621(.data_in(wire_d36_20),.data_out(wire_d36_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373622(.data_in(wire_d36_21),.data_out(wire_d36_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373623(.data_in(wire_d36_22),.data_out(wire_d36_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373624(.data_in(wire_d36_23),.data_out(wire_d36_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373625(.data_in(wire_d36_24),.data_out(wire_d36_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373626(.data_in(wire_d36_25),.data_out(wire_d36_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373627(.data_in(wire_d36_26),.data_out(wire_d36_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373628(.data_in(wire_d36_27),.data_out(wire_d36_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373629(.data_in(wire_d36_28),.data_out(wire_d36_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373630(.data_in(wire_d36_29),.data_out(wire_d36_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373631(.data_in(wire_d36_30),.data_out(wire_d36_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373632(.data_in(wire_d36_31),.data_out(wire_d36_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373633(.data_in(wire_d36_32),.data_out(wire_d36_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373634(.data_in(wire_d36_33),.data_out(wire_d36_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373635(.data_in(wire_d36_34),.data_out(wire_d36_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373636(.data_in(wire_d36_35),.data_out(wire_d36_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373637(.data_in(wire_d36_36),.data_out(wire_d36_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373638(.data_in(wire_d36_37),.data_out(wire_d36_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373639(.data_in(wire_d36_38),.data_out(wire_d36_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373640(.data_in(wire_d36_39),.data_out(wire_d36_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373641(.data_in(wire_d36_40),.data_out(wire_d36_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373642(.data_in(wire_d36_41),.data_out(wire_d36_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373643(.data_in(wire_d36_42),.data_out(wire_d36_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373644(.data_in(wire_d36_43),.data_out(wire_d36_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373645(.data_in(wire_d36_44),.data_out(wire_d36_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373646(.data_in(wire_d36_45),.data_out(wire_d36_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373647(.data_in(wire_d36_46),.data_out(wire_d36_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373648(.data_in(wire_d36_47),.data_out(wire_d36_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373649(.data_in(wire_d36_48),.data_out(wire_d36_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373650(.data_in(wire_d36_49),.data_out(wire_d36_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373651(.data_in(wire_d36_50),.data_out(wire_d36_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373652(.data_in(wire_d36_51),.data_out(wire_d36_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373653(.data_in(wire_d36_52),.data_out(wire_d36_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373654(.data_in(wire_d36_53),.data_out(wire_d36_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373655(.data_in(wire_d36_54),.data_out(wire_d36_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373656(.data_in(wire_d36_55),.data_out(wire_d36_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373657(.data_in(wire_d36_56),.data_out(wire_d36_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373658(.data_in(wire_d36_57),.data_out(wire_d36_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373659(.data_in(wire_d36_58),.data_out(wire_d36_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373660(.data_in(wire_d36_59),.data_out(wire_d36_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373661(.data_in(wire_d36_60),.data_out(wire_d36_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373662(.data_in(wire_d36_61),.data_out(wire_d36_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373663(.data_in(wire_d36_62),.data_out(wire_d36_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373664(.data_in(wire_d36_63),.data_out(wire_d36_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373665(.data_in(wire_d36_64),.data_out(wire_d36_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373666(.data_in(wire_d36_65),.data_out(wire_d36_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373667(.data_in(wire_d36_66),.data_out(wire_d36_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373668(.data_in(wire_d36_67),.data_out(wire_d36_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373669(.data_in(wire_d36_68),.data_out(wire_d36_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373670(.data_in(wire_d36_69),.data_out(wire_d36_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373671(.data_in(wire_d36_70),.data_out(wire_d36_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373672(.data_in(wire_d36_71),.data_out(wire_d36_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373673(.data_in(wire_d36_72),.data_out(wire_d36_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373674(.data_in(wire_d36_73),.data_out(wire_d36_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373675(.data_in(wire_d36_74),.data_out(wire_d36_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373676(.data_in(wire_d36_75),.data_out(wire_d36_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373677(.data_in(wire_d36_76),.data_out(wire_d36_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373678(.data_in(wire_d36_77),.data_out(wire_d36_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373679(.data_in(wire_d36_78),.data_out(wire_d36_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373680(.data_in(wire_d36_79),.data_out(wire_d36_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373681(.data_in(wire_d36_80),.data_out(wire_d36_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373682(.data_in(wire_d36_81),.data_out(wire_d36_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373683(.data_in(wire_d36_82),.data_out(wire_d36_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373684(.data_in(wire_d36_83),.data_out(wire_d36_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373685(.data_in(wire_d36_84),.data_out(wire_d36_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373686(.data_in(wire_d36_85),.data_out(wire_d36_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373687(.data_in(wire_d36_86),.data_out(wire_d36_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373688(.data_in(wire_d36_87),.data_out(wire_d36_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373689(.data_in(wire_d36_88),.data_out(wire_d36_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373690(.data_in(wire_d36_89),.data_out(wire_d36_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373691(.data_in(wire_d36_90),.data_out(wire_d36_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373692(.data_in(wire_d36_91),.data_out(wire_d36_92),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373693(.data_in(wire_d36_92),.data_out(wire_d36_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373694(.data_in(wire_d36_93),.data_out(wire_d36_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373695(.data_in(wire_d36_94),.data_out(wire_d36_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373696(.data_in(wire_d36_95),.data_out(wire_d36_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373697(.data_in(wire_d36_96),.data_out(wire_d36_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373698(.data_in(wire_d36_97),.data_out(wire_d36_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373699(.data_in(wire_d36_98),.data_out(d_out36),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance38370(.data_in(d_in37),.data_out(wire_d37_0),.clk(clk),.rst(rst));            //channel 38
	encoder #(.WIDTH(WIDTH)) encoder_instance38371(.data_in(wire_d37_0),.data_out(wire_d37_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance38372(.data_in(wire_d37_1),.data_out(wire_d37_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance38373(.data_in(wire_d37_2),.data_out(wire_d37_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance38374(.data_in(wire_d37_3),.data_out(wire_d37_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance38375(.data_in(wire_d37_4),.data_out(wire_d37_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance38376(.data_in(wire_d37_5),.data_out(wire_d37_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance38377(.data_in(wire_d37_6),.data_out(wire_d37_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance38378(.data_in(wire_d37_7),.data_out(wire_d37_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance38379(.data_in(wire_d37_8),.data_out(wire_d37_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383710(.data_in(wire_d37_9),.data_out(wire_d37_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383711(.data_in(wire_d37_10),.data_out(wire_d37_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383712(.data_in(wire_d37_11),.data_out(wire_d37_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383713(.data_in(wire_d37_12),.data_out(wire_d37_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383714(.data_in(wire_d37_13),.data_out(wire_d37_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383715(.data_in(wire_d37_14),.data_out(wire_d37_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383716(.data_in(wire_d37_15),.data_out(wire_d37_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383717(.data_in(wire_d37_16),.data_out(wire_d37_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383718(.data_in(wire_d37_17),.data_out(wire_d37_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383719(.data_in(wire_d37_18),.data_out(wire_d37_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383720(.data_in(wire_d37_19),.data_out(wire_d37_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383721(.data_in(wire_d37_20),.data_out(wire_d37_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383722(.data_in(wire_d37_21),.data_out(wire_d37_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383723(.data_in(wire_d37_22),.data_out(wire_d37_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383724(.data_in(wire_d37_23),.data_out(wire_d37_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383725(.data_in(wire_d37_24),.data_out(wire_d37_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383726(.data_in(wire_d37_25),.data_out(wire_d37_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383727(.data_in(wire_d37_26),.data_out(wire_d37_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383728(.data_in(wire_d37_27),.data_out(wire_d37_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383729(.data_in(wire_d37_28),.data_out(wire_d37_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383730(.data_in(wire_d37_29),.data_out(wire_d37_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383731(.data_in(wire_d37_30),.data_out(wire_d37_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383732(.data_in(wire_d37_31),.data_out(wire_d37_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383733(.data_in(wire_d37_32),.data_out(wire_d37_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383734(.data_in(wire_d37_33),.data_out(wire_d37_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383735(.data_in(wire_d37_34),.data_out(wire_d37_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383736(.data_in(wire_d37_35),.data_out(wire_d37_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383737(.data_in(wire_d37_36),.data_out(wire_d37_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383738(.data_in(wire_d37_37),.data_out(wire_d37_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383739(.data_in(wire_d37_38),.data_out(wire_d37_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383740(.data_in(wire_d37_39),.data_out(wire_d37_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383741(.data_in(wire_d37_40),.data_out(wire_d37_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383742(.data_in(wire_d37_41),.data_out(wire_d37_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383743(.data_in(wire_d37_42),.data_out(wire_d37_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383744(.data_in(wire_d37_43),.data_out(wire_d37_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383745(.data_in(wire_d37_44),.data_out(wire_d37_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383746(.data_in(wire_d37_45),.data_out(wire_d37_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383747(.data_in(wire_d37_46),.data_out(wire_d37_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383748(.data_in(wire_d37_47),.data_out(wire_d37_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383749(.data_in(wire_d37_48),.data_out(wire_d37_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383750(.data_in(wire_d37_49),.data_out(wire_d37_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383751(.data_in(wire_d37_50),.data_out(wire_d37_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383752(.data_in(wire_d37_51),.data_out(wire_d37_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383753(.data_in(wire_d37_52),.data_out(wire_d37_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383754(.data_in(wire_d37_53),.data_out(wire_d37_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383755(.data_in(wire_d37_54),.data_out(wire_d37_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383756(.data_in(wire_d37_55),.data_out(wire_d37_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383757(.data_in(wire_d37_56),.data_out(wire_d37_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383758(.data_in(wire_d37_57),.data_out(wire_d37_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383759(.data_in(wire_d37_58),.data_out(wire_d37_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383760(.data_in(wire_d37_59),.data_out(wire_d37_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383761(.data_in(wire_d37_60),.data_out(wire_d37_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383762(.data_in(wire_d37_61),.data_out(wire_d37_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383763(.data_in(wire_d37_62),.data_out(wire_d37_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383764(.data_in(wire_d37_63),.data_out(wire_d37_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383765(.data_in(wire_d37_64),.data_out(wire_d37_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383766(.data_in(wire_d37_65),.data_out(wire_d37_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383767(.data_in(wire_d37_66),.data_out(wire_d37_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383768(.data_in(wire_d37_67),.data_out(wire_d37_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383769(.data_in(wire_d37_68),.data_out(wire_d37_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383770(.data_in(wire_d37_69),.data_out(wire_d37_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383771(.data_in(wire_d37_70),.data_out(wire_d37_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383772(.data_in(wire_d37_71),.data_out(wire_d37_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383773(.data_in(wire_d37_72),.data_out(wire_d37_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383774(.data_in(wire_d37_73),.data_out(wire_d37_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383775(.data_in(wire_d37_74),.data_out(wire_d37_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383776(.data_in(wire_d37_75),.data_out(wire_d37_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383777(.data_in(wire_d37_76),.data_out(wire_d37_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383778(.data_in(wire_d37_77),.data_out(wire_d37_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383779(.data_in(wire_d37_78),.data_out(wire_d37_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383780(.data_in(wire_d37_79),.data_out(wire_d37_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383781(.data_in(wire_d37_80),.data_out(wire_d37_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383782(.data_in(wire_d37_81),.data_out(wire_d37_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383783(.data_in(wire_d37_82),.data_out(wire_d37_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383784(.data_in(wire_d37_83),.data_out(wire_d37_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383785(.data_in(wire_d37_84),.data_out(wire_d37_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383786(.data_in(wire_d37_85),.data_out(wire_d37_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383787(.data_in(wire_d37_86),.data_out(wire_d37_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383788(.data_in(wire_d37_87),.data_out(wire_d37_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383789(.data_in(wire_d37_88),.data_out(wire_d37_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383790(.data_in(wire_d37_89),.data_out(wire_d37_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383791(.data_in(wire_d37_90),.data_out(wire_d37_91),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383792(.data_in(wire_d37_91),.data_out(wire_d37_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383793(.data_in(wire_d37_92),.data_out(wire_d37_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383794(.data_in(wire_d37_93),.data_out(wire_d37_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383795(.data_in(wire_d37_94),.data_out(wire_d37_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383796(.data_in(wire_d37_95),.data_out(wire_d37_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383797(.data_in(wire_d37_96),.data_out(wire_d37_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383798(.data_in(wire_d37_97),.data_out(wire_d37_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383799(.data_in(wire_d37_98),.data_out(d_out37),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance39380(.data_in(d_in38),.data_out(wire_d38_0),.clk(clk),.rst(rst));            //channel 39
	large_mux #(.WIDTH(WIDTH)) large_mux_instance39381(.data_in(wire_d38_0),.data_out(wire_d38_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance39382(.data_in(wire_d38_1),.data_out(wire_d38_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance39383(.data_in(wire_d38_2),.data_out(wire_d38_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance39384(.data_in(wire_d38_3),.data_out(wire_d38_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance39385(.data_in(wire_d38_4),.data_out(wire_d38_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance39386(.data_in(wire_d38_5),.data_out(wire_d38_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance39387(.data_in(wire_d38_6),.data_out(wire_d38_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance39388(.data_in(wire_d38_7),.data_out(wire_d38_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance39389(.data_in(wire_d38_8),.data_out(wire_d38_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393810(.data_in(wire_d38_9),.data_out(wire_d38_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393811(.data_in(wire_d38_10),.data_out(wire_d38_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393812(.data_in(wire_d38_11),.data_out(wire_d38_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393813(.data_in(wire_d38_12),.data_out(wire_d38_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393814(.data_in(wire_d38_13),.data_out(wire_d38_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393815(.data_in(wire_d38_14),.data_out(wire_d38_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393816(.data_in(wire_d38_15),.data_out(wire_d38_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393817(.data_in(wire_d38_16),.data_out(wire_d38_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393818(.data_in(wire_d38_17),.data_out(wire_d38_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393819(.data_in(wire_d38_18),.data_out(wire_d38_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393820(.data_in(wire_d38_19),.data_out(wire_d38_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393821(.data_in(wire_d38_20),.data_out(wire_d38_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393822(.data_in(wire_d38_21),.data_out(wire_d38_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393823(.data_in(wire_d38_22),.data_out(wire_d38_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393824(.data_in(wire_d38_23),.data_out(wire_d38_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393825(.data_in(wire_d38_24),.data_out(wire_d38_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393826(.data_in(wire_d38_25),.data_out(wire_d38_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393827(.data_in(wire_d38_26),.data_out(wire_d38_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393828(.data_in(wire_d38_27),.data_out(wire_d38_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393829(.data_in(wire_d38_28),.data_out(wire_d38_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393830(.data_in(wire_d38_29),.data_out(wire_d38_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393831(.data_in(wire_d38_30),.data_out(wire_d38_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393832(.data_in(wire_d38_31),.data_out(wire_d38_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393833(.data_in(wire_d38_32),.data_out(wire_d38_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393834(.data_in(wire_d38_33),.data_out(wire_d38_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393835(.data_in(wire_d38_34),.data_out(wire_d38_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393836(.data_in(wire_d38_35),.data_out(wire_d38_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393837(.data_in(wire_d38_36),.data_out(wire_d38_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393838(.data_in(wire_d38_37),.data_out(wire_d38_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393839(.data_in(wire_d38_38),.data_out(wire_d38_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393840(.data_in(wire_d38_39),.data_out(wire_d38_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393841(.data_in(wire_d38_40),.data_out(wire_d38_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393842(.data_in(wire_d38_41),.data_out(wire_d38_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393843(.data_in(wire_d38_42),.data_out(wire_d38_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393844(.data_in(wire_d38_43),.data_out(wire_d38_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393845(.data_in(wire_d38_44),.data_out(wire_d38_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393846(.data_in(wire_d38_45),.data_out(wire_d38_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393847(.data_in(wire_d38_46),.data_out(wire_d38_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393848(.data_in(wire_d38_47),.data_out(wire_d38_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393849(.data_in(wire_d38_48),.data_out(wire_d38_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393850(.data_in(wire_d38_49),.data_out(wire_d38_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393851(.data_in(wire_d38_50),.data_out(wire_d38_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393852(.data_in(wire_d38_51),.data_out(wire_d38_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393853(.data_in(wire_d38_52),.data_out(wire_d38_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393854(.data_in(wire_d38_53),.data_out(wire_d38_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393855(.data_in(wire_d38_54),.data_out(wire_d38_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393856(.data_in(wire_d38_55),.data_out(wire_d38_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393857(.data_in(wire_d38_56),.data_out(wire_d38_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393858(.data_in(wire_d38_57),.data_out(wire_d38_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393859(.data_in(wire_d38_58),.data_out(wire_d38_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393860(.data_in(wire_d38_59),.data_out(wire_d38_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393861(.data_in(wire_d38_60),.data_out(wire_d38_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393862(.data_in(wire_d38_61),.data_out(wire_d38_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393863(.data_in(wire_d38_62),.data_out(wire_d38_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393864(.data_in(wire_d38_63),.data_out(wire_d38_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393865(.data_in(wire_d38_64),.data_out(wire_d38_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393866(.data_in(wire_d38_65),.data_out(wire_d38_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393867(.data_in(wire_d38_66),.data_out(wire_d38_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393868(.data_in(wire_d38_67),.data_out(wire_d38_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393869(.data_in(wire_d38_68),.data_out(wire_d38_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393870(.data_in(wire_d38_69),.data_out(wire_d38_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393871(.data_in(wire_d38_70),.data_out(wire_d38_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393872(.data_in(wire_d38_71),.data_out(wire_d38_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393873(.data_in(wire_d38_72),.data_out(wire_d38_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393874(.data_in(wire_d38_73),.data_out(wire_d38_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393875(.data_in(wire_d38_74),.data_out(wire_d38_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393876(.data_in(wire_d38_75),.data_out(wire_d38_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393877(.data_in(wire_d38_76),.data_out(wire_d38_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393878(.data_in(wire_d38_77),.data_out(wire_d38_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393879(.data_in(wire_d38_78),.data_out(wire_d38_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393880(.data_in(wire_d38_79),.data_out(wire_d38_80),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393881(.data_in(wire_d38_80),.data_out(wire_d38_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393882(.data_in(wire_d38_81),.data_out(wire_d38_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393883(.data_in(wire_d38_82),.data_out(wire_d38_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393884(.data_in(wire_d38_83),.data_out(wire_d38_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393885(.data_in(wire_d38_84),.data_out(wire_d38_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393886(.data_in(wire_d38_85),.data_out(wire_d38_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393887(.data_in(wire_d38_86),.data_out(wire_d38_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393888(.data_in(wire_d38_87),.data_out(wire_d38_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393889(.data_in(wire_d38_88),.data_out(wire_d38_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393890(.data_in(wire_d38_89),.data_out(wire_d38_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393891(.data_in(wire_d38_90),.data_out(wire_d38_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393892(.data_in(wire_d38_91),.data_out(wire_d38_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393893(.data_in(wire_d38_92),.data_out(wire_d38_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393894(.data_in(wire_d38_93),.data_out(wire_d38_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393895(.data_in(wire_d38_94),.data_out(wire_d38_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393896(.data_in(wire_d38_95),.data_out(wire_d38_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393897(.data_in(wire_d38_96),.data_out(wire_d38_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393898(.data_in(wire_d38_97),.data_out(wire_d38_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393899(.data_in(wire_d38_98),.data_out(d_out38),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance40390(.data_in(d_in39),.data_out(wire_d39_0),.clk(clk),.rst(rst));            //channel 40
	encoder #(.WIDTH(WIDTH)) encoder_instance40391(.data_in(wire_d39_0),.data_out(wire_d39_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance40392(.data_in(wire_d39_1),.data_out(wire_d39_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance40393(.data_in(wire_d39_2),.data_out(wire_d39_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance40394(.data_in(wire_d39_3),.data_out(wire_d39_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance40395(.data_in(wire_d39_4),.data_out(wire_d39_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance40396(.data_in(wire_d39_5),.data_out(wire_d39_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance40397(.data_in(wire_d39_6),.data_out(wire_d39_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance40398(.data_in(wire_d39_7),.data_out(wire_d39_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance40399(.data_in(wire_d39_8),.data_out(wire_d39_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403910(.data_in(wire_d39_9),.data_out(wire_d39_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403911(.data_in(wire_d39_10),.data_out(wire_d39_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403912(.data_in(wire_d39_11),.data_out(wire_d39_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403913(.data_in(wire_d39_12),.data_out(wire_d39_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403914(.data_in(wire_d39_13),.data_out(wire_d39_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403915(.data_in(wire_d39_14),.data_out(wire_d39_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403916(.data_in(wire_d39_15),.data_out(wire_d39_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403917(.data_in(wire_d39_16),.data_out(wire_d39_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403918(.data_in(wire_d39_17),.data_out(wire_d39_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403919(.data_in(wire_d39_18),.data_out(wire_d39_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403920(.data_in(wire_d39_19),.data_out(wire_d39_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403921(.data_in(wire_d39_20),.data_out(wire_d39_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403922(.data_in(wire_d39_21),.data_out(wire_d39_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403923(.data_in(wire_d39_22),.data_out(wire_d39_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403924(.data_in(wire_d39_23),.data_out(wire_d39_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403925(.data_in(wire_d39_24),.data_out(wire_d39_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403926(.data_in(wire_d39_25),.data_out(wire_d39_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403927(.data_in(wire_d39_26),.data_out(wire_d39_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403928(.data_in(wire_d39_27),.data_out(wire_d39_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403929(.data_in(wire_d39_28),.data_out(wire_d39_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403930(.data_in(wire_d39_29),.data_out(wire_d39_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403931(.data_in(wire_d39_30),.data_out(wire_d39_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403932(.data_in(wire_d39_31),.data_out(wire_d39_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403933(.data_in(wire_d39_32),.data_out(wire_d39_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403934(.data_in(wire_d39_33),.data_out(wire_d39_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403935(.data_in(wire_d39_34),.data_out(wire_d39_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403936(.data_in(wire_d39_35),.data_out(wire_d39_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403937(.data_in(wire_d39_36),.data_out(wire_d39_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403938(.data_in(wire_d39_37),.data_out(wire_d39_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403939(.data_in(wire_d39_38),.data_out(wire_d39_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403940(.data_in(wire_d39_39),.data_out(wire_d39_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403941(.data_in(wire_d39_40),.data_out(wire_d39_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403942(.data_in(wire_d39_41),.data_out(wire_d39_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403943(.data_in(wire_d39_42),.data_out(wire_d39_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403944(.data_in(wire_d39_43),.data_out(wire_d39_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403945(.data_in(wire_d39_44),.data_out(wire_d39_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403946(.data_in(wire_d39_45),.data_out(wire_d39_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403947(.data_in(wire_d39_46),.data_out(wire_d39_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403948(.data_in(wire_d39_47),.data_out(wire_d39_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403949(.data_in(wire_d39_48),.data_out(wire_d39_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403950(.data_in(wire_d39_49),.data_out(wire_d39_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403951(.data_in(wire_d39_50),.data_out(wire_d39_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403952(.data_in(wire_d39_51),.data_out(wire_d39_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403953(.data_in(wire_d39_52),.data_out(wire_d39_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403954(.data_in(wire_d39_53),.data_out(wire_d39_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403955(.data_in(wire_d39_54),.data_out(wire_d39_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403956(.data_in(wire_d39_55),.data_out(wire_d39_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403957(.data_in(wire_d39_56),.data_out(wire_d39_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403958(.data_in(wire_d39_57),.data_out(wire_d39_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403959(.data_in(wire_d39_58),.data_out(wire_d39_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403960(.data_in(wire_d39_59),.data_out(wire_d39_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403961(.data_in(wire_d39_60),.data_out(wire_d39_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403962(.data_in(wire_d39_61),.data_out(wire_d39_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403963(.data_in(wire_d39_62),.data_out(wire_d39_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403964(.data_in(wire_d39_63),.data_out(wire_d39_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403965(.data_in(wire_d39_64),.data_out(wire_d39_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403966(.data_in(wire_d39_65),.data_out(wire_d39_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403967(.data_in(wire_d39_66),.data_out(wire_d39_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403968(.data_in(wire_d39_67),.data_out(wire_d39_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403969(.data_in(wire_d39_68),.data_out(wire_d39_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403970(.data_in(wire_d39_69),.data_out(wire_d39_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403971(.data_in(wire_d39_70),.data_out(wire_d39_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403972(.data_in(wire_d39_71),.data_out(wire_d39_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403973(.data_in(wire_d39_72),.data_out(wire_d39_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403974(.data_in(wire_d39_73),.data_out(wire_d39_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403975(.data_in(wire_d39_74),.data_out(wire_d39_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403976(.data_in(wire_d39_75),.data_out(wire_d39_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403977(.data_in(wire_d39_76),.data_out(wire_d39_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403978(.data_in(wire_d39_77),.data_out(wire_d39_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403979(.data_in(wire_d39_78),.data_out(wire_d39_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403980(.data_in(wire_d39_79),.data_out(wire_d39_80),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403981(.data_in(wire_d39_80),.data_out(wire_d39_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403982(.data_in(wire_d39_81),.data_out(wire_d39_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403983(.data_in(wire_d39_82),.data_out(wire_d39_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403984(.data_in(wire_d39_83),.data_out(wire_d39_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403985(.data_in(wire_d39_84),.data_out(wire_d39_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403986(.data_in(wire_d39_85),.data_out(wire_d39_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403987(.data_in(wire_d39_86),.data_out(wire_d39_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403988(.data_in(wire_d39_87),.data_out(wire_d39_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403989(.data_in(wire_d39_88),.data_out(wire_d39_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403990(.data_in(wire_d39_89),.data_out(wire_d39_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403991(.data_in(wire_d39_90),.data_out(wire_d39_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403992(.data_in(wire_d39_91),.data_out(wire_d39_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403993(.data_in(wire_d39_92),.data_out(wire_d39_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403994(.data_in(wire_d39_93),.data_out(wire_d39_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403995(.data_in(wire_d39_94),.data_out(wire_d39_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403996(.data_in(wire_d39_95),.data_out(wire_d39_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403997(.data_in(wire_d39_96),.data_out(wire_d39_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403998(.data_in(wire_d39_97),.data_out(wire_d39_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403999(.data_in(wire_d39_98),.data_out(d_out39),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance41400(.data_in(d_in40),.data_out(wire_d40_0),.clk(clk),.rst(rst));            //channel 41
	invertion #(.WIDTH(WIDTH)) invertion_instance41401(.data_in(wire_d40_0),.data_out(wire_d40_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance41402(.data_in(wire_d40_1),.data_out(wire_d40_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance41403(.data_in(wire_d40_2),.data_out(wire_d40_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance41404(.data_in(wire_d40_3),.data_out(wire_d40_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance41405(.data_in(wire_d40_4),.data_out(wire_d40_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance41406(.data_in(wire_d40_5),.data_out(wire_d40_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance41407(.data_in(wire_d40_6),.data_out(wire_d40_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance41408(.data_in(wire_d40_7),.data_out(wire_d40_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance41409(.data_in(wire_d40_8),.data_out(wire_d40_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414010(.data_in(wire_d40_9),.data_out(wire_d40_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414011(.data_in(wire_d40_10),.data_out(wire_d40_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414012(.data_in(wire_d40_11),.data_out(wire_d40_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414013(.data_in(wire_d40_12),.data_out(wire_d40_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414014(.data_in(wire_d40_13),.data_out(wire_d40_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414015(.data_in(wire_d40_14),.data_out(wire_d40_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414016(.data_in(wire_d40_15),.data_out(wire_d40_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414017(.data_in(wire_d40_16),.data_out(wire_d40_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414018(.data_in(wire_d40_17),.data_out(wire_d40_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414019(.data_in(wire_d40_18),.data_out(wire_d40_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414020(.data_in(wire_d40_19),.data_out(wire_d40_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414021(.data_in(wire_d40_20),.data_out(wire_d40_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414022(.data_in(wire_d40_21),.data_out(wire_d40_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414023(.data_in(wire_d40_22),.data_out(wire_d40_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414024(.data_in(wire_d40_23),.data_out(wire_d40_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414025(.data_in(wire_d40_24),.data_out(wire_d40_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414026(.data_in(wire_d40_25),.data_out(wire_d40_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414027(.data_in(wire_d40_26),.data_out(wire_d40_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414028(.data_in(wire_d40_27),.data_out(wire_d40_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414029(.data_in(wire_d40_28),.data_out(wire_d40_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414030(.data_in(wire_d40_29),.data_out(wire_d40_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414031(.data_in(wire_d40_30),.data_out(wire_d40_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414032(.data_in(wire_d40_31),.data_out(wire_d40_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414033(.data_in(wire_d40_32),.data_out(wire_d40_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414034(.data_in(wire_d40_33),.data_out(wire_d40_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414035(.data_in(wire_d40_34),.data_out(wire_d40_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414036(.data_in(wire_d40_35),.data_out(wire_d40_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414037(.data_in(wire_d40_36),.data_out(wire_d40_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414038(.data_in(wire_d40_37),.data_out(wire_d40_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414039(.data_in(wire_d40_38),.data_out(wire_d40_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414040(.data_in(wire_d40_39),.data_out(wire_d40_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414041(.data_in(wire_d40_40),.data_out(wire_d40_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414042(.data_in(wire_d40_41),.data_out(wire_d40_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414043(.data_in(wire_d40_42),.data_out(wire_d40_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414044(.data_in(wire_d40_43),.data_out(wire_d40_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414045(.data_in(wire_d40_44),.data_out(wire_d40_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414046(.data_in(wire_d40_45),.data_out(wire_d40_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414047(.data_in(wire_d40_46),.data_out(wire_d40_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414048(.data_in(wire_d40_47),.data_out(wire_d40_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414049(.data_in(wire_d40_48),.data_out(wire_d40_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414050(.data_in(wire_d40_49),.data_out(wire_d40_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414051(.data_in(wire_d40_50),.data_out(wire_d40_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414052(.data_in(wire_d40_51),.data_out(wire_d40_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414053(.data_in(wire_d40_52),.data_out(wire_d40_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414054(.data_in(wire_d40_53),.data_out(wire_d40_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414055(.data_in(wire_d40_54),.data_out(wire_d40_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414056(.data_in(wire_d40_55),.data_out(wire_d40_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414057(.data_in(wire_d40_56),.data_out(wire_d40_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414058(.data_in(wire_d40_57),.data_out(wire_d40_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414059(.data_in(wire_d40_58),.data_out(wire_d40_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414060(.data_in(wire_d40_59),.data_out(wire_d40_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414061(.data_in(wire_d40_60),.data_out(wire_d40_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414062(.data_in(wire_d40_61),.data_out(wire_d40_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414063(.data_in(wire_d40_62),.data_out(wire_d40_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414064(.data_in(wire_d40_63),.data_out(wire_d40_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414065(.data_in(wire_d40_64),.data_out(wire_d40_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414066(.data_in(wire_d40_65),.data_out(wire_d40_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414067(.data_in(wire_d40_66),.data_out(wire_d40_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414068(.data_in(wire_d40_67),.data_out(wire_d40_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414069(.data_in(wire_d40_68),.data_out(wire_d40_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414070(.data_in(wire_d40_69),.data_out(wire_d40_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414071(.data_in(wire_d40_70),.data_out(wire_d40_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414072(.data_in(wire_d40_71),.data_out(wire_d40_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414073(.data_in(wire_d40_72),.data_out(wire_d40_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414074(.data_in(wire_d40_73),.data_out(wire_d40_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414075(.data_in(wire_d40_74),.data_out(wire_d40_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414076(.data_in(wire_d40_75),.data_out(wire_d40_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414077(.data_in(wire_d40_76),.data_out(wire_d40_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414078(.data_in(wire_d40_77),.data_out(wire_d40_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414079(.data_in(wire_d40_78),.data_out(wire_d40_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414080(.data_in(wire_d40_79),.data_out(wire_d40_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414081(.data_in(wire_d40_80),.data_out(wire_d40_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414082(.data_in(wire_d40_81),.data_out(wire_d40_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414083(.data_in(wire_d40_82),.data_out(wire_d40_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414084(.data_in(wire_d40_83),.data_out(wire_d40_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414085(.data_in(wire_d40_84),.data_out(wire_d40_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414086(.data_in(wire_d40_85),.data_out(wire_d40_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414087(.data_in(wire_d40_86),.data_out(wire_d40_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414088(.data_in(wire_d40_87),.data_out(wire_d40_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414089(.data_in(wire_d40_88),.data_out(wire_d40_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414090(.data_in(wire_d40_89),.data_out(wire_d40_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414091(.data_in(wire_d40_90),.data_out(wire_d40_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414092(.data_in(wire_d40_91),.data_out(wire_d40_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414093(.data_in(wire_d40_92),.data_out(wire_d40_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414094(.data_in(wire_d40_93),.data_out(wire_d40_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414095(.data_in(wire_d40_94),.data_out(wire_d40_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414096(.data_in(wire_d40_95),.data_out(wire_d40_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414097(.data_in(wire_d40_96),.data_out(wire_d40_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414098(.data_in(wire_d40_97),.data_out(wire_d40_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414099(.data_in(wire_d40_98),.data_out(d_out40),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance42410(.data_in(d_in41),.data_out(wire_d41_0),.clk(clk),.rst(rst));            //channel 42
	invertion #(.WIDTH(WIDTH)) invertion_instance42411(.data_in(wire_d41_0),.data_out(wire_d41_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance42412(.data_in(wire_d41_1),.data_out(wire_d41_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance42413(.data_in(wire_d41_2),.data_out(wire_d41_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance42414(.data_in(wire_d41_3),.data_out(wire_d41_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance42415(.data_in(wire_d41_4),.data_out(wire_d41_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance42416(.data_in(wire_d41_5),.data_out(wire_d41_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance42417(.data_in(wire_d41_6),.data_out(wire_d41_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance42418(.data_in(wire_d41_7),.data_out(wire_d41_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance42419(.data_in(wire_d41_8),.data_out(wire_d41_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424110(.data_in(wire_d41_9),.data_out(wire_d41_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424111(.data_in(wire_d41_10),.data_out(wire_d41_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424112(.data_in(wire_d41_11),.data_out(wire_d41_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424113(.data_in(wire_d41_12),.data_out(wire_d41_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424114(.data_in(wire_d41_13),.data_out(wire_d41_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424115(.data_in(wire_d41_14),.data_out(wire_d41_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424116(.data_in(wire_d41_15),.data_out(wire_d41_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424117(.data_in(wire_d41_16),.data_out(wire_d41_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424118(.data_in(wire_d41_17),.data_out(wire_d41_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424119(.data_in(wire_d41_18),.data_out(wire_d41_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424120(.data_in(wire_d41_19),.data_out(wire_d41_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424121(.data_in(wire_d41_20),.data_out(wire_d41_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424122(.data_in(wire_d41_21),.data_out(wire_d41_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424123(.data_in(wire_d41_22),.data_out(wire_d41_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424124(.data_in(wire_d41_23),.data_out(wire_d41_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424125(.data_in(wire_d41_24),.data_out(wire_d41_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424126(.data_in(wire_d41_25),.data_out(wire_d41_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424127(.data_in(wire_d41_26),.data_out(wire_d41_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424128(.data_in(wire_d41_27),.data_out(wire_d41_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424129(.data_in(wire_d41_28),.data_out(wire_d41_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424130(.data_in(wire_d41_29),.data_out(wire_d41_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424131(.data_in(wire_d41_30),.data_out(wire_d41_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424132(.data_in(wire_d41_31),.data_out(wire_d41_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424133(.data_in(wire_d41_32),.data_out(wire_d41_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424134(.data_in(wire_d41_33),.data_out(wire_d41_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424135(.data_in(wire_d41_34),.data_out(wire_d41_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424136(.data_in(wire_d41_35),.data_out(wire_d41_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424137(.data_in(wire_d41_36),.data_out(wire_d41_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424138(.data_in(wire_d41_37),.data_out(wire_d41_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424139(.data_in(wire_d41_38),.data_out(wire_d41_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424140(.data_in(wire_d41_39),.data_out(wire_d41_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424141(.data_in(wire_d41_40),.data_out(wire_d41_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424142(.data_in(wire_d41_41),.data_out(wire_d41_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424143(.data_in(wire_d41_42),.data_out(wire_d41_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424144(.data_in(wire_d41_43),.data_out(wire_d41_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424145(.data_in(wire_d41_44),.data_out(wire_d41_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424146(.data_in(wire_d41_45),.data_out(wire_d41_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424147(.data_in(wire_d41_46),.data_out(wire_d41_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424148(.data_in(wire_d41_47),.data_out(wire_d41_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424149(.data_in(wire_d41_48),.data_out(wire_d41_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424150(.data_in(wire_d41_49),.data_out(wire_d41_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424151(.data_in(wire_d41_50),.data_out(wire_d41_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424152(.data_in(wire_d41_51),.data_out(wire_d41_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424153(.data_in(wire_d41_52),.data_out(wire_d41_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424154(.data_in(wire_d41_53),.data_out(wire_d41_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424155(.data_in(wire_d41_54),.data_out(wire_d41_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424156(.data_in(wire_d41_55),.data_out(wire_d41_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424157(.data_in(wire_d41_56),.data_out(wire_d41_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424158(.data_in(wire_d41_57),.data_out(wire_d41_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424159(.data_in(wire_d41_58),.data_out(wire_d41_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424160(.data_in(wire_d41_59),.data_out(wire_d41_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424161(.data_in(wire_d41_60),.data_out(wire_d41_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424162(.data_in(wire_d41_61),.data_out(wire_d41_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424163(.data_in(wire_d41_62),.data_out(wire_d41_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424164(.data_in(wire_d41_63),.data_out(wire_d41_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424165(.data_in(wire_d41_64),.data_out(wire_d41_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424166(.data_in(wire_d41_65),.data_out(wire_d41_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424167(.data_in(wire_d41_66),.data_out(wire_d41_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424168(.data_in(wire_d41_67),.data_out(wire_d41_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424169(.data_in(wire_d41_68),.data_out(wire_d41_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424170(.data_in(wire_d41_69),.data_out(wire_d41_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424171(.data_in(wire_d41_70),.data_out(wire_d41_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424172(.data_in(wire_d41_71),.data_out(wire_d41_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424173(.data_in(wire_d41_72),.data_out(wire_d41_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424174(.data_in(wire_d41_73),.data_out(wire_d41_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424175(.data_in(wire_d41_74),.data_out(wire_d41_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424176(.data_in(wire_d41_75),.data_out(wire_d41_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424177(.data_in(wire_d41_76),.data_out(wire_d41_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424178(.data_in(wire_d41_77),.data_out(wire_d41_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424179(.data_in(wire_d41_78),.data_out(wire_d41_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424180(.data_in(wire_d41_79),.data_out(wire_d41_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424181(.data_in(wire_d41_80),.data_out(wire_d41_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424182(.data_in(wire_d41_81),.data_out(wire_d41_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424183(.data_in(wire_d41_82),.data_out(wire_d41_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424184(.data_in(wire_d41_83),.data_out(wire_d41_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424185(.data_in(wire_d41_84),.data_out(wire_d41_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424186(.data_in(wire_d41_85),.data_out(wire_d41_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424187(.data_in(wire_d41_86),.data_out(wire_d41_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424188(.data_in(wire_d41_87),.data_out(wire_d41_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424189(.data_in(wire_d41_88),.data_out(wire_d41_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424190(.data_in(wire_d41_89),.data_out(wire_d41_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424191(.data_in(wire_d41_90),.data_out(wire_d41_91),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424192(.data_in(wire_d41_91),.data_out(wire_d41_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424193(.data_in(wire_d41_92),.data_out(wire_d41_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424194(.data_in(wire_d41_93),.data_out(wire_d41_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424195(.data_in(wire_d41_94),.data_out(wire_d41_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424196(.data_in(wire_d41_95),.data_out(wire_d41_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424197(.data_in(wire_d41_96),.data_out(wire_d41_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424198(.data_in(wire_d41_97),.data_out(wire_d41_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424199(.data_in(wire_d41_98),.data_out(d_out41),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance43420(.data_in(d_in42),.data_out(wire_d42_0),.clk(clk),.rst(rst));            //channel 43
	large_mux #(.WIDTH(WIDTH)) large_mux_instance43421(.data_in(wire_d42_0),.data_out(wire_d42_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43422(.data_in(wire_d42_1),.data_out(wire_d42_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance43423(.data_in(wire_d42_2),.data_out(wire_d42_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance43424(.data_in(wire_d42_3),.data_out(wire_d42_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance43425(.data_in(wire_d42_4),.data_out(wire_d42_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43426(.data_in(wire_d42_5),.data_out(wire_d42_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43427(.data_in(wire_d42_6),.data_out(wire_d42_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43428(.data_in(wire_d42_7),.data_out(wire_d42_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance43429(.data_in(wire_d42_8),.data_out(wire_d42_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434210(.data_in(wire_d42_9),.data_out(wire_d42_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434211(.data_in(wire_d42_10),.data_out(wire_d42_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434212(.data_in(wire_d42_11),.data_out(wire_d42_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434213(.data_in(wire_d42_12),.data_out(wire_d42_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434214(.data_in(wire_d42_13),.data_out(wire_d42_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434215(.data_in(wire_d42_14),.data_out(wire_d42_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434216(.data_in(wire_d42_15),.data_out(wire_d42_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434217(.data_in(wire_d42_16),.data_out(wire_d42_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434218(.data_in(wire_d42_17),.data_out(wire_d42_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434219(.data_in(wire_d42_18),.data_out(wire_d42_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434220(.data_in(wire_d42_19),.data_out(wire_d42_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434221(.data_in(wire_d42_20),.data_out(wire_d42_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434222(.data_in(wire_d42_21),.data_out(wire_d42_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434223(.data_in(wire_d42_22),.data_out(wire_d42_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434224(.data_in(wire_d42_23),.data_out(wire_d42_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434225(.data_in(wire_d42_24),.data_out(wire_d42_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434226(.data_in(wire_d42_25),.data_out(wire_d42_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434227(.data_in(wire_d42_26),.data_out(wire_d42_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434228(.data_in(wire_d42_27),.data_out(wire_d42_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434229(.data_in(wire_d42_28),.data_out(wire_d42_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434230(.data_in(wire_d42_29),.data_out(wire_d42_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434231(.data_in(wire_d42_30),.data_out(wire_d42_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434232(.data_in(wire_d42_31),.data_out(wire_d42_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434233(.data_in(wire_d42_32),.data_out(wire_d42_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434234(.data_in(wire_d42_33),.data_out(wire_d42_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434235(.data_in(wire_d42_34),.data_out(wire_d42_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434236(.data_in(wire_d42_35),.data_out(wire_d42_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434237(.data_in(wire_d42_36),.data_out(wire_d42_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434238(.data_in(wire_d42_37),.data_out(wire_d42_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434239(.data_in(wire_d42_38),.data_out(wire_d42_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434240(.data_in(wire_d42_39),.data_out(wire_d42_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434241(.data_in(wire_d42_40),.data_out(wire_d42_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434242(.data_in(wire_d42_41),.data_out(wire_d42_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434243(.data_in(wire_d42_42),.data_out(wire_d42_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434244(.data_in(wire_d42_43),.data_out(wire_d42_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434245(.data_in(wire_d42_44),.data_out(wire_d42_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434246(.data_in(wire_d42_45),.data_out(wire_d42_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434247(.data_in(wire_d42_46),.data_out(wire_d42_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434248(.data_in(wire_d42_47),.data_out(wire_d42_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434249(.data_in(wire_d42_48),.data_out(wire_d42_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434250(.data_in(wire_d42_49),.data_out(wire_d42_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434251(.data_in(wire_d42_50),.data_out(wire_d42_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434252(.data_in(wire_d42_51),.data_out(wire_d42_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434253(.data_in(wire_d42_52),.data_out(wire_d42_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434254(.data_in(wire_d42_53),.data_out(wire_d42_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434255(.data_in(wire_d42_54),.data_out(wire_d42_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434256(.data_in(wire_d42_55),.data_out(wire_d42_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434257(.data_in(wire_d42_56),.data_out(wire_d42_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434258(.data_in(wire_d42_57),.data_out(wire_d42_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434259(.data_in(wire_d42_58),.data_out(wire_d42_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434260(.data_in(wire_d42_59),.data_out(wire_d42_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434261(.data_in(wire_d42_60),.data_out(wire_d42_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434262(.data_in(wire_d42_61),.data_out(wire_d42_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434263(.data_in(wire_d42_62),.data_out(wire_d42_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434264(.data_in(wire_d42_63),.data_out(wire_d42_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434265(.data_in(wire_d42_64),.data_out(wire_d42_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434266(.data_in(wire_d42_65),.data_out(wire_d42_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434267(.data_in(wire_d42_66),.data_out(wire_d42_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434268(.data_in(wire_d42_67),.data_out(wire_d42_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434269(.data_in(wire_d42_68),.data_out(wire_d42_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434270(.data_in(wire_d42_69),.data_out(wire_d42_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434271(.data_in(wire_d42_70),.data_out(wire_d42_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434272(.data_in(wire_d42_71),.data_out(wire_d42_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434273(.data_in(wire_d42_72),.data_out(wire_d42_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434274(.data_in(wire_d42_73),.data_out(wire_d42_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434275(.data_in(wire_d42_74),.data_out(wire_d42_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434276(.data_in(wire_d42_75),.data_out(wire_d42_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434277(.data_in(wire_d42_76),.data_out(wire_d42_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434278(.data_in(wire_d42_77),.data_out(wire_d42_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434279(.data_in(wire_d42_78),.data_out(wire_d42_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434280(.data_in(wire_d42_79),.data_out(wire_d42_80),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434281(.data_in(wire_d42_80),.data_out(wire_d42_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434282(.data_in(wire_d42_81),.data_out(wire_d42_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434283(.data_in(wire_d42_82),.data_out(wire_d42_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434284(.data_in(wire_d42_83),.data_out(wire_d42_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434285(.data_in(wire_d42_84),.data_out(wire_d42_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434286(.data_in(wire_d42_85),.data_out(wire_d42_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434287(.data_in(wire_d42_86),.data_out(wire_d42_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434288(.data_in(wire_d42_87),.data_out(wire_d42_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434289(.data_in(wire_d42_88),.data_out(wire_d42_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434290(.data_in(wire_d42_89),.data_out(wire_d42_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434291(.data_in(wire_d42_90),.data_out(wire_d42_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434292(.data_in(wire_d42_91),.data_out(wire_d42_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434293(.data_in(wire_d42_92),.data_out(wire_d42_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434294(.data_in(wire_d42_93),.data_out(wire_d42_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434295(.data_in(wire_d42_94),.data_out(wire_d42_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434296(.data_in(wire_d42_95),.data_out(wire_d42_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434297(.data_in(wire_d42_96),.data_out(wire_d42_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434298(.data_in(wire_d42_97),.data_out(wire_d42_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434299(.data_in(wire_d42_98),.data_out(d_out42),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance44430(.data_in(d_in43),.data_out(wire_d43_0),.clk(clk),.rst(rst));            //channel 44
	encoder #(.WIDTH(WIDTH)) encoder_instance44431(.data_in(wire_d43_0),.data_out(wire_d43_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance44432(.data_in(wire_d43_1),.data_out(wire_d43_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance44433(.data_in(wire_d43_2),.data_out(wire_d43_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance44434(.data_in(wire_d43_3),.data_out(wire_d43_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance44435(.data_in(wire_d43_4),.data_out(wire_d43_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance44436(.data_in(wire_d43_5),.data_out(wire_d43_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance44437(.data_in(wire_d43_6),.data_out(wire_d43_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance44438(.data_in(wire_d43_7),.data_out(wire_d43_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance44439(.data_in(wire_d43_8),.data_out(wire_d43_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444310(.data_in(wire_d43_9),.data_out(wire_d43_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444311(.data_in(wire_d43_10),.data_out(wire_d43_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444312(.data_in(wire_d43_11),.data_out(wire_d43_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444313(.data_in(wire_d43_12),.data_out(wire_d43_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444314(.data_in(wire_d43_13),.data_out(wire_d43_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444315(.data_in(wire_d43_14),.data_out(wire_d43_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444316(.data_in(wire_d43_15),.data_out(wire_d43_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444317(.data_in(wire_d43_16),.data_out(wire_d43_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444318(.data_in(wire_d43_17),.data_out(wire_d43_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444319(.data_in(wire_d43_18),.data_out(wire_d43_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444320(.data_in(wire_d43_19),.data_out(wire_d43_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444321(.data_in(wire_d43_20),.data_out(wire_d43_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444322(.data_in(wire_d43_21),.data_out(wire_d43_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444323(.data_in(wire_d43_22),.data_out(wire_d43_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444324(.data_in(wire_d43_23),.data_out(wire_d43_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444325(.data_in(wire_d43_24),.data_out(wire_d43_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444326(.data_in(wire_d43_25),.data_out(wire_d43_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444327(.data_in(wire_d43_26),.data_out(wire_d43_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444328(.data_in(wire_d43_27),.data_out(wire_d43_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444329(.data_in(wire_d43_28),.data_out(wire_d43_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444330(.data_in(wire_d43_29),.data_out(wire_d43_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444331(.data_in(wire_d43_30),.data_out(wire_d43_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444332(.data_in(wire_d43_31),.data_out(wire_d43_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444333(.data_in(wire_d43_32),.data_out(wire_d43_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444334(.data_in(wire_d43_33),.data_out(wire_d43_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444335(.data_in(wire_d43_34),.data_out(wire_d43_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444336(.data_in(wire_d43_35),.data_out(wire_d43_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444337(.data_in(wire_d43_36),.data_out(wire_d43_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444338(.data_in(wire_d43_37),.data_out(wire_d43_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444339(.data_in(wire_d43_38),.data_out(wire_d43_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444340(.data_in(wire_d43_39),.data_out(wire_d43_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444341(.data_in(wire_d43_40),.data_out(wire_d43_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444342(.data_in(wire_d43_41),.data_out(wire_d43_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444343(.data_in(wire_d43_42),.data_out(wire_d43_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444344(.data_in(wire_d43_43),.data_out(wire_d43_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444345(.data_in(wire_d43_44),.data_out(wire_d43_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444346(.data_in(wire_d43_45),.data_out(wire_d43_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444347(.data_in(wire_d43_46),.data_out(wire_d43_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444348(.data_in(wire_d43_47),.data_out(wire_d43_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444349(.data_in(wire_d43_48),.data_out(wire_d43_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444350(.data_in(wire_d43_49),.data_out(wire_d43_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444351(.data_in(wire_d43_50),.data_out(wire_d43_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444352(.data_in(wire_d43_51),.data_out(wire_d43_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444353(.data_in(wire_d43_52),.data_out(wire_d43_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444354(.data_in(wire_d43_53),.data_out(wire_d43_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444355(.data_in(wire_d43_54),.data_out(wire_d43_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444356(.data_in(wire_d43_55),.data_out(wire_d43_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444357(.data_in(wire_d43_56),.data_out(wire_d43_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444358(.data_in(wire_d43_57),.data_out(wire_d43_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444359(.data_in(wire_d43_58),.data_out(wire_d43_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444360(.data_in(wire_d43_59),.data_out(wire_d43_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444361(.data_in(wire_d43_60),.data_out(wire_d43_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444362(.data_in(wire_d43_61),.data_out(wire_d43_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444363(.data_in(wire_d43_62),.data_out(wire_d43_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444364(.data_in(wire_d43_63),.data_out(wire_d43_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444365(.data_in(wire_d43_64),.data_out(wire_d43_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444366(.data_in(wire_d43_65),.data_out(wire_d43_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444367(.data_in(wire_d43_66),.data_out(wire_d43_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444368(.data_in(wire_d43_67),.data_out(wire_d43_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444369(.data_in(wire_d43_68),.data_out(wire_d43_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444370(.data_in(wire_d43_69),.data_out(wire_d43_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444371(.data_in(wire_d43_70),.data_out(wire_d43_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444372(.data_in(wire_d43_71),.data_out(wire_d43_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444373(.data_in(wire_d43_72),.data_out(wire_d43_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444374(.data_in(wire_d43_73),.data_out(wire_d43_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444375(.data_in(wire_d43_74),.data_out(wire_d43_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444376(.data_in(wire_d43_75),.data_out(wire_d43_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444377(.data_in(wire_d43_76),.data_out(wire_d43_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444378(.data_in(wire_d43_77),.data_out(wire_d43_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444379(.data_in(wire_d43_78),.data_out(wire_d43_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444380(.data_in(wire_d43_79),.data_out(wire_d43_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444381(.data_in(wire_d43_80),.data_out(wire_d43_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444382(.data_in(wire_d43_81),.data_out(wire_d43_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444383(.data_in(wire_d43_82),.data_out(wire_d43_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444384(.data_in(wire_d43_83),.data_out(wire_d43_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444385(.data_in(wire_d43_84),.data_out(wire_d43_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444386(.data_in(wire_d43_85),.data_out(wire_d43_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444387(.data_in(wire_d43_86),.data_out(wire_d43_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444388(.data_in(wire_d43_87),.data_out(wire_d43_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444389(.data_in(wire_d43_88),.data_out(wire_d43_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444390(.data_in(wire_d43_89),.data_out(wire_d43_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444391(.data_in(wire_d43_90),.data_out(wire_d43_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444392(.data_in(wire_d43_91),.data_out(wire_d43_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444393(.data_in(wire_d43_92),.data_out(wire_d43_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444394(.data_in(wire_d43_93),.data_out(wire_d43_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444395(.data_in(wire_d43_94),.data_out(wire_d43_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444396(.data_in(wire_d43_95),.data_out(wire_d43_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444397(.data_in(wire_d43_96),.data_out(wire_d43_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444398(.data_in(wire_d43_97),.data_out(wire_d43_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444399(.data_in(wire_d43_98),.data_out(d_out43),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance45440(.data_in(d_in44),.data_out(wire_d44_0),.clk(clk),.rst(rst));            //channel 45
	large_mux #(.WIDTH(WIDTH)) large_mux_instance45441(.data_in(wire_d44_0),.data_out(wire_d44_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance45442(.data_in(wire_d44_1),.data_out(wire_d44_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance45443(.data_in(wire_d44_2),.data_out(wire_d44_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance45444(.data_in(wire_d44_3),.data_out(wire_d44_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance45445(.data_in(wire_d44_4),.data_out(wire_d44_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance45446(.data_in(wire_d44_5),.data_out(wire_d44_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance45447(.data_in(wire_d44_6),.data_out(wire_d44_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance45448(.data_in(wire_d44_7),.data_out(wire_d44_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance45449(.data_in(wire_d44_8),.data_out(wire_d44_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454410(.data_in(wire_d44_9),.data_out(wire_d44_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454411(.data_in(wire_d44_10),.data_out(wire_d44_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454412(.data_in(wire_d44_11),.data_out(wire_d44_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454413(.data_in(wire_d44_12),.data_out(wire_d44_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454414(.data_in(wire_d44_13),.data_out(wire_d44_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454415(.data_in(wire_d44_14),.data_out(wire_d44_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454416(.data_in(wire_d44_15),.data_out(wire_d44_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454417(.data_in(wire_d44_16),.data_out(wire_d44_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454418(.data_in(wire_d44_17),.data_out(wire_d44_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454419(.data_in(wire_d44_18),.data_out(wire_d44_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454420(.data_in(wire_d44_19),.data_out(wire_d44_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454421(.data_in(wire_d44_20),.data_out(wire_d44_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454422(.data_in(wire_d44_21),.data_out(wire_d44_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454423(.data_in(wire_d44_22),.data_out(wire_d44_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454424(.data_in(wire_d44_23),.data_out(wire_d44_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454425(.data_in(wire_d44_24),.data_out(wire_d44_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454426(.data_in(wire_d44_25),.data_out(wire_d44_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454427(.data_in(wire_d44_26),.data_out(wire_d44_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454428(.data_in(wire_d44_27),.data_out(wire_d44_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454429(.data_in(wire_d44_28),.data_out(wire_d44_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454430(.data_in(wire_d44_29),.data_out(wire_d44_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454431(.data_in(wire_d44_30),.data_out(wire_d44_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454432(.data_in(wire_d44_31),.data_out(wire_d44_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454433(.data_in(wire_d44_32),.data_out(wire_d44_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454434(.data_in(wire_d44_33),.data_out(wire_d44_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454435(.data_in(wire_d44_34),.data_out(wire_d44_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454436(.data_in(wire_d44_35),.data_out(wire_d44_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454437(.data_in(wire_d44_36),.data_out(wire_d44_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454438(.data_in(wire_d44_37),.data_out(wire_d44_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454439(.data_in(wire_d44_38),.data_out(wire_d44_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454440(.data_in(wire_d44_39),.data_out(wire_d44_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454441(.data_in(wire_d44_40),.data_out(wire_d44_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454442(.data_in(wire_d44_41),.data_out(wire_d44_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454443(.data_in(wire_d44_42),.data_out(wire_d44_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454444(.data_in(wire_d44_43),.data_out(wire_d44_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454445(.data_in(wire_d44_44),.data_out(wire_d44_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454446(.data_in(wire_d44_45),.data_out(wire_d44_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454447(.data_in(wire_d44_46),.data_out(wire_d44_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454448(.data_in(wire_d44_47),.data_out(wire_d44_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454449(.data_in(wire_d44_48),.data_out(wire_d44_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454450(.data_in(wire_d44_49),.data_out(wire_d44_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454451(.data_in(wire_d44_50),.data_out(wire_d44_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454452(.data_in(wire_d44_51),.data_out(wire_d44_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454453(.data_in(wire_d44_52),.data_out(wire_d44_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454454(.data_in(wire_d44_53),.data_out(wire_d44_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454455(.data_in(wire_d44_54),.data_out(wire_d44_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454456(.data_in(wire_d44_55),.data_out(wire_d44_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454457(.data_in(wire_d44_56),.data_out(wire_d44_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454458(.data_in(wire_d44_57),.data_out(wire_d44_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454459(.data_in(wire_d44_58),.data_out(wire_d44_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454460(.data_in(wire_d44_59),.data_out(wire_d44_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454461(.data_in(wire_d44_60),.data_out(wire_d44_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454462(.data_in(wire_d44_61),.data_out(wire_d44_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454463(.data_in(wire_d44_62),.data_out(wire_d44_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454464(.data_in(wire_d44_63),.data_out(wire_d44_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454465(.data_in(wire_d44_64),.data_out(wire_d44_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454466(.data_in(wire_d44_65),.data_out(wire_d44_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454467(.data_in(wire_d44_66),.data_out(wire_d44_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454468(.data_in(wire_d44_67),.data_out(wire_d44_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454469(.data_in(wire_d44_68),.data_out(wire_d44_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454470(.data_in(wire_d44_69),.data_out(wire_d44_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454471(.data_in(wire_d44_70),.data_out(wire_d44_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454472(.data_in(wire_d44_71),.data_out(wire_d44_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454473(.data_in(wire_d44_72),.data_out(wire_d44_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454474(.data_in(wire_d44_73),.data_out(wire_d44_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454475(.data_in(wire_d44_74),.data_out(wire_d44_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454476(.data_in(wire_d44_75),.data_out(wire_d44_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454477(.data_in(wire_d44_76),.data_out(wire_d44_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454478(.data_in(wire_d44_77),.data_out(wire_d44_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454479(.data_in(wire_d44_78),.data_out(wire_d44_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454480(.data_in(wire_d44_79),.data_out(wire_d44_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454481(.data_in(wire_d44_80),.data_out(wire_d44_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454482(.data_in(wire_d44_81),.data_out(wire_d44_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454483(.data_in(wire_d44_82),.data_out(wire_d44_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454484(.data_in(wire_d44_83),.data_out(wire_d44_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454485(.data_in(wire_d44_84),.data_out(wire_d44_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454486(.data_in(wire_d44_85),.data_out(wire_d44_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454487(.data_in(wire_d44_86),.data_out(wire_d44_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454488(.data_in(wire_d44_87),.data_out(wire_d44_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454489(.data_in(wire_d44_88),.data_out(wire_d44_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454490(.data_in(wire_d44_89),.data_out(wire_d44_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454491(.data_in(wire_d44_90),.data_out(wire_d44_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454492(.data_in(wire_d44_91),.data_out(wire_d44_92),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454493(.data_in(wire_d44_92),.data_out(wire_d44_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454494(.data_in(wire_d44_93),.data_out(wire_d44_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454495(.data_in(wire_d44_94),.data_out(wire_d44_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454496(.data_in(wire_d44_95),.data_out(wire_d44_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454497(.data_in(wire_d44_96),.data_out(wire_d44_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454498(.data_in(wire_d44_97),.data_out(wire_d44_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454499(.data_in(wire_d44_98),.data_out(d_out44),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance46450(.data_in(d_in45),.data_out(wire_d45_0),.clk(clk),.rst(rst));            //channel 46
	invertion #(.WIDTH(WIDTH)) invertion_instance46451(.data_in(wire_d45_0),.data_out(wire_d45_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance46452(.data_in(wire_d45_1),.data_out(wire_d45_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance46453(.data_in(wire_d45_2),.data_out(wire_d45_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance46454(.data_in(wire_d45_3),.data_out(wire_d45_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance46455(.data_in(wire_d45_4),.data_out(wire_d45_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance46456(.data_in(wire_d45_5),.data_out(wire_d45_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance46457(.data_in(wire_d45_6),.data_out(wire_d45_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance46458(.data_in(wire_d45_7),.data_out(wire_d45_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance46459(.data_in(wire_d45_8),.data_out(wire_d45_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464510(.data_in(wire_d45_9),.data_out(wire_d45_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464511(.data_in(wire_d45_10),.data_out(wire_d45_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464512(.data_in(wire_d45_11),.data_out(wire_d45_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464513(.data_in(wire_d45_12),.data_out(wire_d45_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464514(.data_in(wire_d45_13),.data_out(wire_d45_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464515(.data_in(wire_d45_14),.data_out(wire_d45_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464516(.data_in(wire_d45_15),.data_out(wire_d45_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464517(.data_in(wire_d45_16),.data_out(wire_d45_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464518(.data_in(wire_d45_17),.data_out(wire_d45_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464519(.data_in(wire_d45_18),.data_out(wire_d45_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464520(.data_in(wire_d45_19),.data_out(wire_d45_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464521(.data_in(wire_d45_20),.data_out(wire_d45_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464522(.data_in(wire_d45_21),.data_out(wire_d45_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464523(.data_in(wire_d45_22),.data_out(wire_d45_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464524(.data_in(wire_d45_23),.data_out(wire_d45_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464525(.data_in(wire_d45_24),.data_out(wire_d45_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464526(.data_in(wire_d45_25),.data_out(wire_d45_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464527(.data_in(wire_d45_26),.data_out(wire_d45_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464528(.data_in(wire_d45_27),.data_out(wire_d45_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464529(.data_in(wire_d45_28),.data_out(wire_d45_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464530(.data_in(wire_d45_29),.data_out(wire_d45_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464531(.data_in(wire_d45_30),.data_out(wire_d45_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464532(.data_in(wire_d45_31),.data_out(wire_d45_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464533(.data_in(wire_d45_32),.data_out(wire_d45_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464534(.data_in(wire_d45_33),.data_out(wire_d45_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464535(.data_in(wire_d45_34),.data_out(wire_d45_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464536(.data_in(wire_d45_35),.data_out(wire_d45_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464537(.data_in(wire_d45_36),.data_out(wire_d45_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464538(.data_in(wire_d45_37),.data_out(wire_d45_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464539(.data_in(wire_d45_38),.data_out(wire_d45_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464540(.data_in(wire_d45_39),.data_out(wire_d45_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464541(.data_in(wire_d45_40),.data_out(wire_d45_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464542(.data_in(wire_d45_41),.data_out(wire_d45_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464543(.data_in(wire_d45_42),.data_out(wire_d45_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464544(.data_in(wire_d45_43),.data_out(wire_d45_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464545(.data_in(wire_d45_44),.data_out(wire_d45_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464546(.data_in(wire_d45_45),.data_out(wire_d45_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464547(.data_in(wire_d45_46),.data_out(wire_d45_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464548(.data_in(wire_d45_47),.data_out(wire_d45_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464549(.data_in(wire_d45_48),.data_out(wire_d45_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464550(.data_in(wire_d45_49),.data_out(wire_d45_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464551(.data_in(wire_d45_50),.data_out(wire_d45_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464552(.data_in(wire_d45_51),.data_out(wire_d45_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464553(.data_in(wire_d45_52),.data_out(wire_d45_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464554(.data_in(wire_d45_53),.data_out(wire_d45_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464555(.data_in(wire_d45_54),.data_out(wire_d45_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464556(.data_in(wire_d45_55),.data_out(wire_d45_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464557(.data_in(wire_d45_56),.data_out(wire_d45_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464558(.data_in(wire_d45_57),.data_out(wire_d45_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464559(.data_in(wire_d45_58),.data_out(wire_d45_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464560(.data_in(wire_d45_59),.data_out(wire_d45_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464561(.data_in(wire_d45_60),.data_out(wire_d45_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464562(.data_in(wire_d45_61),.data_out(wire_d45_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464563(.data_in(wire_d45_62),.data_out(wire_d45_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464564(.data_in(wire_d45_63),.data_out(wire_d45_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464565(.data_in(wire_d45_64),.data_out(wire_d45_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464566(.data_in(wire_d45_65),.data_out(wire_d45_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464567(.data_in(wire_d45_66),.data_out(wire_d45_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464568(.data_in(wire_d45_67),.data_out(wire_d45_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464569(.data_in(wire_d45_68),.data_out(wire_d45_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464570(.data_in(wire_d45_69),.data_out(wire_d45_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464571(.data_in(wire_d45_70),.data_out(wire_d45_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464572(.data_in(wire_d45_71),.data_out(wire_d45_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464573(.data_in(wire_d45_72),.data_out(wire_d45_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464574(.data_in(wire_d45_73),.data_out(wire_d45_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464575(.data_in(wire_d45_74),.data_out(wire_d45_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464576(.data_in(wire_d45_75),.data_out(wire_d45_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464577(.data_in(wire_d45_76),.data_out(wire_d45_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464578(.data_in(wire_d45_77),.data_out(wire_d45_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464579(.data_in(wire_d45_78),.data_out(wire_d45_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464580(.data_in(wire_d45_79),.data_out(wire_d45_80),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464581(.data_in(wire_d45_80),.data_out(wire_d45_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464582(.data_in(wire_d45_81),.data_out(wire_d45_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464583(.data_in(wire_d45_82),.data_out(wire_d45_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464584(.data_in(wire_d45_83),.data_out(wire_d45_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464585(.data_in(wire_d45_84),.data_out(wire_d45_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464586(.data_in(wire_d45_85),.data_out(wire_d45_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464587(.data_in(wire_d45_86),.data_out(wire_d45_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464588(.data_in(wire_d45_87),.data_out(wire_d45_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464589(.data_in(wire_d45_88),.data_out(wire_d45_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464590(.data_in(wire_d45_89),.data_out(wire_d45_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464591(.data_in(wire_d45_90),.data_out(wire_d45_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464592(.data_in(wire_d45_91),.data_out(wire_d45_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464593(.data_in(wire_d45_92),.data_out(wire_d45_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464594(.data_in(wire_d45_93),.data_out(wire_d45_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464595(.data_in(wire_d45_94),.data_out(wire_d45_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464596(.data_in(wire_d45_95),.data_out(wire_d45_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464597(.data_in(wire_d45_96),.data_out(wire_d45_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464598(.data_in(wire_d45_97),.data_out(wire_d45_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464599(.data_in(wire_d45_98),.data_out(d_out45),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance47460(.data_in(d_in46),.data_out(wire_d46_0),.clk(clk),.rst(rst));            //channel 47
	register #(.WIDTH(WIDTH)) register_instance47461(.data_in(wire_d46_0),.data_out(wire_d46_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance47462(.data_in(wire_d46_1),.data_out(wire_d46_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance47463(.data_in(wire_d46_2),.data_out(wire_d46_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance47464(.data_in(wire_d46_3),.data_out(wire_d46_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance47465(.data_in(wire_d46_4),.data_out(wire_d46_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance47466(.data_in(wire_d46_5),.data_out(wire_d46_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance47467(.data_in(wire_d46_6),.data_out(wire_d46_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance47468(.data_in(wire_d46_7),.data_out(wire_d46_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance47469(.data_in(wire_d46_8),.data_out(wire_d46_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474610(.data_in(wire_d46_9),.data_out(wire_d46_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474611(.data_in(wire_d46_10),.data_out(wire_d46_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474612(.data_in(wire_d46_11),.data_out(wire_d46_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474613(.data_in(wire_d46_12),.data_out(wire_d46_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474614(.data_in(wire_d46_13),.data_out(wire_d46_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474615(.data_in(wire_d46_14),.data_out(wire_d46_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474616(.data_in(wire_d46_15),.data_out(wire_d46_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474617(.data_in(wire_d46_16),.data_out(wire_d46_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474618(.data_in(wire_d46_17),.data_out(wire_d46_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474619(.data_in(wire_d46_18),.data_out(wire_d46_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474620(.data_in(wire_d46_19),.data_out(wire_d46_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474621(.data_in(wire_d46_20),.data_out(wire_d46_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474622(.data_in(wire_d46_21),.data_out(wire_d46_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474623(.data_in(wire_d46_22),.data_out(wire_d46_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474624(.data_in(wire_d46_23),.data_out(wire_d46_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474625(.data_in(wire_d46_24),.data_out(wire_d46_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474626(.data_in(wire_d46_25),.data_out(wire_d46_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474627(.data_in(wire_d46_26),.data_out(wire_d46_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474628(.data_in(wire_d46_27),.data_out(wire_d46_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474629(.data_in(wire_d46_28),.data_out(wire_d46_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474630(.data_in(wire_d46_29),.data_out(wire_d46_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474631(.data_in(wire_d46_30),.data_out(wire_d46_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474632(.data_in(wire_d46_31),.data_out(wire_d46_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474633(.data_in(wire_d46_32),.data_out(wire_d46_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474634(.data_in(wire_d46_33),.data_out(wire_d46_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474635(.data_in(wire_d46_34),.data_out(wire_d46_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474636(.data_in(wire_d46_35),.data_out(wire_d46_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474637(.data_in(wire_d46_36),.data_out(wire_d46_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474638(.data_in(wire_d46_37),.data_out(wire_d46_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474639(.data_in(wire_d46_38),.data_out(wire_d46_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474640(.data_in(wire_d46_39),.data_out(wire_d46_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474641(.data_in(wire_d46_40),.data_out(wire_d46_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474642(.data_in(wire_d46_41),.data_out(wire_d46_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474643(.data_in(wire_d46_42),.data_out(wire_d46_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474644(.data_in(wire_d46_43),.data_out(wire_d46_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474645(.data_in(wire_d46_44),.data_out(wire_d46_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474646(.data_in(wire_d46_45),.data_out(wire_d46_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474647(.data_in(wire_d46_46),.data_out(wire_d46_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474648(.data_in(wire_d46_47),.data_out(wire_d46_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474649(.data_in(wire_d46_48),.data_out(wire_d46_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474650(.data_in(wire_d46_49),.data_out(wire_d46_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474651(.data_in(wire_d46_50),.data_out(wire_d46_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474652(.data_in(wire_d46_51),.data_out(wire_d46_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474653(.data_in(wire_d46_52),.data_out(wire_d46_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474654(.data_in(wire_d46_53),.data_out(wire_d46_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474655(.data_in(wire_d46_54),.data_out(wire_d46_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474656(.data_in(wire_d46_55),.data_out(wire_d46_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474657(.data_in(wire_d46_56),.data_out(wire_d46_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474658(.data_in(wire_d46_57),.data_out(wire_d46_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474659(.data_in(wire_d46_58),.data_out(wire_d46_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474660(.data_in(wire_d46_59),.data_out(wire_d46_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474661(.data_in(wire_d46_60),.data_out(wire_d46_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474662(.data_in(wire_d46_61),.data_out(wire_d46_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474663(.data_in(wire_d46_62),.data_out(wire_d46_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474664(.data_in(wire_d46_63),.data_out(wire_d46_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474665(.data_in(wire_d46_64),.data_out(wire_d46_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474666(.data_in(wire_d46_65),.data_out(wire_d46_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474667(.data_in(wire_d46_66),.data_out(wire_d46_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474668(.data_in(wire_d46_67),.data_out(wire_d46_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474669(.data_in(wire_d46_68),.data_out(wire_d46_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474670(.data_in(wire_d46_69),.data_out(wire_d46_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474671(.data_in(wire_d46_70),.data_out(wire_d46_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474672(.data_in(wire_d46_71),.data_out(wire_d46_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474673(.data_in(wire_d46_72),.data_out(wire_d46_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474674(.data_in(wire_d46_73),.data_out(wire_d46_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474675(.data_in(wire_d46_74),.data_out(wire_d46_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474676(.data_in(wire_d46_75),.data_out(wire_d46_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474677(.data_in(wire_d46_76),.data_out(wire_d46_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474678(.data_in(wire_d46_77),.data_out(wire_d46_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474679(.data_in(wire_d46_78),.data_out(wire_d46_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474680(.data_in(wire_d46_79),.data_out(wire_d46_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474681(.data_in(wire_d46_80),.data_out(wire_d46_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474682(.data_in(wire_d46_81),.data_out(wire_d46_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474683(.data_in(wire_d46_82),.data_out(wire_d46_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474684(.data_in(wire_d46_83),.data_out(wire_d46_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474685(.data_in(wire_d46_84),.data_out(wire_d46_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474686(.data_in(wire_d46_85),.data_out(wire_d46_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474687(.data_in(wire_d46_86),.data_out(wire_d46_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474688(.data_in(wire_d46_87),.data_out(wire_d46_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474689(.data_in(wire_d46_88),.data_out(wire_d46_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474690(.data_in(wire_d46_89),.data_out(wire_d46_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474691(.data_in(wire_d46_90),.data_out(wire_d46_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474692(.data_in(wire_d46_91),.data_out(wire_d46_92),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474693(.data_in(wire_d46_92),.data_out(wire_d46_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474694(.data_in(wire_d46_93),.data_out(wire_d46_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474695(.data_in(wire_d46_94),.data_out(wire_d46_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474696(.data_in(wire_d46_95),.data_out(wire_d46_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474697(.data_in(wire_d46_96),.data_out(wire_d46_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474698(.data_in(wire_d46_97),.data_out(wire_d46_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474699(.data_in(wire_d46_98),.data_out(d_out46),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance48470(.data_in(d_in47),.data_out(wire_d47_0),.clk(clk),.rst(rst));            //channel 48
	register #(.WIDTH(WIDTH)) register_instance48471(.data_in(wire_d47_0),.data_out(wire_d47_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance48472(.data_in(wire_d47_1),.data_out(wire_d47_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance48473(.data_in(wire_d47_2),.data_out(wire_d47_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance48474(.data_in(wire_d47_3),.data_out(wire_d47_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance48475(.data_in(wire_d47_4),.data_out(wire_d47_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance48476(.data_in(wire_d47_5),.data_out(wire_d47_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance48477(.data_in(wire_d47_6),.data_out(wire_d47_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance48478(.data_in(wire_d47_7),.data_out(wire_d47_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance48479(.data_in(wire_d47_8),.data_out(wire_d47_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484710(.data_in(wire_d47_9),.data_out(wire_d47_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484711(.data_in(wire_d47_10),.data_out(wire_d47_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484712(.data_in(wire_d47_11),.data_out(wire_d47_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484713(.data_in(wire_d47_12),.data_out(wire_d47_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484714(.data_in(wire_d47_13),.data_out(wire_d47_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484715(.data_in(wire_d47_14),.data_out(wire_d47_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484716(.data_in(wire_d47_15),.data_out(wire_d47_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484717(.data_in(wire_d47_16),.data_out(wire_d47_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484718(.data_in(wire_d47_17),.data_out(wire_d47_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484719(.data_in(wire_d47_18),.data_out(wire_d47_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484720(.data_in(wire_d47_19),.data_out(wire_d47_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484721(.data_in(wire_d47_20),.data_out(wire_d47_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484722(.data_in(wire_d47_21),.data_out(wire_d47_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484723(.data_in(wire_d47_22),.data_out(wire_d47_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484724(.data_in(wire_d47_23),.data_out(wire_d47_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484725(.data_in(wire_d47_24),.data_out(wire_d47_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484726(.data_in(wire_d47_25),.data_out(wire_d47_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484727(.data_in(wire_d47_26),.data_out(wire_d47_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484728(.data_in(wire_d47_27),.data_out(wire_d47_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484729(.data_in(wire_d47_28),.data_out(wire_d47_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484730(.data_in(wire_d47_29),.data_out(wire_d47_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484731(.data_in(wire_d47_30),.data_out(wire_d47_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484732(.data_in(wire_d47_31),.data_out(wire_d47_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484733(.data_in(wire_d47_32),.data_out(wire_d47_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484734(.data_in(wire_d47_33),.data_out(wire_d47_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484735(.data_in(wire_d47_34),.data_out(wire_d47_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484736(.data_in(wire_d47_35),.data_out(wire_d47_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484737(.data_in(wire_d47_36),.data_out(wire_d47_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484738(.data_in(wire_d47_37),.data_out(wire_d47_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484739(.data_in(wire_d47_38),.data_out(wire_d47_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484740(.data_in(wire_d47_39),.data_out(wire_d47_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484741(.data_in(wire_d47_40),.data_out(wire_d47_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484742(.data_in(wire_d47_41),.data_out(wire_d47_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484743(.data_in(wire_d47_42),.data_out(wire_d47_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484744(.data_in(wire_d47_43),.data_out(wire_d47_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484745(.data_in(wire_d47_44),.data_out(wire_d47_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484746(.data_in(wire_d47_45),.data_out(wire_d47_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484747(.data_in(wire_d47_46),.data_out(wire_d47_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484748(.data_in(wire_d47_47),.data_out(wire_d47_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484749(.data_in(wire_d47_48),.data_out(wire_d47_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484750(.data_in(wire_d47_49),.data_out(wire_d47_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484751(.data_in(wire_d47_50),.data_out(wire_d47_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484752(.data_in(wire_d47_51),.data_out(wire_d47_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484753(.data_in(wire_d47_52),.data_out(wire_d47_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484754(.data_in(wire_d47_53),.data_out(wire_d47_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484755(.data_in(wire_d47_54),.data_out(wire_d47_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484756(.data_in(wire_d47_55),.data_out(wire_d47_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484757(.data_in(wire_d47_56),.data_out(wire_d47_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484758(.data_in(wire_d47_57),.data_out(wire_d47_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484759(.data_in(wire_d47_58),.data_out(wire_d47_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484760(.data_in(wire_d47_59),.data_out(wire_d47_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484761(.data_in(wire_d47_60),.data_out(wire_d47_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484762(.data_in(wire_d47_61),.data_out(wire_d47_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484763(.data_in(wire_d47_62),.data_out(wire_d47_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484764(.data_in(wire_d47_63),.data_out(wire_d47_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484765(.data_in(wire_d47_64),.data_out(wire_d47_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484766(.data_in(wire_d47_65),.data_out(wire_d47_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484767(.data_in(wire_d47_66),.data_out(wire_d47_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484768(.data_in(wire_d47_67),.data_out(wire_d47_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484769(.data_in(wire_d47_68),.data_out(wire_d47_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484770(.data_in(wire_d47_69),.data_out(wire_d47_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484771(.data_in(wire_d47_70),.data_out(wire_d47_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484772(.data_in(wire_d47_71),.data_out(wire_d47_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484773(.data_in(wire_d47_72),.data_out(wire_d47_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484774(.data_in(wire_d47_73),.data_out(wire_d47_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484775(.data_in(wire_d47_74),.data_out(wire_d47_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484776(.data_in(wire_d47_75),.data_out(wire_d47_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484777(.data_in(wire_d47_76),.data_out(wire_d47_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484778(.data_in(wire_d47_77),.data_out(wire_d47_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484779(.data_in(wire_d47_78),.data_out(wire_d47_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484780(.data_in(wire_d47_79),.data_out(wire_d47_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484781(.data_in(wire_d47_80),.data_out(wire_d47_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484782(.data_in(wire_d47_81),.data_out(wire_d47_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484783(.data_in(wire_d47_82),.data_out(wire_d47_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484784(.data_in(wire_d47_83),.data_out(wire_d47_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484785(.data_in(wire_d47_84),.data_out(wire_d47_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484786(.data_in(wire_d47_85),.data_out(wire_d47_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484787(.data_in(wire_d47_86),.data_out(wire_d47_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484788(.data_in(wire_d47_87),.data_out(wire_d47_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484789(.data_in(wire_d47_88),.data_out(wire_d47_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484790(.data_in(wire_d47_89),.data_out(wire_d47_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484791(.data_in(wire_d47_90),.data_out(wire_d47_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484792(.data_in(wire_d47_91),.data_out(wire_d47_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484793(.data_in(wire_d47_92),.data_out(wire_d47_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484794(.data_in(wire_d47_93),.data_out(wire_d47_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484795(.data_in(wire_d47_94),.data_out(wire_d47_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484796(.data_in(wire_d47_95),.data_out(wire_d47_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484797(.data_in(wire_d47_96),.data_out(wire_d47_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484798(.data_in(wire_d47_97),.data_out(wire_d47_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484799(.data_in(wire_d47_98),.data_out(d_out47),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance49480(.data_in(d_in48),.data_out(wire_d48_0),.clk(clk),.rst(rst));            //channel 49
	register #(.WIDTH(WIDTH)) register_instance49481(.data_in(wire_d48_0),.data_out(wire_d48_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance49482(.data_in(wire_d48_1),.data_out(wire_d48_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance49483(.data_in(wire_d48_2),.data_out(wire_d48_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance49484(.data_in(wire_d48_3),.data_out(wire_d48_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance49485(.data_in(wire_d48_4),.data_out(wire_d48_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance49486(.data_in(wire_d48_5),.data_out(wire_d48_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance49487(.data_in(wire_d48_6),.data_out(wire_d48_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance49488(.data_in(wire_d48_7),.data_out(wire_d48_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance49489(.data_in(wire_d48_8),.data_out(wire_d48_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494810(.data_in(wire_d48_9),.data_out(wire_d48_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494811(.data_in(wire_d48_10),.data_out(wire_d48_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494812(.data_in(wire_d48_11),.data_out(wire_d48_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494813(.data_in(wire_d48_12),.data_out(wire_d48_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494814(.data_in(wire_d48_13),.data_out(wire_d48_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494815(.data_in(wire_d48_14),.data_out(wire_d48_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494816(.data_in(wire_d48_15),.data_out(wire_d48_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494817(.data_in(wire_d48_16),.data_out(wire_d48_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494818(.data_in(wire_d48_17),.data_out(wire_d48_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494819(.data_in(wire_d48_18),.data_out(wire_d48_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494820(.data_in(wire_d48_19),.data_out(wire_d48_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494821(.data_in(wire_d48_20),.data_out(wire_d48_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494822(.data_in(wire_d48_21),.data_out(wire_d48_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494823(.data_in(wire_d48_22),.data_out(wire_d48_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494824(.data_in(wire_d48_23),.data_out(wire_d48_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494825(.data_in(wire_d48_24),.data_out(wire_d48_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494826(.data_in(wire_d48_25),.data_out(wire_d48_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494827(.data_in(wire_d48_26),.data_out(wire_d48_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494828(.data_in(wire_d48_27),.data_out(wire_d48_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494829(.data_in(wire_d48_28),.data_out(wire_d48_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494830(.data_in(wire_d48_29),.data_out(wire_d48_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494831(.data_in(wire_d48_30),.data_out(wire_d48_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494832(.data_in(wire_d48_31),.data_out(wire_d48_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494833(.data_in(wire_d48_32),.data_out(wire_d48_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494834(.data_in(wire_d48_33),.data_out(wire_d48_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494835(.data_in(wire_d48_34),.data_out(wire_d48_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494836(.data_in(wire_d48_35),.data_out(wire_d48_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494837(.data_in(wire_d48_36),.data_out(wire_d48_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494838(.data_in(wire_d48_37),.data_out(wire_d48_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494839(.data_in(wire_d48_38),.data_out(wire_d48_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494840(.data_in(wire_d48_39),.data_out(wire_d48_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494841(.data_in(wire_d48_40),.data_out(wire_d48_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494842(.data_in(wire_d48_41),.data_out(wire_d48_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494843(.data_in(wire_d48_42),.data_out(wire_d48_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494844(.data_in(wire_d48_43),.data_out(wire_d48_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494845(.data_in(wire_d48_44),.data_out(wire_d48_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494846(.data_in(wire_d48_45),.data_out(wire_d48_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494847(.data_in(wire_d48_46),.data_out(wire_d48_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494848(.data_in(wire_d48_47),.data_out(wire_d48_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494849(.data_in(wire_d48_48),.data_out(wire_d48_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494850(.data_in(wire_d48_49),.data_out(wire_d48_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494851(.data_in(wire_d48_50),.data_out(wire_d48_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494852(.data_in(wire_d48_51),.data_out(wire_d48_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494853(.data_in(wire_d48_52),.data_out(wire_d48_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494854(.data_in(wire_d48_53),.data_out(wire_d48_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494855(.data_in(wire_d48_54),.data_out(wire_d48_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494856(.data_in(wire_d48_55),.data_out(wire_d48_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494857(.data_in(wire_d48_56),.data_out(wire_d48_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494858(.data_in(wire_d48_57),.data_out(wire_d48_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494859(.data_in(wire_d48_58),.data_out(wire_d48_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494860(.data_in(wire_d48_59),.data_out(wire_d48_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494861(.data_in(wire_d48_60),.data_out(wire_d48_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494862(.data_in(wire_d48_61),.data_out(wire_d48_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494863(.data_in(wire_d48_62),.data_out(wire_d48_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494864(.data_in(wire_d48_63),.data_out(wire_d48_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494865(.data_in(wire_d48_64),.data_out(wire_d48_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494866(.data_in(wire_d48_65),.data_out(wire_d48_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494867(.data_in(wire_d48_66),.data_out(wire_d48_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494868(.data_in(wire_d48_67),.data_out(wire_d48_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494869(.data_in(wire_d48_68),.data_out(wire_d48_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494870(.data_in(wire_d48_69),.data_out(wire_d48_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494871(.data_in(wire_d48_70),.data_out(wire_d48_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494872(.data_in(wire_d48_71),.data_out(wire_d48_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494873(.data_in(wire_d48_72),.data_out(wire_d48_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494874(.data_in(wire_d48_73),.data_out(wire_d48_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494875(.data_in(wire_d48_74),.data_out(wire_d48_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494876(.data_in(wire_d48_75),.data_out(wire_d48_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494877(.data_in(wire_d48_76),.data_out(wire_d48_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494878(.data_in(wire_d48_77),.data_out(wire_d48_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494879(.data_in(wire_d48_78),.data_out(wire_d48_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494880(.data_in(wire_d48_79),.data_out(wire_d48_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494881(.data_in(wire_d48_80),.data_out(wire_d48_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494882(.data_in(wire_d48_81),.data_out(wire_d48_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494883(.data_in(wire_d48_82),.data_out(wire_d48_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494884(.data_in(wire_d48_83),.data_out(wire_d48_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494885(.data_in(wire_d48_84),.data_out(wire_d48_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494886(.data_in(wire_d48_85),.data_out(wire_d48_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494887(.data_in(wire_d48_86),.data_out(wire_d48_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494888(.data_in(wire_d48_87),.data_out(wire_d48_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494889(.data_in(wire_d48_88),.data_out(wire_d48_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494890(.data_in(wire_d48_89),.data_out(wire_d48_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494891(.data_in(wire_d48_90),.data_out(wire_d48_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494892(.data_in(wire_d48_91),.data_out(wire_d48_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494893(.data_in(wire_d48_92),.data_out(wire_d48_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494894(.data_in(wire_d48_93),.data_out(wire_d48_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494895(.data_in(wire_d48_94),.data_out(wire_d48_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494896(.data_in(wire_d48_95),.data_out(wire_d48_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494897(.data_in(wire_d48_96),.data_out(wire_d48_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494898(.data_in(wire_d48_97),.data_out(wire_d48_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494899(.data_in(wire_d48_98),.data_out(d_out48),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance50490(.data_in(d_in49),.data_out(wire_d49_0),.clk(clk),.rst(rst));            //channel 50
	large_mux #(.WIDTH(WIDTH)) large_mux_instance50491(.data_in(wire_d49_0),.data_out(wire_d49_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance50492(.data_in(wire_d49_1),.data_out(wire_d49_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance50493(.data_in(wire_d49_2),.data_out(wire_d49_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance50494(.data_in(wire_d49_3),.data_out(wire_d49_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance50495(.data_in(wire_d49_4),.data_out(wire_d49_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance50496(.data_in(wire_d49_5),.data_out(wire_d49_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance50497(.data_in(wire_d49_6),.data_out(wire_d49_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance50498(.data_in(wire_d49_7),.data_out(wire_d49_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance50499(.data_in(wire_d49_8),.data_out(wire_d49_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504910(.data_in(wire_d49_9),.data_out(wire_d49_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504911(.data_in(wire_d49_10),.data_out(wire_d49_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504912(.data_in(wire_d49_11),.data_out(wire_d49_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504913(.data_in(wire_d49_12),.data_out(wire_d49_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504914(.data_in(wire_d49_13),.data_out(wire_d49_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504915(.data_in(wire_d49_14),.data_out(wire_d49_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504916(.data_in(wire_d49_15),.data_out(wire_d49_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504917(.data_in(wire_d49_16),.data_out(wire_d49_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504918(.data_in(wire_d49_17),.data_out(wire_d49_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504919(.data_in(wire_d49_18),.data_out(wire_d49_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504920(.data_in(wire_d49_19),.data_out(wire_d49_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504921(.data_in(wire_d49_20),.data_out(wire_d49_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504922(.data_in(wire_d49_21),.data_out(wire_d49_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504923(.data_in(wire_d49_22),.data_out(wire_d49_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504924(.data_in(wire_d49_23),.data_out(wire_d49_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504925(.data_in(wire_d49_24),.data_out(wire_d49_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504926(.data_in(wire_d49_25),.data_out(wire_d49_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504927(.data_in(wire_d49_26),.data_out(wire_d49_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504928(.data_in(wire_d49_27),.data_out(wire_d49_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504929(.data_in(wire_d49_28),.data_out(wire_d49_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504930(.data_in(wire_d49_29),.data_out(wire_d49_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504931(.data_in(wire_d49_30),.data_out(wire_d49_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504932(.data_in(wire_d49_31),.data_out(wire_d49_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504933(.data_in(wire_d49_32),.data_out(wire_d49_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504934(.data_in(wire_d49_33),.data_out(wire_d49_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504935(.data_in(wire_d49_34),.data_out(wire_d49_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504936(.data_in(wire_d49_35),.data_out(wire_d49_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504937(.data_in(wire_d49_36),.data_out(wire_d49_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504938(.data_in(wire_d49_37),.data_out(wire_d49_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504939(.data_in(wire_d49_38),.data_out(wire_d49_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504940(.data_in(wire_d49_39),.data_out(wire_d49_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504941(.data_in(wire_d49_40),.data_out(wire_d49_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504942(.data_in(wire_d49_41),.data_out(wire_d49_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504943(.data_in(wire_d49_42),.data_out(wire_d49_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504944(.data_in(wire_d49_43),.data_out(wire_d49_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504945(.data_in(wire_d49_44),.data_out(wire_d49_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504946(.data_in(wire_d49_45),.data_out(wire_d49_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504947(.data_in(wire_d49_46),.data_out(wire_d49_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504948(.data_in(wire_d49_47),.data_out(wire_d49_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504949(.data_in(wire_d49_48),.data_out(wire_d49_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504950(.data_in(wire_d49_49),.data_out(wire_d49_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504951(.data_in(wire_d49_50),.data_out(wire_d49_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504952(.data_in(wire_d49_51),.data_out(wire_d49_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504953(.data_in(wire_d49_52),.data_out(wire_d49_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504954(.data_in(wire_d49_53),.data_out(wire_d49_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504955(.data_in(wire_d49_54),.data_out(wire_d49_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504956(.data_in(wire_d49_55),.data_out(wire_d49_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504957(.data_in(wire_d49_56),.data_out(wire_d49_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504958(.data_in(wire_d49_57),.data_out(wire_d49_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504959(.data_in(wire_d49_58),.data_out(wire_d49_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504960(.data_in(wire_d49_59),.data_out(wire_d49_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504961(.data_in(wire_d49_60),.data_out(wire_d49_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504962(.data_in(wire_d49_61),.data_out(wire_d49_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504963(.data_in(wire_d49_62),.data_out(wire_d49_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504964(.data_in(wire_d49_63),.data_out(wire_d49_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504965(.data_in(wire_d49_64),.data_out(wire_d49_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504966(.data_in(wire_d49_65),.data_out(wire_d49_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504967(.data_in(wire_d49_66),.data_out(wire_d49_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504968(.data_in(wire_d49_67),.data_out(wire_d49_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504969(.data_in(wire_d49_68),.data_out(wire_d49_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504970(.data_in(wire_d49_69),.data_out(wire_d49_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504971(.data_in(wire_d49_70),.data_out(wire_d49_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504972(.data_in(wire_d49_71),.data_out(wire_d49_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504973(.data_in(wire_d49_72),.data_out(wire_d49_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504974(.data_in(wire_d49_73),.data_out(wire_d49_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504975(.data_in(wire_d49_74),.data_out(wire_d49_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504976(.data_in(wire_d49_75),.data_out(wire_d49_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504977(.data_in(wire_d49_76),.data_out(wire_d49_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504978(.data_in(wire_d49_77),.data_out(wire_d49_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504979(.data_in(wire_d49_78),.data_out(wire_d49_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504980(.data_in(wire_d49_79),.data_out(wire_d49_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504981(.data_in(wire_d49_80),.data_out(wire_d49_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504982(.data_in(wire_d49_81),.data_out(wire_d49_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504983(.data_in(wire_d49_82),.data_out(wire_d49_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504984(.data_in(wire_d49_83),.data_out(wire_d49_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504985(.data_in(wire_d49_84),.data_out(wire_d49_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504986(.data_in(wire_d49_85),.data_out(wire_d49_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504987(.data_in(wire_d49_86),.data_out(wire_d49_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504988(.data_in(wire_d49_87),.data_out(wire_d49_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504989(.data_in(wire_d49_88),.data_out(wire_d49_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504990(.data_in(wire_d49_89),.data_out(wire_d49_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504991(.data_in(wire_d49_90),.data_out(wire_d49_91),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504992(.data_in(wire_d49_91),.data_out(wire_d49_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504993(.data_in(wire_d49_92),.data_out(wire_d49_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504994(.data_in(wire_d49_93),.data_out(wire_d49_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504995(.data_in(wire_d49_94),.data_out(wire_d49_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504996(.data_in(wire_d49_95),.data_out(wire_d49_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504997(.data_in(wire_d49_96),.data_out(wire_d49_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504998(.data_in(wire_d49_97),.data_out(wire_d49_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504999(.data_in(wire_d49_98),.data_out(d_out49),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance51500(.data_in(d_in50),.data_out(wire_d50_0),.clk(clk),.rst(rst));            //channel 51
	large_mux #(.WIDTH(WIDTH)) large_mux_instance51501(.data_in(wire_d50_0),.data_out(wire_d50_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance51502(.data_in(wire_d50_1),.data_out(wire_d50_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance51503(.data_in(wire_d50_2),.data_out(wire_d50_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance51504(.data_in(wire_d50_3),.data_out(wire_d50_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance51505(.data_in(wire_d50_4),.data_out(wire_d50_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance51506(.data_in(wire_d50_5),.data_out(wire_d50_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance51507(.data_in(wire_d50_6),.data_out(wire_d50_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance51508(.data_in(wire_d50_7),.data_out(wire_d50_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance51509(.data_in(wire_d50_8),.data_out(wire_d50_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515010(.data_in(wire_d50_9),.data_out(wire_d50_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515011(.data_in(wire_d50_10),.data_out(wire_d50_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515012(.data_in(wire_d50_11),.data_out(wire_d50_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance515013(.data_in(wire_d50_12),.data_out(wire_d50_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515014(.data_in(wire_d50_13),.data_out(wire_d50_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515015(.data_in(wire_d50_14),.data_out(wire_d50_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515016(.data_in(wire_d50_15),.data_out(wire_d50_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515017(.data_in(wire_d50_16),.data_out(wire_d50_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515018(.data_in(wire_d50_17),.data_out(wire_d50_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515019(.data_in(wire_d50_18),.data_out(wire_d50_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515020(.data_in(wire_d50_19),.data_out(wire_d50_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515021(.data_in(wire_d50_20),.data_out(wire_d50_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance515022(.data_in(wire_d50_21),.data_out(wire_d50_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515023(.data_in(wire_d50_22),.data_out(wire_d50_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance515024(.data_in(wire_d50_23),.data_out(wire_d50_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance515025(.data_in(wire_d50_24),.data_out(wire_d50_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515026(.data_in(wire_d50_25),.data_out(wire_d50_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance515027(.data_in(wire_d50_26),.data_out(wire_d50_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515028(.data_in(wire_d50_27),.data_out(wire_d50_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515029(.data_in(wire_d50_28),.data_out(wire_d50_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance515030(.data_in(wire_d50_29),.data_out(wire_d50_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515031(.data_in(wire_d50_30),.data_out(wire_d50_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515032(.data_in(wire_d50_31),.data_out(wire_d50_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance515033(.data_in(wire_d50_32),.data_out(wire_d50_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515034(.data_in(wire_d50_33),.data_out(wire_d50_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515035(.data_in(wire_d50_34),.data_out(wire_d50_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515036(.data_in(wire_d50_35),.data_out(wire_d50_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515037(.data_in(wire_d50_36),.data_out(wire_d50_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515038(.data_in(wire_d50_37),.data_out(wire_d50_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515039(.data_in(wire_d50_38),.data_out(wire_d50_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515040(.data_in(wire_d50_39),.data_out(wire_d50_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515041(.data_in(wire_d50_40),.data_out(wire_d50_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515042(.data_in(wire_d50_41),.data_out(wire_d50_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515043(.data_in(wire_d50_42),.data_out(wire_d50_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance515044(.data_in(wire_d50_43),.data_out(wire_d50_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515045(.data_in(wire_d50_44),.data_out(wire_d50_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515046(.data_in(wire_d50_45),.data_out(wire_d50_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance515047(.data_in(wire_d50_46),.data_out(wire_d50_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515048(.data_in(wire_d50_47),.data_out(wire_d50_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance515049(.data_in(wire_d50_48),.data_out(wire_d50_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance515050(.data_in(wire_d50_49),.data_out(wire_d50_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515051(.data_in(wire_d50_50),.data_out(wire_d50_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515052(.data_in(wire_d50_51),.data_out(wire_d50_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance515053(.data_in(wire_d50_52),.data_out(wire_d50_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515054(.data_in(wire_d50_53),.data_out(wire_d50_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515055(.data_in(wire_d50_54),.data_out(wire_d50_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance515056(.data_in(wire_d50_55),.data_out(wire_d50_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515057(.data_in(wire_d50_56),.data_out(wire_d50_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515058(.data_in(wire_d50_57),.data_out(wire_d50_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance515059(.data_in(wire_d50_58),.data_out(wire_d50_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance515060(.data_in(wire_d50_59),.data_out(wire_d50_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515061(.data_in(wire_d50_60),.data_out(wire_d50_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515062(.data_in(wire_d50_61),.data_out(wire_d50_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515063(.data_in(wire_d50_62),.data_out(wire_d50_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515064(.data_in(wire_d50_63),.data_out(wire_d50_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515065(.data_in(wire_d50_64),.data_out(wire_d50_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515066(.data_in(wire_d50_65),.data_out(wire_d50_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515067(.data_in(wire_d50_66),.data_out(wire_d50_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance515068(.data_in(wire_d50_67),.data_out(wire_d50_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance515069(.data_in(wire_d50_68),.data_out(wire_d50_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515070(.data_in(wire_d50_69),.data_out(wire_d50_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance515071(.data_in(wire_d50_70),.data_out(wire_d50_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515072(.data_in(wire_d50_71),.data_out(wire_d50_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515073(.data_in(wire_d50_72),.data_out(wire_d50_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515074(.data_in(wire_d50_73),.data_out(wire_d50_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515075(.data_in(wire_d50_74),.data_out(wire_d50_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515076(.data_in(wire_d50_75),.data_out(wire_d50_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515077(.data_in(wire_d50_76),.data_out(wire_d50_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515078(.data_in(wire_d50_77),.data_out(wire_d50_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515079(.data_in(wire_d50_78),.data_out(wire_d50_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515080(.data_in(wire_d50_79),.data_out(wire_d50_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515081(.data_in(wire_d50_80),.data_out(wire_d50_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515082(.data_in(wire_d50_81),.data_out(wire_d50_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515083(.data_in(wire_d50_82),.data_out(wire_d50_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515084(.data_in(wire_d50_83),.data_out(wire_d50_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515085(.data_in(wire_d50_84),.data_out(wire_d50_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515086(.data_in(wire_d50_85),.data_out(wire_d50_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515087(.data_in(wire_d50_86),.data_out(wire_d50_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance515088(.data_in(wire_d50_87),.data_out(wire_d50_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance515089(.data_in(wire_d50_88),.data_out(wire_d50_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515090(.data_in(wire_d50_89),.data_out(wire_d50_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515091(.data_in(wire_d50_90),.data_out(wire_d50_91),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance515092(.data_in(wire_d50_91),.data_out(wire_d50_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515093(.data_in(wire_d50_92),.data_out(wire_d50_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515094(.data_in(wire_d50_93),.data_out(wire_d50_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515095(.data_in(wire_d50_94),.data_out(wire_d50_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance515096(.data_in(wire_d50_95),.data_out(wire_d50_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515097(.data_in(wire_d50_96),.data_out(wire_d50_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515098(.data_in(wire_d50_97),.data_out(wire_d50_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance515099(.data_in(wire_d50_98),.data_out(d_out50),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance52510(.data_in(d_in51),.data_out(wire_d51_0),.clk(clk),.rst(rst));            //channel 52
	large_mux #(.WIDTH(WIDTH)) large_mux_instance52511(.data_in(wire_d51_0),.data_out(wire_d51_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance52512(.data_in(wire_d51_1),.data_out(wire_d51_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance52513(.data_in(wire_d51_2),.data_out(wire_d51_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance52514(.data_in(wire_d51_3),.data_out(wire_d51_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance52515(.data_in(wire_d51_4),.data_out(wire_d51_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance52516(.data_in(wire_d51_5),.data_out(wire_d51_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance52517(.data_in(wire_d51_6),.data_out(wire_d51_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance52518(.data_in(wire_d51_7),.data_out(wire_d51_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance52519(.data_in(wire_d51_8),.data_out(wire_d51_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525110(.data_in(wire_d51_9),.data_out(wire_d51_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525111(.data_in(wire_d51_10),.data_out(wire_d51_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525112(.data_in(wire_d51_11),.data_out(wire_d51_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance525113(.data_in(wire_d51_12),.data_out(wire_d51_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525114(.data_in(wire_d51_13),.data_out(wire_d51_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance525115(.data_in(wire_d51_14),.data_out(wire_d51_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525116(.data_in(wire_d51_15),.data_out(wire_d51_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance525117(.data_in(wire_d51_16),.data_out(wire_d51_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance525118(.data_in(wire_d51_17),.data_out(wire_d51_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525119(.data_in(wire_d51_18),.data_out(wire_d51_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525120(.data_in(wire_d51_19),.data_out(wire_d51_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance525121(.data_in(wire_d51_20),.data_out(wire_d51_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525122(.data_in(wire_d51_21),.data_out(wire_d51_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525123(.data_in(wire_d51_22),.data_out(wire_d51_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525124(.data_in(wire_d51_23),.data_out(wire_d51_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525125(.data_in(wire_d51_24),.data_out(wire_d51_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525126(.data_in(wire_d51_25),.data_out(wire_d51_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance525127(.data_in(wire_d51_26),.data_out(wire_d51_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525128(.data_in(wire_d51_27),.data_out(wire_d51_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525129(.data_in(wire_d51_28),.data_out(wire_d51_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525130(.data_in(wire_d51_29),.data_out(wire_d51_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525131(.data_in(wire_d51_30),.data_out(wire_d51_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525132(.data_in(wire_d51_31),.data_out(wire_d51_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525133(.data_in(wire_d51_32),.data_out(wire_d51_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525134(.data_in(wire_d51_33),.data_out(wire_d51_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525135(.data_in(wire_d51_34),.data_out(wire_d51_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525136(.data_in(wire_d51_35),.data_out(wire_d51_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525137(.data_in(wire_d51_36),.data_out(wire_d51_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525138(.data_in(wire_d51_37),.data_out(wire_d51_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance525139(.data_in(wire_d51_38),.data_out(wire_d51_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525140(.data_in(wire_d51_39),.data_out(wire_d51_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525141(.data_in(wire_d51_40),.data_out(wire_d51_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525142(.data_in(wire_d51_41),.data_out(wire_d51_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525143(.data_in(wire_d51_42),.data_out(wire_d51_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525144(.data_in(wire_d51_43),.data_out(wire_d51_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525145(.data_in(wire_d51_44),.data_out(wire_d51_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525146(.data_in(wire_d51_45),.data_out(wire_d51_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance525147(.data_in(wire_d51_46),.data_out(wire_d51_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525148(.data_in(wire_d51_47),.data_out(wire_d51_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525149(.data_in(wire_d51_48),.data_out(wire_d51_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525150(.data_in(wire_d51_49),.data_out(wire_d51_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance525151(.data_in(wire_d51_50),.data_out(wire_d51_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525152(.data_in(wire_d51_51),.data_out(wire_d51_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525153(.data_in(wire_d51_52),.data_out(wire_d51_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance525154(.data_in(wire_d51_53),.data_out(wire_d51_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance525155(.data_in(wire_d51_54),.data_out(wire_d51_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525156(.data_in(wire_d51_55),.data_out(wire_d51_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525157(.data_in(wire_d51_56),.data_out(wire_d51_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525158(.data_in(wire_d51_57),.data_out(wire_d51_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance525159(.data_in(wire_d51_58),.data_out(wire_d51_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance525160(.data_in(wire_d51_59),.data_out(wire_d51_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525161(.data_in(wire_d51_60),.data_out(wire_d51_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525162(.data_in(wire_d51_61),.data_out(wire_d51_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525163(.data_in(wire_d51_62),.data_out(wire_d51_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525164(.data_in(wire_d51_63),.data_out(wire_d51_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525165(.data_in(wire_d51_64),.data_out(wire_d51_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525166(.data_in(wire_d51_65),.data_out(wire_d51_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525167(.data_in(wire_d51_66),.data_out(wire_d51_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525168(.data_in(wire_d51_67),.data_out(wire_d51_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525169(.data_in(wire_d51_68),.data_out(wire_d51_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance525170(.data_in(wire_d51_69),.data_out(wire_d51_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525171(.data_in(wire_d51_70),.data_out(wire_d51_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525172(.data_in(wire_d51_71),.data_out(wire_d51_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance525173(.data_in(wire_d51_72),.data_out(wire_d51_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525174(.data_in(wire_d51_73),.data_out(wire_d51_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525175(.data_in(wire_d51_74),.data_out(wire_d51_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525176(.data_in(wire_d51_75),.data_out(wire_d51_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525177(.data_in(wire_d51_76),.data_out(wire_d51_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525178(.data_in(wire_d51_77),.data_out(wire_d51_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525179(.data_in(wire_d51_78),.data_out(wire_d51_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525180(.data_in(wire_d51_79),.data_out(wire_d51_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525181(.data_in(wire_d51_80),.data_out(wire_d51_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525182(.data_in(wire_d51_81),.data_out(wire_d51_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance525183(.data_in(wire_d51_82),.data_out(wire_d51_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525184(.data_in(wire_d51_83),.data_out(wire_d51_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance525185(.data_in(wire_d51_84),.data_out(wire_d51_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525186(.data_in(wire_d51_85),.data_out(wire_d51_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525187(.data_in(wire_d51_86),.data_out(wire_d51_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525188(.data_in(wire_d51_87),.data_out(wire_d51_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525189(.data_in(wire_d51_88),.data_out(wire_d51_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance525190(.data_in(wire_d51_89),.data_out(wire_d51_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525191(.data_in(wire_d51_90),.data_out(wire_d51_91),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525192(.data_in(wire_d51_91),.data_out(wire_d51_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525193(.data_in(wire_d51_92),.data_out(wire_d51_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525194(.data_in(wire_d51_93),.data_out(wire_d51_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance525195(.data_in(wire_d51_94),.data_out(wire_d51_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525196(.data_in(wire_d51_95),.data_out(wire_d51_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance525197(.data_in(wire_d51_96),.data_out(wire_d51_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance525198(.data_in(wire_d51_97),.data_out(wire_d51_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance525199(.data_in(wire_d51_98),.data_out(d_out51),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance53520(.data_in(d_in52),.data_out(wire_d52_0),.clk(clk),.rst(rst));            //channel 53
	large_mux #(.WIDTH(WIDTH)) large_mux_instance53521(.data_in(wire_d52_0),.data_out(wire_d52_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance53522(.data_in(wire_d52_1),.data_out(wire_d52_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance53523(.data_in(wire_d52_2),.data_out(wire_d52_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance53524(.data_in(wire_d52_3),.data_out(wire_d52_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance53525(.data_in(wire_d52_4),.data_out(wire_d52_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance53526(.data_in(wire_d52_5),.data_out(wire_d52_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance53527(.data_in(wire_d52_6),.data_out(wire_d52_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance53528(.data_in(wire_d52_7),.data_out(wire_d52_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance53529(.data_in(wire_d52_8),.data_out(wire_d52_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535210(.data_in(wire_d52_9),.data_out(wire_d52_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535211(.data_in(wire_d52_10),.data_out(wire_d52_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535212(.data_in(wire_d52_11),.data_out(wire_d52_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535213(.data_in(wire_d52_12),.data_out(wire_d52_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance535214(.data_in(wire_d52_13),.data_out(wire_d52_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535215(.data_in(wire_d52_14),.data_out(wire_d52_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535216(.data_in(wire_d52_15),.data_out(wire_d52_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance535217(.data_in(wire_d52_16),.data_out(wire_d52_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance535218(.data_in(wire_d52_17),.data_out(wire_d52_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535219(.data_in(wire_d52_18),.data_out(wire_d52_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance535220(.data_in(wire_d52_19),.data_out(wire_d52_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance535221(.data_in(wire_d52_20),.data_out(wire_d52_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535222(.data_in(wire_d52_21),.data_out(wire_d52_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance535223(.data_in(wire_d52_22),.data_out(wire_d52_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535224(.data_in(wire_d52_23),.data_out(wire_d52_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance535225(.data_in(wire_d52_24),.data_out(wire_d52_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance535226(.data_in(wire_d52_25),.data_out(wire_d52_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance535227(.data_in(wire_d52_26),.data_out(wire_d52_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535228(.data_in(wire_d52_27),.data_out(wire_d52_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535229(.data_in(wire_d52_28),.data_out(wire_d52_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance535230(.data_in(wire_d52_29),.data_out(wire_d52_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535231(.data_in(wire_d52_30),.data_out(wire_d52_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535232(.data_in(wire_d52_31),.data_out(wire_d52_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535233(.data_in(wire_d52_32),.data_out(wire_d52_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance535234(.data_in(wire_d52_33),.data_out(wire_d52_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535235(.data_in(wire_d52_34),.data_out(wire_d52_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance535236(.data_in(wire_d52_35),.data_out(wire_d52_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance535237(.data_in(wire_d52_36),.data_out(wire_d52_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance535238(.data_in(wire_d52_37),.data_out(wire_d52_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance535239(.data_in(wire_d52_38),.data_out(wire_d52_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535240(.data_in(wire_d52_39),.data_out(wire_d52_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535241(.data_in(wire_d52_40),.data_out(wire_d52_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535242(.data_in(wire_d52_41),.data_out(wire_d52_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance535243(.data_in(wire_d52_42),.data_out(wire_d52_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance535244(.data_in(wire_d52_43),.data_out(wire_d52_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance535245(.data_in(wire_d52_44),.data_out(wire_d52_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535246(.data_in(wire_d52_45),.data_out(wire_d52_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance535247(.data_in(wire_d52_46),.data_out(wire_d52_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535248(.data_in(wire_d52_47),.data_out(wire_d52_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance535249(.data_in(wire_d52_48),.data_out(wire_d52_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance535250(.data_in(wire_d52_49),.data_out(wire_d52_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535251(.data_in(wire_d52_50),.data_out(wire_d52_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535252(.data_in(wire_d52_51),.data_out(wire_d52_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance535253(.data_in(wire_d52_52),.data_out(wire_d52_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance535254(.data_in(wire_d52_53),.data_out(wire_d52_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535255(.data_in(wire_d52_54),.data_out(wire_d52_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535256(.data_in(wire_d52_55),.data_out(wire_d52_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance535257(.data_in(wire_d52_56),.data_out(wire_d52_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535258(.data_in(wire_d52_57),.data_out(wire_d52_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535259(.data_in(wire_d52_58),.data_out(wire_d52_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance535260(.data_in(wire_d52_59),.data_out(wire_d52_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance535261(.data_in(wire_d52_60),.data_out(wire_d52_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535262(.data_in(wire_d52_61),.data_out(wire_d52_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance535263(.data_in(wire_d52_62),.data_out(wire_d52_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance535264(.data_in(wire_d52_63),.data_out(wire_d52_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance535265(.data_in(wire_d52_64),.data_out(wire_d52_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535266(.data_in(wire_d52_65),.data_out(wire_d52_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535267(.data_in(wire_d52_66),.data_out(wire_d52_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance535268(.data_in(wire_d52_67),.data_out(wire_d52_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance535269(.data_in(wire_d52_68),.data_out(wire_d52_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535270(.data_in(wire_d52_69),.data_out(wire_d52_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535271(.data_in(wire_d52_70),.data_out(wire_d52_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance535272(.data_in(wire_d52_71),.data_out(wire_d52_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535273(.data_in(wire_d52_72),.data_out(wire_d52_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance535274(.data_in(wire_d52_73),.data_out(wire_d52_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance535275(.data_in(wire_d52_74),.data_out(wire_d52_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535276(.data_in(wire_d52_75),.data_out(wire_d52_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535277(.data_in(wire_d52_76),.data_out(wire_d52_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535278(.data_in(wire_d52_77),.data_out(wire_d52_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535279(.data_in(wire_d52_78),.data_out(wire_d52_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535280(.data_in(wire_d52_79),.data_out(wire_d52_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance535281(.data_in(wire_d52_80),.data_out(wire_d52_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance535282(.data_in(wire_d52_81),.data_out(wire_d52_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535283(.data_in(wire_d52_82),.data_out(wire_d52_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535284(.data_in(wire_d52_83),.data_out(wire_d52_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance535285(.data_in(wire_d52_84),.data_out(wire_d52_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535286(.data_in(wire_d52_85),.data_out(wire_d52_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance535287(.data_in(wire_d52_86),.data_out(wire_d52_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535288(.data_in(wire_d52_87),.data_out(wire_d52_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535289(.data_in(wire_d52_88),.data_out(wire_d52_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance535290(.data_in(wire_d52_89),.data_out(wire_d52_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance535291(.data_in(wire_d52_90),.data_out(wire_d52_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535292(.data_in(wire_d52_91),.data_out(wire_d52_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535293(.data_in(wire_d52_92),.data_out(wire_d52_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance535294(.data_in(wire_d52_93),.data_out(wire_d52_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance535295(.data_in(wire_d52_94),.data_out(wire_d52_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535296(.data_in(wire_d52_95),.data_out(wire_d52_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance535297(.data_in(wire_d52_96),.data_out(wire_d52_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance535298(.data_in(wire_d52_97),.data_out(wire_d52_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance535299(.data_in(wire_d52_98),.data_out(d_out52),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance54530(.data_in(d_in53),.data_out(wire_d53_0),.clk(clk),.rst(rst));            //channel 54
	register #(.WIDTH(WIDTH)) register_instance54531(.data_in(wire_d53_0),.data_out(wire_d53_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance54532(.data_in(wire_d53_1),.data_out(wire_d53_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54533(.data_in(wire_d53_2),.data_out(wire_d53_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance54534(.data_in(wire_d53_3),.data_out(wire_d53_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance54535(.data_in(wire_d53_4),.data_out(wire_d53_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54536(.data_in(wire_d53_5),.data_out(wire_d53_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54537(.data_in(wire_d53_6),.data_out(wire_d53_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54538(.data_in(wire_d53_7),.data_out(wire_d53_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance54539(.data_in(wire_d53_8),.data_out(wire_d53_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545310(.data_in(wire_d53_9),.data_out(wire_d53_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545311(.data_in(wire_d53_10),.data_out(wire_d53_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545312(.data_in(wire_d53_11),.data_out(wire_d53_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545313(.data_in(wire_d53_12),.data_out(wire_d53_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545314(.data_in(wire_d53_13),.data_out(wire_d53_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545315(.data_in(wire_d53_14),.data_out(wire_d53_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545316(.data_in(wire_d53_15),.data_out(wire_d53_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545317(.data_in(wire_d53_16),.data_out(wire_d53_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545318(.data_in(wire_d53_17),.data_out(wire_d53_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545319(.data_in(wire_d53_18),.data_out(wire_d53_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545320(.data_in(wire_d53_19),.data_out(wire_d53_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545321(.data_in(wire_d53_20),.data_out(wire_d53_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545322(.data_in(wire_d53_21),.data_out(wire_d53_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545323(.data_in(wire_d53_22),.data_out(wire_d53_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545324(.data_in(wire_d53_23),.data_out(wire_d53_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545325(.data_in(wire_d53_24),.data_out(wire_d53_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545326(.data_in(wire_d53_25),.data_out(wire_d53_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545327(.data_in(wire_d53_26),.data_out(wire_d53_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545328(.data_in(wire_d53_27),.data_out(wire_d53_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545329(.data_in(wire_d53_28),.data_out(wire_d53_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545330(.data_in(wire_d53_29),.data_out(wire_d53_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545331(.data_in(wire_d53_30),.data_out(wire_d53_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545332(.data_in(wire_d53_31),.data_out(wire_d53_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545333(.data_in(wire_d53_32),.data_out(wire_d53_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545334(.data_in(wire_d53_33),.data_out(wire_d53_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545335(.data_in(wire_d53_34),.data_out(wire_d53_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545336(.data_in(wire_d53_35),.data_out(wire_d53_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545337(.data_in(wire_d53_36),.data_out(wire_d53_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545338(.data_in(wire_d53_37),.data_out(wire_d53_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545339(.data_in(wire_d53_38),.data_out(wire_d53_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545340(.data_in(wire_d53_39),.data_out(wire_d53_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545341(.data_in(wire_d53_40),.data_out(wire_d53_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545342(.data_in(wire_d53_41),.data_out(wire_d53_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545343(.data_in(wire_d53_42),.data_out(wire_d53_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545344(.data_in(wire_d53_43),.data_out(wire_d53_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545345(.data_in(wire_d53_44),.data_out(wire_d53_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545346(.data_in(wire_d53_45),.data_out(wire_d53_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545347(.data_in(wire_d53_46),.data_out(wire_d53_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545348(.data_in(wire_d53_47),.data_out(wire_d53_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545349(.data_in(wire_d53_48),.data_out(wire_d53_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545350(.data_in(wire_d53_49),.data_out(wire_d53_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545351(.data_in(wire_d53_50),.data_out(wire_d53_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545352(.data_in(wire_d53_51),.data_out(wire_d53_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545353(.data_in(wire_d53_52),.data_out(wire_d53_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545354(.data_in(wire_d53_53),.data_out(wire_d53_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545355(.data_in(wire_d53_54),.data_out(wire_d53_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545356(.data_in(wire_d53_55),.data_out(wire_d53_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545357(.data_in(wire_d53_56),.data_out(wire_d53_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545358(.data_in(wire_d53_57),.data_out(wire_d53_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545359(.data_in(wire_d53_58),.data_out(wire_d53_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545360(.data_in(wire_d53_59),.data_out(wire_d53_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545361(.data_in(wire_d53_60),.data_out(wire_d53_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545362(.data_in(wire_d53_61),.data_out(wire_d53_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545363(.data_in(wire_d53_62),.data_out(wire_d53_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545364(.data_in(wire_d53_63),.data_out(wire_d53_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545365(.data_in(wire_d53_64),.data_out(wire_d53_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545366(.data_in(wire_d53_65),.data_out(wire_d53_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545367(.data_in(wire_d53_66),.data_out(wire_d53_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545368(.data_in(wire_d53_67),.data_out(wire_d53_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545369(.data_in(wire_d53_68),.data_out(wire_d53_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545370(.data_in(wire_d53_69),.data_out(wire_d53_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545371(.data_in(wire_d53_70),.data_out(wire_d53_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545372(.data_in(wire_d53_71),.data_out(wire_d53_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545373(.data_in(wire_d53_72),.data_out(wire_d53_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545374(.data_in(wire_d53_73),.data_out(wire_d53_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545375(.data_in(wire_d53_74),.data_out(wire_d53_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545376(.data_in(wire_d53_75),.data_out(wire_d53_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545377(.data_in(wire_d53_76),.data_out(wire_d53_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545378(.data_in(wire_d53_77),.data_out(wire_d53_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545379(.data_in(wire_d53_78),.data_out(wire_d53_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545380(.data_in(wire_d53_79),.data_out(wire_d53_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545381(.data_in(wire_d53_80),.data_out(wire_d53_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545382(.data_in(wire_d53_81),.data_out(wire_d53_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545383(.data_in(wire_d53_82),.data_out(wire_d53_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545384(.data_in(wire_d53_83),.data_out(wire_d53_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545385(.data_in(wire_d53_84),.data_out(wire_d53_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545386(.data_in(wire_d53_85),.data_out(wire_d53_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545387(.data_in(wire_d53_86),.data_out(wire_d53_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545388(.data_in(wire_d53_87),.data_out(wire_d53_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545389(.data_in(wire_d53_88),.data_out(wire_d53_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545390(.data_in(wire_d53_89),.data_out(wire_d53_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545391(.data_in(wire_d53_90),.data_out(wire_d53_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545392(.data_in(wire_d53_91),.data_out(wire_d53_92),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545393(.data_in(wire_d53_92),.data_out(wire_d53_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545394(.data_in(wire_d53_93),.data_out(wire_d53_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545395(.data_in(wire_d53_94),.data_out(wire_d53_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545396(.data_in(wire_d53_95),.data_out(wire_d53_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545397(.data_in(wire_d53_96),.data_out(wire_d53_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545398(.data_in(wire_d53_97),.data_out(wire_d53_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance545399(.data_in(wire_d53_98),.data_out(d_out53),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance55540(.data_in(d_in54),.data_out(wire_d54_0),.clk(clk),.rst(rst));            //channel 55
	invertion #(.WIDTH(WIDTH)) invertion_instance55541(.data_in(wire_d54_0),.data_out(wire_d54_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance55542(.data_in(wire_d54_1),.data_out(wire_d54_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance55543(.data_in(wire_d54_2),.data_out(wire_d54_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance55544(.data_in(wire_d54_3),.data_out(wire_d54_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance55545(.data_in(wire_d54_4),.data_out(wire_d54_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance55546(.data_in(wire_d54_5),.data_out(wire_d54_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance55547(.data_in(wire_d54_6),.data_out(wire_d54_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance55548(.data_in(wire_d54_7),.data_out(wire_d54_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance55549(.data_in(wire_d54_8),.data_out(wire_d54_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance555410(.data_in(wire_d54_9),.data_out(wire_d54_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555411(.data_in(wire_d54_10),.data_out(wire_d54_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555412(.data_in(wire_d54_11),.data_out(wire_d54_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555413(.data_in(wire_d54_12),.data_out(wire_d54_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555414(.data_in(wire_d54_13),.data_out(wire_d54_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance555415(.data_in(wire_d54_14),.data_out(wire_d54_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555416(.data_in(wire_d54_15),.data_out(wire_d54_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555417(.data_in(wire_d54_16),.data_out(wire_d54_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555418(.data_in(wire_d54_17),.data_out(wire_d54_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555419(.data_in(wire_d54_18),.data_out(wire_d54_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance555420(.data_in(wire_d54_19),.data_out(wire_d54_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance555421(.data_in(wire_d54_20),.data_out(wire_d54_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555422(.data_in(wire_d54_21),.data_out(wire_d54_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555423(.data_in(wire_d54_22),.data_out(wire_d54_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance555424(.data_in(wire_d54_23),.data_out(wire_d54_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555425(.data_in(wire_d54_24),.data_out(wire_d54_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance555426(.data_in(wire_d54_25),.data_out(wire_d54_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance555427(.data_in(wire_d54_26),.data_out(wire_d54_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance555428(.data_in(wire_d54_27),.data_out(wire_d54_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555429(.data_in(wire_d54_28),.data_out(wire_d54_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555430(.data_in(wire_d54_29),.data_out(wire_d54_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555431(.data_in(wire_d54_30),.data_out(wire_d54_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555432(.data_in(wire_d54_31),.data_out(wire_d54_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555433(.data_in(wire_d54_32),.data_out(wire_d54_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance555434(.data_in(wire_d54_33),.data_out(wire_d54_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555435(.data_in(wire_d54_34),.data_out(wire_d54_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance555436(.data_in(wire_d54_35),.data_out(wire_d54_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555437(.data_in(wire_d54_36),.data_out(wire_d54_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555438(.data_in(wire_d54_37),.data_out(wire_d54_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555439(.data_in(wire_d54_38),.data_out(wire_d54_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance555440(.data_in(wire_d54_39),.data_out(wire_d54_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance555441(.data_in(wire_d54_40),.data_out(wire_d54_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555442(.data_in(wire_d54_41),.data_out(wire_d54_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance555443(.data_in(wire_d54_42),.data_out(wire_d54_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance555444(.data_in(wire_d54_43),.data_out(wire_d54_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance555445(.data_in(wire_d54_44),.data_out(wire_d54_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555446(.data_in(wire_d54_45),.data_out(wire_d54_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance555447(.data_in(wire_d54_46),.data_out(wire_d54_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance555448(.data_in(wire_d54_47),.data_out(wire_d54_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance555449(.data_in(wire_d54_48),.data_out(wire_d54_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance555450(.data_in(wire_d54_49),.data_out(wire_d54_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555451(.data_in(wire_d54_50),.data_out(wire_d54_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance555452(.data_in(wire_d54_51),.data_out(wire_d54_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance555453(.data_in(wire_d54_52),.data_out(wire_d54_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555454(.data_in(wire_d54_53),.data_out(wire_d54_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555455(.data_in(wire_d54_54),.data_out(wire_d54_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555456(.data_in(wire_d54_55),.data_out(wire_d54_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555457(.data_in(wire_d54_56),.data_out(wire_d54_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance555458(.data_in(wire_d54_57),.data_out(wire_d54_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555459(.data_in(wire_d54_58),.data_out(wire_d54_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance555460(.data_in(wire_d54_59),.data_out(wire_d54_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance555461(.data_in(wire_d54_60),.data_out(wire_d54_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance555462(.data_in(wire_d54_61),.data_out(wire_d54_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555463(.data_in(wire_d54_62),.data_out(wire_d54_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance555464(.data_in(wire_d54_63),.data_out(wire_d54_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance555465(.data_in(wire_d54_64),.data_out(wire_d54_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555466(.data_in(wire_d54_65),.data_out(wire_d54_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555467(.data_in(wire_d54_66),.data_out(wire_d54_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance555468(.data_in(wire_d54_67),.data_out(wire_d54_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance555469(.data_in(wire_d54_68),.data_out(wire_d54_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555470(.data_in(wire_d54_69),.data_out(wire_d54_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555471(.data_in(wire_d54_70),.data_out(wire_d54_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555472(.data_in(wire_d54_71),.data_out(wire_d54_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance555473(.data_in(wire_d54_72),.data_out(wire_d54_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555474(.data_in(wire_d54_73),.data_out(wire_d54_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance555475(.data_in(wire_d54_74),.data_out(wire_d54_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance555476(.data_in(wire_d54_75),.data_out(wire_d54_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555477(.data_in(wire_d54_76),.data_out(wire_d54_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance555478(.data_in(wire_d54_77),.data_out(wire_d54_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance555479(.data_in(wire_d54_78),.data_out(wire_d54_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance555480(.data_in(wire_d54_79),.data_out(wire_d54_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555481(.data_in(wire_d54_80),.data_out(wire_d54_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance555482(.data_in(wire_d54_81),.data_out(wire_d54_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555483(.data_in(wire_d54_82),.data_out(wire_d54_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance555484(.data_in(wire_d54_83),.data_out(wire_d54_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555485(.data_in(wire_d54_84),.data_out(wire_d54_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555486(.data_in(wire_d54_85),.data_out(wire_d54_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555487(.data_in(wire_d54_86),.data_out(wire_d54_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance555488(.data_in(wire_d54_87),.data_out(wire_d54_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance555489(.data_in(wire_d54_88),.data_out(wire_d54_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance555490(.data_in(wire_d54_89),.data_out(wire_d54_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance555491(.data_in(wire_d54_90),.data_out(wire_d54_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555492(.data_in(wire_d54_91),.data_out(wire_d54_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance555493(.data_in(wire_d54_92),.data_out(wire_d54_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555494(.data_in(wire_d54_93),.data_out(wire_d54_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555495(.data_in(wire_d54_94),.data_out(wire_d54_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555496(.data_in(wire_d54_95),.data_out(wire_d54_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555497(.data_in(wire_d54_96),.data_out(wire_d54_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance555498(.data_in(wire_d54_97),.data_out(wire_d54_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance555499(.data_in(wire_d54_98),.data_out(d_out54),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance56550(.data_in(d_in55),.data_out(wire_d55_0),.clk(clk),.rst(rst));            //channel 56
	invertion #(.WIDTH(WIDTH)) invertion_instance56551(.data_in(wire_d55_0),.data_out(wire_d55_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance56552(.data_in(wire_d55_1),.data_out(wire_d55_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance56553(.data_in(wire_d55_2),.data_out(wire_d55_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance56554(.data_in(wire_d55_3),.data_out(wire_d55_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance56555(.data_in(wire_d55_4),.data_out(wire_d55_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance56556(.data_in(wire_d55_5),.data_out(wire_d55_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance56557(.data_in(wire_d55_6),.data_out(wire_d55_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance56558(.data_in(wire_d55_7),.data_out(wire_d55_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance56559(.data_in(wire_d55_8),.data_out(wire_d55_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565510(.data_in(wire_d55_9),.data_out(wire_d55_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565511(.data_in(wire_d55_10),.data_out(wire_d55_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565512(.data_in(wire_d55_11),.data_out(wire_d55_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance565513(.data_in(wire_d55_12),.data_out(wire_d55_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565514(.data_in(wire_d55_13),.data_out(wire_d55_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance565515(.data_in(wire_d55_14),.data_out(wire_d55_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance565516(.data_in(wire_d55_15),.data_out(wire_d55_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565517(.data_in(wire_d55_16),.data_out(wire_d55_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance565518(.data_in(wire_d55_17),.data_out(wire_d55_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565519(.data_in(wire_d55_18),.data_out(wire_d55_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565520(.data_in(wire_d55_19),.data_out(wire_d55_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance565521(.data_in(wire_d55_20),.data_out(wire_d55_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565522(.data_in(wire_d55_21),.data_out(wire_d55_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565523(.data_in(wire_d55_22),.data_out(wire_d55_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565524(.data_in(wire_d55_23),.data_out(wire_d55_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565525(.data_in(wire_d55_24),.data_out(wire_d55_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance565526(.data_in(wire_d55_25),.data_out(wire_d55_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565527(.data_in(wire_d55_26),.data_out(wire_d55_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance565528(.data_in(wire_d55_27),.data_out(wire_d55_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance565529(.data_in(wire_d55_28),.data_out(wire_d55_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565530(.data_in(wire_d55_29),.data_out(wire_d55_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance565531(.data_in(wire_d55_30),.data_out(wire_d55_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance565532(.data_in(wire_d55_31),.data_out(wire_d55_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565533(.data_in(wire_d55_32),.data_out(wire_d55_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance565534(.data_in(wire_d55_33),.data_out(wire_d55_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance565535(.data_in(wire_d55_34),.data_out(wire_d55_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565536(.data_in(wire_d55_35),.data_out(wire_d55_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance565537(.data_in(wire_d55_36),.data_out(wire_d55_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565538(.data_in(wire_d55_37),.data_out(wire_d55_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance565539(.data_in(wire_d55_38),.data_out(wire_d55_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565540(.data_in(wire_d55_39),.data_out(wire_d55_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565541(.data_in(wire_d55_40),.data_out(wire_d55_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565542(.data_in(wire_d55_41),.data_out(wire_d55_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565543(.data_in(wire_d55_42),.data_out(wire_d55_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565544(.data_in(wire_d55_43),.data_out(wire_d55_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565545(.data_in(wire_d55_44),.data_out(wire_d55_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565546(.data_in(wire_d55_45),.data_out(wire_d55_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565547(.data_in(wire_d55_46),.data_out(wire_d55_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance565548(.data_in(wire_d55_47),.data_out(wire_d55_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565549(.data_in(wire_d55_48),.data_out(wire_d55_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565550(.data_in(wire_d55_49),.data_out(wire_d55_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565551(.data_in(wire_d55_50),.data_out(wire_d55_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565552(.data_in(wire_d55_51),.data_out(wire_d55_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565553(.data_in(wire_d55_52),.data_out(wire_d55_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565554(.data_in(wire_d55_53),.data_out(wire_d55_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565555(.data_in(wire_d55_54),.data_out(wire_d55_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565556(.data_in(wire_d55_55),.data_out(wire_d55_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance565557(.data_in(wire_d55_56),.data_out(wire_d55_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance565558(.data_in(wire_d55_57),.data_out(wire_d55_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance565559(.data_in(wire_d55_58),.data_out(wire_d55_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance565560(.data_in(wire_d55_59),.data_out(wire_d55_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565561(.data_in(wire_d55_60),.data_out(wire_d55_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance565562(.data_in(wire_d55_61),.data_out(wire_d55_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance565563(.data_in(wire_d55_62),.data_out(wire_d55_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance565564(.data_in(wire_d55_63),.data_out(wire_d55_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565565(.data_in(wire_d55_64),.data_out(wire_d55_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565566(.data_in(wire_d55_65),.data_out(wire_d55_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565567(.data_in(wire_d55_66),.data_out(wire_d55_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance565568(.data_in(wire_d55_67),.data_out(wire_d55_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565569(.data_in(wire_d55_68),.data_out(wire_d55_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance565570(.data_in(wire_d55_69),.data_out(wire_d55_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance565571(.data_in(wire_d55_70),.data_out(wire_d55_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance565572(.data_in(wire_d55_71),.data_out(wire_d55_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance565573(.data_in(wire_d55_72),.data_out(wire_d55_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565574(.data_in(wire_d55_73),.data_out(wire_d55_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565575(.data_in(wire_d55_74),.data_out(wire_d55_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance565576(.data_in(wire_d55_75),.data_out(wire_d55_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565577(.data_in(wire_d55_76),.data_out(wire_d55_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565578(.data_in(wire_d55_77),.data_out(wire_d55_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance565579(.data_in(wire_d55_78),.data_out(wire_d55_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565580(.data_in(wire_d55_79),.data_out(wire_d55_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance565581(.data_in(wire_d55_80),.data_out(wire_d55_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance565582(.data_in(wire_d55_81),.data_out(wire_d55_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance565583(.data_in(wire_d55_82),.data_out(wire_d55_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance565584(.data_in(wire_d55_83),.data_out(wire_d55_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565585(.data_in(wire_d55_84),.data_out(wire_d55_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance565586(.data_in(wire_d55_85),.data_out(wire_d55_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance565587(.data_in(wire_d55_86),.data_out(wire_d55_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565588(.data_in(wire_d55_87),.data_out(wire_d55_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance565589(.data_in(wire_d55_88),.data_out(wire_d55_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance565590(.data_in(wire_d55_89),.data_out(wire_d55_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance565591(.data_in(wire_d55_90),.data_out(wire_d55_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565592(.data_in(wire_d55_91),.data_out(wire_d55_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance565593(.data_in(wire_d55_92),.data_out(wire_d55_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance565594(.data_in(wire_d55_93),.data_out(wire_d55_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance565595(.data_in(wire_d55_94),.data_out(wire_d55_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance565596(.data_in(wire_d55_95),.data_out(wire_d55_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance565597(.data_in(wire_d55_96),.data_out(wire_d55_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance565598(.data_in(wire_d55_97),.data_out(wire_d55_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance565599(.data_in(wire_d55_98),.data_out(d_out55),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance57560(.data_in(d_in56),.data_out(wire_d56_0),.clk(clk),.rst(rst));            //channel 57
	invertion #(.WIDTH(WIDTH)) invertion_instance57561(.data_in(wire_d56_0),.data_out(wire_d56_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance57562(.data_in(wire_d56_1),.data_out(wire_d56_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance57563(.data_in(wire_d56_2),.data_out(wire_d56_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance57564(.data_in(wire_d56_3),.data_out(wire_d56_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance57565(.data_in(wire_d56_4),.data_out(wire_d56_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance57566(.data_in(wire_d56_5),.data_out(wire_d56_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance57567(.data_in(wire_d56_6),.data_out(wire_d56_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance57568(.data_in(wire_d56_7),.data_out(wire_d56_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance57569(.data_in(wire_d56_8),.data_out(wire_d56_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance575610(.data_in(wire_d56_9),.data_out(wire_d56_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575611(.data_in(wire_d56_10),.data_out(wire_d56_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance575612(.data_in(wire_d56_11),.data_out(wire_d56_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance575613(.data_in(wire_d56_12),.data_out(wire_d56_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance575614(.data_in(wire_d56_13),.data_out(wire_d56_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575615(.data_in(wire_d56_14),.data_out(wire_d56_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575616(.data_in(wire_d56_15),.data_out(wire_d56_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575617(.data_in(wire_d56_16),.data_out(wire_d56_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575618(.data_in(wire_d56_17),.data_out(wire_d56_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance575619(.data_in(wire_d56_18),.data_out(wire_d56_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575620(.data_in(wire_d56_19),.data_out(wire_d56_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance575621(.data_in(wire_d56_20),.data_out(wire_d56_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575622(.data_in(wire_d56_21),.data_out(wire_d56_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance575623(.data_in(wire_d56_22),.data_out(wire_d56_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575624(.data_in(wire_d56_23),.data_out(wire_d56_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575625(.data_in(wire_d56_24),.data_out(wire_d56_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575626(.data_in(wire_d56_25),.data_out(wire_d56_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance575627(.data_in(wire_d56_26),.data_out(wire_d56_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance575628(.data_in(wire_d56_27),.data_out(wire_d56_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance575629(.data_in(wire_d56_28),.data_out(wire_d56_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575630(.data_in(wire_d56_29),.data_out(wire_d56_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575631(.data_in(wire_d56_30),.data_out(wire_d56_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance575632(.data_in(wire_d56_31),.data_out(wire_d56_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance575633(.data_in(wire_d56_32),.data_out(wire_d56_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575634(.data_in(wire_d56_33),.data_out(wire_d56_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance575635(.data_in(wire_d56_34),.data_out(wire_d56_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575636(.data_in(wire_d56_35),.data_out(wire_d56_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance575637(.data_in(wire_d56_36),.data_out(wire_d56_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575638(.data_in(wire_d56_37),.data_out(wire_d56_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance575639(.data_in(wire_d56_38),.data_out(wire_d56_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575640(.data_in(wire_d56_39),.data_out(wire_d56_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance575641(.data_in(wire_d56_40),.data_out(wire_d56_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance575642(.data_in(wire_d56_41),.data_out(wire_d56_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575643(.data_in(wire_d56_42),.data_out(wire_d56_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575644(.data_in(wire_d56_43),.data_out(wire_d56_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575645(.data_in(wire_d56_44),.data_out(wire_d56_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575646(.data_in(wire_d56_45),.data_out(wire_d56_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance575647(.data_in(wire_d56_46),.data_out(wire_d56_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575648(.data_in(wire_d56_47),.data_out(wire_d56_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance575649(.data_in(wire_d56_48),.data_out(wire_d56_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance575650(.data_in(wire_d56_49),.data_out(wire_d56_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance575651(.data_in(wire_d56_50),.data_out(wire_d56_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575652(.data_in(wire_d56_51),.data_out(wire_d56_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance575653(.data_in(wire_d56_52),.data_out(wire_d56_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575654(.data_in(wire_d56_53),.data_out(wire_d56_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance575655(.data_in(wire_d56_54),.data_out(wire_d56_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance575656(.data_in(wire_d56_55),.data_out(wire_d56_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575657(.data_in(wire_d56_56),.data_out(wire_d56_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance575658(.data_in(wire_d56_57),.data_out(wire_d56_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575659(.data_in(wire_d56_58),.data_out(wire_d56_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575660(.data_in(wire_d56_59),.data_out(wire_d56_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575661(.data_in(wire_d56_60),.data_out(wire_d56_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575662(.data_in(wire_d56_61),.data_out(wire_d56_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance575663(.data_in(wire_d56_62),.data_out(wire_d56_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance575664(.data_in(wire_d56_63),.data_out(wire_d56_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance575665(.data_in(wire_d56_64),.data_out(wire_d56_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575666(.data_in(wire_d56_65),.data_out(wire_d56_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance575667(.data_in(wire_d56_66),.data_out(wire_d56_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance575668(.data_in(wire_d56_67),.data_out(wire_d56_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance575669(.data_in(wire_d56_68),.data_out(wire_d56_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575670(.data_in(wire_d56_69),.data_out(wire_d56_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575671(.data_in(wire_d56_70),.data_out(wire_d56_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575672(.data_in(wire_d56_71),.data_out(wire_d56_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575673(.data_in(wire_d56_72),.data_out(wire_d56_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575674(.data_in(wire_d56_73),.data_out(wire_d56_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575675(.data_in(wire_d56_74),.data_out(wire_d56_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575676(.data_in(wire_d56_75),.data_out(wire_d56_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575677(.data_in(wire_d56_76),.data_out(wire_d56_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575678(.data_in(wire_d56_77),.data_out(wire_d56_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575679(.data_in(wire_d56_78),.data_out(wire_d56_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance575680(.data_in(wire_d56_79),.data_out(wire_d56_80),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance575681(.data_in(wire_d56_80),.data_out(wire_d56_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575682(.data_in(wire_d56_81),.data_out(wire_d56_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575683(.data_in(wire_d56_82),.data_out(wire_d56_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575684(.data_in(wire_d56_83),.data_out(wire_d56_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance575685(.data_in(wire_d56_84),.data_out(wire_d56_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575686(.data_in(wire_d56_85),.data_out(wire_d56_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance575687(.data_in(wire_d56_86),.data_out(wire_d56_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575688(.data_in(wire_d56_87),.data_out(wire_d56_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance575689(.data_in(wire_d56_88),.data_out(wire_d56_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575690(.data_in(wire_d56_89),.data_out(wire_d56_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575691(.data_in(wire_d56_90),.data_out(wire_d56_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575692(.data_in(wire_d56_91),.data_out(wire_d56_92),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance575693(.data_in(wire_d56_92),.data_out(wire_d56_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance575694(.data_in(wire_d56_93),.data_out(wire_d56_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance575695(.data_in(wire_d56_94),.data_out(wire_d56_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance575696(.data_in(wire_d56_95),.data_out(wire_d56_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance575697(.data_in(wire_d56_96),.data_out(wire_d56_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance575698(.data_in(wire_d56_97),.data_out(wire_d56_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance575699(.data_in(wire_d56_98),.data_out(d_out56),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance58570(.data_in(d_in57),.data_out(wire_d57_0),.clk(clk),.rst(rst));            //channel 58
	encoder #(.WIDTH(WIDTH)) encoder_instance58571(.data_in(wire_d57_0),.data_out(wire_d57_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance58572(.data_in(wire_d57_1),.data_out(wire_d57_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance58573(.data_in(wire_d57_2),.data_out(wire_d57_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance58574(.data_in(wire_d57_3),.data_out(wire_d57_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance58575(.data_in(wire_d57_4),.data_out(wire_d57_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance58576(.data_in(wire_d57_5),.data_out(wire_d57_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance58577(.data_in(wire_d57_6),.data_out(wire_d57_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance58578(.data_in(wire_d57_7),.data_out(wire_d57_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance58579(.data_in(wire_d57_8),.data_out(wire_d57_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585710(.data_in(wire_d57_9),.data_out(wire_d57_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance585711(.data_in(wire_d57_10),.data_out(wire_d57_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance585712(.data_in(wire_d57_11),.data_out(wire_d57_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance585713(.data_in(wire_d57_12),.data_out(wire_d57_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance585714(.data_in(wire_d57_13),.data_out(wire_d57_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585715(.data_in(wire_d57_14),.data_out(wire_d57_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585716(.data_in(wire_d57_15),.data_out(wire_d57_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585717(.data_in(wire_d57_16),.data_out(wire_d57_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585718(.data_in(wire_d57_17),.data_out(wire_d57_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance585719(.data_in(wire_d57_18),.data_out(wire_d57_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585720(.data_in(wire_d57_19),.data_out(wire_d57_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585721(.data_in(wire_d57_20),.data_out(wire_d57_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585722(.data_in(wire_d57_21),.data_out(wire_d57_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance585723(.data_in(wire_d57_22),.data_out(wire_d57_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance585724(.data_in(wire_d57_23),.data_out(wire_d57_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585725(.data_in(wire_d57_24),.data_out(wire_d57_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance585726(.data_in(wire_d57_25),.data_out(wire_d57_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585727(.data_in(wire_d57_26),.data_out(wire_d57_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585728(.data_in(wire_d57_27),.data_out(wire_d57_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance585729(.data_in(wire_d57_28),.data_out(wire_d57_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585730(.data_in(wire_d57_29),.data_out(wire_d57_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585731(.data_in(wire_d57_30),.data_out(wire_d57_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance585732(.data_in(wire_d57_31),.data_out(wire_d57_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance585733(.data_in(wire_d57_32),.data_out(wire_d57_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance585734(.data_in(wire_d57_33),.data_out(wire_d57_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance585735(.data_in(wire_d57_34),.data_out(wire_d57_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance585736(.data_in(wire_d57_35),.data_out(wire_d57_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance585737(.data_in(wire_d57_36),.data_out(wire_d57_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance585738(.data_in(wire_d57_37),.data_out(wire_d57_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585739(.data_in(wire_d57_38),.data_out(wire_d57_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585740(.data_in(wire_d57_39),.data_out(wire_d57_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585741(.data_in(wire_d57_40),.data_out(wire_d57_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585742(.data_in(wire_d57_41),.data_out(wire_d57_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585743(.data_in(wire_d57_42),.data_out(wire_d57_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585744(.data_in(wire_d57_43),.data_out(wire_d57_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585745(.data_in(wire_d57_44),.data_out(wire_d57_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance585746(.data_in(wire_d57_45),.data_out(wire_d57_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance585747(.data_in(wire_d57_46),.data_out(wire_d57_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance585748(.data_in(wire_d57_47),.data_out(wire_d57_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585749(.data_in(wire_d57_48),.data_out(wire_d57_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance585750(.data_in(wire_d57_49),.data_out(wire_d57_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585751(.data_in(wire_d57_50),.data_out(wire_d57_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585752(.data_in(wire_d57_51),.data_out(wire_d57_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance585753(.data_in(wire_d57_52),.data_out(wire_d57_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance585754(.data_in(wire_d57_53),.data_out(wire_d57_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585755(.data_in(wire_d57_54),.data_out(wire_d57_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585756(.data_in(wire_d57_55),.data_out(wire_d57_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance585757(.data_in(wire_d57_56),.data_out(wire_d57_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585758(.data_in(wire_d57_57),.data_out(wire_d57_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585759(.data_in(wire_d57_58),.data_out(wire_d57_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance585760(.data_in(wire_d57_59),.data_out(wire_d57_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance585761(.data_in(wire_d57_60),.data_out(wire_d57_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585762(.data_in(wire_d57_61),.data_out(wire_d57_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585763(.data_in(wire_d57_62),.data_out(wire_d57_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance585764(.data_in(wire_d57_63),.data_out(wire_d57_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585765(.data_in(wire_d57_64),.data_out(wire_d57_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance585766(.data_in(wire_d57_65),.data_out(wire_d57_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance585767(.data_in(wire_d57_66),.data_out(wire_d57_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance585768(.data_in(wire_d57_67),.data_out(wire_d57_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585769(.data_in(wire_d57_68),.data_out(wire_d57_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance585770(.data_in(wire_d57_69),.data_out(wire_d57_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585771(.data_in(wire_d57_70),.data_out(wire_d57_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585772(.data_in(wire_d57_71),.data_out(wire_d57_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance585773(.data_in(wire_d57_72),.data_out(wire_d57_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585774(.data_in(wire_d57_73),.data_out(wire_d57_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585775(.data_in(wire_d57_74),.data_out(wire_d57_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance585776(.data_in(wire_d57_75),.data_out(wire_d57_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585777(.data_in(wire_d57_76),.data_out(wire_d57_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585778(.data_in(wire_d57_77),.data_out(wire_d57_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance585779(.data_in(wire_d57_78),.data_out(wire_d57_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance585780(.data_in(wire_d57_79),.data_out(wire_d57_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance585781(.data_in(wire_d57_80),.data_out(wire_d57_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance585782(.data_in(wire_d57_81),.data_out(wire_d57_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance585783(.data_in(wire_d57_82),.data_out(wire_d57_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance585784(.data_in(wire_d57_83),.data_out(wire_d57_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585785(.data_in(wire_d57_84),.data_out(wire_d57_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585786(.data_in(wire_d57_85),.data_out(wire_d57_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585787(.data_in(wire_d57_86),.data_out(wire_d57_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585788(.data_in(wire_d57_87),.data_out(wire_d57_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance585789(.data_in(wire_d57_88),.data_out(wire_d57_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585790(.data_in(wire_d57_89),.data_out(wire_d57_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance585791(.data_in(wire_d57_90),.data_out(wire_d57_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance585792(.data_in(wire_d57_91),.data_out(wire_d57_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585793(.data_in(wire_d57_92),.data_out(wire_d57_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance585794(.data_in(wire_d57_93),.data_out(wire_d57_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585795(.data_in(wire_d57_94),.data_out(wire_d57_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585796(.data_in(wire_d57_95),.data_out(wire_d57_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance585797(.data_in(wire_d57_96),.data_out(wire_d57_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance585798(.data_in(wire_d57_97),.data_out(wire_d57_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance585799(.data_in(wire_d57_98),.data_out(d_out57),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance59580(.data_in(d_in58),.data_out(wire_d58_0),.clk(clk),.rst(rst));            //channel 59
	encoder #(.WIDTH(WIDTH)) encoder_instance59581(.data_in(wire_d58_0),.data_out(wire_d58_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance59582(.data_in(wire_d58_1),.data_out(wire_d58_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance59583(.data_in(wire_d58_2),.data_out(wire_d58_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance59584(.data_in(wire_d58_3),.data_out(wire_d58_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance59585(.data_in(wire_d58_4),.data_out(wire_d58_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance59586(.data_in(wire_d58_5),.data_out(wire_d58_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance59587(.data_in(wire_d58_6),.data_out(wire_d58_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance59588(.data_in(wire_d58_7),.data_out(wire_d58_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance59589(.data_in(wire_d58_8),.data_out(wire_d58_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595810(.data_in(wire_d58_9),.data_out(wire_d58_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595811(.data_in(wire_d58_10),.data_out(wire_d58_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595812(.data_in(wire_d58_11),.data_out(wire_d58_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance595813(.data_in(wire_d58_12),.data_out(wire_d58_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595814(.data_in(wire_d58_13),.data_out(wire_d58_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance595815(.data_in(wire_d58_14),.data_out(wire_d58_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595816(.data_in(wire_d58_15),.data_out(wire_d58_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595817(.data_in(wire_d58_16),.data_out(wire_d58_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595818(.data_in(wire_d58_17),.data_out(wire_d58_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance595819(.data_in(wire_d58_18),.data_out(wire_d58_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595820(.data_in(wire_d58_19),.data_out(wire_d58_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595821(.data_in(wire_d58_20),.data_out(wire_d58_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595822(.data_in(wire_d58_21),.data_out(wire_d58_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595823(.data_in(wire_d58_22),.data_out(wire_d58_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance595824(.data_in(wire_d58_23),.data_out(wire_d58_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595825(.data_in(wire_d58_24),.data_out(wire_d58_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance595826(.data_in(wire_d58_25),.data_out(wire_d58_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595827(.data_in(wire_d58_26),.data_out(wire_d58_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595828(.data_in(wire_d58_27),.data_out(wire_d58_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance595829(.data_in(wire_d58_28),.data_out(wire_d58_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance595830(.data_in(wire_d58_29),.data_out(wire_d58_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595831(.data_in(wire_d58_30),.data_out(wire_d58_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595832(.data_in(wire_d58_31),.data_out(wire_d58_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595833(.data_in(wire_d58_32),.data_out(wire_d58_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance595834(.data_in(wire_d58_33),.data_out(wire_d58_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595835(.data_in(wire_d58_34),.data_out(wire_d58_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595836(.data_in(wire_d58_35),.data_out(wire_d58_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595837(.data_in(wire_d58_36),.data_out(wire_d58_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595838(.data_in(wire_d58_37),.data_out(wire_d58_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595839(.data_in(wire_d58_38),.data_out(wire_d58_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance595840(.data_in(wire_d58_39),.data_out(wire_d58_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595841(.data_in(wire_d58_40),.data_out(wire_d58_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595842(.data_in(wire_d58_41),.data_out(wire_d58_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595843(.data_in(wire_d58_42),.data_out(wire_d58_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595844(.data_in(wire_d58_43),.data_out(wire_d58_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595845(.data_in(wire_d58_44),.data_out(wire_d58_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595846(.data_in(wire_d58_45),.data_out(wire_d58_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance595847(.data_in(wire_d58_46),.data_out(wire_d58_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595848(.data_in(wire_d58_47),.data_out(wire_d58_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595849(.data_in(wire_d58_48),.data_out(wire_d58_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance595850(.data_in(wire_d58_49),.data_out(wire_d58_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595851(.data_in(wire_d58_50),.data_out(wire_d58_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595852(.data_in(wire_d58_51),.data_out(wire_d58_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595853(.data_in(wire_d58_52),.data_out(wire_d58_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595854(.data_in(wire_d58_53),.data_out(wire_d58_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595855(.data_in(wire_d58_54),.data_out(wire_d58_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595856(.data_in(wire_d58_55),.data_out(wire_d58_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance595857(.data_in(wire_d58_56),.data_out(wire_d58_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595858(.data_in(wire_d58_57),.data_out(wire_d58_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595859(.data_in(wire_d58_58),.data_out(wire_d58_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance595860(.data_in(wire_d58_59),.data_out(wire_d58_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595861(.data_in(wire_d58_60),.data_out(wire_d58_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595862(.data_in(wire_d58_61),.data_out(wire_d58_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595863(.data_in(wire_d58_62),.data_out(wire_d58_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595864(.data_in(wire_d58_63),.data_out(wire_d58_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595865(.data_in(wire_d58_64),.data_out(wire_d58_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595866(.data_in(wire_d58_65),.data_out(wire_d58_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595867(.data_in(wire_d58_66),.data_out(wire_d58_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance595868(.data_in(wire_d58_67),.data_out(wire_d58_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance595869(.data_in(wire_d58_68),.data_out(wire_d58_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595870(.data_in(wire_d58_69),.data_out(wire_d58_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance595871(.data_in(wire_d58_70),.data_out(wire_d58_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance595872(.data_in(wire_d58_71),.data_out(wire_d58_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595873(.data_in(wire_d58_72),.data_out(wire_d58_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595874(.data_in(wire_d58_73),.data_out(wire_d58_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595875(.data_in(wire_d58_74),.data_out(wire_d58_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595876(.data_in(wire_d58_75),.data_out(wire_d58_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595877(.data_in(wire_d58_76),.data_out(wire_d58_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595878(.data_in(wire_d58_77),.data_out(wire_d58_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595879(.data_in(wire_d58_78),.data_out(wire_d58_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595880(.data_in(wire_d58_79),.data_out(wire_d58_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595881(.data_in(wire_d58_80),.data_out(wire_d58_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595882(.data_in(wire_d58_81),.data_out(wire_d58_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance595883(.data_in(wire_d58_82),.data_out(wire_d58_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance595884(.data_in(wire_d58_83),.data_out(wire_d58_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595885(.data_in(wire_d58_84),.data_out(wire_d58_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595886(.data_in(wire_d58_85),.data_out(wire_d58_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595887(.data_in(wire_d58_86),.data_out(wire_d58_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595888(.data_in(wire_d58_87),.data_out(wire_d58_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595889(.data_in(wire_d58_88),.data_out(wire_d58_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595890(.data_in(wire_d58_89),.data_out(wire_d58_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595891(.data_in(wire_d58_90),.data_out(wire_d58_91),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595892(.data_in(wire_d58_91),.data_out(wire_d58_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595893(.data_in(wire_d58_92),.data_out(wire_d58_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance595894(.data_in(wire_d58_93),.data_out(wire_d58_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance595895(.data_in(wire_d58_94),.data_out(wire_d58_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595896(.data_in(wire_d58_95),.data_out(wire_d58_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595897(.data_in(wire_d58_96),.data_out(wire_d58_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance595898(.data_in(wire_d58_97),.data_out(wire_d58_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance595899(.data_in(wire_d58_98),.data_out(d_out58),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance60590(.data_in(d_in59),.data_out(wire_d59_0),.clk(clk),.rst(rst));            //channel 60
	large_mux #(.WIDTH(WIDTH)) large_mux_instance60591(.data_in(wire_d59_0),.data_out(wire_d59_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance60592(.data_in(wire_d59_1),.data_out(wire_d59_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance60593(.data_in(wire_d59_2),.data_out(wire_d59_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance60594(.data_in(wire_d59_3),.data_out(wire_d59_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance60595(.data_in(wire_d59_4),.data_out(wire_d59_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance60596(.data_in(wire_d59_5),.data_out(wire_d59_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance60597(.data_in(wire_d59_6),.data_out(wire_d59_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance60598(.data_in(wire_d59_7),.data_out(wire_d59_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance60599(.data_in(wire_d59_8),.data_out(wire_d59_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605910(.data_in(wire_d59_9),.data_out(wire_d59_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance605911(.data_in(wire_d59_10),.data_out(wire_d59_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605912(.data_in(wire_d59_11),.data_out(wire_d59_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance605913(.data_in(wire_d59_12),.data_out(wire_d59_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605914(.data_in(wire_d59_13),.data_out(wire_d59_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance605915(.data_in(wire_d59_14),.data_out(wire_d59_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance605916(.data_in(wire_d59_15),.data_out(wire_d59_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605917(.data_in(wire_d59_16),.data_out(wire_d59_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605918(.data_in(wire_d59_17),.data_out(wire_d59_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605919(.data_in(wire_d59_18),.data_out(wire_d59_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605920(.data_in(wire_d59_19),.data_out(wire_d59_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance605921(.data_in(wire_d59_20),.data_out(wire_d59_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance605922(.data_in(wire_d59_21),.data_out(wire_d59_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605923(.data_in(wire_d59_22),.data_out(wire_d59_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605924(.data_in(wire_d59_23),.data_out(wire_d59_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance605925(.data_in(wire_d59_24),.data_out(wire_d59_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605926(.data_in(wire_d59_25),.data_out(wire_d59_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605927(.data_in(wire_d59_26),.data_out(wire_d59_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605928(.data_in(wire_d59_27),.data_out(wire_d59_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605929(.data_in(wire_d59_28),.data_out(wire_d59_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605930(.data_in(wire_d59_29),.data_out(wire_d59_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605931(.data_in(wire_d59_30),.data_out(wire_d59_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605932(.data_in(wire_d59_31),.data_out(wire_d59_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605933(.data_in(wire_d59_32),.data_out(wire_d59_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605934(.data_in(wire_d59_33),.data_out(wire_d59_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance605935(.data_in(wire_d59_34),.data_out(wire_d59_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605936(.data_in(wire_d59_35),.data_out(wire_d59_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605937(.data_in(wire_d59_36),.data_out(wire_d59_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605938(.data_in(wire_d59_37),.data_out(wire_d59_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605939(.data_in(wire_d59_38),.data_out(wire_d59_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605940(.data_in(wire_d59_39),.data_out(wire_d59_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605941(.data_in(wire_d59_40),.data_out(wire_d59_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605942(.data_in(wire_d59_41),.data_out(wire_d59_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605943(.data_in(wire_d59_42),.data_out(wire_d59_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605944(.data_in(wire_d59_43),.data_out(wire_d59_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605945(.data_in(wire_d59_44),.data_out(wire_d59_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605946(.data_in(wire_d59_45),.data_out(wire_d59_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance605947(.data_in(wire_d59_46),.data_out(wire_d59_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605948(.data_in(wire_d59_47),.data_out(wire_d59_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605949(.data_in(wire_d59_48),.data_out(wire_d59_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605950(.data_in(wire_d59_49),.data_out(wire_d59_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605951(.data_in(wire_d59_50),.data_out(wire_d59_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605952(.data_in(wire_d59_51),.data_out(wire_d59_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605953(.data_in(wire_d59_52),.data_out(wire_d59_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance605954(.data_in(wire_d59_53),.data_out(wire_d59_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605955(.data_in(wire_d59_54),.data_out(wire_d59_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605956(.data_in(wire_d59_55),.data_out(wire_d59_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605957(.data_in(wire_d59_56),.data_out(wire_d59_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance605958(.data_in(wire_d59_57),.data_out(wire_d59_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605959(.data_in(wire_d59_58),.data_out(wire_d59_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance605960(.data_in(wire_d59_59),.data_out(wire_d59_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605961(.data_in(wire_d59_60),.data_out(wire_d59_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605962(.data_in(wire_d59_61),.data_out(wire_d59_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605963(.data_in(wire_d59_62),.data_out(wire_d59_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605964(.data_in(wire_d59_63),.data_out(wire_d59_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605965(.data_in(wire_d59_64),.data_out(wire_d59_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605966(.data_in(wire_d59_65),.data_out(wire_d59_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605967(.data_in(wire_d59_66),.data_out(wire_d59_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605968(.data_in(wire_d59_67),.data_out(wire_d59_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605969(.data_in(wire_d59_68),.data_out(wire_d59_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605970(.data_in(wire_d59_69),.data_out(wire_d59_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605971(.data_in(wire_d59_70),.data_out(wire_d59_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605972(.data_in(wire_d59_71),.data_out(wire_d59_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605973(.data_in(wire_d59_72),.data_out(wire_d59_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605974(.data_in(wire_d59_73),.data_out(wire_d59_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance605975(.data_in(wire_d59_74),.data_out(wire_d59_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605976(.data_in(wire_d59_75),.data_out(wire_d59_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605977(.data_in(wire_d59_76),.data_out(wire_d59_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605978(.data_in(wire_d59_77),.data_out(wire_d59_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605979(.data_in(wire_d59_78),.data_out(wire_d59_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance605980(.data_in(wire_d59_79),.data_out(wire_d59_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605981(.data_in(wire_d59_80),.data_out(wire_d59_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance605982(.data_in(wire_d59_81),.data_out(wire_d59_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance605983(.data_in(wire_d59_82),.data_out(wire_d59_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance605984(.data_in(wire_d59_83),.data_out(wire_d59_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605985(.data_in(wire_d59_84),.data_out(wire_d59_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605986(.data_in(wire_d59_85),.data_out(wire_d59_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605987(.data_in(wire_d59_86),.data_out(wire_d59_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance605988(.data_in(wire_d59_87),.data_out(wire_d59_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605989(.data_in(wire_d59_88),.data_out(wire_d59_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605990(.data_in(wire_d59_89),.data_out(wire_d59_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance605991(.data_in(wire_d59_90),.data_out(wire_d59_91),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605992(.data_in(wire_d59_91),.data_out(wire_d59_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance605993(.data_in(wire_d59_92),.data_out(wire_d59_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605994(.data_in(wire_d59_93),.data_out(wire_d59_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605995(.data_in(wire_d59_94),.data_out(wire_d59_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance605996(.data_in(wire_d59_95),.data_out(wire_d59_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance605997(.data_in(wire_d59_96),.data_out(wire_d59_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605998(.data_in(wire_d59_97),.data_out(wire_d59_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance605999(.data_in(wire_d59_98),.data_out(d_out59),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance61600(.data_in(d_in60),.data_out(wire_d60_0),.clk(clk),.rst(rst));            //channel 61
	register #(.WIDTH(WIDTH)) register_instance61601(.data_in(wire_d60_0),.data_out(wire_d60_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance61602(.data_in(wire_d60_1),.data_out(wire_d60_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance61603(.data_in(wire_d60_2),.data_out(wire_d60_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance61604(.data_in(wire_d60_3),.data_out(wire_d60_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance61605(.data_in(wire_d60_4),.data_out(wire_d60_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance61606(.data_in(wire_d60_5),.data_out(wire_d60_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance61607(.data_in(wire_d60_6),.data_out(wire_d60_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance61608(.data_in(wire_d60_7),.data_out(wire_d60_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance61609(.data_in(wire_d60_8),.data_out(wire_d60_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance616010(.data_in(wire_d60_9),.data_out(wire_d60_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616011(.data_in(wire_d60_10),.data_out(wire_d60_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616012(.data_in(wire_d60_11),.data_out(wire_d60_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance616013(.data_in(wire_d60_12),.data_out(wire_d60_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance616014(.data_in(wire_d60_13),.data_out(wire_d60_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616015(.data_in(wire_d60_14),.data_out(wire_d60_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616016(.data_in(wire_d60_15),.data_out(wire_d60_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance616017(.data_in(wire_d60_16),.data_out(wire_d60_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616018(.data_in(wire_d60_17),.data_out(wire_d60_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616019(.data_in(wire_d60_18),.data_out(wire_d60_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance616020(.data_in(wire_d60_19),.data_out(wire_d60_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616021(.data_in(wire_d60_20),.data_out(wire_d60_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance616022(.data_in(wire_d60_21),.data_out(wire_d60_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance616023(.data_in(wire_d60_22),.data_out(wire_d60_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance616024(.data_in(wire_d60_23),.data_out(wire_d60_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance616025(.data_in(wire_d60_24),.data_out(wire_d60_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616026(.data_in(wire_d60_25),.data_out(wire_d60_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616027(.data_in(wire_d60_26),.data_out(wire_d60_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616028(.data_in(wire_d60_27),.data_out(wire_d60_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616029(.data_in(wire_d60_28),.data_out(wire_d60_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616030(.data_in(wire_d60_29),.data_out(wire_d60_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance616031(.data_in(wire_d60_30),.data_out(wire_d60_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance616032(.data_in(wire_d60_31),.data_out(wire_d60_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616033(.data_in(wire_d60_32),.data_out(wire_d60_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance616034(.data_in(wire_d60_33),.data_out(wire_d60_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616035(.data_in(wire_d60_34),.data_out(wire_d60_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616036(.data_in(wire_d60_35),.data_out(wire_d60_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616037(.data_in(wire_d60_36),.data_out(wire_d60_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616038(.data_in(wire_d60_37),.data_out(wire_d60_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616039(.data_in(wire_d60_38),.data_out(wire_d60_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616040(.data_in(wire_d60_39),.data_out(wire_d60_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance616041(.data_in(wire_d60_40),.data_out(wire_d60_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance616042(.data_in(wire_d60_41),.data_out(wire_d60_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616043(.data_in(wire_d60_42),.data_out(wire_d60_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616044(.data_in(wire_d60_43),.data_out(wire_d60_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance616045(.data_in(wire_d60_44),.data_out(wire_d60_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance616046(.data_in(wire_d60_45),.data_out(wire_d60_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance616047(.data_in(wire_d60_46),.data_out(wire_d60_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616048(.data_in(wire_d60_47),.data_out(wire_d60_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance616049(.data_in(wire_d60_48),.data_out(wire_d60_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616050(.data_in(wire_d60_49),.data_out(wire_d60_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616051(.data_in(wire_d60_50),.data_out(wire_d60_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance616052(.data_in(wire_d60_51),.data_out(wire_d60_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance616053(.data_in(wire_d60_52),.data_out(wire_d60_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616054(.data_in(wire_d60_53),.data_out(wire_d60_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance616055(.data_in(wire_d60_54),.data_out(wire_d60_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance616056(.data_in(wire_d60_55),.data_out(wire_d60_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance616057(.data_in(wire_d60_56),.data_out(wire_d60_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance616058(.data_in(wire_d60_57),.data_out(wire_d60_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616059(.data_in(wire_d60_58),.data_out(wire_d60_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616060(.data_in(wire_d60_59),.data_out(wire_d60_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616061(.data_in(wire_d60_60),.data_out(wire_d60_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616062(.data_in(wire_d60_61),.data_out(wire_d60_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance616063(.data_in(wire_d60_62),.data_out(wire_d60_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance616064(.data_in(wire_d60_63),.data_out(wire_d60_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616065(.data_in(wire_d60_64),.data_out(wire_d60_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance616066(.data_in(wire_d60_65),.data_out(wire_d60_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616067(.data_in(wire_d60_66),.data_out(wire_d60_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance616068(.data_in(wire_d60_67),.data_out(wire_d60_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance616069(.data_in(wire_d60_68),.data_out(wire_d60_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance616070(.data_in(wire_d60_69),.data_out(wire_d60_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance616071(.data_in(wire_d60_70),.data_out(wire_d60_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616072(.data_in(wire_d60_71),.data_out(wire_d60_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance616073(.data_in(wire_d60_72),.data_out(wire_d60_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance616074(.data_in(wire_d60_73),.data_out(wire_d60_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616075(.data_in(wire_d60_74),.data_out(wire_d60_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance616076(.data_in(wire_d60_75),.data_out(wire_d60_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616077(.data_in(wire_d60_76),.data_out(wire_d60_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616078(.data_in(wire_d60_77),.data_out(wire_d60_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance616079(.data_in(wire_d60_78),.data_out(wire_d60_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance616080(.data_in(wire_d60_79),.data_out(wire_d60_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616081(.data_in(wire_d60_80),.data_out(wire_d60_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616082(.data_in(wire_d60_81),.data_out(wire_d60_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance616083(.data_in(wire_d60_82),.data_out(wire_d60_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616084(.data_in(wire_d60_83),.data_out(wire_d60_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616085(.data_in(wire_d60_84),.data_out(wire_d60_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616086(.data_in(wire_d60_85),.data_out(wire_d60_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616087(.data_in(wire_d60_86),.data_out(wire_d60_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616088(.data_in(wire_d60_87),.data_out(wire_d60_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616089(.data_in(wire_d60_88),.data_out(wire_d60_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance616090(.data_in(wire_d60_89),.data_out(wire_d60_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616091(.data_in(wire_d60_90),.data_out(wire_d60_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616092(.data_in(wire_d60_91),.data_out(wire_d60_92),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance616093(.data_in(wire_d60_92),.data_out(wire_d60_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance616094(.data_in(wire_d60_93),.data_out(wire_d60_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance616095(.data_in(wire_d60_94),.data_out(wire_d60_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616096(.data_in(wire_d60_95),.data_out(wire_d60_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616097(.data_in(wire_d60_96),.data_out(wire_d60_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance616098(.data_in(wire_d60_97),.data_out(wire_d60_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance616099(.data_in(wire_d60_98),.data_out(d_out60),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance62610(.data_in(d_in61),.data_out(wire_d61_0),.clk(clk),.rst(rst));            //channel 62
	encoder #(.WIDTH(WIDTH)) encoder_instance62611(.data_in(wire_d61_0),.data_out(wire_d61_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance62612(.data_in(wire_d61_1),.data_out(wire_d61_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance62613(.data_in(wire_d61_2),.data_out(wire_d61_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance62614(.data_in(wire_d61_3),.data_out(wire_d61_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance62615(.data_in(wire_d61_4),.data_out(wire_d61_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance62616(.data_in(wire_d61_5),.data_out(wire_d61_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance62617(.data_in(wire_d61_6),.data_out(wire_d61_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance62618(.data_in(wire_d61_7),.data_out(wire_d61_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance62619(.data_in(wire_d61_8),.data_out(wire_d61_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626110(.data_in(wire_d61_9),.data_out(wire_d61_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance626111(.data_in(wire_d61_10),.data_out(wire_d61_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance626112(.data_in(wire_d61_11),.data_out(wire_d61_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626113(.data_in(wire_d61_12),.data_out(wire_d61_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance626114(.data_in(wire_d61_13),.data_out(wire_d61_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance626115(.data_in(wire_d61_14),.data_out(wire_d61_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626116(.data_in(wire_d61_15),.data_out(wire_d61_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance626117(.data_in(wire_d61_16),.data_out(wire_d61_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626118(.data_in(wire_d61_17),.data_out(wire_d61_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626119(.data_in(wire_d61_18),.data_out(wire_d61_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626120(.data_in(wire_d61_19),.data_out(wire_d61_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626121(.data_in(wire_d61_20),.data_out(wire_d61_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626122(.data_in(wire_d61_21),.data_out(wire_d61_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626123(.data_in(wire_d61_22),.data_out(wire_d61_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626124(.data_in(wire_d61_23),.data_out(wire_d61_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626125(.data_in(wire_d61_24),.data_out(wire_d61_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance626126(.data_in(wire_d61_25),.data_out(wire_d61_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance626127(.data_in(wire_d61_26),.data_out(wire_d61_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626128(.data_in(wire_d61_27),.data_out(wire_d61_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance626129(.data_in(wire_d61_28),.data_out(wire_d61_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626130(.data_in(wire_d61_29),.data_out(wire_d61_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626131(.data_in(wire_d61_30),.data_out(wire_d61_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance626132(.data_in(wire_d61_31),.data_out(wire_d61_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance626133(.data_in(wire_d61_32),.data_out(wire_d61_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance626134(.data_in(wire_d61_33),.data_out(wire_d61_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626135(.data_in(wire_d61_34),.data_out(wire_d61_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance626136(.data_in(wire_d61_35),.data_out(wire_d61_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626137(.data_in(wire_d61_36),.data_out(wire_d61_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626138(.data_in(wire_d61_37),.data_out(wire_d61_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626139(.data_in(wire_d61_38),.data_out(wire_d61_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626140(.data_in(wire_d61_39),.data_out(wire_d61_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626141(.data_in(wire_d61_40),.data_out(wire_d61_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance626142(.data_in(wire_d61_41),.data_out(wire_d61_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626143(.data_in(wire_d61_42),.data_out(wire_d61_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance626144(.data_in(wire_d61_43),.data_out(wire_d61_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance626145(.data_in(wire_d61_44),.data_out(wire_d61_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626146(.data_in(wire_d61_45),.data_out(wire_d61_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626147(.data_in(wire_d61_46),.data_out(wire_d61_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626148(.data_in(wire_d61_47),.data_out(wire_d61_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626149(.data_in(wire_d61_48),.data_out(wire_d61_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626150(.data_in(wire_d61_49),.data_out(wire_d61_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626151(.data_in(wire_d61_50),.data_out(wire_d61_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance626152(.data_in(wire_d61_51),.data_out(wire_d61_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626153(.data_in(wire_d61_52),.data_out(wire_d61_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626154(.data_in(wire_d61_53),.data_out(wire_d61_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance626155(.data_in(wire_d61_54),.data_out(wire_d61_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance626156(.data_in(wire_d61_55),.data_out(wire_d61_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance626157(.data_in(wire_d61_56),.data_out(wire_d61_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626158(.data_in(wire_d61_57),.data_out(wire_d61_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626159(.data_in(wire_d61_58),.data_out(wire_d61_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626160(.data_in(wire_d61_59),.data_out(wire_d61_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626161(.data_in(wire_d61_60),.data_out(wire_d61_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626162(.data_in(wire_d61_61),.data_out(wire_d61_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance626163(.data_in(wire_d61_62),.data_out(wire_d61_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626164(.data_in(wire_d61_63),.data_out(wire_d61_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance626165(.data_in(wire_d61_64),.data_out(wire_d61_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance626166(.data_in(wire_d61_65),.data_out(wire_d61_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626167(.data_in(wire_d61_66),.data_out(wire_d61_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance626168(.data_in(wire_d61_67),.data_out(wire_d61_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance626169(.data_in(wire_d61_68),.data_out(wire_d61_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance626170(.data_in(wire_d61_69),.data_out(wire_d61_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626171(.data_in(wire_d61_70),.data_out(wire_d61_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance626172(.data_in(wire_d61_71),.data_out(wire_d61_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance626173(.data_in(wire_d61_72),.data_out(wire_d61_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626174(.data_in(wire_d61_73),.data_out(wire_d61_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626175(.data_in(wire_d61_74),.data_out(wire_d61_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626176(.data_in(wire_d61_75),.data_out(wire_d61_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance626177(.data_in(wire_d61_76),.data_out(wire_d61_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626178(.data_in(wire_d61_77),.data_out(wire_d61_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance626179(.data_in(wire_d61_78),.data_out(wire_d61_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626180(.data_in(wire_d61_79),.data_out(wire_d61_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626181(.data_in(wire_d61_80),.data_out(wire_d61_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626182(.data_in(wire_d61_81),.data_out(wire_d61_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance626183(.data_in(wire_d61_82),.data_out(wire_d61_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance626184(.data_in(wire_d61_83),.data_out(wire_d61_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626185(.data_in(wire_d61_84),.data_out(wire_d61_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626186(.data_in(wire_d61_85),.data_out(wire_d61_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance626187(.data_in(wire_d61_86),.data_out(wire_d61_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance626188(.data_in(wire_d61_87),.data_out(wire_d61_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance626189(.data_in(wire_d61_88),.data_out(wire_d61_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance626190(.data_in(wire_d61_89),.data_out(wire_d61_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance626191(.data_in(wire_d61_90),.data_out(wire_d61_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance626192(.data_in(wire_d61_91),.data_out(wire_d61_92),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance626193(.data_in(wire_d61_92),.data_out(wire_d61_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance626194(.data_in(wire_d61_93),.data_out(wire_d61_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626195(.data_in(wire_d61_94),.data_out(wire_d61_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance626196(.data_in(wire_d61_95),.data_out(wire_d61_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance626197(.data_in(wire_d61_96),.data_out(wire_d61_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance626198(.data_in(wire_d61_97),.data_out(wire_d61_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance626199(.data_in(wire_d61_98),.data_out(d_out61),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance63620(.data_in(d_in62),.data_out(wire_d62_0),.clk(clk),.rst(rst));            //channel 63
	register #(.WIDTH(WIDTH)) register_instance63621(.data_in(wire_d62_0),.data_out(wire_d62_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance63622(.data_in(wire_d62_1),.data_out(wire_d62_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance63623(.data_in(wire_d62_2),.data_out(wire_d62_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance63624(.data_in(wire_d62_3),.data_out(wire_d62_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance63625(.data_in(wire_d62_4),.data_out(wire_d62_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance63626(.data_in(wire_d62_5),.data_out(wire_d62_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance63627(.data_in(wire_d62_6),.data_out(wire_d62_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance63628(.data_in(wire_d62_7),.data_out(wire_d62_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance63629(.data_in(wire_d62_8),.data_out(wire_d62_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636210(.data_in(wire_d62_9),.data_out(wire_d62_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance636211(.data_in(wire_d62_10),.data_out(wire_d62_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636212(.data_in(wire_d62_11),.data_out(wire_d62_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636213(.data_in(wire_d62_12),.data_out(wire_d62_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance636214(.data_in(wire_d62_13),.data_out(wire_d62_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636215(.data_in(wire_d62_14),.data_out(wire_d62_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance636216(.data_in(wire_d62_15),.data_out(wire_d62_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance636217(.data_in(wire_d62_16),.data_out(wire_d62_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance636218(.data_in(wire_d62_17),.data_out(wire_d62_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance636219(.data_in(wire_d62_18),.data_out(wire_d62_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance636220(.data_in(wire_d62_19),.data_out(wire_d62_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636221(.data_in(wire_d62_20),.data_out(wire_d62_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance636222(.data_in(wire_d62_21),.data_out(wire_d62_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance636223(.data_in(wire_d62_22),.data_out(wire_d62_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636224(.data_in(wire_d62_23),.data_out(wire_d62_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance636225(.data_in(wire_d62_24),.data_out(wire_d62_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance636226(.data_in(wire_d62_25),.data_out(wire_d62_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance636227(.data_in(wire_d62_26),.data_out(wire_d62_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636228(.data_in(wire_d62_27),.data_out(wire_d62_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance636229(.data_in(wire_d62_28),.data_out(wire_d62_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance636230(.data_in(wire_d62_29),.data_out(wire_d62_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance636231(.data_in(wire_d62_30),.data_out(wire_d62_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance636232(.data_in(wire_d62_31),.data_out(wire_d62_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance636233(.data_in(wire_d62_32),.data_out(wire_d62_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636234(.data_in(wire_d62_33),.data_out(wire_d62_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance636235(.data_in(wire_d62_34),.data_out(wire_d62_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance636236(.data_in(wire_d62_35),.data_out(wire_d62_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance636237(.data_in(wire_d62_36),.data_out(wire_d62_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance636238(.data_in(wire_d62_37),.data_out(wire_d62_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance636239(.data_in(wire_d62_38),.data_out(wire_d62_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance636240(.data_in(wire_d62_39),.data_out(wire_d62_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance636241(.data_in(wire_d62_40),.data_out(wire_d62_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636242(.data_in(wire_d62_41),.data_out(wire_d62_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance636243(.data_in(wire_d62_42),.data_out(wire_d62_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance636244(.data_in(wire_d62_43),.data_out(wire_d62_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance636245(.data_in(wire_d62_44),.data_out(wire_d62_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636246(.data_in(wire_d62_45),.data_out(wire_d62_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance636247(.data_in(wire_d62_46),.data_out(wire_d62_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance636248(.data_in(wire_d62_47),.data_out(wire_d62_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance636249(.data_in(wire_d62_48),.data_out(wire_d62_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636250(.data_in(wire_d62_49),.data_out(wire_d62_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance636251(.data_in(wire_d62_50),.data_out(wire_d62_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636252(.data_in(wire_d62_51),.data_out(wire_d62_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance636253(.data_in(wire_d62_52),.data_out(wire_d62_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636254(.data_in(wire_d62_53),.data_out(wire_d62_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636255(.data_in(wire_d62_54),.data_out(wire_d62_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636256(.data_in(wire_d62_55),.data_out(wire_d62_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance636257(.data_in(wire_d62_56),.data_out(wire_d62_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance636258(.data_in(wire_d62_57),.data_out(wire_d62_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance636259(.data_in(wire_d62_58),.data_out(wire_d62_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance636260(.data_in(wire_d62_59),.data_out(wire_d62_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance636261(.data_in(wire_d62_60),.data_out(wire_d62_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance636262(.data_in(wire_d62_61),.data_out(wire_d62_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance636263(.data_in(wire_d62_62),.data_out(wire_d62_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance636264(.data_in(wire_d62_63),.data_out(wire_d62_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636265(.data_in(wire_d62_64),.data_out(wire_d62_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance636266(.data_in(wire_d62_65),.data_out(wire_d62_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636267(.data_in(wire_d62_66),.data_out(wire_d62_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance636268(.data_in(wire_d62_67),.data_out(wire_d62_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance636269(.data_in(wire_d62_68),.data_out(wire_d62_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance636270(.data_in(wire_d62_69),.data_out(wire_d62_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance636271(.data_in(wire_d62_70),.data_out(wire_d62_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636272(.data_in(wire_d62_71),.data_out(wire_d62_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636273(.data_in(wire_d62_72),.data_out(wire_d62_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance636274(.data_in(wire_d62_73),.data_out(wire_d62_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance636275(.data_in(wire_d62_74),.data_out(wire_d62_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance636276(.data_in(wire_d62_75),.data_out(wire_d62_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance636277(.data_in(wire_d62_76),.data_out(wire_d62_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636278(.data_in(wire_d62_77),.data_out(wire_d62_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance636279(.data_in(wire_d62_78),.data_out(wire_d62_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance636280(.data_in(wire_d62_79),.data_out(wire_d62_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance636281(.data_in(wire_d62_80),.data_out(wire_d62_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance636282(.data_in(wire_d62_81),.data_out(wire_d62_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance636283(.data_in(wire_d62_82),.data_out(wire_d62_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance636284(.data_in(wire_d62_83),.data_out(wire_d62_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance636285(.data_in(wire_d62_84),.data_out(wire_d62_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636286(.data_in(wire_d62_85),.data_out(wire_d62_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance636287(.data_in(wire_d62_86),.data_out(wire_d62_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance636288(.data_in(wire_d62_87),.data_out(wire_d62_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636289(.data_in(wire_d62_88),.data_out(wire_d62_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance636290(.data_in(wire_d62_89),.data_out(wire_d62_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance636291(.data_in(wire_d62_90),.data_out(wire_d62_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance636292(.data_in(wire_d62_91),.data_out(wire_d62_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance636293(.data_in(wire_d62_92),.data_out(wire_d62_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636294(.data_in(wire_d62_93),.data_out(wire_d62_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance636295(.data_in(wire_d62_94),.data_out(wire_d62_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance636296(.data_in(wire_d62_95),.data_out(wire_d62_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance636297(.data_in(wire_d62_96),.data_out(wire_d62_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance636298(.data_in(wire_d62_97),.data_out(wire_d62_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance636299(.data_in(wire_d62_98),.data_out(d_out62),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance64630(.data_in(d_in63),.data_out(wire_d63_0),.clk(clk),.rst(rst));            //channel 64
	register #(.WIDTH(WIDTH)) register_instance64631(.data_in(wire_d63_0),.data_out(wire_d63_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance64632(.data_in(wire_d63_1),.data_out(wire_d63_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance64633(.data_in(wire_d63_2),.data_out(wire_d63_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance64634(.data_in(wire_d63_3),.data_out(wire_d63_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance64635(.data_in(wire_d63_4),.data_out(wire_d63_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance64636(.data_in(wire_d63_5),.data_out(wire_d63_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance64637(.data_in(wire_d63_6),.data_out(wire_d63_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance64638(.data_in(wire_d63_7),.data_out(wire_d63_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance64639(.data_in(wire_d63_8),.data_out(wire_d63_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance646310(.data_in(wire_d63_9),.data_out(wire_d63_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646311(.data_in(wire_d63_10),.data_out(wire_d63_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646312(.data_in(wire_d63_11),.data_out(wire_d63_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance646313(.data_in(wire_d63_12),.data_out(wire_d63_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646314(.data_in(wire_d63_13),.data_out(wire_d63_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646315(.data_in(wire_d63_14),.data_out(wire_d63_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance646316(.data_in(wire_d63_15),.data_out(wire_d63_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646317(.data_in(wire_d63_16),.data_out(wire_d63_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646318(.data_in(wire_d63_17),.data_out(wire_d63_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646319(.data_in(wire_d63_18),.data_out(wire_d63_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance646320(.data_in(wire_d63_19),.data_out(wire_d63_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646321(.data_in(wire_d63_20),.data_out(wire_d63_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance646322(.data_in(wire_d63_21),.data_out(wire_d63_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646323(.data_in(wire_d63_22),.data_out(wire_d63_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646324(.data_in(wire_d63_23),.data_out(wire_d63_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646325(.data_in(wire_d63_24),.data_out(wire_d63_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance646326(.data_in(wire_d63_25),.data_out(wire_d63_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646327(.data_in(wire_d63_26),.data_out(wire_d63_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646328(.data_in(wire_d63_27),.data_out(wire_d63_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646329(.data_in(wire_d63_28),.data_out(wire_d63_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646330(.data_in(wire_d63_29),.data_out(wire_d63_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646331(.data_in(wire_d63_30),.data_out(wire_d63_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646332(.data_in(wire_d63_31),.data_out(wire_d63_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646333(.data_in(wire_d63_32),.data_out(wire_d63_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance646334(.data_in(wire_d63_33),.data_out(wire_d63_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646335(.data_in(wire_d63_34),.data_out(wire_d63_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646336(.data_in(wire_d63_35),.data_out(wire_d63_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646337(.data_in(wire_d63_36),.data_out(wire_d63_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646338(.data_in(wire_d63_37),.data_out(wire_d63_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance646339(.data_in(wire_d63_38),.data_out(wire_d63_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646340(.data_in(wire_d63_39),.data_out(wire_d63_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646341(.data_in(wire_d63_40),.data_out(wire_d63_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646342(.data_in(wire_d63_41),.data_out(wire_d63_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646343(.data_in(wire_d63_42),.data_out(wire_d63_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646344(.data_in(wire_d63_43),.data_out(wire_d63_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646345(.data_in(wire_d63_44),.data_out(wire_d63_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646346(.data_in(wire_d63_45),.data_out(wire_d63_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646347(.data_in(wire_d63_46),.data_out(wire_d63_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646348(.data_in(wire_d63_47),.data_out(wire_d63_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646349(.data_in(wire_d63_48),.data_out(wire_d63_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646350(.data_in(wire_d63_49),.data_out(wire_d63_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646351(.data_in(wire_d63_50),.data_out(wire_d63_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646352(.data_in(wire_d63_51),.data_out(wire_d63_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646353(.data_in(wire_d63_52),.data_out(wire_d63_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance646354(.data_in(wire_d63_53),.data_out(wire_d63_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646355(.data_in(wire_d63_54),.data_out(wire_d63_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646356(.data_in(wire_d63_55),.data_out(wire_d63_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646357(.data_in(wire_d63_56),.data_out(wire_d63_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646358(.data_in(wire_d63_57),.data_out(wire_d63_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646359(.data_in(wire_d63_58),.data_out(wire_d63_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646360(.data_in(wire_d63_59),.data_out(wire_d63_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance646361(.data_in(wire_d63_60),.data_out(wire_d63_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646362(.data_in(wire_d63_61),.data_out(wire_d63_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646363(.data_in(wire_d63_62),.data_out(wire_d63_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance646364(.data_in(wire_d63_63),.data_out(wire_d63_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646365(.data_in(wire_d63_64),.data_out(wire_d63_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646366(.data_in(wire_d63_65),.data_out(wire_d63_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646367(.data_in(wire_d63_66),.data_out(wire_d63_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646368(.data_in(wire_d63_67),.data_out(wire_d63_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646369(.data_in(wire_d63_68),.data_out(wire_d63_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance646370(.data_in(wire_d63_69),.data_out(wire_d63_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646371(.data_in(wire_d63_70),.data_out(wire_d63_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646372(.data_in(wire_d63_71),.data_out(wire_d63_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646373(.data_in(wire_d63_72),.data_out(wire_d63_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance646374(.data_in(wire_d63_73),.data_out(wire_d63_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance646375(.data_in(wire_d63_74),.data_out(wire_d63_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646376(.data_in(wire_d63_75),.data_out(wire_d63_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646377(.data_in(wire_d63_76),.data_out(wire_d63_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance646378(.data_in(wire_d63_77),.data_out(wire_d63_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646379(.data_in(wire_d63_78),.data_out(wire_d63_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646380(.data_in(wire_d63_79),.data_out(wire_d63_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance646381(.data_in(wire_d63_80),.data_out(wire_d63_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646382(.data_in(wire_d63_81),.data_out(wire_d63_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646383(.data_in(wire_d63_82),.data_out(wire_d63_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646384(.data_in(wire_d63_83),.data_out(wire_d63_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance646385(.data_in(wire_d63_84),.data_out(wire_d63_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance646386(.data_in(wire_d63_85),.data_out(wire_d63_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646387(.data_in(wire_d63_86),.data_out(wire_d63_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance646388(.data_in(wire_d63_87),.data_out(wire_d63_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646389(.data_in(wire_d63_88),.data_out(wire_d63_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646390(.data_in(wire_d63_89),.data_out(wire_d63_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646391(.data_in(wire_d63_90),.data_out(wire_d63_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646392(.data_in(wire_d63_91),.data_out(wire_d63_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance646393(.data_in(wire_d63_92),.data_out(wire_d63_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance646394(.data_in(wire_d63_93),.data_out(wire_d63_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646395(.data_in(wire_d63_94),.data_out(wire_d63_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646396(.data_in(wire_d63_95),.data_out(wire_d63_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance646397(.data_in(wire_d63_96),.data_out(wire_d63_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance646398(.data_in(wire_d63_97),.data_out(wire_d63_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance646399(.data_in(wire_d63_98),.data_out(d_out63),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance65640(.data_in(d_in64),.data_out(wire_d64_0),.clk(clk),.rst(rst));            //channel 65
	encoder #(.WIDTH(WIDTH)) encoder_instance65641(.data_in(wire_d64_0),.data_out(wire_d64_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance65642(.data_in(wire_d64_1),.data_out(wire_d64_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65643(.data_in(wire_d64_2),.data_out(wire_d64_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance65644(.data_in(wire_d64_3),.data_out(wire_d64_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance65645(.data_in(wire_d64_4),.data_out(wire_d64_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance65646(.data_in(wire_d64_5),.data_out(wire_d64_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance65647(.data_in(wire_d64_6),.data_out(wire_d64_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance65648(.data_in(wire_d64_7),.data_out(wire_d64_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65649(.data_in(wire_d64_8),.data_out(wire_d64_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance656410(.data_in(wire_d64_9),.data_out(wire_d64_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656411(.data_in(wire_d64_10),.data_out(wire_d64_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656412(.data_in(wire_d64_11),.data_out(wire_d64_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656413(.data_in(wire_d64_12),.data_out(wire_d64_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance656414(.data_in(wire_d64_13),.data_out(wire_d64_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656415(.data_in(wire_d64_14),.data_out(wire_d64_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656416(.data_in(wire_d64_15),.data_out(wire_d64_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656417(.data_in(wire_d64_16),.data_out(wire_d64_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656418(.data_in(wire_d64_17),.data_out(wire_d64_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656419(.data_in(wire_d64_18),.data_out(wire_d64_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656420(.data_in(wire_d64_19),.data_out(wire_d64_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656421(.data_in(wire_d64_20),.data_out(wire_d64_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance656422(.data_in(wire_d64_21),.data_out(wire_d64_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance656423(.data_in(wire_d64_22),.data_out(wire_d64_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656424(.data_in(wire_d64_23),.data_out(wire_d64_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656425(.data_in(wire_d64_24),.data_out(wire_d64_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656426(.data_in(wire_d64_25),.data_out(wire_d64_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656427(.data_in(wire_d64_26),.data_out(wire_d64_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656428(.data_in(wire_d64_27),.data_out(wire_d64_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656429(.data_in(wire_d64_28),.data_out(wire_d64_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656430(.data_in(wire_d64_29),.data_out(wire_d64_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance656431(.data_in(wire_d64_30),.data_out(wire_d64_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656432(.data_in(wire_d64_31),.data_out(wire_d64_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656433(.data_in(wire_d64_32),.data_out(wire_d64_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656434(.data_in(wire_d64_33),.data_out(wire_d64_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656435(.data_in(wire_d64_34),.data_out(wire_d64_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656436(.data_in(wire_d64_35),.data_out(wire_d64_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656437(.data_in(wire_d64_36),.data_out(wire_d64_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656438(.data_in(wire_d64_37),.data_out(wire_d64_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656439(.data_in(wire_d64_38),.data_out(wire_d64_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656440(.data_in(wire_d64_39),.data_out(wire_d64_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance656441(.data_in(wire_d64_40),.data_out(wire_d64_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656442(.data_in(wire_d64_41),.data_out(wire_d64_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656443(.data_in(wire_d64_42),.data_out(wire_d64_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656444(.data_in(wire_d64_43),.data_out(wire_d64_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance656445(.data_in(wire_d64_44),.data_out(wire_d64_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656446(.data_in(wire_d64_45),.data_out(wire_d64_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656447(.data_in(wire_d64_46),.data_out(wire_d64_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656448(.data_in(wire_d64_47),.data_out(wire_d64_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656449(.data_in(wire_d64_48),.data_out(wire_d64_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656450(.data_in(wire_d64_49),.data_out(wire_d64_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656451(.data_in(wire_d64_50),.data_out(wire_d64_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656452(.data_in(wire_d64_51),.data_out(wire_d64_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance656453(.data_in(wire_d64_52),.data_out(wire_d64_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance656454(.data_in(wire_d64_53),.data_out(wire_d64_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656455(.data_in(wire_d64_54),.data_out(wire_d64_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance656456(.data_in(wire_d64_55),.data_out(wire_d64_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656457(.data_in(wire_d64_56),.data_out(wire_d64_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656458(.data_in(wire_d64_57),.data_out(wire_d64_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656459(.data_in(wire_d64_58),.data_out(wire_d64_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance656460(.data_in(wire_d64_59),.data_out(wire_d64_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656461(.data_in(wire_d64_60),.data_out(wire_d64_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656462(.data_in(wire_d64_61),.data_out(wire_d64_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656463(.data_in(wire_d64_62),.data_out(wire_d64_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance656464(.data_in(wire_d64_63),.data_out(wire_d64_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656465(.data_in(wire_d64_64),.data_out(wire_d64_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656466(.data_in(wire_d64_65),.data_out(wire_d64_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance656467(.data_in(wire_d64_66),.data_out(wire_d64_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656468(.data_in(wire_d64_67),.data_out(wire_d64_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance656469(.data_in(wire_d64_68),.data_out(wire_d64_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656470(.data_in(wire_d64_69),.data_out(wire_d64_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656471(.data_in(wire_d64_70),.data_out(wire_d64_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656472(.data_in(wire_d64_71),.data_out(wire_d64_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656473(.data_in(wire_d64_72),.data_out(wire_d64_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656474(.data_in(wire_d64_73),.data_out(wire_d64_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656475(.data_in(wire_d64_74),.data_out(wire_d64_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance656476(.data_in(wire_d64_75),.data_out(wire_d64_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance656477(.data_in(wire_d64_76),.data_out(wire_d64_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656478(.data_in(wire_d64_77),.data_out(wire_d64_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656479(.data_in(wire_d64_78),.data_out(wire_d64_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656480(.data_in(wire_d64_79),.data_out(wire_d64_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656481(.data_in(wire_d64_80),.data_out(wire_d64_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656482(.data_in(wire_d64_81),.data_out(wire_d64_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656483(.data_in(wire_d64_82),.data_out(wire_d64_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656484(.data_in(wire_d64_83),.data_out(wire_d64_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656485(.data_in(wire_d64_84),.data_out(wire_d64_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656486(.data_in(wire_d64_85),.data_out(wire_d64_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance656487(.data_in(wire_d64_86),.data_out(wire_d64_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656488(.data_in(wire_d64_87),.data_out(wire_d64_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance656489(.data_in(wire_d64_88),.data_out(wire_d64_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656490(.data_in(wire_d64_89),.data_out(wire_d64_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656491(.data_in(wire_d64_90),.data_out(wire_d64_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656492(.data_in(wire_d64_91),.data_out(wire_d64_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance656493(.data_in(wire_d64_92),.data_out(wire_d64_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance656494(.data_in(wire_d64_93),.data_out(wire_d64_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance656495(.data_in(wire_d64_94),.data_out(wire_d64_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656496(.data_in(wire_d64_95),.data_out(wire_d64_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656497(.data_in(wire_d64_96),.data_out(wire_d64_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656498(.data_in(wire_d64_97),.data_out(wire_d64_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance656499(.data_in(wire_d64_98),.data_out(d_out64),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance66650(.data_in(d_in65),.data_out(wire_d65_0),.clk(clk),.rst(rst));            //channel 66
	large_mux #(.WIDTH(WIDTH)) large_mux_instance66651(.data_in(wire_d65_0),.data_out(wire_d65_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance66652(.data_in(wire_d65_1),.data_out(wire_d65_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance66653(.data_in(wire_d65_2),.data_out(wire_d65_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance66654(.data_in(wire_d65_3),.data_out(wire_d65_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance66655(.data_in(wire_d65_4),.data_out(wire_d65_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance66656(.data_in(wire_d65_5),.data_out(wire_d65_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance66657(.data_in(wire_d65_6),.data_out(wire_d65_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance66658(.data_in(wire_d65_7),.data_out(wire_d65_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance66659(.data_in(wire_d65_8),.data_out(wire_d65_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666510(.data_in(wire_d65_9),.data_out(wire_d65_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance666511(.data_in(wire_d65_10),.data_out(wire_d65_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666512(.data_in(wire_d65_11),.data_out(wire_d65_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance666513(.data_in(wire_d65_12),.data_out(wire_d65_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666514(.data_in(wire_d65_13),.data_out(wire_d65_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666515(.data_in(wire_d65_14),.data_out(wire_d65_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance666516(.data_in(wire_d65_15),.data_out(wire_d65_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666517(.data_in(wire_d65_16),.data_out(wire_d65_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance666518(.data_in(wire_d65_17),.data_out(wire_d65_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666519(.data_in(wire_d65_18),.data_out(wire_d65_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666520(.data_in(wire_d65_19),.data_out(wire_d65_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666521(.data_in(wire_d65_20),.data_out(wire_d65_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666522(.data_in(wire_d65_21),.data_out(wire_d65_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance666523(.data_in(wire_d65_22),.data_out(wire_d65_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance666524(.data_in(wire_d65_23),.data_out(wire_d65_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance666525(.data_in(wire_d65_24),.data_out(wire_d65_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance666526(.data_in(wire_d65_25),.data_out(wire_d65_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666527(.data_in(wire_d65_26),.data_out(wire_d65_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance666528(.data_in(wire_d65_27),.data_out(wire_d65_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance666529(.data_in(wire_d65_28),.data_out(wire_d65_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666530(.data_in(wire_d65_29),.data_out(wire_d65_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666531(.data_in(wire_d65_30),.data_out(wire_d65_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance666532(.data_in(wire_d65_31),.data_out(wire_d65_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance666533(.data_in(wire_d65_32),.data_out(wire_d65_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance666534(.data_in(wire_d65_33),.data_out(wire_d65_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance666535(.data_in(wire_d65_34),.data_out(wire_d65_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666536(.data_in(wire_d65_35),.data_out(wire_d65_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666537(.data_in(wire_d65_36),.data_out(wire_d65_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance666538(.data_in(wire_d65_37),.data_out(wire_d65_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666539(.data_in(wire_d65_38),.data_out(wire_d65_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance666540(.data_in(wire_d65_39),.data_out(wire_d65_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance666541(.data_in(wire_d65_40),.data_out(wire_d65_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance666542(.data_in(wire_d65_41),.data_out(wire_d65_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666543(.data_in(wire_d65_42),.data_out(wire_d65_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance666544(.data_in(wire_d65_43),.data_out(wire_d65_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666545(.data_in(wire_d65_44),.data_out(wire_d65_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance666546(.data_in(wire_d65_45),.data_out(wire_d65_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance666547(.data_in(wire_d65_46),.data_out(wire_d65_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666548(.data_in(wire_d65_47),.data_out(wire_d65_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance666549(.data_in(wire_d65_48),.data_out(wire_d65_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance666550(.data_in(wire_d65_49),.data_out(wire_d65_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666551(.data_in(wire_d65_50),.data_out(wire_d65_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance666552(.data_in(wire_d65_51),.data_out(wire_d65_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666553(.data_in(wire_d65_52),.data_out(wire_d65_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance666554(.data_in(wire_d65_53),.data_out(wire_d65_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666555(.data_in(wire_d65_54),.data_out(wire_d65_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance666556(.data_in(wire_d65_55),.data_out(wire_d65_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666557(.data_in(wire_d65_56),.data_out(wire_d65_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666558(.data_in(wire_d65_57),.data_out(wire_d65_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance666559(.data_in(wire_d65_58),.data_out(wire_d65_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666560(.data_in(wire_d65_59),.data_out(wire_d65_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666561(.data_in(wire_d65_60),.data_out(wire_d65_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666562(.data_in(wire_d65_61),.data_out(wire_d65_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance666563(.data_in(wire_d65_62),.data_out(wire_d65_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance666564(.data_in(wire_d65_63),.data_out(wire_d65_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666565(.data_in(wire_d65_64),.data_out(wire_d65_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance666566(.data_in(wire_d65_65),.data_out(wire_d65_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666567(.data_in(wire_d65_66),.data_out(wire_d65_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666568(.data_in(wire_d65_67),.data_out(wire_d65_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666569(.data_in(wire_d65_68),.data_out(wire_d65_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance666570(.data_in(wire_d65_69),.data_out(wire_d65_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666571(.data_in(wire_d65_70),.data_out(wire_d65_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666572(.data_in(wire_d65_71),.data_out(wire_d65_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance666573(.data_in(wire_d65_72),.data_out(wire_d65_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance666574(.data_in(wire_d65_73),.data_out(wire_d65_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666575(.data_in(wire_d65_74),.data_out(wire_d65_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance666576(.data_in(wire_d65_75),.data_out(wire_d65_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance666577(.data_in(wire_d65_76),.data_out(wire_d65_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance666578(.data_in(wire_d65_77),.data_out(wire_d65_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance666579(.data_in(wire_d65_78),.data_out(wire_d65_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance666580(.data_in(wire_d65_79),.data_out(wire_d65_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance666581(.data_in(wire_d65_80),.data_out(wire_d65_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance666582(.data_in(wire_d65_81),.data_out(wire_d65_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666583(.data_in(wire_d65_82),.data_out(wire_d65_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666584(.data_in(wire_d65_83),.data_out(wire_d65_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666585(.data_in(wire_d65_84),.data_out(wire_d65_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666586(.data_in(wire_d65_85),.data_out(wire_d65_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666587(.data_in(wire_d65_86),.data_out(wire_d65_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666588(.data_in(wire_d65_87),.data_out(wire_d65_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666589(.data_in(wire_d65_88),.data_out(wire_d65_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666590(.data_in(wire_d65_89),.data_out(wire_d65_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666591(.data_in(wire_d65_90),.data_out(wire_d65_91),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666592(.data_in(wire_d65_91),.data_out(wire_d65_92),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666593(.data_in(wire_d65_92),.data_out(wire_d65_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666594(.data_in(wire_d65_93),.data_out(wire_d65_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666595(.data_in(wire_d65_94),.data_out(wire_d65_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance666596(.data_in(wire_d65_95),.data_out(wire_d65_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance666597(.data_in(wire_d65_96),.data_out(wire_d65_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance666598(.data_in(wire_d65_97),.data_out(wire_d65_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance666599(.data_in(wire_d65_98),.data_out(d_out65),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance67660(.data_in(d_in66),.data_out(wire_d66_0),.clk(clk),.rst(rst));            //channel 67
	invertion #(.WIDTH(WIDTH)) invertion_instance67661(.data_in(wire_d66_0),.data_out(wire_d66_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance67662(.data_in(wire_d66_1),.data_out(wire_d66_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance67663(.data_in(wire_d66_2),.data_out(wire_d66_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance67664(.data_in(wire_d66_3),.data_out(wire_d66_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance67665(.data_in(wire_d66_4),.data_out(wire_d66_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance67666(.data_in(wire_d66_5),.data_out(wire_d66_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance67667(.data_in(wire_d66_6),.data_out(wire_d66_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance67668(.data_in(wire_d66_7),.data_out(wire_d66_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance67669(.data_in(wire_d66_8),.data_out(wire_d66_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance676610(.data_in(wire_d66_9),.data_out(wire_d66_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance676611(.data_in(wire_d66_10),.data_out(wire_d66_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676612(.data_in(wire_d66_11),.data_out(wire_d66_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676613(.data_in(wire_d66_12),.data_out(wire_d66_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676614(.data_in(wire_d66_13),.data_out(wire_d66_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676615(.data_in(wire_d66_14),.data_out(wire_d66_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676616(.data_in(wire_d66_15),.data_out(wire_d66_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance676617(.data_in(wire_d66_16),.data_out(wire_d66_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance676618(.data_in(wire_d66_17),.data_out(wire_d66_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676619(.data_in(wire_d66_18),.data_out(wire_d66_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676620(.data_in(wire_d66_19),.data_out(wire_d66_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance676621(.data_in(wire_d66_20),.data_out(wire_d66_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676622(.data_in(wire_d66_21),.data_out(wire_d66_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance676623(.data_in(wire_d66_22),.data_out(wire_d66_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance676624(.data_in(wire_d66_23),.data_out(wire_d66_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676625(.data_in(wire_d66_24),.data_out(wire_d66_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676626(.data_in(wire_d66_25),.data_out(wire_d66_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance676627(.data_in(wire_d66_26),.data_out(wire_d66_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676628(.data_in(wire_d66_27),.data_out(wire_d66_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance676629(.data_in(wire_d66_28),.data_out(wire_d66_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676630(.data_in(wire_d66_29),.data_out(wire_d66_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676631(.data_in(wire_d66_30),.data_out(wire_d66_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676632(.data_in(wire_d66_31),.data_out(wire_d66_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance676633(.data_in(wire_d66_32),.data_out(wire_d66_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676634(.data_in(wire_d66_33),.data_out(wire_d66_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance676635(.data_in(wire_d66_34),.data_out(wire_d66_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance676636(.data_in(wire_d66_35),.data_out(wire_d66_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance676637(.data_in(wire_d66_36),.data_out(wire_d66_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance676638(.data_in(wire_d66_37),.data_out(wire_d66_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676639(.data_in(wire_d66_38),.data_out(wire_d66_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676640(.data_in(wire_d66_39),.data_out(wire_d66_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676641(.data_in(wire_d66_40),.data_out(wire_d66_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance676642(.data_in(wire_d66_41),.data_out(wire_d66_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance676643(.data_in(wire_d66_42),.data_out(wire_d66_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676644(.data_in(wire_d66_43),.data_out(wire_d66_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676645(.data_in(wire_d66_44),.data_out(wire_d66_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance676646(.data_in(wire_d66_45),.data_out(wire_d66_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance676647(.data_in(wire_d66_46),.data_out(wire_d66_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance676648(.data_in(wire_d66_47),.data_out(wire_d66_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance676649(.data_in(wire_d66_48),.data_out(wire_d66_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance676650(.data_in(wire_d66_49),.data_out(wire_d66_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676651(.data_in(wire_d66_50),.data_out(wire_d66_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676652(.data_in(wire_d66_51),.data_out(wire_d66_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676653(.data_in(wire_d66_52),.data_out(wire_d66_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676654(.data_in(wire_d66_53),.data_out(wire_d66_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676655(.data_in(wire_d66_54),.data_out(wire_d66_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676656(.data_in(wire_d66_55),.data_out(wire_d66_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676657(.data_in(wire_d66_56),.data_out(wire_d66_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance676658(.data_in(wire_d66_57),.data_out(wire_d66_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance676659(.data_in(wire_d66_58),.data_out(wire_d66_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance676660(.data_in(wire_d66_59),.data_out(wire_d66_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676661(.data_in(wire_d66_60),.data_out(wire_d66_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance676662(.data_in(wire_d66_61),.data_out(wire_d66_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676663(.data_in(wire_d66_62),.data_out(wire_d66_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance676664(.data_in(wire_d66_63),.data_out(wire_d66_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance676665(.data_in(wire_d66_64),.data_out(wire_d66_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676666(.data_in(wire_d66_65),.data_out(wire_d66_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance676667(.data_in(wire_d66_66),.data_out(wire_d66_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance676668(.data_in(wire_d66_67),.data_out(wire_d66_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance676669(.data_in(wire_d66_68),.data_out(wire_d66_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676670(.data_in(wire_d66_69),.data_out(wire_d66_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676671(.data_in(wire_d66_70),.data_out(wire_d66_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676672(.data_in(wire_d66_71),.data_out(wire_d66_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance676673(.data_in(wire_d66_72),.data_out(wire_d66_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676674(.data_in(wire_d66_73),.data_out(wire_d66_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676675(.data_in(wire_d66_74),.data_out(wire_d66_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676676(.data_in(wire_d66_75),.data_out(wire_d66_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance676677(.data_in(wire_d66_76),.data_out(wire_d66_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676678(.data_in(wire_d66_77),.data_out(wire_d66_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676679(.data_in(wire_d66_78),.data_out(wire_d66_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676680(.data_in(wire_d66_79),.data_out(wire_d66_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance676681(.data_in(wire_d66_80),.data_out(wire_d66_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676682(.data_in(wire_d66_81),.data_out(wire_d66_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676683(.data_in(wire_d66_82),.data_out(wire_d66_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance676684(.data_in(wire_d66_83),.data_out(wire_d66_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance676685(.data_in(wire_d66_84),.data_out(wire_d66_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance676686(.data_in(wire_d66_85),.data_out(wire_d66_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676687(.data_in(wire_d66_86),.data_out(wire_d66_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance676688(.data_in(wire_d66_87),.data_out(wire_d66_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676689(.data_in(wire_d66_88),.data_out(wire_d66_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance676690(.data_in(wire_d66_89),.data_out(wire_d66_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance676691(.data_in(wire_d66_90),.data_out(wire_d66_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676692(.data_in(wire_d66_91),.data_out(wire_d66_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance676693(.data_in(wire_d66_92),.data_out(wire_d66_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676694(.data_in(wire_d66_93),.data_out(wire_d66_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676695(.data_in(wire_d66_94),.data_out(wire_d66_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance676696(.data_in(wire_d66_95),.data_out(wire_d66_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance676697(.data_in(wire_d66_96),.data_out(wire_d66_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance676698(.data_in(wire_d66_97),.data_out(wire_d66_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance676699(.data_in(wire_d66_98),.data_out(d_out66),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance68670(.data_in(d_in67),.data_out(wire_d67_0),.clk(clk),.rst(rst));            //channel 68
	invertion #(.WIDTH(WIDTH)) invertion_instance68671(.data_in(wire_d67_0),.data_out(wire_d67_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance68672(.data_in(wire_d67_1),.data_out(wire_d67_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance68673(.data_in(wire_d67_2),.data_out(wire_d67_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance68674(.data_in(wire_d67_3),.data_out(wire_d67_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance68675(.data_in(wire_d67_4),.data_out(wire_d67_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance68676(.data_in(wire_d67_5),.data_out(wire_d67_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance68677(.data_in(wire_d67_6),.data_out(wire_d67_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance68678(.data_in(wire_d67_7),.data_out(wire_d67_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance68679(.data_in(wire_d67_8),.data_out(wire_d67_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance686710(.data_in(wire_d67_9),.data_out(wire_d67_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686711(.data_in(wire_d67_10),.data_out(wire_d67_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686712(.data_in(wire_d67_11),.data_out(wire_d67_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686713(.data_in(wire_d67_12),.data_out(wire_d67_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance686714(.data_in(wire_d67_13),.data_out(wire_d67_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686715(.data_in(wire_d67_14),.data_out(wire_d67_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686716(.data_in(wire_d67_15),.data_out(wire_d67_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686717(.data_in(wire_d67_16),.data_out(wire_d67_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686718(.data_in(wire_d67_17),.data_out(wire_d67_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance686719(.data_in(wire_d67_18),.data_out(wire_d67_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance686720(.data_in(wire_d67_19),.data_out(wire_d67_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance686721(.data_in(wire_d67_20),.data_out(wire_d67_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686722(.data_in(wire_d67_21),.data_out(wire_d67_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance686723(.data_in(wire_d67_22),.data_out(wire_d67_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance686724(.data_in(wire_d67_23),.data_out(wire_d67_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686725(.data_in(wire_d67_24),.data_out(wire_d67_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686726(.data_in(wire_d67_25),.data_out(wire_d67_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686727(.data_in(wire_d67_26),.data_out(wire_d67_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686728(.data_in(wire_d67_27),.data_out(wire_d67_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686729(.data_in(wire_d67_28),.data_out(wire_d67_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance686730(.data_in(wire_d67_29),.data_out(wire_d67_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686731(.data_in(wire_d67_30),.data_out(wire_d67_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686732(.data_in(wire_d67_31),.data_out(wire_d67_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance686733(.data_in(wire_d67_32),.data_out(wire_d67_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance686734(.data_in(wire_d67_33),.data_out(wire_d67_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance686735(.data_in(wire_d67_34),.data_out(wire_d67_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance686736(.data_in(wire_d67_35),.data_out(wire_d67_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686737(.data_in(wire_d67_36),.data_out(wire_d67_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686738(.data_in(wire_d67_37),.data_out(wire_d67_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance686739(.data_in(wire_d67_38),.data_out(wire_d67_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance686740(.data_in(wire_d67_39),.data_out(wire_d67_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686741(.data_in(wire_d67_40),.data_out(wire_d67_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686742(.data_in(wire_d67_41),.data_out(wire_d67_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686743(.data_in(wire_d67_42),.data_out(wire_d67_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance686744(.data_in(wire_d67_43),.data_out(wire_d67_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance686745(.data_in(wire_d67_44),.data_out(wire_d67_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance686746(.data_in(wire_d67_45),.data_out(wire_d67_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686747(.data_in(wire_d67_46),.data_out(wire_d67_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686748(.data_in(wire_d67_47),.data_out(wire_d67_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance686749(.data_in(wire_d67_48),.data_out(wire_d67_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance686750(.data_in(wire_d67_49),.data_out(wire_d67_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance686751(.data_in(wire_d67_50),.data_out(wire_d67_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance686752(.data_in(wire_d67_51),.data_out(wire_d67_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686753(.data_in(wire_d67_52),.data_out(wire_d67_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686754(.data_in(wire_d67_53),.data_out(wire_d67_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686755(.data_in(wire_d67_54),.data_out(wire_d67_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance686756(.data_in(wire_d67_55),.data_out(wire_d67_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance686757(.data_in(wire_d67_56),.data_out(wire_d67_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686758(.data_in(wire_d67_57),.data_out(wire_d67_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance686759(.data_in(wire_d67_58),.data_out(wire_d67_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance686760(.data_in(wire_d67_59),.data_out(wire_d67_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance686761(.data_in(wire_d67_60),.data_out(wire_d67_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance686762(.data_in(wire_d67_61),.data_out(wire_d67_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance686763(.data_in(wire_d67_62),.data_out(wire_d67_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686764(.data_in(wire_d67_63),.data_out(wire_d67_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance686765(.data_in(wire_d67_64),.data_out(wire_d67_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686766(.data_in(wire_d67_65),.data_out(wire_d67_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686767(.data_in(wire_d67_66),.data_out(wire_d67_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686768(.data_in(wire_d67_67),.data_out(wire_d67_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance686769(.data_in(wire_d67_68),.data_out(wire_d67_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance686770(.data_in(wire_d67_69),.data_out(wire_d67_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance686771(.data_in(wire_d67_70),.data_out(wire_d67_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance686772(.data_in(wire_d67_71),.data_out(wire_d67_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686773(.data_in(wire_d67_72),.data_out(wire_d67_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686774(.data_in(wire_d67_73),.data_out(wire_d67_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686775(.data_in(wire_d67_74),.data_out(wire_d67_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance686776(.data_in(wire_d67_75),.data_out(wire_d67_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686777(.data_in(wire_d67_76),.data_out(wire_d67_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686778(.data_in(wire_d67_77),.data_out(wire_d67_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686779(.data_in(wire_d67_78),.data_out(wire_d67_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance686780(.data_in(wire_d67_79),.data_out(wire_d67_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686781(.data_in(wire_d67_80),.data_out(wire_d67_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance686782(.data_in(wire_d67_81),.data_out(wire_d67_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686783(.data_in(wire_d67_82),.data_out(wire_d67_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance686784(.data_in(wire_d67_83),.data_out(wire_d67_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance686785(.data_in(wire_d67_84),.data_out(wire_d67_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686786(.data_in(wire_d67_85),.data_out(wire_d67_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686787(.data_in(wire_d67_86),.data_out(wire_d67_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance686788(.data_in(wire_d67_87),.data_out(wire_d67_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686789(.data_in(wire_d67_88),.data_out(wire_d67_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance686790(.data_in(wire_d67_89),.data_out(wire_d67_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686791(.data_in(wire_d67_90),.data_out(wire_d67_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686792(.data_in(wire_d67_91),.data_out(wire_d67_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance686793(.data_in(wire_d67_92),.data_out(wire_d67_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance686794(.data_in(wire_d67_93),.data_out(wire_d67_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance686795(.data_in(wire_d67_94),.data_out(wire_d67_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686796(.data_in(wire_d67_95),.data_out(wire_d67_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance686797(.data_in(wire_d67_96),.data_out(wire_d67_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance686798(.data_in(wire_d67_97),.data_out(wire_d67_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance686799(.data_in(wire_d67_98),.data_out(d_out67),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance69680(.data_in(d_in68),.data_out(wire_d68_0),.clk(clk),.rst(rst));            //channel 69
	large_mux #(.WIDTH(WIDTH)) large_mux_instance69681(.data_in(wire_d68_0),.data_out(wire_d68_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance69682(.data_in(wire_d68_1),.data_out(wire_d68_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance69683(.data_in(wire_d68_2),.data_out(wire_d68_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance69684(.data_in(wire_d68_3),.data_out(wire_d68_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance69685(.data_in(wire_d68_4),.data_out(wire_d68_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance69686(.data_in(wire_d68_5),.data_out(wire_d68_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance69687(.data_in(wire_d68_6),.data_out(wire_d68_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance69688(.data_in(wire_d68_7),.data_out(wire_d68_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance69689(.data_in(wire_d68_8),.data_out(wire_d68_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696810(.data_in(wire_d68_9),.data_out(wire_d68_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696811(.data_in(wire_d68_10),.data_out(wire_d68_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696812(.data_in(wire_d68_11),.data_out(wire_d68_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance696813(.data_in(wire_d68_12),.data_out(wire_d68_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance696814(.data_in(wire_d68_13),.data_out(wire_d68_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance696815(.data_in(wire_d68_14),.data_out(wire_d68_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696816(.data_in(wire_d68_15),.data_out(wire_d68_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696817(.data_in(wire_d68_16),.data_out(wire_d68_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696818(.data_in(wire_d68_17),.data_out(wire_d68_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance696819(.data_in(wire_d68_18),.data_out(wire_d68_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696820(.data_in(wire_d68_19),.data_out(wire_d68_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696821(.data_in(wire_d68_20),.data_out(wire_d68_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance696822(.data_in(wire_d68_21),.data_out(wire_d68_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance696823(.data_in(wire_d68_22),.data_out(wire_d68_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance696824(.data_in(wire_d68_23),.data_out(wire_d68_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696825(.data_in(wire_d68_24),.data_out(wire_d68_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance696826(.data_in(wire_d68_25),.data_out(wire_d68_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696827(.data_in(wire_d68_26),.data_out(wire_d68_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance696828(.data_in(wire_d68_27),.data_out(wire_d68_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance696829(.data_in(wire_d68_28),.data_out(wire_d68_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696830(.data_in(wire_d68_29),.data_out(wire_d68_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance696831(.data_in(wire_d68_30),.data_out(wire_d68_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance696832(.data_in(wire_d68_31),.data_out(wire_d68_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance696833(.data_in(wire_d68_32),.data_out(wire_d68_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696834(.data_in(wire_d68_33),.data_out(wire_d68_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696835(.data_in(wire_d68_34),.data_out(wire_d68_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance696836(.data_in(wire_d68_35),.data_out(wire_d68_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696837(.data_in(wire_d68_36),.data_out(wire_d68_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696838(.data_in(wire_d68_37),.data_out(wire_d68_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance696839(.data_in(wire_d68_38),.data_out(wire_d68_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696840(.data_in(wire_d68_39),.data_out(wire_d68_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696841(.data_in(wire_d68_40),.data_out(wire_d68_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696842(.data_in(wire_d68_41),.data_out(wire_d68_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696843(.data_in(wire_d68_42),.data_out(wire_d68_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696844(.data_in(wire_d68_43),.data_out(wire_d68_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance696845(.data_in(wire_d68_44),.data_out(wire_d68_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696846(.data_in(wire_d68_45),.data_out(wire_d68_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance696847(.data_in(wire_d68_46),.data_out(wire_d68_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696848(.data_in(wire_d68_47),.data_out(wire_d68_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696849(.data_in(wire_d68_48),.data_out(wire_d68_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696850(.data_in(wire_d68_49),.data_out(wire_d68_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696851(.data_in(wire_d68_50),.data_out(wire_d68_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance696852(.data_in(wire_d68_51),.data_out(wire_d68_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance696853(.data_in(wire_d68_52),.data_out(wire_d68_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance696854(.data_in(wire_d68_53),.data_out(wire_d68_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance696855(.data_in(wire_d68_54),.data_out(wire_d68_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance696856(.data_in(wire_d68_55),.data_out(wire_d68_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696857(.data_in(wire_d68_56),.data_out(wire_d68_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696858(.data_in(wire_d68_57),.data_out(wire_d68_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance696859(.data_in(wire_d68_58),.data_out(wire_d68_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance696860(.data_in(wire_d68_59),.data_out(wire_d68_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance696861(.data_in(wire_d68_60),.data_out(wire_d68_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696862(.data_in(wire_d68_61),.data_out(wire_d68_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696863(.data_in(wire_d68_62),.data_out(wire_d68_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696864(.data_in(wire_d68_63),.data_out(wire_d68_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696865(.data_in(wire_d68_64),.data_out(wire_d68_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696866(.data_in(wire_d68_65),.data_out(wire_d68_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696867(.data_in(wire_d68_66),.data_out(wire_d68_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696868(.data_in(wire_d68_67),.data_out(wire_d68_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance696869(.data_in(wire_d68_68),.data_out(wire_d68_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance696870(.data_in(wire_d68_69),.data_out(wire_d68_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696871(.data_in(wire_d68_70),.data_out(wire_d68_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance696872(.data_in(wire_d68_71),.data_out(wire_d68_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696873(.data_in(wire_d68_72),.data_out(wire_d68_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696874(.data_in(wire_d68_73),.data_out(wire_d68_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696875(.data_in(wire_d68_74),.data_out(wire_d68_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance696876(.data_in(wire_d68_75),.data_out(wire_d68_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696877(.data_in(wire_d68_76),.data_out(wire_d68_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696878(.data_in(wire_d68_77),.data_out(wire_d68_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance696879(.data_in(wire_d68_78),.data_out(wire_d68_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696880(.data_in(wire_d68_79),.data_out(wire_d68_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696881(.data_in(wire_d68_80),.data_out(wire_d68_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696882(.data_in(wire_d68_81),.data_out(wire_d68_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance696883(.data_in(wire_d68_82),.data_out(wire_d68_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance696884(.data_in(wire_d68_83),.data_out(wire_d68_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696885(.data_in(wire_d68_84),.data_out(wire_d68_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance696886(.data_in(wire_d68_85),.data_out(wire_d68_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance696887(.data_in(wire_d68_86),.data_out(wire_d68_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance696888(.data_in(wire_d68_87),.data_out(wire_d68_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696889(.data_in(wire_d68_88),.data_out(wire_d68_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance696890(.data_in(wire_d68_89),.data_out(wire_d68_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance696891(.data_in(wire_d68_90),.data_out(wire_d68_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance696892(.data_in(wire_d68_91),.data_out(wire_d68_92),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696893(.data_in(wire_d68_92),.data_out(wire_d68_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance696894(.data_in(wire_d68_93),.data_out(wire_d68_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance696895(.data_in(wire_d68_94),.data_out(wire_d68_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance696896(.data_in(wire_d68_95),.data_out(wire_d68_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance696897(.data_in(wire_d68_96),.data_out(wire_d68_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance696898(.data_in(wire_d68_97),.data_out(wire_d68_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance696899(.data_in(wire_d68_98),.data_out(d_out68),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance70690(.data_in(d_in69),.data_out(wire_d69_0),.clk(clk),.rst(rst));            //channel 70
	register #(.WIDTH(WIDTH)) register_instance70691(.data_in(wire_d69_0),.data_out(wire_d69_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance70692(.data_in(wire_d69_1),.data_out(wire_d69_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance70693(.data_in(wire_d69_2),.data_out(wire_d69_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance70694(.data_in(wire_d69_3),.data_out(wire_d69_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance70695(.data_in(wire_d69_4),.data_out(wire_d69_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance70696(.data_in(wire_d69_5),.data_out(wire_d69_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance70697(.data_in(wire_d69_6),.data_out(wire_d69_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance70698(.data_in(wire_d69_7),.data_out(wire_d69_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance70699(.data_in(wire_d69_8),.data_out(wire_d69_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706910(.data_in(wire_d69_9),.data_out(wire_d69_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance706911(.data_in(wire_d69_10),.data_out(wire_d69_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706912(.data_in(wire_d69_11),.data_out(wire_d69_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706913(.data_in(wire_d69_12),.data_out(wire_d69_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance706914(.data_in(wire_d69_13),.data_out(wire_d69_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706915(.data_in(wire_d69_14),.data_out(wire_d69_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706916(.data_in(wire_d69_15),.data_out(wire_d69_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706917(.data_in(wire_d69_16),.data_out(wire_d69_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance706918(.data_in(wire_d69_17),.data_out(wire_d69_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance706919(.data_in(wire_d69_18),.data_out(wire_d69_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance706920(.data_in(wire_d69_19),.data_out(wire_d69_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance706921(.data_in(wire_d69_20),.data_out(wire_d69_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance706922(.data_in(wire_d69_21),.data_out(wire_d69_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance706923(.data_in(wire_d69_22),.data_out(wire_d69_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706924(.data_in(wire_d69_23),.data_out(wire_d69_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance706925(.data_in(wire_d69_24),.data_out(wire_d69_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance706926(.data_in(wire_d69_25),.data_out(wire_d69_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706927(.data_in(wire_d69_26),.data_out(wire_d69_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706928(.data_in(wire_d69_27),.data_out(wire_d69_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance706929(.data_in(wire_d69_28),.data_out(wire_d69_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706930(.data_in(wire_d69_29),.data_out(wire_d69_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706931(.data_in(wire_d69_30),.data_out(wire_d69_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706932(.data_in(wire_d69_31),.data_out(wire_d69_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance706933(.data_in(wire_d69_32),.data_out(wire_d69_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance706934(.data_in(wire_d69_33),.data_out(wire_d69_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance706935(.data_in(wire_d69_34),.data_out(wire_d69_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706936(.data_in(wire_d69_35),.data_out(wire_d69_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706937(.data_in(wire_d69_36),.data_out(wire_d69_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance706938(.data_in(wire_d69_37),.data_out(wire_d69_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance706939(.data_in(wire_d69_38),.data_out(wire_d69_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance706940(.data_in(wire_d69_39),.data_out(wire_d69_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706941(.data_in(wire_d69_40),.data_out(wire_d69_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706942(.data_in(wire_d69_41),.data_out(wire_d69_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706943(.data_in(wire_d69_42),.data_out(wire_d69_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706944(.data_in(wire_d69_43),.data_out(wire_d69_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance706945(.data_in(wire_d69_44),.data_out(wire_d69_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance706946(.data_in(wire_d69_45),.data_out(wire_d69_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706947(.data_in(wire_d69_46),.data_out(wire_d69_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706948(.data_in(wire_d69_47),.data_out(wire_d69_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance706949(.data_in(wire_d69_48),.data_out(wire_d69_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance706950(.data_in(wire_d69_49),.data_out(wire_d69_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706951(.data_in(wire_d69_50),.data_out(wire_d69_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706952(.data_in(wire_d69_51),.data_out(wire_d69_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance706953(.data_in(wire_d69_52),.data_out(wire_d69_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706954(.data_in(wire_d69_53),.data_out(wire_d69_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706955(.data_in(wire_d69_54),.data_out(wire_d69_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706956(.data_in(wire_d69_55),.data_out(wire_d69_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706957(.data_in(wire_d69_56),.data_out(wire_d69_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706958(.data_in(wire_d69_57),.data_out(wire_d69_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance706959(.data_in(wire_d69_58),.data_out(wire_d69_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706960(.data_in(wire_d69_59),.data_out(wire_d69_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance706961(.data_in(wire_d69_60),.data_out(wire_d69_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706962(.data_in(wire_d69_61),.data_out(wire_d69_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance706963(.data_in(wire_d69_62),.data_out(wire_d69_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706964(.data_in(wire_d69_63),.data_out(wire_d69_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance706965(.data_in(wire_d69_64),.data_out(wire_d69_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance706966(.data_in(wire_d69_65),.data_out(wire_d69_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706967(.data_in(wire_d69_66),.data_out(wire_d69_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance706968(.data_in(wire_d69_67),.data_out(wire_d69_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706969(.data_in(wire_d69_68),.data_out(wire_d69_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance706970(.data_in(wire_d69_69),.data_out(wire_d69_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance706971(.data_in(wire_d69_70),.data_out(wire_d69_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706972(.data_in(wire_d69_71),.data_out(wire_d69_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance706973(.data_in(wire_d69_72),.data_out(wire_d69_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance706974(.data_in(wire_d69_73),.data_out(wire_d69_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance706975(.data_in(wire_d69_74),.data_out(wire_d69_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706976(.data_in(wire_d69_75),.data_out(wire_d69_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706977(.data_in(wire_d69_76),.data_out(wire_d69_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance706978(.data_in(wire_d69_77),.data_out(wire_d69_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706979(.data_in(wire_d69_78),.data_out(wire_d69_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706980(.data_in(wire_d69_79),.data_out(wire_d69_80),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706981(.data_in(wire_d69_80),.data_out(wire_d69_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706982(.data_in(wire_d69_81),.data_out(wire_d69_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance706983(.data_in(wire_d69_82),.data_out(wire_d69_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance706984(.data_in(wire_d69_83),.data_out(wire_d69_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance706985(.data_in(wire_d69_84),.data_out(wire_d69_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706986(.data_in(wire_d69_85),.data_out(wire_d69_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance706987(.data_in(wire_d69_86),.data_out(wire_d69_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706988(.data_in(wire_d69_87),.data_out(wire_d69_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance706989(.data_in(wire_d69_88),.data_out(wire_d69_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance706990(.data_in(wire_d69_89),.data_out(wire_d69_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706991(.data_in(wire_d69_90),.data_out(wire_d69_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706992(.data_in(wire_d69_91),.data_out(wire_d69_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance706993(.data_in(wire_d69_92),.data_out(wire_d69_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance706994(.data_in(wire_d69_93),.data_out(wire_d69_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706995(.data_in(wire_d69_94),.data_out(wire_d69_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance706996(.data_in(wire_d69_95),.data_out(wire_d69_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706997(.data_in(wire_d69_96),.data_out(wire_d69_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance706998(.data_in(wire_d69_97),.data_out(wire_d69_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance706999(.data_in(wire_d69_98),.data_out(d_out69),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance71700(.data_in(d_in70),.data_out(wire_d70_0),.clk(clk),.rst(rst));            //channel 71
	large_mux #(.WIDTH(WIDTH)) large_mux_instance71701(.data_in(wire_d70_0),.data_out(wire_d70_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance71702(.data_in(wire_d70_1),.data_out(wire_d70_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance71703(.data_in(wire_d70_2),.data_out(wire_d70_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance71704(.data_in(wire_d70_3),.data_out(wire_d70_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance71705(.data_in(wire_d70_4),.data_out(wire_d70_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance71706(.data_in(wire_d70_5),.data_out(wire_d70_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance71707(.data_in(wire_d70_6),.data_out(wire_d70_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance71708(.data_in(wire_d70_7),.data_out(wire_d70_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance71709(.data_in(wire_d70_8),.data_out(wire_d70_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance717010(.data_in(wire_d70_9),.data_out(wire_d70_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717011(.data_in(wire_d70_10),.data_out(wire_d70_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717012(.data_in(wire_d70_11),.data_out(wire_d70_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717013(.data_in(wire_d70_12),.data_out(wire_d70_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717014(.data_in(wire_d70_13),.data_out(wire_d70_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance717015(.data_in(wire_d70_14),.data_out(wire_d70_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance717016(.data_in(wire_d70_15),.data_out(wire_d70_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717017(.data_in(wire_d70_16),.data_out(wire_d70_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance717018(.data_in(wire_d70_17),.data_out(wire_d70_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717019(.data_in(wire_d70_18),.data_out(wire_d70_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance717020(.data_in(wire_d70_19),.data_out(wire_d70_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717021(.data_in(wire_d70_20),.data_out(wire_d70_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717022(.data_in(wire_d70_21),.data_out(wire_d70_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717023(.data_in(wire_d70_22),.data_out(wire_d70_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717024(.data_in(wire_d70_23),.data_out(wire_d70_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717025(.data_in(wire_d70_24),.data_out(wire_d70_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717026(.data_in(wire_d70_25),.data_out(wire_d70_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance717027(.data_in(wire_d70_26),.data_out(wire_d70_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717028(.data_in(wire_d70_27),.data_out(wire_d70_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717029(.data_in(wire_d70_28),.data_out(wire_d70_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717030(.data_in(wire_d70_29),.data_out(wire_d70_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717031(.data_in(wire_d70_30),.data_out(wire_d70_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717032(.data_in(wire_d70_31),.data_out(wire_d70_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717033(.data_in(wire_d70_32),.data_out(wire_d70_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717034(.data_in(wire_d70_33),.data_out(wire_d70_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717035(.data_in(wire_d70_34),.data_out(wire_d70_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717036(.data_in(wire_d70_35),.data_out(wire_d70_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717037(.data_in(wire_d70_36),.data_out(wire_d70_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717038(.data_in(wire_d70_37),.data_out(wire_d70_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717039(.data_in(wire_d70_38),.data_out(wire_d70_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717040(.data_in(wire_d70_39),.data_out(wire_d70_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717041(.data_in(wire_d70_40),.data_out(wire_d70_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717042(.data_in(wire_d70_41),.data_out(wire_d70_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717043(.data_in(wire_d70_42),.data_out(wire_d70_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance717044(.data_in(wire_d70_43),.data_out(wire_d70_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717045(.data_in(wire_d70_44),.data_out(wire_d70_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717046(.data_in(wire_d70_45),.data_out(wire_d70_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance717047(.data_in(wire_d70_46),.data_out(wire_d70_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717048(.data_in(wire_d70_47),.data_out(wire_d70_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717049(.data_in(wire_d70_48),.data_out(wire_d70_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717050(.data_in(wire_d70_49),.data_out(wire_d70_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717051(.data_in(wire_d70_50),.data_out(wire_d70_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717052(.data_in(wire_d70_51),.data_out(wire_d70_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance717053(.data_in(wire_d70_52),.data_out(wire_d70_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717054(.data_in(wire_d70_53),.data_out(wire_d70_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance717055(.data_in(wire_d70_54),.data_out(wire_d70_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717056(.data_in(wire_d70_55),.data_out(wire_d70_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717057(.data_in(wire_d70_56),.data_out(wire_d70_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717058(.data_in(wire_d70_57),.data_out(wire_d70_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717059(.data_in(wire_d70_58),.data_out(wire_d70_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance717060(.data_in(wire_d70_59),.data_out(wire_d70_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717061(.data_in(wire_d70_60),.data_out(wire_d70_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717062(.data_in(wire_d70_61),.data_out(wire_d70_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717063(.data_in(wire_d70_62),.data_out(wire_d70_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717064(.data_in(wire_d70_63),.data_out(wire_d70_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717065(.data_in(wire_d70_64),.data_out(wire_d70_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance717066(.data_in(wire_d70_65),.data_out(wire_d70_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717067(.data_in(wire_d70_66),.data_out(wire_d70_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717068(.data_in(wire_d70_67),.data_out(wire_d70_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717069(.data_in(wire_d70_68),.data_out(wire_d70_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717070(.data_in(wire_d70_69),.data_out(wire_d70_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance717071(.data_in(wire_d70_70),.data_out(wire_d70_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717072(.data_in(wire_d70_71),.data_out(wire_d70_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717073(.data_in(wire_d70_72),.data_out(wire_d70_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717074(.data_in(wire_d70_73),.data_out(wire_d70_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance717075(.data_in(wire_d70_74),.data_out(wire_d70_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance717076(.data_in(wire_d70_75),.data_out(wire_d70_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717077(.data_in(wire_d70_76),.data_out(wire_d70_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717078(.data_in(wire_d70_77),.data_out(wire_d70_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717079(.data_in(wire_d70_78),.data_out(wire_d70_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717080(.data_in(wire_d70_79),.data_out(wire_d70_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717081(.data_in(wire_d70_80),.data_out(wire_d70_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance717082(.data_in(wire_d70_81),.data_out(wire_d70_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance717083(.data_in(wire_d70_82),.data_out(wire_d70_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance717084(.data_in(wire_d70_83),.data_out(wire_d70_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717085(.data_in(wire_d70_84),.data_out(wire_d70_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717086(.data_in(wire_d70_85),.data_out(wire_d70_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717087(.data_in(wire_d70_86),.data_out(wire_d70_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717088(.data_in(wire_d70_87),.data_out(wire_d70_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717089(.data_in(wire_d70_88),.data_out(wire_d70_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717090(.data_in(wire_d70_89),.data_out(wire_d70_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717091(.data_in(wire_d70_90),.data_out(wire_d70_91),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance717092(.data_in(wire_d70_91),.data_out(wire_d70_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance717093(.data_in(wire_d70_92),.data_out(wire_d70_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717094(.data_in(wire_d70_93),.data_out(wire_d70_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717095(.data_in(wire_d70_94),.data_out(wire_d70_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717096(.data_in(wire_d70_95),.data_out(wire_d70_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717097(.data_in(wire_d70_96),.data_out(wire_d70_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance717098(.data_in(wire_d70_97),.data_out(wire_d70_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance717099(.data_in(wire_d70_98),.data_out(d_out70),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance72710(.data_in(d_in71),.data_out(wire_d71_0),.clk(clk),.rst(rst));            //channel 72
	encoder #(.WIDTH(WIDTH)) encoder_instance72711(.data_in(wire_d71_0),.data_out(wire_d71_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance72712(.data_in(wire_d71_1),.data_out(wire_d71_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance72713(.data_in(wire_d71_2),.data_out(wire_d71_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance72714(.data_in(wire_d71_3),.data_out(wire_d71_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance72715(.data_in(wire_d71_4),.data_out(wire_d71_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance72716(.data_in(wire_d71_5),.data_out(wire_d71_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance72717(.data_in(wire_d71_6),.data_out(wire_d71_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance72718(.data_in(wire_d71_7),.data_out(wire_d71_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance72719(.data_in(wire_d71_8),.data_out(wire_d71_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727110(.data_in(wire_d71_9),.data_out(wire_d71_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance727111(.data_in(wire_d71_10),.data_out(wire_d71_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance727112(.data_in(wire_d71_11),.data_out(wire_d71_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727113(.data_in(wire_d71_12),.data_out(wire_d71_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727114(.data_in(wire_d71_13),.data_out(wire_d71_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727115(.data_in(wire_d71_14),.data_out(wire_d71_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727116(.data_in(wire_d71_15),.data_out(wire_d71_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727117(.data_in(wire_d71_16),.data_out(wire_d71_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727118(.data_in(wire_d71_17),.data_out(wire_d71_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727119(.data_in(wire_d71_18),.data_out(wire_d71_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727120(.data_in(wire_d71_19),.data_out(wire_d71_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727121(.data_in(wire_d71_20),.data_out(wire_d71_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727122(.data_in(wire_d71_21),.data_out(wire_d71_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727123(.data_in(wire_d71_22),.data_out(wire_d71_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727124(.data_in(wire_d71_23),.data_out(wire_d71_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance727125(.data_in(wire_d71_24),.data_out(wire_d71_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance727126(.data_in(wire_d71_25),.data_out(wire_d71_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727127(.data_in(wire_d71_26),.data_out(wire_d71_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727128(.data_in(wire_d71_27),.data_out(wire_d71_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727129(.data_in(wire_d71_28),.data_out(wire_d71_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727130(.data_in(wire_d71_29),.data_out(wire_d71_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727131(.data_in(wire_d71_30),.data_out(wire_d71_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727132(.data_in(wire_d71_31),.data_out(wire_d71_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727133(.data_in(wire_d71_32),.data_out(wire_d71_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance727134(.data_in(wire_d71_33),.data_out(wire_d71_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance727135(.data_in(wire_d71_34),.data_out(wire_d71_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727136(.data_in(wire_d71_35),.data_out(wire_d71_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance727137(.data_in(wire_d71_36),.data_out(wire_d71_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance727138(.data_in(wire_d71_37),.data_out(wire_d71_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727139(.data_in(wire_d71_38),.data_out(wire_d71_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance727140(.data_in(wire_d71_39),.data_out(wire_d71_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727141(.data_in(wire_d71_40),.data_out(wire_d71_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727142(.data_in(wire_d71_41),.data_out(wire_d71_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727143(.data_in(wire_d71_42),.data_out(wire_d71_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727144(.data_in(wire_d71_43),.data_out(wire_d71_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727145(.data_in(wire_d71_44),.data_out(wire_d71_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance727146(.data_in(wire_d71_45),.data_out(wire_d71_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance727147(.data_in(wire_d71_46),.data_out(wire_d71_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance727148(.data_in(wire_d71_47),.data_out(wire_d71_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727149(.data_in(wire_d71_48),.data_out(wire_d71_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727150(.data_in(wire_d71_49),.data_out(wire_d71_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727151(.data_in(wire_d71_50),.data_out(wire_d71_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727152(.data_in(wire_d71_51),.data_out(wire_d71_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance727153(.data_in(wire_d71_52),.data_out(wire_d71_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727154(.data_in(wire_d71_53),.data_out(wire_d71_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727155(.data_in(wire_d71_54),.data_out(wire_d71_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727156(.data_in(wire_d71_55),.data_out(wire_d71_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727157(.data_in(wire_d71_56),.data_out(wire_d71_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727158(.data_in(wire_d71_57),.data_out(wire_d71_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727159(.data_in(wire_d71_58),.data_out(wire_d71_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727160(.data_in(wire_d71_59),.data_out(wire_d71_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727161(.data_in(wire_d71_60),.data_out(wire_d71_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727162(.data_in(wire_d71_61),.data_out(wire_d71_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727163(.data_in(wire_d71_62),.data_out(wire_d71_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727164(.data_in(wire_d71_63),.data_out(wire_d71_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727165(.data_in(wire_d71_64),.data_out(wire_d71_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727166(.data_in(wire_d71_65),.data_out(wire_d71_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727167(.data_in(wire_d71_66),.data_out(wire_d71_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727168(.data_in(wire_d71_67),.data_out(wire_d71_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727169(.data_in(wire_d71_68),.data_out(wire_d71_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727170(.data_in(wire_d71_69),.data_out(wire_d71_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727171(.data_in(wire_d71_70),.data_out(wire_d71_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727172(.data_in(wire_d71_71),.data_out(wire_d71_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance727173(.data_in(wire_d71_72),.data_out(wire_d71_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727174(.data_in(wire_d71_73),.data_out(wire_d71_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727175(.data_in(wire_d71_74),.data_out(wire_d71_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727176(.data_in(wire_d71_75),.data_out(wire_d71_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727177(.data_in(wire_d71_76),.data_out(wire_d71_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727178(.data_in(wire_d71_77),.data_out(wire_d71_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727179(.data_in(wire_d71_78),.data_out(wire_d71_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727180(.data_in(wire_d71_79),.data_out(wire_d71_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance727181(.data_in(wire_d71_80),.data_out(wire_d71_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance727182(.data_in(wire_d71_81),.data_out(wire_d71_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727183(.data_in(wire_d71_82),.data_out(wire_d71_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727184(.data_in(wire_d71_83),.data_out(wire_d71_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727185(.data_in(wire_d71_84),.data_out(wire_d71_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727186(.data_in(wire_d71_85),.data_out(wire_d71_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727187(.data_in(wire_d71_86),.data_out(wire_d71_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727188(.data_in(wire_d71_87),.data_out(wire_d71_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance727189(.data_in(wire_d71_88),.data_out(wire_d71_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727190(.data_in(wire_d71_89),.data_out(wire_d71_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance727191(.data_in(wire_d71_90),.data_out(wire_d71_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727192(.data_in(wire_d71_91),.data_out(wire_d71_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727193(.data_in(wire_d71_92),.data_out(wire_d71_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727194(.data_in(wire_d71_93),.data_out(wire_d71_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance727195(.data_in(wire_d71_94),.data_out(wire_d71_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727196(.data_in(wire_d71_95),.data_out(wire_d71_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance727197(.data_in(wire_d71_96),.data_out(wire_d71_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance727198(.data_in(wire_d71_97),.data_out(wire_d71_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance727199(.data_in(wire_d71_98),.data_out(d_out71),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance73720(.data_in(d_in72),.data_out(wire_d72_0),.clk(clk),.rst(rst));            //channel 73
	register #(.WIDTH(WIDTH)) register_instance73721(.data_in(wire_d72_0),.data_out(wire_d72_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance73722(.data_in(wire_d72_1),.data_out(wire_d72_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance73723(.data_in(wire_d72_2),.data_out(wire_d72_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance73724(.data_in(wire_d72_3),.data_out(wire_d72_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance73725(.data_in(wire_d72_4),.data_out(wire_d72_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance73726(.data_in(wire_d72_5),.data_out(wire_d72_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance73727(.data_in(wire_d72_6),.data_out(wire_d72_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance73728(.data_in(wire_d72_7),.data_out(wire_d72_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance73729(.data_in(wire_d72_8),.data_out(wire_d72_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance737210(.data_in(wire_d72_9),.data_out(wire_d72_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737211(.data_in(wire_d72_10),.data_out(wire_d72_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737212(.data_in(wire_d72_11),.data_out(wire_d72_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737213(.data_in(wire_d72_12),.data_out(wire_d72_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737214(.data_in(wire_d72_13),.data_out(wire_d72_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737215(.data_in(wire_d72_14),.data_out(wire_d72_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737216(.data_in(wire_d72_15),.data_out(wire_d72_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737217(.data_in(wire_d72_16),.data_out(wire_d72_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance737218(.data_in(wire_d72_17),.data_out(wire_d72_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737219(.data_in(wire_d72_18),.data_out(wire_d72_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737220(.data_in(wire_d72_19),.data_out(wire_d72_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance737221(.data_in(wire_d72_20),.data_out(wire_d72_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance737222(.data_in(wire_d72_21),.data_out(wire_d72_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737223(.data_in(wire_d72_22),.data_out(wire_d72_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737224(.data_in(wire_d72_23),.data_out(wire_d72_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance737225(.data_in(wire_d72_24),.data_out(wire_d72_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737226(.data_in(wire_d72_25),.data_out(wire_d72_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737227(.data_in(wire_d72_26),.data_out(wire_d72_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737228(.data_in(wire_d72_27),.data_out(wire_d72_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance737229(.data_in(wire_d72_28),.data_out(wire_d72_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance737230(.data_in(wire_d72_29),.data_out(wire_d72_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737231(.data_in(wire_d72_30),.data_out(wire_d72_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance737232(.data_in(wire_d72_31),.data_out(wire_d72_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737233(.data_in(wire_d72_32),.data_out(wire_d72_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance737234(.data_in(wire_d72_33),.data_out(wire_d72_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance737235(.data_in(wire_d72_34),.data_out(wire_d72_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance737236(.data_in(wire_d72_35),.data_out(wire_d72_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance737237(.data_in(wire_d72_36),.data_out(wire_d72_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737238(.data_in(wire_d72_37),.data_out(wire_d72_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737239(.data_in(wire_d72_38),.data_out(wire_d72_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737240(.data_in(wire_d72_39),.data_out(wire_d72_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737241(.data_in(wire_d72_40),.data_out(wire_d72_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737242(.data_in(wire_d72_41),.data_out(wire_d72_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance737243(.data_in(wire_d72_42),.data_out(wire_d72_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance737244(.data_in(wire_d72_43),.data_out(wire_d72_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737245(.data_in(wire_d72_44),.data_out(wire_d72_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance737246(.data_in(wire_d72_45),.data_out(wire_d72_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737247(.data_in(wire_d72_46),.data_out(wire_d72_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance737248(.data_in(wire_d72_47),.data_out(wire_d72_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737249(.data_in(wire_d72_48),.data_out(wire_d72_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance737250(.data_in(wire_d72_49),.data_out(wire_d72_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737251(.data_in(wire_d72_50),.data_out(wire_d72_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737252(.data_in(wire_d72_51),.data_out(wire_d72_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance737253(.data_in(wire_d72_52),.data_out(wire_d72_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance737254(.data_in(wire_d72_53),.data_out(wire_d72_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737255(.data_in(wire_d72_54),.data_out(wire_d72_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance737256(.data_in(wire_d72_55),.data_out(wire_d72_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance737257(.data_in(wire_d72_56),.data_out(wire_d72_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737258(.data_in(wire_d72_57),.data_out(wire_d72_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737259(.data_in(wire_d72_58),.data_out(wire_d72_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance737260(.data_in(wire_d72_59),.data_out(wire_d72_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance737261(.data_in(wire_d72_60),.data_out(wire_d72_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737262(.data_in(wire_d72_61),.data_out(wire_d72_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737263(.data_in(wire_d72_62),.data_out(wire_d72_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance737264(.data_in(wire_d72_63),.data_out(wire_d72_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance737265(.data_in(wire_d72_64),.data_out(wire_d72_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance737266(.data_in(wire_d72_65),.data_out(wire_d72_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance737267(.data_in(wire_d72_66),.data_out(wire_d72_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737268(.data_in(wire_d72_67),.data_out(wire_d72_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737269(.data_in(wire_d72_68),.data_out(wire_d72_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737270(.data_in(wire_d72_69),.data_out(wire_d72_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737271(.data_in(wire_d72_70),.data_out(wire_d72_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737272(.data_in(wire_d72_71),.data_out(wire_d72_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance737273(.data_in(wire_d72_72),.data_out(wire_d72_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance737274(.data_in(wire_d72_73),.data_out(wire_d72_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance737275(.data_in(wire_d72_74),.data_out(wire_d72_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737276(.data_in(wire_d72_75),.data_out(wire_d72_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737277(.data_in(wire_d72_76),.data_out(wire_d72_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance737278(.data_in(wire_d72_77),.data_out(wire_d72_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance737279(.data_in(wire_d72_78),.data_out(wire_d72_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance737280(.data_in(wire_d72_79),.data_out(wire_d72_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance737281(.data_in(wire_d72_80),.data_out(wire_d72_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance737282(.data_in(wire_d72_81),.data_out(wire_d72_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737283(.data_in(wire_d72_82),.data_out(wire_d72_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737284(.data_in(wire_d72_83),.data_out(wire_d72_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737285(.data_in(wire_d72_84),.data_out(wire_d72_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance737286(.data_in(wire_d72_85),.data_out(wire_d72_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737287(.data_in(wire_d72_86),.data_out(wire_d72_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance737288(.data_in(wire_d72_87),.data_out(wire_d72_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737289(.data_in(wire_d72_88),.data_out(wire_d72_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance737290(.data_in(wire_d72_89),.data_out(wire_d72_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737291(.data_in(wire_d72_90),.data_out(wire_d72_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance737292(.data_in(wire_d72_91),.data_out(wire_d72_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance737293(.data_in(wire_d72_92),.data_out(wire_d72_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737294(.data_in(wire_d72_93),.data_out(wire_d72_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance737295(.data_in(wire_d72_94),.data_out(wire_d72_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance737296(.data_in(wire_d72_95),.data_out(wire_d72_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance737297(.data_in(wire_d72_96),.data_out(wire_d72_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance737298(.data_in(wire_d72_97),.data_out(wire_d72_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance737299(.data_in(wire_d72_98),.data_out(d_out72),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance74730(.data_in(d_in73),.data_out(wire_d73_0),.clk(clk),.rst(rst));            //channel 74
	register #(.WIDTH(WIDTH)) register_instance74731(.data_in(wire_d73_0),.data_out(wire_d73_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance74732(.data_in(wire_d73_1),.data_out(wire_d73_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance74733(.data_in(wire_d73_2),.data_out(wire_d73_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance74734(.data_in(wire_d73_3),.data_out(wire_d73_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance74735(.data_in(wire_d73_4),.data_out(wire_d73_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance74736(.data_in(wire_d73_5),.data_out(wire_d73_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance74737(.data_in(wire_d73_6),.data_out(wire_d73_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance74738(.data_in(wire_d73_7),.data_out(wire_d73_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance74739(.data_in(wire_d73_8),.data_out(wire_d73_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747310(.data_in(wire_d73_9),.data_out(wire_d73_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance747311(.data_in(wire_d73_10),.data_out(wire_d73_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747312(.data_in(wire_d73_11),.data_out(wire_d73_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance747313(.data_in(wire_d73_12),.data_out(wire_d73_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747314(.data_in(wire_d73_13),.data_out(wire_d73_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance747315(.data_in(wire_d73_14),.data_out(wire_d73_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747316(.data_in(wire_d73_15),.data_out(wire_d73_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance747317(.data_in(wire_d73_16),.data_out(wire_d73_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance747318(.data_in(wire_d73_17),.data_out(wire_d73_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance747319(.data_in(wire_d73_18),.data_out(wire_d73_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747320(.data_in(wire_d73_19),.data_out(wire_d73_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance747321(.data_in(wire_d73_20),.data_out(wire_d73_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance747322(.data_in(wire_d73_21),.data_out(wire_d73_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance747323(.data_in(wire_d73_22),.data_out(wire_d73_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance747324(.data_in(wire_d73_23),.data_out(wire_d73_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747325(.data_in(wire_d73_24),.data_out(wire_d73_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747326(.data_in(wire_d73_25),.data_out(wire_d73_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance747327(.data_in(wire_d73_26),.data_out(wire_d73_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747328(.data_in(wire_d73_27),.data_out(wire_d73_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747329(.data_in(wire_d73_28),.data_out(wire_d73_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747330(.data_in(wire_d73_29),.data_out(wire_d73_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance747331(.data_in(wire_d73_30),.data_out(wire_d73_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747332(.data_in(wire_d73_31),.data_out(wire_d73_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747333(.data_in(wire_d73_32),.data_out(wire_d73_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance747334(.data_in(wire_d73_33),.data_out(wire_d73_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747335(.data_in(wire_d73_34),.data_out(wire_d73_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance747336(.data_in(wire_d73_35),.data_out(wire_d73_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance747337(.data_in(wire_d73_36),.data_out(wire_d73_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747338(.data_in(wire_d73_37),.data_out(wire_d73_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747339(.data_in(wire_d73_38),.data_out(wire_d73_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747340(.data_in(wire_d73_39),.data_out(wire_d73_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747341(.data_in(wire_d73_40),.data_out(wire_d73_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance747342(.data_in(wire_d73_41),.data_out(wire_d73_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance747343(.data_in(wire_d73_42),.data_out(wire_d73_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance747344(.data_in(wire_d73_43),.data_out(wire_d73_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747345(.data_in(wire_d73_44),.data_out(wire_d73_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance747346(.data_in(wire_d73_45),.data_out(wire_d73_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance747347(.data_in(wire_d73_46),.data_out(wire_d73_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747348(.data_in(wire_d73_47),.data_out(wire_d73_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747349(.data_in(wire_d73_48),.data_out(wire_d73_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747350(.data_in(wire_d73_49),.data_out(wire_d73_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747351(.data_in(wire_d73_50),.data_out(wire_d73_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance747352(.data_in(wire_d73_51),.data_out(wire_d73_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance747353(.data_in(wire_d73_52),.data_out(wire_d73_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747354(.data_in(wire_d73_53),.data_out(wire_d73_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747355(.data_in(wire_d73_54),.data_out(wire_d73_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance747356(.data_in(wire_d73_55),.data_out(wire_d73_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance747357(.data_in(wire_d73_56),.data_out(wire_d73_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747358(.data_in(wire_d73_57),.data_out(wire_d73_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747359(.data_in(wire_d73_58),.data_out(wire_d73_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance747360(.data_in(wire_d73_59),.data_out(wire_d73_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747361(.data_in(wire_d73_60),.data_out(wire_d73_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747362(.data_in(wire_d73_61),.data_out(wire_d73_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747363(.data_in(wire_d73_62),.data_out(wire_d73_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747364(.data_in(wire_d73_63),.data_out(wire_d73_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747365(.data_in(wire_d73_64),.data_out(wire_d73_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance747366(.data_in(wire_d73_65),.data_out(wire_d73_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance747367(.data_in(wire_d73_66),.data_out(wire_d73_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747368(.data_in(wire_d73_67),.data_out(wire_d73_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance747369(.data_in(wire_d73_68),.data_out(wire_d73_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747370(.data_in(wire_d73_69),.data_out(wire_d73_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747371(.data_in(wire_d73_70),.data_out(wire_d73_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747372(.data_in(wire_d73_71),.data_out(wire_d73_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747373(.data_in(wire_d73_72),.data_out(wire_d73_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance747374(.data_in(wire_d73_73),.data_out(wire_d73_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance747375(.data_in(wire_d73_74),.data_out(wire_d73_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747376(.data_in(wire_d73_75),.data_out(wire_d73_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747377(.data_in(wire_d73_76),.data_out(wire_d73_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance747378(.data_in(wire_d73_77),.data_out(wire_d73_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747379(.data_in(wire_d73_78),.data_out(wire_d73_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance747380(.data_in(wire_d73_79),.data_out(wire_d73_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance747381(.data_in(wire_d73_80),.data_out(wire_d73_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance747382(.data_in(wire_d73_81),.data_out(wire_d73_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747383(.data_in(wire_d73_82),.data_out(wire_d73_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance747384(.data_in(wire_d73_83),.data_out(wire_d73_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance747385(.data_in(wire_d73_84),.data_out(wire_d73_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747386(.data_in(wire_d73_85),.data_out(wire_d73_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance747387(.data_in(wire_d73_86),.data_out(wire_d73_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747388(.data_in(wire_d73_87),.data_out(wire_d73_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance747389(.data_in(wire_d73_88),.data_out(wire_d73_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747390(.data_in(wire_d73_89),.data_out(wire_d73_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747391(.data_in(wire_d73_90),.data_out(wire_d73_91),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747392(.data_in(wire_d73_91),.data_out(wire_d73_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747393(.data_in(wire_d73_92),.data_out(wire_d73_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance747394(.data_in(wire_d73_93),.data_out(wire_d73_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance747395(.data_in(wire_d73_94),.data_out(wire_d73_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance747396(.data_in(wire_d73_95),.data_out(wire_d73_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance747397(.data_in(wire_d73_96),.data_out(wire_d73_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance747398(.data_in(wire_d73_97),.data_out(wire_d73_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance747399(.data_in(wire_d73_98),.data_out(d_out73),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance75740(.data_in(d_in74),.data_out(wire_d74_0),.clk(clk),.rst(rst));            //channel 75
	register #(.WIDTH(WIDTH)) register_instance75741(.data_in(wire_d74_0),.data_out(wire_d74_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance75742(.data_in(wire_d74_1),.data_out(wire_d74_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance75743(.data_in(wire_d74_2),.data_out(wire_d74_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance75744(.data_in(wire_d74_3),.data_out(wire_d74_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance75745(.data_in(wire_d74_4),.data_out(wire_d74_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance75746(.data_in(wire_d74_5),.data_out(wire_d74_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance75747(.data_in(wire_d74_6),.data_out(wire_d74_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance75748(.data_in(wire_d74_7),.data_out(wire_d74_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance75749(.data_in(wire_d74_8),.data_out(wire_d74_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757410(.data_in(wire_d74_9),.data_out(wire_d74_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757411(.data_in(wire_d74_10),.data_out(wire_d74_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757412(.data_in(wire_d74_11),.data_out(wire_d74_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757413(.data_in(wire_d74_12),.data_out(wire_d74_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757414(.data_in(wire_d74_13),.data_out(wire_d74_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757415(.data_in(wire_d74_14),.data_out(wire_d74_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance757416(.data_in(wire_d74_15),.data_out(wire_d74_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757417(.data_in(wire_d74_16),.data_out(wire_d74_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757418(.data_in(wire_d74_17),.data_out(wire_d74_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance757419(.data_in(wire_d74_18),.data_out(wire_d74_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757420(.data_in(wire_d74_19),.data_out(wire_d74_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance757421(.data_in(wire_d74_20),.data_out(wire_d74_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757422(.data_in(wire_d74_21),.data_out(wire_d74_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757423(.data_in(wire_d74_22),.data_out(wire_d74_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757424(.data_in(wire_d74_23),.data_out(wire_d74_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757425(.data_in(wire_d74_24),.data_out(wire_d74_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757426(.data_in(wire_d74_25),.data_out(wire_d74_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757427(.data_in(wire_d74_26),.data_out(wire_d74_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757428(.data_in(wire_d74_27),.data_out(wire_d74_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757429(.data_in(wire_d74_28),.data_out(wire_d74_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757430(.data_in(wire_d74_29),.data_out(wire_d74_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757431(.data_in(wire_d74_30),.data_out(wire_d74_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757432(.data_in(wire_d74_31),.data_out(wire_d74_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757433(.data_in(wire_d74_32),.data_out(wire_d74_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757434(.data_in(wire_d74_33),.data_out(wire_d74_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance757435(.data_in(wire_d74_34),.data_out(wire_d74_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757436(.data_in(wire_d74_35),.data_out(wire_d74_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757437(.data_in(wire_d74_36),.data_out(wire_d74_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757438(.data_in(wire_d74_37),.data_out(wire_d74_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757439(.data_in(wire_d74_38),.data_out(wire_d74_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757440(.data_in(wire_d74_39),.data_out(wire_d74_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance757441(.data_in(wire_d74_40),.data_out(wire_d74_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance757442(.data_in(wire_d74_41),.data_out(wire_d74_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757443(.data_in(wire_d74_42),.data_out(wire_d74_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757444(.data_in(wire_d74_43),.data_out(wire_d74_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757445(.data_in(wire_d74_44),.data_out(wire_d74_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757446(.data_in(wire_d74_45),.data_out(wire_d74_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757447(.data_in(wire_d74_46),.data_out(wire_d74_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance757448(.data_in(wire_d74_47),.data_out(wire_d74_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757449(.data_in(wire_d74_48),.data_out(wire_d74_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance757450(.data_in(wire_d74_49),.data_out(wire_d74_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757451(.data_in(wire_d74_50),.data_out(wire_d74_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757452(.data_in(wire_d74_51),.data_out(wire_d74_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance757453(.data_in(wire_d74_52),.data_out(wire_d74_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757454(.data_in(wire_d74_53),.data_out(wire_d74_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757455(.data_in(wire_d74_54),.data_out(wire_d74_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757456(.data_in(wire_d74_55),.data_out(wire_d74_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757457(.data_in(wire_d74_56),.data_out(wire_d74_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757458(.data_in(wire_d74_57),.data_out(wire_d74_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance757459(.data_in(wire_d74_58),.data_out(wire_d74_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757460(.data_in(wire_d74_59),.data_out(wire_d74_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance757461(.data_in(wire_d74_60),.data_out(wire_d74_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757462(.data_in(wire_d74_61),.data_out(wire_d74_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757463(.data_in(wire_d74_62),.data_out(wire_d74_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757464(.data_in(wire_d74_63),.data_out(wire_d74_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757465(.data_in(wire_d74_64),.data_out(wire_d74_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance757466(.data_in(wire_d74_65),.data_out(wire_d74_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance757467(.data_in(wire_d74_66),.data_out(wire_d74_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance757468(.data_in(wire_d74_67),.data_out(wire_d74_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757469(.data_in(wire_d74_68),.data_out(wire_d74_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757470(.data_in(wire_d74_69),.data_out(wire_d74_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757471(.data_in(wire_d74_70),.data_out(wire_d74_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757472(.data_in(wire_d74_71),.data_out(wire_d74_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757473(.data_in(wire_d74_72),.data_out(wire_d74_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757474(.data_in(wire_d74_73),.data_out(wire_d74_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757475(.data_in(wire_d74_74),.data_out(wire_d74_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757476(.data_in(wire_d74_75),.data_out(wire_d74_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757477(.data_in(wire_d74_76),.data_out(wire_d74_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757478(.data_in(wire_d74_77),.data_out(wire_d74_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757479(.data_in(wire_d74_78),.data_out(wire_d74_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance757480(.data_in(wire_d74_79),.data_out(wire_d74_80),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757481(.data_in(wire_d74_80),.data_out(wire_d74_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757482(.data_in(wire_d74_81),.data_out(wire_d74_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757483(.data_in(wire_d74_82),.data_out(wire_d74_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance757484(.data_in(wire_d74_83),.data_out(wire_d74_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance757485(.data_in(wire_d74_84),.data_out(wire_d74_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757486(.data_in(wire_d74_85),.data_out(wire_d74_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance757487(.data_in(wire_d74_86),.data_out(wire_d74_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance757488(.data_in(wire_d74_87),.data_out(wire_d74_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757489(.data_in(wire_d74_88),.data_out(wire_d74_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance757490(.data_in(wire_d74_89),.data_out(wire_d74_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757491(.data_in(wire_d74_90),.data_out(wire_d74_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757492(.data_in(wire_d74_91),.data_out(wire_d74_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757493(.data_in(wire_d74_92),.data_out(wire_d74_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance757494(.data_in(wire_d74_93),.data_out(wire_d74_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757495(.data_in(wire_d74_94),.data_out(wire_d74_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance757496(.data_in(wire_d74_95),.data_out(wire_d74_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance757497(.data_in(wire_d74_96),.data_out(wire_d74_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757498(.data_in(wire_d74_97),.data_out(wire_d74_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance757499(.data_in(wire_d74_98),.data_out(d_out74),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance76750(.data_in(d_in75),.data_out(wire_d75_0),.clk(clk),.rst(rst));            //channel 76
	invertion #(.WIDTH(WIDTH)) invertion_instance76751(.data_in(wire_d75_0),.data_out(wire_d75_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance76752(.data_in(wire_d75_1),.data_out(wire_d75_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance76753(.data_in(wire_d75_2),.data_out(wire_d75_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance76754(.data_in(wire_d75_3),.data_out(wire_d75_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance76755(.data_in(wire_d75_4),.data_out(wire_d75_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance76756(.data_in(wire_d75_5),.data_out(wire_d75_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance76757(.data_in(wire_d75_6),.data_out(wire_d75_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance76758(.data_in(wire_d75_7),.data_out(wire_d75_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76759(.data_in(wire_d75_8),.data_out(wire_d75_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767510(.data_in(wire_d75_9),.data_out(wire_d75_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767511(.data_in(wire_d75_10),.data_out(wire_d75_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767512(.data_in(wire_d75_11),.data_out(wire_d75_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767513(.data_in(wire_d75_12),.data_out(wire_d75_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance767514(.data_in(wire_d75_13),.data_out(wire_d75_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance767515(.data_in(wire_d75_14),.data_out(wire_d75_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767516(.data_in(wire_d75_15),.data_out(wire_d75_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance767517(.data_in(wire_d75_16),.data_out(wire_d75_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767518(.data_in(wire_d75_17),.data_out(wire_d75_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance767519(.data_in(wire_d75_18),.data_out(wire_d75_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767520(.data_in(wire_d75_19),.data_out(wire_d75_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767521(.data_in(wire_d75_20),.data_out(wire_d75_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767522(.data_in(wire_d75_21),.data_out(wire_d75_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767523(.data_in(wire_d75_22),.data_out(wire_d75_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767524(.data_in(wire_d75_23),.data_out(wire_d75_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767525(.data_in(wire_d75_24),.data_out(wire_d75_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767526(.data_in(wire_d75_25),.data_out(wire_d75_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance767527(.data_in(wire_d75_26),.data_out(wire_d75_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance767528(.data_in(wire_d75_27),.data_out(wire_d75_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance767529(.data_in(wire_d75_28),.data_out(wire_d75_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767530(.data_in(wire_d75_29),.data_out(wire_d75_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767531(.data_in(wire_d75_30),.data_out(wire_d75_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767532(.data_in(wire_d75_31),.data_out(wire_d75_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767533(.data_in(wire_d75_32),.data_out(wire_d75_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance767534(.data_in(wire_d75_33),.data_out(wire_d75_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767535(.data_in(wire_d75_34),.data_out(wire_d75_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767536(.data_in(wire_d75_35),.data_out(wire_d75_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767537(.data_in(wire_d75_36),.data_out(wire_d75_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767538(.data_in(wire_d75_37),.data_out(wire_d75_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767539(.data_in(wire_d75_38),.data_out(wire_d75_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767540(.data_in(wire_d75_39),.data_out(wire_d75_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767541(.data_in(wire_d75_40),.data_out(wire_d75_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance767542(.data_in(wire_d75_41),.data_out(wire_d75_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767543(.data_in(wire_d75_42),.data_out(wire_d75_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767544(.data_in(wire_d75_43),.data_out(wire_d75_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767545(.data_in(wire_d75_44),.data_out(wire_d75_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance767546(.data_in(wire_d75_45),.data_out(wire_d75_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767547(.data_in(wire_d75_46),.data_out(wire_d75_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767548(.data_in(wire_d75_47),.data_out(wire_d75_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767549(.data_in(wire_d75_48),.data_out(wire_d75_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767550(.data_in(wire_d75_49),.data_out(wire_d75_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767551(.data_in(wire_d75_50),.data_out(wire_d75_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767552(.data_in(wire_d75_51),.data_out(wire_d75_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance767553(.data_in(wire_d75_52),.data_out(wire_d75_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767554(.data_in(wire_d75_53),.data_out(wire_d75_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767555(.data_in(wire_d75_54),.data_out(wire_d75_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767556(.data_in(wire_d75_55),.data_out(wire_d75_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767557(.data_in(wire_d75_56),.data_out(wire_d75_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767558(.data_in(wire_d75_57),.data_out(wire_d75_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance767559(.data_in(wire_d75_58),.data_out(wire_d75_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767560(.data_in(wire_d75_59),.data_out(wire_d75_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767561(.data_in(wire_d75_60),.data_out(wire_d75_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767562(.data_in(wire_d75_61),.data_out(wire_d75_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance767563(.data_in(wire_d75_62),.data_out(wire_d75_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767564(.data_in(wire_d75_63),.data_out(wire_d75_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance767565(.data_in(wire_d75_64),.data_out(wire_d75_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767566(.data_in(wire_d75_65),.data_out(wire_d75_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767567(.data_in(wire_d75_66),.data_out(wire_d75_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767568(.data_in(wire_d75_67),.data_out(wire_d75_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767569(.data_in(wire_d75_68),.data_out(wire_d75_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767570(.data_in(wire_d75_69),.data_out(wire_d75_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767571(.data_in(wire_d75_70),.data_out(wire_d75_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767572(.data_in(wire_d75_71),.data_out(wire_d75_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767573(.data_in(wire_d75_72),.data_out(wire_d75_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767574(.data_in(wire_d75_73),.data_out(wire_d75_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767575(.data_in(wire_d75_74),.data_out(wire_d75_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767576(.data_in(wire_d75_75),.data_out(wire_d75_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767577(.data_in(wire_d75_76),.data_out(wire_d75_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767578(.data_in(wire_d75_77),.data_out(wire_d75_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767579(.data_in(wire_d75_78),.data_out(wire_d75_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance767580(.data_in(wire_d75_79),.data_out(wire_d75_80),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance767581(.data_in(wire_d75_80),.data_out(wire_d75_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance767582(.data_in(wire_d75_81),.data_out(wire_d75_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767583(.data_in(wire_d75_82),.data_out(wire_d75_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767584(.data_in(wire_d75_83),.data_out(wire_d75_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance767585(.data_in(wire_d75_84),.data_out(wire_d75_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767586(.data_in(wire_d75_85),.data_out(wire_d75_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767587(.data_in(wire_d75_86),.data_out(wire_d75_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance767588(.data_in(wire_d75_87),.data_out(wire_d75_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767589(.data_in(wire_d75_88),.data_out(wire_d75_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767590(.data_in(wire_d75_89),.data_out(wire_d75_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance767591(.data_in(wire_d75_90),.data_out(wire_d75_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767592(.data_in(wire_d75_91),.data_out(wire_d75_92),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance767593(.data_in(wire_d75_92),.data_out(wire_d75_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767594(.data_in(wire_d75_93),.data_out(wire_d75_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767595(.data_in(wire_d75_94),.data_out(wire_d75_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767596(.data_in(wire_d75_95),.data_out(wire_d75_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance767597(.data_in(wire_d75_96),.data_out(wire_d75_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767598(.data_in(wire_d75_97),.data_out(wire_d75_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767599(.data_in(wire_d75_98),.data_out(d_out75),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance77760(.data_in(d_in76),.data_out(wire_d76_0),.clk(clk),.rst(rst));            //channel 77
	large_mux #(.WIDTH(WIDTH)) large_mux_instance77761(.data_in(wire_d76_0),.data_out(wire_d76_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance77762(.data_in(wire_d76_1),.data_out(wire_d76_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance77763(.data_in(wire_d76_2),.data_out(wire_d76_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance77764(.data_in(wire_d76_3),.data_out(wire_d76_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance77765(.data_in(wire_d76_4),.data_out(wire_d76_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance77766(.data_in(wire_d76_5),.data_out(wire_d76_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance77767(.data_in(wire_d76_6),.data_out(wire_d76_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance77768(.data_in(wire_d76_7),.data_out(wire_d76_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance77769(.data_in(wire_d76_8),.data_out(wire_d76_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777610(.data_in(wire_d76_9),.data_out(wire_d76_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777611(.data_in(wire_d76_10),.data_out(wire_d76_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777612(.data_in(wire_d76_11),.data_out(wire_d76_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance777613(.data_in(wire_d76_12),.data_out(wire_d76_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance777614(.data_in(wire_d76_13),.data_out(wire_d76_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance777615(.data_in(wire_d76_14),.data_out(wire_d76_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance777616(.data_in(wire_d76_15),.data_out(wire_d76_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777617(.data_in(wire_d76_16),.data_out(wire_d76_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777618(.data_in(wire_d76_17),.data_out(wire_d76_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777619(.data_in(wire_d76_18),.data_out(wire_d76_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777620(.data_in(wire_d76_19),.data_out(wire_d76_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777621(.data_in(wire_d76_20),.data_out(wire_d76_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777622(.data_in(wire_d76_21),.data_out(wire_d76_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance777623(.data_in(wire_d76_22),.data_out(wire_d76_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance777624(.data_in(wire_d76_23),.data_out(wire_d76_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777625(.data_in(wire_d76_24),.data_out(wire_d76_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777626(.data_in(wire_d76_25),.data_out(wire_d76_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777627(.data_in(wire_d76_26),.data_out(wire_d76_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777628(.data_in(wire_d76_27),.data_out(wire_d76_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance777629(.data_in(wire_d76_28),.data_out(wire_d76_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777630(.data_in(wire_d76_29),.data_out(wire_d76_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777631(.data_in(wire_d76_30),.data_out(wire_d76_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777632(.data_in(wire_d76_31),.data_out(wire_d76_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777633(.data_in(wire_d76_32),.data_out(wire_d76_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777634(.data_in(wire_d76_33),.data_out(wire_d76_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777635(.data_in(wire_d76_34),.data_out(wire_d76_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777636(.data_in(wire_d76_35),.data_out(wire_d76_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777637(.data_in(wire_d76_36),.data_out(wire_d76_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777638(.data_in(wire_d76_37),.data_out(wire_d76_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777639(.data_in(wire_d76_38),.data_out(wire_d76_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance777640(.data_in(wire_d76_39),.data_out(wire_d76_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777641(.data_in(wire_d76_40),.data_out(wire_d76_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance777642(.data_in(wire_d76_41),.data_out(wire_d76_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777643(.data_in(wire_d76_42),.data_out(wire_d76_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance777644(.data_in(wire_d76_43),.data_out(wire_d76_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777645(.data_in(wire_d76_44),.data_out(wire_d76_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777646(.data_in(wire_d76_45),.data_out(wire_d76_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777647(.data_in(wire_d76_46),.data_out(wire_d76_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777648(.data_in(wire_d76_47),.data_out(wire_d76_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777649(.data_in(wire_d76_48),.data_out(wire_d76_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance777650(.data_in(wire_d76_49),.data_out(wire_d76_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance777651(.data_in(wire_d76_50),.data_out(wire_d76_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777652(.data_in(wire_d76_51),.data_out(wire_d76_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777653(.data_in(wire_d76_52),.data_out(wire_d76_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777654(.data_in(wire_d76_53),.data_out(wire_d76_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777655(.data_in(wire_d76_54),.data_out(wire_d76_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777656(.data_in(wire_d76_55),.data_out(wire_d76_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777657(.data_in(wire_d76_56),.data_out(wire_d76_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777658(.data_in(wire_d76_57),.data_out(wire_d76_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777659(.data_in(wire_d76_58),.data_out(wire_d76_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777660(.data_in(wire_d76_59),.data_out(wire_d76_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777661(.data_in(wire_d76_60),.data_out(wire_d76_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777662(.data_in(wire_d76_61),.data_out(wire_d76_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777663(.data_in(wire_d76_62),.data_out(wire_d76_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777664(.data_in(wire_d76_63),.data_out(wire_d76_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777665(.data_in(wire_d76_64),.data_out(wire_d76_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance777666(.data_in(wire_d76_65),.data_out(wire_d76_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance777667(.data_in(wire_d76_66),.data_out(wire_d76_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777668(.data_in(wire_d76_67),.data_out(wire_d76_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777669(.data_in(wire_d76_68),.data_out(wire_d76_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777670(.data_in(wire_d76_69),.data_out(wire_d76_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777671(.data_in(wire_d76_70),.data_out(wire_d76_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance777672(.data_in(wire_d76_71),.data_out(wire_d76_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777673(.data_in(wire_d76_72),.data_out(wire_d76_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777674(.data_in(wire_d76_73),.data_out(wire_d76_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777675(.data_in(wire_d76_74),.data_out(wire_d76_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777676(.data_in(wire_d76_75),.data_out(wire_d76_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777677(.data_in(wire_d76_76),.data_out(wire_d76_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance777678(.data_in(wire_d76_77),.data_out(wire_d76_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777679(.data_in(wire_d76_78),.data_out(wire_d76_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777680(.data_in(wire_d76_79),.data_out(wire_d76_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance777681(.data_in(wire_d76_80),.data_out(wire_d76_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777682(.data_in(wire_d76_81),.data_out(wire_d76_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777683(.data_in(wire_d76_82),.data_out(wire_d76_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777684(.data_in(wire_d76_83),.data_out(wire_d76_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance777685(.data_in(wire_d76_84),.data_out(wire_d76_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777686(.data_in(wire_d76_85),.data_out(wire_d76_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777687(.data_in(wire_d76_86),.data_out(wire_d76_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777688(.data_in(wire_d76_87),.data_out(wire_d76_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance777689(.data_in(wire_d76_88),.data_out(wire_d76_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance777690(.data_in(wire_d76_89),.data_out(wire_d76_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777691(.data_in(wire_d76_90),.data_out(wire_d76_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance777692(.data_in(wire_d76_91),.data_out(wire_d76_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777693(.data_in(wire_d76_92),.data_out(wire_d76_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777694(.data_in(wire_d76_93),.data_out(wire_d76_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance777695(.data_in(wire_d76_94),.data_out(wire_d76_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777696(.data_in(wire_d76_95),.data_out(wire_d76_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777697(.data_in(wire_d76_96),.data_out(wire_d76_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance777698(.data_in(wire_d76_97),.data_out(wire_d76_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance777699(.data_in(wire_d76_98),.data_out(d_out76),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance78770(.data_in(d_in77),.data_out(wire_d77_0),.clk(clk),.rst(rst));            //channel 78
	register #(.WIDTH(WIDTH)) register_instance78771(.data_in(wire_d77_0),.data_out(wire_d77_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance78772(.data_in(wire_d77_1),.data_out(wire_d77_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance78773(.data_in(wire_d77_2),.data_out(wire_d77_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance78774(.data_in(wire_d77_3),.data_out(wire_d77_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance78775(.data_in(wire_d77_4),.data_out(wire_d77_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance78776(.data_in(wire_d77_5),.data_out(wire_d77_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance78777(.data_in(wire_d77_6),.data_out(wire_d77_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance78778(.data_in(wire_d77_7),.data_out(wire_d77_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance78779(.data_in(wire_d77_8),.data_out(wire_d77_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787710(.data_in(wire_d77_9),.data_out(wire_d77_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787711(.data_in(wire_d77_10),.data_out(wire_d77_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787712(.data_in(wire_d77_11),.data_out(wire_d77_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787713(.data_in(wire_d77_12),.data_out(wire_d77_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787714(.data_in(wire_d77_13),.data_out(wire_d77_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787715(.data_in(wire_d77_14),.data_out(wire_d77_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance787716(.data_in(wire_d77_15),.data_out(wire_d77_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787717(.data_in(wire_d77_16),.data_out(wire_d77_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787718(.data_in(wire_d77_17),.data_out(wire_d77_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787719(.data_in(wire_d77_18),.data_out(wire_d77_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787720(.data_in(wire_d77_19),.data_out(wire_d77_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787721(.data_in(wire_d77_20),.data_out(wire_d77_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787722(.data_in(wire_d77_21),.data_out(wire_d77_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance787723(.data_in(wire_d77_22),.data_out(wire_d77_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787724(.data_in(wire_d77_23),.data_out(wire_d77_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787725(.data_in(wire_d77_24),.data_out(wire_d77_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787726(.data_in(wire_d77_25),.data_out(wire_d77_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787727(.data_in(wire_d77_26),.data_out(wire_d77_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance787728(.data_in(wire_d77_27),.data_out(wire_d77_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787729(.data_in(wire_d77_28),.data_out(wire_d77_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787730(.data_in(wire_d77_29),.data_out(wire_d77_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787731(.data_in(wire_d77_30),.data_out(wire_d77_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance787732(.data_in(wire_d77_31),.data_out(wire_d77_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787733(.data_in(wire_d77_32),.data_out(wire_d77_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787734(.data_in(wire_d77_33),.data_out(wire_d77_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787735(.data_in(wire_d77_34),.data_out(wire_d77_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787736(.data_in(wire_d77_35),.data_out(wire_d77_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787737(.data_in(wire_d77_36),.data_out(wire_d77_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787738(.data_in(wire_d77_37),.data_out(wire_d77_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787739(.data_in(wire_d77_38),.data_out(wire_d77_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787740(.data_in(wire_d77_39),.data_out(wire_d77_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787741(.data_in(wire_d77_40),.data_out(wire_d77_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance787742(.data_in(wire_d77_41),.data_out(wire_d77_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787743(.data_in(wire_d77_42),.data_out(wire_d77_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787744(.data_in(wire_d77_43),.data_out(wire_d77_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance787745(.data_in(wire_d77_44),.data_out(wire_d77_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787746(.data_in(wire_d77_45),.data_out(wire_d77_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787747(.data_in(wire_d77_46),.data_out(wire_d77_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance787748(.data_in(wire_d77_47),.data_out(wire_d77_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787749(.data_in(wire_d77_48),.data_out(wire_d77_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance787750(.data_in(wire_d77_49),.data_out(wire_d77_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787751(.data_in(wire_d77_50),.data_out(wire_d77_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance787752(.data_in(wire_d77_51),.data_out(wire_d77_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787753(.data_in(wire_d77_52),.data_out(wire_d77_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787754(.data_in(wire_d77_53),.data_out(wire_d77_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787755(.data_in(wire_d77_54),.data_out(wire_d77_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787756(.data_in(wire_d77_55),.data_out(wire_d77_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787757(.data_in(wire_d77_56),.data_out(wire_d77_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787758(.data_in(wire_d77_57),.data_out(wire_d77_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787759(.data_in(wire_d77_58),.data_out(wire_d77_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787760(.data_in(wire_d77_59),.data_out(wire_d77_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance787761(.data_in(wire_d77_60),.data_out(wire_d77_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787762(.data_in(wire_d77_61),.data_out(wire_d77_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance787763(.data_in(wire_d77_62),.data_out(wire_d77_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance787764(.data_in(wire_d77_63),.data_out(wire_d77_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787765(.data_in(wire_d77_64),.data_out(wire_d77_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance787766(.data_in(wire_d77_65),.data_out(wire_d77_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance787767(.data_in(wire_d77_66),.data_out(wire_d77_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance787768(.data_in(wire_d77_67),.data_out(wire_d77_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787769(.data_in(wire_d77_68),.data_out(wire_d77_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787770(.data_in(wire_d77_69),.data_out(wire_d77_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787771(.data_in(wire_d77_70),.data_out(wire_d77_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance787772(.data_in(wire_d77_71),.data_out(wire_d77_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787773(.data_in(wire_d77_72),.data_out(wire_d77_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787774(.data_in(wire_d77_73),.data_out(wire_d77_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance787775(.data_in(wire_d77_74),.data_out(wire_d77_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787776(.data_in(wire_d77_75),.data_out(wire_d77_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787777(.data_in(wire_d77_76),.data_out(wire_d77_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787778(.data_in(wire_d77_77),.data_out(wire_d77_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance787779(.data_in(wire_d77_78),.data_out(wire_d77_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787780(.data_in(wire_d77_79),.data_out(wire_d77_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787781(.data_in(wire_d77_80),.data_out(wire_d77_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787782(.data_in(wire_d77_81),.data_out(wire_d77_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787783(.data_in(wire_d77_82),.data_out(wire_d77_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787784(.data_in(wire_d77_83),.data_out(wire_d77_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787785(.data_in(wire_d77_84),.data_out(wire_d77_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787786(.data_in(wire_d77_85),.data_out(wire_d77_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787787(.data_in(wire_d77_86),.data_out(wire_d77_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787788(.data_in(wire_d77_87),.data_out(wire_d77_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787789(.data_in(wire_d77_88),.data_out(wire_d77_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787790(.data_in(wire_d77_89),.data_out(wire_d77_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance787791(.data_in(wire_d77_90),.data_out(wire_d77_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance787792(.data_in(wire_d77_91),.data_out(wire_d77_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance787793(.data_in(wire_d77_92),.data_out(wire_d77_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787794(.data_in(wire_d77_93),.data_out(wire_d77_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787795(.data_in(wire_d77_94),.data_out(wire_d77_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787796(.data_in(wire_d77_95),.data_out(wire_d77_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance787797(.data_in(wire_d77_96),.data_out(wire_d77_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance787798(.data_in(wire_d77_97),.data_out(wire_d77_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance787799(.data_in(wire_d77_98),.data_out(d_out77),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance79780(.data_in(d_in78),.data_out(wire_d78_0),.clk(clk),.rst(rst));            //channel 79
	invertion #(.WIDTH(WIDTH)) invertion_instance79781(.data_in(wire_d78_0),.data_out(wire_d78_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance79782(.data_in(wire_d78_1),.data_out(wire_d78_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance79783(.data_in(wire_d78_2),.data_out(wire_d78_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance79784(.data_in(wire_d78_3),.data_out(wire_d78_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance79785(.data_in(wire_d78_4),.data_out(wire_d78_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance79786(.data_in(wire_d78_5),.data_out(wire_d78_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance79787(.data_in(wire_d78_6),.data_out(wire_d78_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance79788(.data_in(wire_d78_7),.data_out(wire_d78_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance79789(.data_in(wire_d78_8),.data_out(wire_d78_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance797810(.data_in(wire_d78_9),.data_out(wire_d78_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797811(.data_in(wire_d78_10),.data_out(wire_d78_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797812(.data_in(wire_d78_11),.data_out(wire_d78_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797813(.data_in(wire_d78_12),.data_out(wire_d78_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance797814(.data_in(wire_d78_13),.data_out(wire_d78_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance797815(.data_in(wire_d78_14),.data_out(wire_d78_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance797816(.data_in(wire_d78_15),.data_out(wire_d78_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance797817(.data_in(wire_d78_16),.data_out(wire_d78_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance797818(.data_in(wire_d78_17),.data_out(wire_d78_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance797819(.data_in(wire_d78_18),.data_out(wire_d78_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797820(.data_in(wire_d78_19),.data_out(wire_d78_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance797821(.data_in(wire_d78_20),.data_out(wire_d78_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance797822(.data_in(wire_d78_21),.data_out(wire_d78_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797823(.data_in(wire_d78_22),.data_out(wire_d78_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance797824(.data_in(wire_d78_23),.data_out(wire_d78_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance797825(.data_in(wire_d78_24),.data_out(wire_d78_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance797826(.data_in(wire_d78_25),.data_out(wire_d78_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797827(.data_in(wire_d78_26),.data_out(wire_d78_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance797828(.data_in(wire_d78_27),.data_out(wire_d78_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance797829(.data_in(wire_d78_28),.data_out(wire_d78_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797830(.data_in(wire_d78_29),.data_out(wire_d78_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance797831(.data_in(wire_d78_30),.data_out(wire_d78_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance797832(.data_in(wire_d78_31),.data_out(wire_d78_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance797833(.data_in(wire_d78_32),.data_out(wire_d78_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797834(.data_in(wire_d78_33),.data_out(wire_d78_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance797835(.data_in(wire_d78_34),.data_out(wire_d78_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance797836(.data_in(wire_d78_35),.data_out(wire_d78_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance797837(.data_in(wire_d78_36),.data_out(wire_d78_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance797838(.data_in(wire_d78_37),.data_out(wire_d78_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance797839(.data_in(wire_d78_38),.data_out(wire_d78_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance797840(.data_in(wire_d78_39),.data_out(wire_d78_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance797841(.data_in(wire_d78_40),.data_out(wire_d78_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797842(.data_in(wire_d78_41),.data_out(wire_d78_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797843(.data_in(wire_d78_42),.data_out(wire_d78_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance797844(.data_in(wire_d78_43),.data_out(wire_d78_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance797845(.data_in(wire_d78_44),.data_out(wire_d78_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797846(.data_in(wire_d78_45),.data_out(wire_d78_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance797847(.data_in(wire_d78_46),.data_out(wire_d78_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance797848(.data_in(wire_d78_47),.data_out(wire_d78_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797849(.data_in(wire_d78_48),.data_out(wire_d78_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance797850(.data_in(wire_d78_49),.data_out(wire_d78_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance797851(.data_in(wire_d78_50),.data_out(wire_d78_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance797852(.data_in(wire_d78_51),.data_out(wire_d78_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance797853(.data_in(wire_d78_52),.data_out(wire_d78_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797854(.data_in(wire_d78_53),.data_out(wire_d78_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797855(.data_in(wire_d78_54),.data_out(wire_d78_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797856(.data_in(wire_d78_55),.data_out(wire_d78_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance797857(.data_in(wire_d78_56),.data_out(wire_d78_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797858(.data_in(wire_d78_57),.data_out(wire_d78_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797859(.data_in(wire_d78_58),.data_out(wire_d78_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance797860(.data_in(wire_d78_59),.data_out(wire_d78_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance797861(.data_in(wire_d78_60),.data_out(wire_d78_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797862(.data_in(wire_d78_61),.data_out(wire_d78_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance797863(.data_in(wire_d78_62),.data_out(wire_d78_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797864(.data_in(wire_d78_63),.data_out(wire_d78_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797865(.data_in(wire_d78_64),.data_out(wire_d78_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance797866(.data_in(wire_d78_65),.data_out(wire_d78_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance797867(.data_in(wire_d78_66),.data_out(wire_d78_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance797868(.data_in(wire_d78_67),.data_out(wire_d78_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance797869(.data_in(wire_d78_68),.data_out(wire_d78_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797870(.data_in(wire_d78_69),.data_out(wire_d78_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance797871(.data_in(wire_d78_70),.data_out(wire_d78_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance797872(.data_in(wire_d78_71),.data_out(wire_d78_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance797873(.data_in(wire_d78_72),.data_out(wire_d78_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance797874(.data_in(wire_d78_73),.data_out(wire_d78_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance797875(.data_in(wire_d78_74),.data_out(wire_d78_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance797876(.data_in(wire_d78_75),.data_out(wire_d78_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance797877(.data_in(wire_d78_76),.data_out(wire_d78_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance797878(.data_in(wire_d78_77),.data_out(wire_d78_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance797879(.data_in(wire_d78_78),.data_out(wire_d78_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance797880(.data_in(wire_d78_79),.data_out(wire_d78_80),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance797881(.data_in(wire_d78_80),.data_out(wire_d78_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance797882(.data_in(wire_d78_81),.data_out(wire_d78_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance797883(.data_in(wire_d78_82),.data_out(wire_d78_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance797884(.data_in(wire_d78_83),.data_out(wire_d78_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance797885(.data_in(wire_d78_84),.data_out(wire_d78_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance797886(.data_in(wire_d78_85),.data_out(wire_d78_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797887(.data_in(wire_d78_86),.data_out(wire_d78_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance797888(.data_in(wire_d78_87),.data_out(wire_d78_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance797889(.data_in(wire_d78_88),.data_out(wire_d78_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797890(.data_in(wire_d78_89),.data_out(wire_d78_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance797891(.data_in(wire_d78_90),.data_out(wire_d78_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance797892(.data_in(wire_d78_91),.data_out(wire_d78_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance797893(.data_in(wire_d78_92),.data_out(wire_d78_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance797894(.data_in(wire_d78_93),.data_out(wire_d78_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance797895(.data_in(wire_d78_94),.data_out(wire_d78_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance797896(.data_in(wire_d78_95),.data_out(wire_d78_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance797897(.data_in(wire_d78_96),.data_out(wire_d78_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance797898(.data_in(wire_d78_97),.data_out(wire_d78_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance797899(.data_in(wire_d78_98),.data_out(d_out78),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance80790(.data_in(d_in79),.data_out(wire_d79_0),.clk(clk),.rst(rst));            //channel 80
	register #(.WIDTH(WIDTH)) register_instance80791(.data_in(wire_d79_0),.data_out(wire_d79_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance80792(.data_in(wire_d79_1),.data_out(wire_d79_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance80793(.data_in(wire_d79_2),.data_out(wire_d79_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance80794(.data_in(wire_d79_3),.data_out(wire_d79_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance80795(.data_in(wire_d79_4),.data_out(wire_d79_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance80796(.data_in(wire_d79_5),.data_out(wire_d79_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance80797(.data_in(wire_d79_6),.data_out(wire_d79_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance80798(.data_in(wire_d79_7),.data_out(wire_d79_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance80799(.data_in(wire_d79_8),.data_out(wire_d79_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807910(.data_in(wire_d79_9),.data_out(wire_d79_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807911(.data_in(wire_d79_10),.data_out(wire_d79_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance807912(.data_in(wire_d79_11),.data_out(wire_d79_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807913(.data_in(wire_d79_12),.data_out(wire_d79_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807914(.data_in(wire_d79_13),.data_out(wire_d79_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance807915(.data_in(wire_d79_14),.data_out(wire_d79_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807916(.data_in(wire_d79_15),.data_out(wire_d79_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance807917(.data_in(wire_d79_16),.data_out(wire_d79_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807918(.data_in(wire_d79_17),.data_out(wire_d79_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance807919(.data_in(wire_d79_18),.data_out(wire_d79_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807920(.data_in(wire_d79_19),.data_out(wire_d79_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807921(.data_in(wire_d79_20),.data_out(wire_d79_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance807922(.data_in(wire_d79_21),.data_out(wire_d79_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807923(.data_in(wire_d79_22),.data_out(wire_d79_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807924(.data_in(wire_d79_23),.data_out(wire_d79_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807925(.data_in(wire_d79_24),.data_out(wire_d79_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807926(.data_in(wire_d79_25),.data_out(wire_d79_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807927(.data_in(wire_d79_26),.data_out(wire_d79_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807928(.data_in(wire_d79_27),.data_out(wire_d79_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance807929(.data_in(wire_d79_28),.data_out(wire_d79_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807930(.data_in(wire_d79_29),.data_out(wire_d79_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807931(.data_in(wire_d79_30),.data_out(wire_d79_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807932(.data_in(wire_d79_31),.data_out(wire_d79_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807933(.data_in(wire_d79_32),.data_out(wire_d79_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance807934(.data_in(wire_d79_33),.data_out(wire_d79_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance807935(.data_in(wire_d79_34),.data_out(wire_d79_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807936(.data_in(wire_d79_35),.data_out(wire_d79_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance807937(.data_in(wire_d79_36),.data_out(wire_d79_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance807938(.data_in(wire_d79_37),.data_out(wire_d79_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance807939(.data_in(wire_d79_38),.data_out(wire_d79_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807940(.data_in(wire_d79_39),.data_out(wire_d79_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807941(.data_in(wire_d79_40),.data_out(wire_d79_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807942(.data_in(wire_d79_41),.data_out(wire_d79_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance807943(.data_in(wire_d79_42),.data_out(wire_d79_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807944(.data_in(wire_d79_43),.data_out(wire_d79_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807945(.data_in(wire_d79_44),.data_out(wire_d79_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807946(.data_in(wire_d79_45),.data_out(wire_d79_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807947(.data_in(wire_d79_46),.data_out(wire_d79_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance807948(.data_in(wire_d79_47),.data_out(wire_d79_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807949(.data_in(wire_d79_48),.data_out(wire_d79_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807950(.data_in(wire_d79_49),.data_out(wire_d79_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance807951(.data_in(wire_d79_50),.data_out(wire_d79_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance807952(.data_in(wire_d79_51),.data_out(wire_d79_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance807953(.data_in(wire_d79_52),.data_out(wire_d79_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance807954(.data_in(wire_d79_53),.data_out(wire_d79_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807955(.data_in(wire_d79_54),.data_out(wire_d79_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance807956(.data_in(wire_d79_55),.data_out(wire_d79_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807957(.data_in(wire_d79_56),.data_out(wire_d79_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807958(.data_in(wire_d79_57),.data_out(wire_d79_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance807959(.data_in(wire_d79_58),.data_out(wire_d79_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance807960(.data_in(wire_d79_59),.data_out(wire_d79_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807961(.data_in(wire_d79_60),.data_out(wire_d79_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807962(.data_in(wire_d79_61),.data_out(wire_d79_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807963(.data_in(wire_d79_62),.data_out(wire_d79_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance807964(.data_in(wire_d79_63),.data_out(wire_d79_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance807965(.data_in(wire_d79_64),.data_out(wire_d79_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807966(.data_in(wire_d79_65),.data_out(wire_d79_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance807967(.data_in(wire_d79_66),.data_out(wire_d79_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807968(.data_in(wire_d79_67),.data_out(wire_d79_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance807969(.data_in(wire_d79_68),.data_out(wire_d79_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807970(.data_in(wire_d79_69),.data_out(wire_d79_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance807971(.data_in(wire_d79_70),.data_out(wire_d79_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance807972(.data_in(wire_d79_71),.data_out(wire_d79_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807973(.data_in(wire_d79_72),.data_out(wire_d79_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance807974(.data_in(wire_d79_73),.data_out(wire_d79_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance807975(.data_in(wire_d79_74),.data_out(wire_d79_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807976(.data_in(wire_d79_75),.data_out(wire_d79_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance807977(.data_in(wire_d79_76),.data_out(wire_d79_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807978(.data_in(wire_d79_77),.data_out(wire_d79_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance807979(.data_in(wire_d79_78),.data_out(wire_d79_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance807980(.data_in(wire_d79_79),.data_out(wire_d79_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807981(.data_in(wire_d79_80),.data_out(wire_d79_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807982(.data_in(wire_d79_81),.data_out(wire_d79_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance807983(.data_in(wire_d79_82),.data_out(wire_d79_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance807984(.data_in(wire_d79_83),.data_out(wire_d79_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807985(.data_in(wire_d79_84),.data_out(wire_d79_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance807986(.data_in(wire_d79_85),.data_out(wire_d79_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance807987(.data_in(wire_d79_86),.data_out(wire_d79_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807988(.data_in(wire_d79_87),.data_out(wire_d79_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807989(.data_in(wire_d79_88),.data_out(wire_d79_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance807990(.data_in(wire_d79_89),.data_out(wire_d79_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807991(.data_in(wire_d79_90),.data_out(wire_d79_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance807992(.data_in(wire_d79_91),.data_out(wire_d79_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance807993(.data_in(wire_d79_92),.data_out(wire_d79_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance807994(.data_in(wire_d79_93),.data_out(wire_d79_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance807995(.data_in(wire_d79_94),.data_out(wire_d79_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance807996(.data_in(wire_d79_95),.data_out(wire_d79_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance807997(.data_in(wire_d79_96),.data_out(wire_d79_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance807998(.data_in(wire_d79_97),.data_out(wire_d79_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance807999(.data_in(wire_d79_98),.data_out(d_out79),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance81800(.data_in(d_in80),.data_out(wire_d80_0),.clk(clk),.rst(rst));            //channel 81
	register #(.WIDTH(WIDTH)) register_instance81801(.data_in(wire_d80_0),.data_out(wire_d80_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance81802(.data_in(wire_d80_1),.data_out(wire_d80_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance81803(.data_in(wire_d80_2),.data_out(wire_d80_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance81804(.data_in(wire_d80_3),.data_out(wire_d80_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance81805(.data_in(wire_d80_4),.data_out(wire_d80_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance81806(.data_in(wire_d80_5),.data_out(wire_d80_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance81807(.data_in(wire_d80_6),.data_out(wire_d80_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance81808(.data_in(wire_d80_7),.data_out(wire_d80_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance81809(.data_in(wire_d80_8),.data_out(wire_d80_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818010(.data_in(wire_d80_9),.data_out(wire_d80_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818011(.data_in(wire_d80_10),.data_out(wire_d80_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818012(.data_in(wire_d80_11),.data_out(wire_d80_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance818013(.data_in(wire_d80_12),.data_out(wire_d80_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818014(.data_in(wire_d80_13),.data_out(wire_d80_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818015(.data_in(wire_d80_14),.data_out(wire_d80_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818016(.data_in(wire_d80_15),.data_out(wire_d80_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818017(.data_in(wire_d80_16),.data_out(wire_d80_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818018(.data_in(wire_d80_17),.data_out(wire_d80_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance818019(.data_in(wire_d80_18),.data_out(wire_d80_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818020(.data_in(wire_d80_19),.data_out(wire_d80_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818021(.data_in(wire_d80_20),.data_out(wire_d80_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance818022(.data_in(wire_d80_21),.data_out(wire_d80_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818023(.data_in(wire_d80_22),.data_out(wire_d80_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance818024(.data_in(wire_d80_23),.data_out(wire_d80_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance818025(.data_in(wire_d80_24),.data_out(wire_d80_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance818026(.data_in(wire_d80_25),.data_out(wire_d80_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818027(.data_in(wire_d80_26),.data_out(wire_d80_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818028(.data_in(wire_d80_27),.data_out(wire_d80_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818029(.data_in(wire_d80_28),.data_out(wire_d80_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance818030(.data_in(wire_d80_29),.data_out(wire_d80_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818031(.data_in(wire_d80_30),.data_out(wire_d80_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818032(.data_in(wire_d80_31),.data_out(wire_d80_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818033(.data_in(wire_d80_32),.data_out(wire_d80_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818034(.data_in(wire_d80_33),.data_out(wire_d80_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818035(.data_in(wire_d80_34),.data_out(wire_d80_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance818036(.data_in(wire_d80_35),.data_out(wire_d80_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818037(.data_in(wire_d80_36),.data_out(wire_d80_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818038(.data_in(wire_d80_37),.data_out(wire_d80_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818039(.data_in(wire_d80_38),.data_out(wire_d80_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818040(.data_in(wire_d80_39),.data_out(wire_d80_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818041(.data_in(wire_d80_40),.data_out(wire_d80_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818042(.data_in(wire_d80_41),.data_out(wire_d80_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance818043(.data_in(wire_d80_42),.data_out(wire_d80_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818044(.data_in(wire_d80_43),.data_out(wire_d80_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance818045(.data_in(wire_d80_44),.data_out(wire_d80_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance818046(.data_in(wire_d80_45),.data_out(wire_d80_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818047(.data_in(wire_d80_46),.data_out(wire_d80_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818048(.data_in(wire_d80_47),.data_out(wire_d80_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818049(.data_in(wire_d80_48),.data_out(wire_d80_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance818050(.data_in(wire_d80_49),.data_out(wire_d80_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance818051(.data_in(wire_d80_50),.data_out(wire_d80_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818052(.data_in(wire_d80_51),.data_out(wire_d80_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818053(.data_in(wire_d80_52),.data_out(wire_d80_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818054(.data_in(wire_d80_53),.data_out(wire_d80_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818055(.data_in(wire_d80_54),.data_out(wire_d80_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818056(.data_in(wire_d80_55),.data_out(wire_d80_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance818057(.data_in(wire_d80_56),.data_out(wire_d80_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818058(.data_in(wire_d80_57),.data_out(wire_d80_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818059(.data_in(wire_d80_58),.data_out(wire_d80_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance818060(.data_in(wire_d80_59),.data_out(wire_d80_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818061(.data_in(wire_d80_60),.data_out(wire_d80_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818062(.data_in(wire_d80_61),.data_out(wire_d80_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818063(.data_in(wire_d80_62),.data_out(wire_d80_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818064(.data_in(wire_d80_63),.data_out(wire_d80_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance818065(.data_in(wire_d80_64),.data_out(wire_d80_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818066(.data_in(wire_d80_65),.data_out(wire_d80_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818067(.data_in(wire_d80_66),.data_out(wire_d80_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818068(.data_in(wire_d80_67),.data_out(wire_d80_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818069(.data_in(wire_d80_68),.data_out(wire_d80_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818070(.data_in(wire_d80_69),.data_out(wire_d80_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance818071(.data_in(wire_d80_70),.data_out(wire_d80_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818072(.data_in(wire_d80_71),.data_out(wire_d80_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818073(.data_in(wire_d80_72),.data_out(wire_d80_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818074(.data_in(wire_d80_73),.data_out(wire_d80_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818075(.data_in(wire_d80_74),.data_out(wire_d80_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818076(.data_in(wire_d80_75),.data_out(wire_d80_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818077(.data_in(wire_d80_76),.data_out(wire_d80_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance818078(.data_in(wire_d80_77),.data_out(wire_d80_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818079(.data_in(wire_d80_78),.data_out(wire_d80_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818080(.data_in(wire_d80_79),.data_out(wire_d80_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818081(.data_in(wire_d80_80),.data_out(wire_d80_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818082(.data_in(wire_d80_81),.data_out(wire_d80_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818083(.data_in(wire_d80_82),.data_out(wire_d80_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818084(.data_in(wire_d80_83),.data_out(wire_d80_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance818085(.data_in(wire_d80_84),.data_out(wire_d80_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818086(.data_in(wire_d80_85),.data_out(wire_d80_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818087(.data_in(wire_d80_86),.data_out(wire_d80_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance818088(.data_in(wire_d80_87),.data_out(wire_d80_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818089(.data_in(wire_d80_88),.data_out(wire_d80_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818090(.data_in(wire_d80_89),.data_out(wire_d80_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818091(.data_in(wire_d80_90),.data_out(wire_d80_91),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818092(.data_in(wire_d80_91),.data_out(wire_d80_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818093(.data_in(wire_d80_92),.data_out(wire_d80_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance818094(.data_in(wire_d80_93),.data_out(wire_d80_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818095(.data_in(wire_d80_94),.data_out(wire_d80_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818096(.data_in(wire_d80_95),.data_out(wire_d80_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance818097(.data_in(wire_d80_96),.data_out(wire_d80_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance818098(.data_in(wire_d80_97),.data_out(wire_d80_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance818099(.data_in(wire_d80_98),.data_out(d_out80),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance82810(.data_in(d_in81),.data_out(wire_d81_0),.clk(clk),.rst(rst));            //channel 82
	large_mux #(.WIDTH(WIDTH)) large_mux_instance82811(.data_in(wire_d81_0),.data_out(wire_d81_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance82812(.data_in(wire_d81_1),.data_out(wire_d81_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance82813(.data_in(wire_d81_2),.data_out(wire_d81_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance82814(.data_in(wire_d81_3),.data_out(wire_d81_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance82815(.data_in(wire_d81_4),.data_out(wire_d81_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance82816(.data_in(wire_d81_5),.data_out(wire_d81_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance82817(.data_in(wire_d81_6),.data_out(wire_d81_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance82818(.data_in(wire_d81_7),.data_out(wire_d81_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance82819(.data_in(wire_d81_8),.data_out(wire_d81_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828110(.data_in(wire_d81_9),.data_out(wire_d81_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828111(.data_in(wire_d81_10),.data_out(wire_d81_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance828112(.data_in(wire_d81_11),.data_out(wire_d81_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828113(.data_in(wire_d81_12),.data_out(wire_d81_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance828114(.data_in(wire_d81_13),.data_out(wire_d81_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance828115(.data_in(wire_d81_14),.data_out(wire_d81_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828116(.data_in(wire_d81_15),.data_out(wire_d81_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828117(.data_in(wire_d81_16),.data_out(wire_d81_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828118(.data_in(wire_d81_17),.data_out(wire_d81_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance828119(.data_in(wire_d81_18),.data_out(wire_d81_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance828120(.data_in(wire_d81_19),.data_out(wire_d81_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828121(.data_in(wire_d81_20),.data_out(wire_d81_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance828122(.data_in(wire_d81_21),.data_out(wire_d81_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828123(.data_in(wire_d81_22),.data_out(wire_d81_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828124(.data_in(wire_d81_23),.data_out(wire_d81_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance828125(.data_in(wire_d81_24),.data_out(wire_d81_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance828126(.data_in(wire_d81_25),.data_out(wire_d81_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance828127(.data_in(wire_d81_26),.data_out(wire_d81_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828128(.data_in(wire_d81_27),.data_out(wire_d81_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance828129(.data_in(wire_d81_28),.data_out(wire_d81_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828130(.data_in(wire_d81_29),.data_out(wire_d81_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance828131(.data_in(wire_d81_30),.data_out(wire_d81_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828132(.data_in(wire_d81_31),.data_out(wire_d81_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance828133(.data_in(wire_d81_32),.data_out(wire_d81_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828134(.data_in(wire_d81_33),.data_out(wire_d81_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance828135(.data_in(wire_d81_34),.data_out(wire_d81_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance828136(.data_in(wire_d81_35),.data_out(wire_d81_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828137(.data_in(wire_d81_36),.data_out(wire_d81_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828138(.data_in(wire_d81_37),.data_out(wire_d81_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828139(.data_in(wire_d81_38),.data_out(wire_d81_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828140(.data_in(wire_d81_39),.data_out(wire_d81_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828141(.data_in(wire_d81_40),.data_out(wire_d81_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828142(.data_in(wire_d81_41),.data_out(wire_d81_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance828143(.data_in(wire_d81_42),.data_out(wire_d81_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828144(.data_in(wire_d81_43),.data_out(wire_d81_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828145(.data_in(wire_d81_44),.data_out(wire_d81_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828146(.data_in(wire_d81_45),.data_out(wire_d81_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828147(.data_in(wire_d81_46),.data_out(wire_d81_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828148(.data_in(wire_d81_47),.data_out(wire_d81_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828149(.data_in(wire_d81_48),.data_out(wire_d81_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828150(.data_in(wire_d81_49),.data_out(wire_d81_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828151(.data_in(wire_d81_50),.data_out(wire_d81_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828152(.data_in(wire_d81_51),.data_out(wire_d81_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance828153(.data_in(wire_d81_52),.data_out(wire_d81_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance828154(.data_in(wire_d81_53),.data_out(wire_d81_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance828155(.data_in(wire_d81_54),.data_out(wire_d81_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828156(.data_in(wire_d81_55),.data_out(wire_d81_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance828157(.data_in(wire_d81_56),.data_out(wire_d81_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance828158(.data_in(wire_d81_57),.data_out(wire_d81_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance828159(.data_in(wire_d81_58),.data_out(wire_d81_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance828160(.data_in(wire_d81_59),.data_out(wire_d81_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance828161(.data_in(wire_d81_60),.data_out(wire_d81_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828162(.data_in(wire_d81_61),.data_out(wire_d81_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828163(.data_in(wire_d81_62),.data_out(wire_d81_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828164(.data_in(wire_d81_63),.data_out(wire_d81_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance828165(.data_in(wire_d81_64),.data_out(wire_d81_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828166(.data_in(wire_d81_65),.data_out(wire_d81_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828167(.data_in(wire_d81_66),.data_out(wire_d81_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828168(.data_in(wire_d81_67),.data_out(wire_d81_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828169(.data_in(wire_d81_68),.data_out(wire_d81_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance828170(.data_in(wire_d81_69),.data_out(wire_d81_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance828171(.data_in(wire_d81_70),.data_out(wire_d81_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance828172(.data_in(wire_d81_71),.data_out(wire_d81_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828173(.data_in(wire_d81_72),.data_out(wire_d81_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance828174(.data_in(wire_d81_73),.data_out(wire_d81_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828175(.data_in(wire_d81_74),.data_out(wire_d81_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828176(.data_in(wire_d81_75),.data_out(wire_d81_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance828177(.data_in(wire_d81_76),.data_out(wire_d81_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance828178(.data_in(wire_d81_77),.data_out(wire_d81_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828179(.data_in(wire_d81_78),.data_out(wire_d81_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance828180(.data_in(wire_d81_79),.data_out(wire_d81_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance828181(.data_in(wire_d81_80),.data_out(wire_d81_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance828182(.data_in(wire_d81_81),.data_out(wire_d81_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance828183(.data_in(wire_d81_82),.data_out(wire_d81_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance828184(.data_in(wire_d81_83),.data_out(wire_d81_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance828185(.data_in(wire_d81_84),.data_out(wire_d81_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance828186(.data_in(wire_d81_85),.data_out(wire_d81_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance828187(.data_in(wire_d81_86),.data_out(wire_d81_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828188(.data_in(wire_d81_87),.data_out(wire_d81_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance828189(.data_in(wire_d81_88),.data_out(wire_d81_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828190(.data_in(wire_d81_89),.data_out(wire_d81_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828191(.data_in(wire_d81_90),.data_out(wire_d81_91),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828192(.data_in(wire_d81_91),.data_out(wire_d81_92),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828193(.data_in(wire_d81_92),.data_out(wire_d81_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance828194(.data_in(wire_d81_93),.data_out(wire_d81_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance828195(.data_in(wire_d81_94),.data_out(wire_d81_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828196(.data_in(wire_d81_95),.data_out(wire_d81_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance828197(.data_in(wire_d81_96),.data_out(wire_d81_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance828198(.data_in(wire_d81_97),.data_out(wire_d81_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance828199(.data_in(wire_d81_98),.data_out(d_out81),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance83820(.data_in(d_in82),.data_out(wire_d82_0),.clk(clk),.rst(rst));            //channel 83
	register #(.WIDTH(WIDTH)) register_instance83821(.data_in(wire_d82_0),.data_out(wire_d82_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance83822(.data_in(wire_d82_1),.data_out(wire_d82_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance83823(.data_in(wire_d82_2),.data_out(wire_d82_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance83824(.data_in(wire_d82_3),.data_out(wire_d82_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance83825(.data_in(wire_d82_4),.data_out(wire_d82_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance83826(.data_in(wire_d82_5),.data_out(wire_d82_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance83827(.data_in(wire_d82_6),.data_out(wire_d82_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance83828(.data_in(wire_d82_7),.data_out(wire_d82_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance83829(.data_in(wire_d82_8),.data_out(wire_d82_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838210(.data_in(wire_d82_9),.data_out(wire_d82_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance838211(.data_in(wire_d82_10),.data_out(wire_d82_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838212(.data_in(wire_d82_11),.data_out(wire_d82_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838213(.data_in(wire_d82_12),.data_out(wire_d82_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance838214(.data_in(wire_d82_13),.data_out(wire_d82_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance838215(.data_in(wire_d82_14),.data_out(wire_d82_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838216(.data_in(wire_d82_15),.data_out(wire_d82_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838217(.data_in(wire_d82_16),.data_out(wire_d82_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance838218(.data_in(wire_d82_17),.data_out(wire_d82_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838219(.data_in(wire_d82_18),.data_out(wire_d82_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance838220(.data_in(wire_d82_19),.data_out(wire_d82_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838221(.data_in(wire_d82_20),.data_out(wire_d82_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance838222(.data_in(wire_d82_21),.data_out(wire_d82_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838223(.data_in(wire_d82_22),.data_out(wire_d82_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance838224(.data_in(wire_d82_23),.data_out(wire_d82_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838225(.data_in(wire_d82_24),.data_out(wire_d82_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838226(.data_in(wire_d82_25),.data_out(wire_d82_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance838227(.data_in(wire_d82_26),.data_out(wire_d82_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838228(.data_in(wire_d82_27),.data_out(wire_d82_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance838229(.data_in(wire_d82_28),.data_out(wire_d82_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838230(.data_in(wire_d82_29),.data_out(wire_d82_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838231(.data_in(wire_d82_30),.data_out(wire_d82_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance838232(.data_in(wire_d82_31),.data_out(wire_d82_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838233(.data_in(wire_d82_32),.data_out(wire_d82_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838234(.data_in(wire_d82_33),.data_out(wire_d82_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838235(.data_in(wire_d82_34),.data_out(wire_d82_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance838236(.data_in(wire_d82_35),.data_out(wire_d82_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance838237(.data_in(wire_d82_36),.data_out(wire_d82_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838238(.data_in(wire_d82_37),.data_out(wire_d82_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838239(.data_in(wire_d82_38),.data_out(wire_d82_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838240(.data_in(wire_d82_39),.data_out(wire_d82_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838241(.data_in(wire_d82_40),.data_out(wire_d82_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838242(.data_in(wire_d82_41),.data_out(wire_d82_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838243(.data_in(wire_d82_42),.data_out(wire_d82_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance838244(.data_in(wire_d82_43),.data_out(wire_d82_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance838245(.data_in(wire_d82_44),.data_out(wire_d82_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance838246(.data_in(wire_d82_45),.data_out(wire_d82_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance838247(.data_in(wire_d82_46),.data_out(wire_d82_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838248(.data_in(wire_d82_47),.data_out(wire_d82_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance838249(.data_in(wire_d82_48),.data_out(wire_d82_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838250(.data_in(wire_d82_49),.data_out(wire_d82_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838251(.data_in(wire_d82_50),.data_out(wire_d82_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838252(.data_in(wire_d82_51),.data_out(wire_d82_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838253(.data_in(wire_d82_52),.data_out(wire_d82_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance838254(.data_in(wire_d82_53),.data_out(wire_d82_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838255(.data_in(wire_d82_54),.data_out(wire_d82_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance838256(.data_in(wire_d82_55),.data_out(wire_d82_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance838257(.data_in(wire_d82_56),.data_out(wire_d82_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance838258(.data_in(wire_d82_57),.data_out(wire_d82_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838259(.data_in(wire_d82_58),.data_out(wire_d82_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance838260(.data_in(wire_d82_59),.data_out(wire_d82_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838261(.data_in(wire_d82_60),.data_out(wire_d82_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance838262(.data_in(wire_d82_61),.data_out(wire_d82_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838263(.data_in(wire_d82_62),.data_out(wire_d82_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838264(.data_in(wire_d82_63),.data_out(wire_d82_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance838265(.data_in(wire_d82_64),.data_out(wire_d82_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838266(.data_in(wire_d82_65),.data_out(wire_d82_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838267(.data_in(wire_d82_66),.data_out(wire_d82_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838268(.data_in(wire_d82_67),.data_out(wire_d82_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance838269(.data_in(wire_d82_68),.data_out(wire_d82_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance838270(.data_in(wire_d82_69),.data_out(wire_d82_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance838271(.data_in(wire_d82_70),.data_out(wire_d82_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838272(.data_in(wire_d82_71),.data_out(wire_d82_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838273(.data_in(wire_d82_72),.data_out(wire_d82_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838274(.data_in(wire_d82_73),.data_out(wire_d82_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance838275(.data_in(wire_d82_74),.data_out(wire_d82_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance838276(.data_in(wire_d82_75),.data_out(wire_d82_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance838277(.data_in(wire_d82_76),.data_out(wire_d82_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838278(.data_in(wire_d82_77),.data_out(wire_d82_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance838279(.data_in(wire_d82_78),.data_out(wire_d82_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance838280(.data_in(wire_d82_79),.data_out(wire_d82_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838281(.data_in(wire_d82_80),.data_out(wire_d82_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance838282(.data_in(wire_d82_81),.data_out(wire_d82_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838283(.data_in(wire_d82_82),.data_out(wire_d82_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838284(.data_in(wire_d82_83),.data_out(wire_d82_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838285(.data_in(wire_d82_84),.data_out(wire_d82_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance838286(.data_in(wire_d82_85),.data_out(wire_d82_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance838287(.data_in(wire_d82_86),.data_out(wire_d82_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance838288(.data_in(wire_d82_87),.data_out(wire_d82_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance838289(.data_in(wire_d82_88),.data_out(wire_d82_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance838290(.data_in(wire_d82_89),.data_out(wire_d82_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance838291(.data_in(wire_d82_90),.data_out(wire_d82_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance838292(.data_in(wire_d82_91),.data_out(wire_d82_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838293(.data_in(wire_d82_92),.data_out(wire_d82_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance838294(.data_in(wire_d82_93),.data_out(wire_d82_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance838295(.data_in(wire_d82_94),.data_out(wire_d82_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838296(.data_in(wire_d82_95),.data_out(wire_d82_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance838297(.data_in(wire_d82_96),.data_out(wire_d82_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance838298(.data_in(wire_d82_97),.data_out(wire_d82_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance838299(.data_in(wire_d82_98),.data_out(d_out82),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance84830(.data_in(d_in83),.data_out(wire_d83_0),.clk(clk),.rst(rst));            //channel 84
	invertion #(.WIDTH(WIDTH)) invertion_instance84831(.data_in(wire_d83_0),.data_out(wire_d83_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance84832(.data_in(wire_d83_1),.data_out(wire_d83_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance84833(.data_in(wire_d83_2),.data_out(wire_d83_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance84834(.data_in(wire_d83_3),.data_out(wire_d83_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance84835(.data_in(wire_d83_4),.data_out(wire_d83_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance84836(.data_in(wire_d83_5),.data_out(wire_d83_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance84837(.data_in(wire_d83_6),.data_out(wire_d83_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance84838(.data_in(wire_d83_7),.data_out(wire_d83_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance84839(.data_in(wire_d83_8),.data_out(wire_d83_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848310(.data_in(wire_d83_9),.data_out(wire_d83_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance848311(.data_in(wire_d83_10),.data_out(wire_d83_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848312(.data_in(wire_d83_11),.data_out(wire_d83_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848313(.data_in(wire_d83_12),.data_out(wire_d83_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance848314(.data_in(wire_d83_13),.data_out(wire_d83_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848315(.data_in(wire_d83_14),.data_out(wire_d83_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance848316(.data_in(wire_d83_15),.data_out(wire_d83_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance848317(.data_in(wire_d83_16),.data_out(wire_d83_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance848318(.data_in(wire_d83_17),.data_out(wire_d83_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848319(.data_in(wire_d83_18),.data_out(wire_d83_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848320(.data_in(wire_d83_19),.data_out(wire_d83_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848321(.data_in(wire_d83_20),.data_out(wire_d83_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance848322(.data_in(wire_d83_21),.data_out(wire_d83_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848323(.data_in(wire_d83_22),.data_out(wire_d83_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance848324(.data_in(wire_d83_23),.data_out(wire_d83_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance848325(.data_in(wire_d83_24),.data_out(wire_d83_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance848326(.data_in(wire_d83_25),.data_out(wire_d83_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848327(.data_in(wire_d83_26),.data_out(wire_d83_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance848328(.data_in(wire_d83_27),.data_out(wire_d83_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848329(.data_in(wire_d83_28),.data_out(wire_d83_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance848330(.data_in(wire_d83_29),.data_out(wire_d83_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848331(.data_in(wire_d83_30),.data_out(wire_d83_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance848332(.data_in(wire_d83_31),.data_out(wire_d83_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848333(.data_in(wire_d83_32),.data_out(wire_d83_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848334(.data_in(wire_d83_33),.data_out(wire_d83_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance848335(.data_in(wire_d83_34),.data_out(wire_d83_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance848336(.data_in(wire_d83_35),.data_out(wire_d83_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance848337(.data_in(wire_d83_36),.data_out(wire_d83_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848338(.data_in(wire_d83_37),.data_out(wire_d83_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance848339(.data_in(wire_d83_38),.data_out(wire_d83_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance848340(.data_in(wire_d83_39),.data_out(wire_d83_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848341(.data_in(wire_d83_40),.data_out(wire_d83_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance848342(.data_in(wire_d83_41),.data_out(wire_d83_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance848343(.data_in(wire_d83_42),.data_out(wire_d83_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848344(.data_in(wire_d83_43),.data_out(wire_d83_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848345(.data_in(wire_d83_44),.data_out(wire_d83_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848346(.data_in(wire_d83_45),.data_out(wire_d83_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance848347(.data_in(wire_d83_46),.data_out(wire_d83_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance848348(.data_in(wire_d83_47),.data_out(wire_d83_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848349(.data_in(wire_d83_48),.data_out(wire_d83_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848350(.data_in(wire_d83_49),.data_out(wire_d83_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance848351(.data_in(wire_d83_50),.data_out(wire_d83_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance848352(.data_in(wire_d83_51),.data_out(wire_d83_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848353(.data_in(wire_d83_52),.data_out(wire_d83_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848354(.data_in(wire_d83_53),.data_out(wire_d83_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance848355(.data_in(wire_d83_54),.data_out(wire_d83_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848356(.data_in(wire_d83_55),.data_out(wire_d83_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848357(.data_in(wire_d83_56),.data_out(wire_d83_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance848358(.data_in(wire_d83_57),.data_out(wire_d83_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance848359(.data_in(wire_d83_58),.data_out(wire_d83_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848360(.data_in(wire_d83_59),.data_out(wire_d83_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance848361(.data_in(wire_d83_60),.data_out(wire_d83_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance848362(.data_in(wire_d83_61),.data_out(wire_d83_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848363(.data_in(wire_d83_62),.data_out(wire_d83_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance848364(.data_in(wire_d83_63),.data_out(wire_d83_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance848365(.data_in(wire_d83_64),.data_out(wire_d83_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance848366(.data_in(wire_d83_65),.data_out(wire_d83_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848367(.data_in(wire_d83_66),.data_out(wire_d83_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848368(.data_in(wire_d83_67),.data_out(wire_d83_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848369(.data_in(wire_d83_68),.data_out(wire_d83_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848370(.data_in(wire_d83_69),.data_out(wire_d83_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance848371(.data_in(wire_d83_70),.data_out(wire_d83_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance848372(.data_in(wire_d83_71),.data_out(wire_d83_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848373(.data_in(wire_d83_72),.data_out(wire_d83_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848374(.data_in(wire_d83_73),.data_out(wire_d83_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848375(.data_in(wire_d83_74),.data_out(wire_d83_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance848376(.data_in(wire_d83_75),.data_out(wire_d83_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848377(.data_in(wire_d83_76),.data_out(wire_d83_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848378(.data_in(wire_d83_77),.data_out(wire_d83_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance848379(.data_in(wire_d83_78),.data_out(wire_d83_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848380(.data_in(wire_d83_79),.data_out(wire_d83_80),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance848381(.data_in(wire_d83_80),.data_out(wire_d83_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance848382(.data_in(wire_d83_81),.data_out(wire_d83_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance848383(.data_in(wire_d83_82),.data_out(wire_d83_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848384(.data_in(wire_d83_83),.data_out(wire_d83_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance848385(.data_in(wire_d83_84),.data_out(wire_d83_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848386(.data_in(wire_d83_85),.data_out(wire_d83_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848387(.data_in(wire_d83_86),.data_out(wire_d83_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance848388(.data_in(wire_d83_87),.data_out(wire_d83_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848389(.data_in(wire_d83_88),.data_out(wire_d83_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance848390(.data_in(wire_d83_89),.data_out(wire_d83_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848391(.data_in(wire_d83_90),.data_out(wire_d83_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance848392(.data_in(wire_d83_91),.data_out(wire_d83_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848393(.data_in(wire_d83_92),.data_out(wire_d83_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance848394(.data_in(wire_d83_93),.data_out(wire_d83_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance848395(.data_in(wire_d83_94),.data_out(wire_d83_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848396(.data_in(wire_d83_95),.data_out(wire_d83_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance848397(.data_in(wire_d83_96),.data_out(wire_d83_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848398(.data_in(wire_d83_97),.data_out(wire_d83_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance848399(.data_in(wire_d83_98),.data_out(d_out83),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance85840(.data_in(d_in84),.data_out(wire_d84_0),.clk(clk),.rst(rst));            //channel 85
	large_mux #(.WIDTH(WIDTH)) large_mux_instance85841(.data_in(wire_d84_0),.data_out(wire_d84_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance85842(.data_in(wire_d84_1),.data_out(wire_d84_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance85843(.data_in(wire_d84_2),.data_out(wire_d84_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance85844(.data_in(wire_d84_3),.data_out(wire_d84_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance85845(.data_in(wire_d84_4),.data_out(wire_d84_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance85846(.data_in(wire_d84_5),.data_out(wire_d84_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance85847(.data_in(wire_d84_6),.data_out(wire_d84_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance85848(.data_in(wire_d84_7),.data_out(wire_d84_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance85849(.data_in(wire_d84_8),.data_out(wire_d84_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance858410(.data_in(wire_d84_9),.data_out(wire_d84_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858411(.data_in(wire_d84_10),.data_out(wire_d84_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance858412(.data_in(wire_d84_11),.data_out(wire_d84_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858413(.data_in(wire_d84_12),.data_out(wire_d84_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858414(.data_in(wire_d84_13),.data_out(wire_d84_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858415(.data_in(wire_d84_14),.data_out(wire_d84_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858416(.data_in(wire_d84_15),.data_out(wire_d84_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858417(.data_in(wire_d84_16),.data_out(wire_d84_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858418(.data_in(wire_d84_17),.data_out(wire_d84_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858419(.data_in(wire_d84_18),.data_out(wire_d84_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance858420(.data_in(wire_d84_19),.data_out(wire_d84_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858421(.data_in(wire_d84_20),.data_out(wire_d84_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance858422(.data_in(wire_d84_21),.data_out(wire_d84_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858423(.data_in(wire_d84_22),.data_out(wire_d84_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858424(.data_in(wire_d84_23),.data_out(wire_d84_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858425(.data_in(wire_d84_24),.data_out(wire_d84_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858426(.data_in(wire_d84_25),.data_out(wire_d84_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858427(.data_in(wire_d84_26),.data_out(wire_d84_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858428(.data_in(wire_d84_27),.data_out(wire_d84_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance858429(.data_in(wire_d84_28),.data_out(wire_d84_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance858430(.data_in(wire_d84_29),.data_out(wire_d84_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858431(.data_in(wire_d84_30),.data_out(wire_d84_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance858432(.data_in(wire_d84_31),.data_out(wire_d84_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858433(.data_in(wire_d84_32),.data_out(wire_d84_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance858434(.data_in(wire_d84_33),.data_out(wire_d84_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance858435(.data_in(wire_d84_34),.data_out(wire_d84_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance858436(.data_in(wire_d84_35),.data_out(wire_d84_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858437(.data_in(wire_d84_36),.data_out(wire_d84_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858438(.data_in(wire_d84_37),.data_out(wire_d84_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858439(.data_in(wire_d84_38),.data_out(wire_d84_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858440(.data_in(wire_d84_39),.data_out(wire_d84_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858441(.data_in(wire_d84_40),.data_out(wire_d84_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858442(.data_in(wire_d84_41),.data_out(wire_d84_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance858443(.data_in(wire_d84_42),.data_out(wire_d84_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858444(.data_in(wire_d84_43),.data_out(wire_d84_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858445(.data_in(wire_d84_44),.data_out(wire_d84_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858446(.data_in(wire_d84_45),.data_out(wire_d84_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858447(.data_in(wire_d84_46),.data_out(wire_d84_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858448(.data_in(wire_d84_47),.data_out(wire_d84_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858449(.data_in(wire_d84_48),.data_out(wire_d84_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance858450(.data_in(wire_d84_49),.data_out(wire_d84_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858451(.data_in(wire_d84_50),.data_out(wire_d84_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858452(.data_in(wire_d84_51),.data_out(wire_d84_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance858453(.data_in(wire_d84_52),.data_out(wire_d84_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance858454(.data_in(wire_d84_53),.data_out(wire_d84_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858455(.data_in(wire_d84_54),.data_out(wire_d84_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858456(.data_in(wire_d84_55),.data_out(wire_d84_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858457(.data_in(wire_d84_56),.data_out(wire_d84_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858458(.data_in(wire_d84_57),.data_out(wire_d84_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance858459(.data_in(wire_d84_58),.data_out(wire_d84_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance858460(.data_in(wire_d84_59),.data_out(wire_d84_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858461(.data_in(wire_d84_60),.data_out(wire_d84_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858462(.data_in(wire_d84_61),.data_out(wire_d84_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858463(.data_in(wire_d84_62),.data_out(wire_d84_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance858464(.data_in(wire_d84_63),.data_out(wire_d84_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858465(.data_in(wire_d84_64),.data_out(wire_d84_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858466(.data_in(wire_d84_65),.data_out(wire_d84_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858467(.data_in(wire_d84_66),.data_out(wire_d84_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858468(.data_in(wire_d84_67),.data_out(wire_d84_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858469(.data_in(wire_d84_68),.data_out(wire_d84_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858470(.data_in(wire_d84_69),.data_out(wire_d84_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance858471(.data_in(wire_d84_70),.data_out(wire_d84_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858472(.data_in(wire_d84_71),.data_out(wire_d84_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858473(.data_in(wire_d84_72),.data_out(wire_d84_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858474(.data_in(wire_d84_73),.data_out(wire_d84_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858475(.data_in(wire_d84_74),.data_out(wire_d84_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858476(.data_in(wire_d84_75),.data_out(wire_d84_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858477(.data_in(wire_d84_76),.data_out(wire_d84_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858478(.data_in(wire_d84_77),.data_out(wire_d84_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance858479(.data_in(wire_d84_78),.data_out(wire_d84_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858480(.data_in(wire_d84_79),.data_out(wire_d84_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858481(.data_in(wire_d84_80),.data_out(wire_d84_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858482(.data_in(wire_d84_81),.data_out(wire_d84_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858483(.data_in(wire_d84_82),.data_out(wire_d84_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858484(.data_in(wire_d84_83),.data_out(wire_d84_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858485(.data_in(wire_d84_84),.data_out(wire_d84_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858486(.data_in(wire_d84_85),.data_out(wire_d84_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858487(.data_in(wire_d84_86),.data_out(wire_d84_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858488(.data_in(wire_d84_87),.data_out(wire_d84_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance858489(.data_in(wire_d84_88),.data_out(wire_d84_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858490(.data_in(wire_d84_89),.data_out(wire_d84_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858491(.data_in(wire_d84_90),.data_out(wire_d84_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858492(.data_in(wire_d84_91),.data_out(wire_d84_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858493(.data_in(wire_d84_92),.data_out(wire_d84_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858494(.data_in(wire_d84_93),.data_out(wire_d84_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858495(.data_in(wire_d84_94),.data_out(wire_d84_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858496(.data_in(wire_d84_95),.data_out(wire_d84_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance858497(.data_in(wire_d84_96),.data_out(wire_d84_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance858498(.data_in(wire_d84_97),.data_out(wire_d84_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance858499(.data_in(wire_d84_98),.data_out(d_out84),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance86850(.data_in(d_in85),.data_out(wire_d85_0),.clk(clk),.rst(rst));            //channel 86
	register #(.WIDTH(WIDTH)) register_instance86851(.data_in(wire_d85_0),.data_out(wire_d85_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance86852(.data_in(wire_d85_1),.data_out(wire_d85_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance86853(.data_in(wire_d85_2),.data_out(wire_d85_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance86854(.data_in(wire_d85_3),.data_out(wire_d85_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance86855(.data_in(wire_d85_4),.data_out(wire_d85_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance86856(.data_in(wire_d85_5),.data_out(wire_d85_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance86857(.data_in(wire_d85_6),.data_out(wire_d85_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance86858(.data_in(wire_d85_7),.data_out(wire_d85_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance86859(.data_in(wire_d85_8),.data_out(wire_d85_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance868510(.data_in(wire_d85_9),.data_out(wire_d85_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868511(.data_in(wire_d85_10),.data_out(wire_d85_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance868512(.data_in(wire_d85_11),.data_out(wire_d85_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868513(.data_in(wire_d85_12),.data_out(wire_d85_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868514(.data_in(wire_d85_13),.data_out(wire_d85_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868515(.data_in(wire_d85_14),.data_out(wire_d85_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868516(.data_in(wire_d85_15),.data_out(wire_d85_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868517(.data_in(wire_d85_16),.data_out(wire_d85_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868518(.data_in(wire_d85_17),.data_out(wire_d85_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance868519(.data_in(wire_d85_18),.data_out(wire_d85_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance868520(.data_in(wire_d85_19),.data_out(wire_d85_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868521(.data_in(wire_d85_20),.data_out(wire_d85_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance868522(.data_in(wire_d85_21),.data_out(wire_d85_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868523(.data_in(wire_d85_22),.data_out(wire_d85_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance868524(.data_in(wire_d85_23),.data_out(wire_d85_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance868525(.data_in(wire_d85_24),.data_out(wire_d85_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868526(.data_in(wire_d85_25),.data_out(wire_d85_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance868527(.data_in(wire_d85_26),.data_out(wire_d85_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868528(.data_in(wire_d85_27),.data_out(wire_d85_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance868529(.data_in(wire_d85_28),.data_out(wire_d85_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance868530(.data_in(wire_d85_29),.data_out(wire_d85_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance868531(.data_in(wire_d85_30),.data_out(wire_d85_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance868532(.data_in(wire_d85_31),.data_out(wire_d85_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868533(.data_in(wire_d85_32),.data_out(wire_d85_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868534(.data_in(wire_d85_33),.data_out(wire_d85_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868535(.data_in(wire_d85_34),.data_out(wire_d85_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance868536(.data_in(wire_d85_35),.data_out(wire_d85_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance868537(.data_in(wire_d85_36),.data_out(wire_d85_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance868538(.data_in(wire_d85_37),.data_out(wire_d85_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance868539(.data_in(wire_d85_38),.data_out(wire_d85_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance868540(.data_in(wire_d85_39),.data_out(wire_d85_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868541(.data_in(wire_d85_40),.data_out(wire_d85_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868542(.data_in(wire_d85_41),.data_out(wire_d85_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868543(.data_in(wire_d85_42),.data_out(wire_d85_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance868544(.data_in(wire_d85_43),.data_out(wire_d85_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868545(.data_in(wire_d85_44),.data_out(wire_d85_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868546(.data_in(wire_d85_45),.data_out(wire_d85_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance868547(.data_in(wire_d85_46),.data_out(wire_d85_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868548(.data_in(wire_d85_47),.data_out(wire_d85_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868549(.data_in(wire_d85_48),.data_out(wire_d85_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance868550(.data_in(wire_d85_49),.data_out(wire_d85_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance868551(.data_in(wire_d85_50),.data_out(wire_d85_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance868552(.data_in(wire_d85_51),.data_out(wire_d85_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance868553(.data_in(wire_d85_52),.data_out(wire_d85_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868554(.data_in(wire_d85_53),.data_out(wire_d85_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868555(.data_in(wire_d85_54),.data_out(wire_d85_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868556(.data_in(wire_d85_55),.data_out(wire_d85_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868557(.data_in(wire_d85_56),.data_out(wire_d85_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance868558(.data_in(wire_d85_57),.data_out(wire_d85_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868559(.data_in(wire_d85_58),.data_out(wire_d85_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868560(.data_in(wire_d85_59),.data_out(wire_d85_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance868561(.data_in(wire_d85_60),.data_out(wire_d85_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance868562(.data_in(wire_d85_61),.data_out(wire_d85_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance868563(.data_in(wire_d85_62),.data_out(wire_d85_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance868564(.data_in(wire_d85_63),.data_out(wire_d85_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868565(.data_in(wire_d85_64),.data_out(wire_d85_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868566(.data_in(wire_d85_65),.data_out(wire_d85_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance868567(.data_in(wire_d85_66),.data_out(wire_d85_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868568(.data_in(wire_d85_67),.data_out(wire_d85_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868569(.data_in(wire_d85_68),.data_out(wire_d85_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance868570(.data_in(wire_d85_69),.data_out(wire_d85_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance868571(.data_in(wire_d85_70),.data_out(wire_d85_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance868572(.data_in(wire_d85_71),.data_out(wire_d85_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance868573(.data_in(wire_d85_72),.data_out(wire_d85_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868574(.data_in(wire_d85_73),.data_out(wire_d85_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868575(.data_in(wire_d85_74),.data_out(wire_d85_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance868576(.data_in(wire_d85_75),.data_out(wire_d85_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance868577(.data_in(wire_d85_76),.data_out(wire_d85_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance868578(.data_in(wire_d85_77),.data_out(wire_d85_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868579(.data_in(wire_d85_78),.data_out(wire_d85_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868580(.data_in(wire_d85_79),.data_out(wire_d85_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868581(.data_in(wire_d85_80),.data_out(wire_d85_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868582(.data_in(wire_d85_81),.data_out(wire_d85_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance868583(.data_in(wire_d85_82),.data_out(wire_d85_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance868584(.data_in(wire_d85_83),.data_out(wire_d85_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868585(.data_in(wire_d85_84),.data_out(wire_d85_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance868586(.data_in(wire_d85_85),.data_out(wire_d85_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868587(.data_in(wire_d85_86),.data_out(wire_d85_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance868588(.data_in(wire_d85_87),.data_out(wire_d85_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868589(.data_in(wire_d85_88),.data_out(wire_d85_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance868590(.data_in(wire_d85_89),.data_out(wire_d85_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868591(.data_in(wire_d85_90),.data_out(wire_d85_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance868592(.data_in(wire_d85_91),.data_out(wire_d85_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868593(.data_in(wire_d85_92),.data_out(wire_d85_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868594(.data_in(wire_d85_93),.data_out(wire_d85_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance868595(.data_in(wire_d85_94),.data_out(wire_d85_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868596(.data_in(wire_d85_95),.data_out(wire_d85_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868597(.data_in(wire_d85_96),.data_out(wire_d85_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance868598(.data_in(wire_d85_97),.data_out(wire_d85_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance868599(.data_in(wire_d85_98),.data_out(d_out85),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance87860(.data_in(d_in86),.data_out(wire_d86_0),.clk(clk),.rst(rst));            //channel 87
	register #(.WIDTH(WIDTH)) register_instance87861(.data_in(wire_d86_0),.data_out(wire_d86_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87862(.data_in(wire_d86_1),.data_out(wire_d86_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance87863(.data_in(wire_d86_2),.data_out(wire_d86_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance87864(.data_in(wire_d86_3),.data_out(wire_d86_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance87865(.data_in(wire_d86_4),.data_out(wire_d86_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance87866(.data_in(wire_d86_5),.data_out(wire_d86_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance87867(.data_in(wire_d86_6),.data_out(wire_d86_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance87868(.data_in(wire_d86_7),.data_out(wire_d86_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance87869(.data_in(wire_d86_8),.data_out(wire_d86_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878610(.data_in(wire_d86_9),.data_out(wire_d86_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878611(.data_in(wire_d86_10),.data_out(wire_d86_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878612(.data_in(wire_d86_11),.data_out(wire_d86_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878613(.data_in(wire_d86_12),.data_out(wire_d86_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878614(.data_in(wire_d86_13),.data_out(wire_d86_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance878615(.data_in(wire_d86_14),.data_out(wire_d86_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878616(.data_in(wire_d86_15),.data_out(wire_d86_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878617(.data_in(wire_d86_16),.data_out(wire_d86_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878618(.data_in(wire_d86_17),.data_out(wire_d86_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance878619(.data_in(wire_d86_18),.data_out(wire_d86_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878620(.data_in(wire_d86_19),.data_out(wire_d86_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878621(.data_in(wire_d86_20),.data_out(wire_d86_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878622(.data_in(wire_d86_21),.data_out(wire_d86_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance878623(.data_in(wire_d86_22),.data_out(wire_d86_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878624(.data_in(wire_d86_23),.data_out(wire_d86_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance878625(.data_in(wire_d86_24),.data_out(wire_d86_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878626(.data_in(wire_d86_25),.data_out(wire_d86_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878627(.data_in(wire_d86_26),.data_out(wire_d86_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878628(.data_in(wire_d86_27),.data_out(wire_d86_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance878629(.data_in(wire_d86_28),.data_out(wire_d86_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878630(.data_in(wire_d86_29),.data_out(wire_d86_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878631(.data_in(wire_d86_30),.data_out(wire_d86_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance878632(.data_in(wire_d86_31),.data_out(wire_d86_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878633(.data_in(wire_d86_32),.data_out(wire_d86_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878634(.data_in(wire_d86_33),.data_out(wire_d86_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878635(.data_in(wire_d86_34),.data_out(wire_d86_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance878636(.data_in(wire_d86_35),.data_out(wire_d86_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878637(.data_in(wire_d86_36),.data_out(wire_d86_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance878638(.data_in(wire_d86_37),.data_out(wire_d86_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance878639(.data_in(wire_d86_38),.data_out(wire_d86_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance878640(.data_in(wire_d86_39),.data_out(wire_d86_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878641(.data_in(wire_d86_40),.data_out(wire_d86_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance878642(.data_in(wire_d86_41),.data_out(wire_d86_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance878643(.data_in(wire_d86_42),.data_out(wire_d86_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878644(.data_in(wire_d86_43),.data_out(wire_d86_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878645(.data_in(wire_d86_44),.data_out(wire_d86_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878646(.data_in(wire_d86_45),.data_out(wire_d86_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance878647(.data_in(wire_d86_46),.data_out(wire_d86_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878648(.data_in(wire_d86_47),.data_out(wire_d86_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878649(.data_in(wire_d86_48),.data_out(wire_d86_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878650(.data_in(wire_d86_49),.data_out(wire_d86_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878651(.data_in(wire_d86_50),.data_out(wire_d86_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878652(.data_in(wire_d86_51),.data_out(wire_d86_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878653(.data_in(wire_d86_52),.data_out(wire_d86_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878654(.data_in(wire_d86_53),.data_out(wire_d86_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878655(.data_in(wire_d86_54),.data_out(wire_d86_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance878656(.data_in(wire_d86_55),.data_out(wire_d86_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance878657(.data_in(wire_d86_56),.data_out(wire_d86_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878658(.data_in(wire_d86_57),.data_out(wire_d86_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878659(.data_in(wire_d86_58),.data_out(wire_d86_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878660(.data_in(wire_d86_59),.data_out(wire_d86_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878661(.data_in(wire_d86_60),.data_out(wire_d86_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance878662(.data_in(wire_d86_61),.data_out(wire_d86_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878663(.data_in(wire_d86_62),.data_out(wire_d86_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878664(.data_in(wire_d86_63),.data_out(wire_d86_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878665(.data_in(wire_d86_64),.data_out(wire_d86_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878666(.data_in(wire_d86_65),.data_out(wire_d86_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878667(.data_in(wire_d86_66),.data_out(wire_d86_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878668(.data_in(wire_d86_67),.data_out(wire_d86_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878669(.data_in(wire_d86_68),.data_out(wire_d86_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878670(.data_in(wire_d86_69),.data_out(wire_d86_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance878671(.data_in(wire_d86_70),.data_out(wire_d86_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878672(.data_in(wire_d86_71),.data_out(wire_d86_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878673(.data_in(wire_d86_72),.data_out(wire_d86_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance878674(.data_in(wire_d86_73),.data_out(wire_d86_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878675(.data_in(wire_d86_74),.data_out(wire_d86_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878676(.data_in(wire_d86_75),.data_out(wire_d86_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance878677(.data_in(wire_d86_76),.data_out(wire_d86_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878678(.data_in(wire_d86_77),.data_out(wire_d86_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878679(.data_in(wire_d86_78),.data_out(wire_d86_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878680(.data_in(wire_d86_79),.data_out(wire_d86_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878681(.data_in(wire_d86_80),.data_out(wire_d86_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878682(.data_in(wire_d86_81),.data_out(wire_d86_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878683(.data_in(wire_d86_82),.data_out(wire_d86_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878684(.data_in(wire_d86_83),.data_out(wire_d86_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878685(.data_in(wire_d86_84),.data_out(wire_d86_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878686(.data_in(wire_d86_85),.data_out(wire_d86_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878687(.data_in(wire_d86_86),.data_out(wire_d86_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878688(.data_in(wire_d86_87),.data_out(wire_d86_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance878689(.data_in(wire_d86_88),.data_out(wire_d86_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878690(.data_in(wire_d86_89),.data_out(wire_d86_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878691(.data_in(wire_d86_90),.data_out(wire_d86_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878692(.data_in(wire_d86_91),.data_out(wire_d86_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878693(.data_in(wire_d86_92),.data_out(wire_d86_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878694(.data_in(wire_d86_93),.data_out(wire_d86_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878695(.data_in(wire_d86_94),.data_out(wire_d86_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance878696(.data_in(wire_d86_95),.data_out(wire_d86_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878697(.data_in(wire_d86_96),.data_out(wire_d86_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878698(.data_in(wire_d86_97),.data_out(wire_d86_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878699(.data_in(wire_d86_98),.data_out(d_out86),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance88870(.data_in(d_in87),.data_out(wire_d87_0),.clk(clk),.rst(rst));            //channel 88
	invertion #(.WIDTH(WIDTH)) invertion_instance88871(.data_in(wire_d87_0),.data_out(wire_d87_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance88872(.data_in(wire_d87_1),.data_out(wire_d87_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance88873(.data_in(wire_d87_2),.data_out(wire_d87_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance88874(.data_in(wire_d87_3),.data_out(wire_d87_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance88875(.data_in(wire_d87_4),.data_out(wire_d87_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance88876(.data_in(wire_d87_5),.data_out(wire_d87_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance88877(.data_in(wire_d87_6),.data_out(wire_d87_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance88878(.data_in(wire_d87_7),.data_out(wire_d87_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance88879(.data_in(wire_d87_8),.data_out(wire_d87_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance888710(.data_in(wire_d87_9),.data_out(wire_d87_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance888711(.data_in(wire_d87_10),.data_out(wire_d87_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance888712(.data_in(wire_d87_11),.data_out(wire_d87_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance888713(.data_in(wire_d87_12),.data_out(wire_d87_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance888714(.data_in(wire_d87_13),.data_out(wire_d87_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance888715(.data_in(wire_d87_14),.data_out(wire_d87_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance888716(.data_in(wire_d87_15),.data_out(wire_d87_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance888717(.data_in(wire_d87_16),.data_out(wire_d87_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance888718(.data_in(wire_d87_17),.data_out(wire_d87_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance888719(.data_in(wire_d87_18),.data_out(wire_d87_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance888720(.data_in(wire_d87_19),.data_out(wire_d87_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance888721(.data_in(wire_d87_20),.data_out(wire_d87_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance888722(.data_in(wire_d87_21),.data_out(wire_d87_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance888723(.data_in(wire_d87_22),.data_out(wire_d87_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888724(.data_in(wire_d87_23),.data_out(wire_d87_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance888725(.data_in(wire_d87_24),.data_out(wire_d87_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance888726(.data_in(wire_d87_25),.data_out(wire_d87_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance888727(.data_in(wire_d87_26),.data_out(wire_d87_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance888728(.data_in(wire_d87_27),.data_out(wire_d87_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance888729(.data_in(wire_d87_28),.data_out(wire_d87_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance888730(.data_in(wire_d87_29),.data_out(wire_d87_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance888731(.data_in(wire_d87_30),.data_out(wire_d87_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888732(.data_in(wire_d87_31),.data_out(wire_d87_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance888733(.data_in(wire_d87_32),.data_out(wire_d87_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance888734(.data_in(wire_d87_33),.data_out(wire_d87_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance888735(.data_in(wire_d87_34),.data_out(wire_d87_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888736(.data_in(wire_d87_35),.data_out(wire_d87_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888737(.data_in(wire_d87_36),.data_out(wire_d87_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888738(.data_in(wire_d87_37),.data_out(wire_d87_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888739(.data_in(wire_d87_38),.data_out(wire_d87_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance888740(.data_in(wire_d87_39),.data_out(wire_d87_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance888741(.data_in(wire_d87_40),.data_out(wire_d87_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888742(.data_in(wire_d87_41),.data_out(wire_d87_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance888743(.data_in(wire_d87_42),.data_out(wire_d87_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance888744(.data_in(wire_d87_43),.data_out(wire_d87_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance888745(.data_in(wire_d87_44),.data_out(wire_d87_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance888746(.data_in(wire_d87_45),.data_out(wire_d87_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance888747(.data_in(wire_d87_46),.data_out(wire_d87_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance888748(.data_in(wire_d87_47),.data_out(wire_d87_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance888749(.data_in(wire_d87_48),.data_out(wire_d87_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888750(.data_in(wire_d87_49),.data_out(wire_d87_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance888751(.data_in(wire_d87_50),.data_out(wire_d87_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance888752(.data_in(wire_d87_51),.data_out(wire_d87_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance888753(.data_in(wire_d87_52),.data_out(wire_d87_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance888754(.data_in(wire_d87_53),.data_out(wire_d87_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888755(.data_in(wire_d87_54),.data_out(wire_d87_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance888756(.data_in(wire_d87_55),.data_out(wire_d87_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance888757(.data_in(wire_d87_56),.data_out(wire_d87_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888758(.data_in(wire_d87_57),.data_out(wire_d87_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance888759(.data_in(wire_d87_58),.data_out(wire_d87_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888760(.data_in(wire_d87_59),.data_out(wire_d87_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888761(.data_in(wire_d87_60),.data_out(wire_d87_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance888762(.data_in(wire_d87_61),.data_out(wire_d87_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance888763(.data_in(wire_d87_62),.data_out(wire_d87_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance888764(.data_in(wire_d87_63),.data_out(wire_d87_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance888765(.data_in(wire_d87_64),.data_out(wire_d87_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance888766(.data_in(wire_d87_65),.data_out(wire_d87_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance888767(.data_in(wire_d87_66),.data_out(wire_d87_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance888768(.data_in(wire_d87_67),.data_out(wire_d87_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888769(.data_in(wire_d87_68),.data_out(wire_d87_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888770(.data_in(wire_d87_69),.data_out(wire_d87_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888771(.data_in(wire_d87_70),.data_out(wire_d87_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance888772(.data_in(wire_d87_71),.data_out(wire_d87_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888773(.data_in(wire_d87_72),.data_out(wire_d87_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance888774(.data_in(wire_d87_73),.data_out(wire_d87_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance888775(.data_in(wire_d87_74),.data_out(wire_d87_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888776(.data_in(wire_d87_75),.data_out(wire_d87_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance888777(.data_in(wire_d87_76),.data_out(wire_d87_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance888778(.data_in(wire_d87_77),.data_out(wire_d87_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888779(.data_in(wire_d87_78),.data_out(wire_d87_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance888780(.data_in(wire_d87_79),.data_out(wire_d87_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888781(.data_in(wire_d87_80),.data_out(wire_d87_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance888782(.data_in(wire_d87_81),.data_out(wire_d87_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888783(.data_in(wire_d87_82),.data_out(wire_d87_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance888784(.data_in(wire_d87_83),.data_out(wire_d87_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance888785(.data_in(wire_d87_84),.data_out(wire_d87_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance888786(.data_in(wire_d87_85),.data_out(wire_d87_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888787(.data_in(wire_d87_86),.data_out(wire_d87_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance888788(.data_in(wire_d87_87),.data_out(wire_d87_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance888789(.data_in(wire_d87_88),.data_out(wire_d87_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance888790(.data_in(wire_d87_89),.data_out(wire_d87_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888791(.data_in(wire_d87_90),.data_out(wire_d87_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance888792(.data_in(wire_d87_91),.data_out(wire_d87_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance888793(.data_in(wire_d87_92),.data_out(wire_d87_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance888794(.data_in(wire_d87_93),.data_out(wire_d87_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance888795(.data_in(wire_d87_94),.data_out(wire_d87_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance888796(.data_in(wire_d87_95),.data_out(wire_d87_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888797(.data_in(wire_d87_96),.data_out(wire_d87_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance888798(.data_in(wire_d87_97),.data_out(wire_d87_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance888799(.data_in(wire_d87_98),.data_out(d_out87),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance89880(.data_in(d_in88),.data_out(wire_d88_0),.clk(clk),.rst(rst));            //channel 89
	large_mux #(.WIDTH(WIDTH)) large_mux_instance89881(.data_in(wire_d88_0),.data_out(wire_d88_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance89882(.data_in(wire_d88_1),.data_out(wire_d88_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance89883(.data_in(wire_d88_2),.data_out(wire_d88_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance89884(.data_in(wire_d88_3),.data_out(wire_d88_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance89885(.data_in(wire_d88_4),.data_out(wire_d88_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance89886(.data_in(wire_d88_5),.data_out(wire_d88_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance89887(.data_in(wire_d88_6),.data_out(wire_d88_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance89888(.data_in(wire_d88_7),.data_out(wire_d88_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance89889(.data_in(wire_d88_8),.data_out(wire_d88_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance898810(.data_in(wire_d88_9),.data_out(wire_d88_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance898811(.data_in(wire_d88_10),.data_out(wire_d88_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898812(.data_in(wire_d88_11),.data_out(wire_d88_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance898813(.data_in(wire_d88_12),.data_out(wire_d88_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898814(.data_in(wire_d88_13),.data_out(wire_d88_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance898815(.data_in(wire_d88_14),.data_out(wire_d88_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance898816(.data_in(wire_d88_15),.data_out(wire_d88_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898817(.data_in(wire_d88_16),.data_out(wire_d88_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance898818(.data_in(wire_d88_17),.data_out(wire_d88_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898819(.data_in(wire_d88_18),.data_out(wire_d88_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance898820(.data_in(wire_d88_19),.data_out(wire_d88_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898821(.data_in(wire_d88_20),.data_out(wire_d88_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance898822(.data_in(wire_d88_21),.data_out(wire_d88_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance898823(.data_in(wire_d88_22),.data_out(wire_d88_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898824(.data_in(wire_d88_23),.data_out(wire_d88_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898825(.data_in(wire_d88_24),.data_out(wire_d88_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance898826(.data_in(wire_d88_25),.data_out(wire_d88_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance898827(.data_in(wire_d88_26),.data_out(wire_d88_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898828(.data_in(wire_d88_27),.data_out(wire_d88_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance898829(.data_in(wire_d88_28),.data_out(wire_d88_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898830(.data_in(wire_d88_29),.data_out(wire_d88_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance898831(.data_in(wire_d88_30),.data_out(wire_d88_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898832(.data_in(wire_d88_31),.data_out(wire_d88_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898833(.data_in(wire_d88_32),.data_out(wire_d88_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance898834(.data_in(wire_d88_33),.data_out(wire_d88_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898835(.data_in(wire_d88_34),.data_out(wire_d88_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance898836(.data_in(wire_d88_35),.data_out(wire_d88_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance898837(.data_in(wire_d88_36),.data_out(wire_d88_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898838(.data_in(wire_d88_37),.data_out(wire_d88_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance898839(.data_in(wire_d88_38),.data_out(wire_d88_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance898840(.data_in(wire_d88_39),.data_out(wire_d88_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance898841(.data_in(wire_d88_40),.data_out(wire_d88_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance898842(.data_in(wire_d88_41),.data_out(wire_d88_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance898843(.data_in(wire_d88_42),.data_out(wire_d88_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance898844(.data_in(wire_d88_43),.data_out(wire_d88_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance898845(.data_in(wire_d88_44),.data_out(wire_d88_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance898846(.data_in(wire_d88_45),.data_out(wire_d88_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898847(.data_in(wire_d88_46),.data_out(wire_d88_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898848(.data_in(wire_d88_47),.data_out(wire_d88_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898849(.data_in(wire_d88_48),.data_out(wire_d88_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance898850(.data_in(wire_d88_49),.data_out(wire_d88_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898851(.data_in(wire_d88_50),.data_out(wire_d88_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898852(.data_in(wire_d88_51),.data_out(wire_d88_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898853(.data_in(wire_d88_52),.data_out(wire_d88_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance898854(.data_in(wire_d88_53),.data_out(wire_d88_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance898855(.data_in(wire_d88_54),.data_out(wire_d88_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898856(.data_in(wire_d88_55),.data_out(wire_d88_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898857(.data_in(wire_d88_56),.data_out(wire_d88_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898858(.data_in(wire_d88_57),.data_out(wire_d88_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898859(.data_in(wire_d88_58),.data_out(wire_d88_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898860(.data_in(wire_d88_59),.data_out(wire_d88_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898861(.data_in(wire_d88_60),.data_out(wire_d88_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance898862(.data_in(wire_d88_61),.data_out(wire_d88_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898863(.data_in(wire_d88_62),.data_out(wire_d88_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance898864(.data_in(wire_d88_63),.data_out(wire_d88_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance898865(.data_in(wire_d88_64),.data_out(wire_d88_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance898866(.data_in(wire_d88_65),.data_out(wire_d88_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898867(.data_in(wire_d88_66),.data_out(wire_d88_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898868(.data_in(wire_d88_67),.data_out(wire_d88_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898869(.data_in(wire_d88_68),.data_out(wire_d88_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898870(.data_in(wire_d88_69),.data_out(wire_d88_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898871(.data_in(wire_d88_70),.data_out(wire_d88_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance898872(.data_in(wire_d88_71),.data_out(wire_d88_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance898873(.data_in(wire_d88_72),.data_out(wire_d88_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance898874(.data_in(wire_d88_73),.data_out(wire_d88_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898875(.data_in(wire_d88_74),.data_out(wire_d88_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898876(.data_in(wire_d88_75),.data_out(wire_d88_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance898877(.data_in(wire_d88_76),.data_out(wire_d88_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance898878(.data_in(wire_d88_77),.data_out(wire_d88_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance898879(.data_in(wire_d88_78),.data_out(wire_d88_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance898880(.data_in(wire_d88_79),.data_out(wire_d88_80),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance898881(.data_in(wire_d88_80),.data_out(wire_d88_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance898882(.data_in(wire_d88_81),.data_out(wire_d88_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance898883(.data_in(wire_d88_82),.data_out(wire_d88_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance898884(.data_in(wire_d88_83),.data_out(wire_d88_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898885(.data_in(wire_d88_84),.data_out(wire_d88_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance898886(.data_in(wire_d88_85),.data_out(wire_d88_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898887(.data_in(wire_d88_86),.data_out(wire_d88_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898888(.data_in(wire_d88_87),.data_out(wire_d88_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898889(.data_in(wire_d88_88),.data_out(wire_d88_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898890(.data_in(wire_d88_89),.data_out(wire_d88_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance898891(.data_in(wire_d88_90),.data_out(wire_d88_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898892(.data_in(wire_d88_91),.data_out(wire_d88_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898893(.data_in(wire_d88_92),.data_out(wire_d88_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance898894(.data_in(wire_d88_93),.data_out(wire_d88_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898895(.data_in(wire_d88_94),.data_out(wire_d88_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898896(.data_in(wire_d88_95),.data_out(wire_d88_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898897(.data_in(wire_d88_96),.data_out(wire_d88_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898898(.data_in(wire_d88_97),.data_out(wire_d88_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance898899(.data_in(wire_d88_98),.data_out(d_out88),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance90890(.data_in(d_in89),.data_out(wire_d89_0),.clk(clk),.rst(rst));            //channel 90
	encoder #(.WIDTH(WIDTH)) encoder_instance90891(.data_in(wire_d89_0),.data_out(wire_d89_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance90892(.data_in(wire_d89_1),.data_out(wire_d89_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance90893(.data_in(wire_d89_2),.data_out(wire_d89_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance90894(.data_in(wire_d89_3),.data_out(wire_d89_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance90895(.data_in(wire_d89_4),.data_out(wire_d89_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance90896(.data_in(wire_d89_5),.data_out(wire_d89_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance90897(.data_in(wire_d89_6),.data_out(wire_d89_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance90898(.data_in(wire_d89_7),.data_out(wire_d89_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance90899(.data_in(wire_d89_8),.data_out(wire_d89_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance908910(.data_in(wire_d89_9),.data_out(wire_d89_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance908911(.data_in(wire_d89_10),.data_out(wire_d89_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908912(.data_in(wire_d89_11),.data_out(wire_d89_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance908913(.data_in(wire_d89_12),.data_out(wire_d89_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908914(.data_in(wire_d89_13),.data_out(wire_d89_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance908915(.data_in(wire_d89_14),.data_out(wire_d89_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908916(.data_in(wire_d89_15),.data_out(wire_d89_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908917(.data_in(wire_d89_16),.data_out(wire_d89_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance908918(.data_in(wire_d89_17),.data_out(wire_d89_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908919(.data_in(wire_d89_18),.data_out(wire_d89_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908920(.data_in(wire_d89_19),.data_out(wire_d89_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance908921(.data_in(wire_d89_20),.data_out(wire_d89_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908922(.data_in(wire_d89_21),.data_out(wire_d89_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance908923(.data_in(wire_d89_22),.data_out(wire_d89_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance908924(.data_in(wire_d89_23),.data_out(wire_d89_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908925(.data_in(wire_d89_24),.data_out(wire_d89_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908926(.data_in(wire_d89_25),.data_out(wire_d89_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance908927(.data_in(wire_d89_26),.data_out(wire_d89_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance908928(.data_in(wire_d89_27),.data_out(wire_d89_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance908929(.data_in(wire_d89_28),.data_out(wire_d89_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908930(.data_in(wire_d89_29),.data_out(wire_d89_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908931(.data_in(wire_d89_30),.data_out(wire_d89_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908932(.data_in(wire_d89_31),.data_out(wire_d89_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908933(.data_in(wire_d89_32),.data_out(wire_d89_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908934(.data_in(wire_d89_33),.data_out(wire_d89_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance908935(.data_in(wire_d89_34),.data_out(wire_d89_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance908936(.data_in(wire_d89_35),.data_out(wire_d89_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908937(.data_in(wire_d89_36),.data_out(wire_d89_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance908938(.data_in(wire_d89_37),.data_out(wire_d89_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908939(.data_in(wire_d89_38),.data_out(wire_d89_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908940(.data_in(wire_d89_39),.data_out(wire_d89_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance908941(.data_in(wire_d89_40),.data_out(wire_d89_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908942(.data_in(wire_d89_41),.data_out(wire_d89_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908943(.data_in(wire_d89_42),.data_out(wire_d89_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance908944(.data_in(wire_d89_43),.data_out(wire_d89_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance908945(.data_in(wire_d89_44),.data_out(wire_d89_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance908946(.data_in(wire_d89_45),.data_out(wire_d89_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908947(.data_in(wire_d89_46),.data_out(wire_d89_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908948(.data_in(wire_d89_47),.data_out(wire_d89_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908949(.data_in(wire_d89_48),.data_out(wire_d89_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance908950(.data_in(wire_d89_49),.data_out(wire_d89_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908951(.data_in(wire_d89_50),.data_out(wire_d89_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance908952(.data_in(wire_d89_51),.data_out(wire_d89_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908953(.data_in(wire_d89_52),.data_out(wire_d89_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908954(.data_in(wire_d89_53),.data_out(wire_d89_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908955(.data_in(wire_d89_54),.data_out(wire_d89_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance908956(.data_in(wire_d89_55),.data_out(wire_d89_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908957(.data_in(wire_d89_56),.data_out(wire_d89_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908958(.data_in(wire_d89_57),.data_out(wire_d89_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908959(.data_in(wire_d89_58),.data_out(wire_d89_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908960(.data_in(wire_d89_59),.data_out(wire_d89_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908961(.data_in(wire_d89_60),.data_out(wire_d89_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908962(.data_in(wire_d89_61),.data_out(wire_d89_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908963(.data_in(wire_d89_62),.data_out(wire_d89_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908964(.data_in(wire_d89_63),.data_out(wire_d89_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance908965(.data_in(wire_d89_64),.data_out(wire_d89_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance908966(.data_in(wire_d89_65),.data_out(wire_d89_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance908967(.data_in(wire_d89_66),.data_out(wire_d89_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance908968(.data_in(wire_d89_67),.data_out(wire_d89_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance908969(.data_in(wire_d89_68),.data_out(wire_d89_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908970(.data_in(wire_d89_69),.data_out(wire_d89_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance908971(.data_in(wire_d89_70),.data_out(wire_d89_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908972(.data_in(wire_d89_71),.data_out(wire_d89_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908973(.data_in(wire_d89_72),.data_out(wire_d89_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance908974(.data_in(wire_d89_73),.data_out(wire_d89_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908975(.data_in(wire_d89_74),.data_out(wire_d89_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908976(.data_in(wire_d89_75),.data_out(wire_d89_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance908977(.data_in(wire_d89_76),.data_out(wire_d89_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance908978(.data_in(wire_d89_77),.data_out(wire_d89_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance908979(.data_in(wire_d89_78),.data_out(wire_d89_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908980(.data_in(wire_d89_79),.data_out(wire_d89_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908981(.data_in(wire_d89_80),.data_out(wire_d89_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908982(.data_in(wire_d89_81),.data_out(wire_d89_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance908983(.data_in(wire_d89_82),.data_out(wire_d89_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908984(.data_in(wire_d89_83),.data_out(wire_d89_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908985(.data_in(wire_d89_84),.data_out(wire_d89_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance908986(.data_in(wire_d89_85),.data_out(wire_d89_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908987(.data_in(wire_d89_86),.data_out(wire_d89_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance908988(.data_in(wire_d89_87),.data_out(wire_d89_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance908989(.data_in(wire_d89_88),.data_out(wire_d89_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance908990(.data_in(wire_d89_89),.data_out(wire_d89_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908991(.data_in(wire_d89_90),.data_out(wire_d89_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance908992(.data_in(wire_d89_91),.data_out(wire_d89_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908993(.data_in(wire_d89_92),.data_out(wire_d89_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance908994(.data_in(wire_d89_93),.data_out(wire_d89_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance908995(.data_in(wire_d89_94),.data_out(wire_d89_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance908996(.data_in(wire_d89_95),.data_out(wire_d89_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance908997(.data_in(wire_d89_96),.data_out(wire_d89_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance908998(.data_in(wire_d89_97),.data_out(wire_d89_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance908999(.data_in(wire_d89_98),.data_out(d_out89),.clk(clk),.rst(rst));


endmodule