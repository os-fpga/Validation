`define P1 32
`define P2 32