module co_sim_matrix_mult_3x3_iverilog;
	reg [143:0] A;
	reg [143:0] B;
	wire [143:0] Result;


	integer mismatch=0;

`ifdef PNR
		matrix_mult_3x3_iverilog inst(
		 A[143] ,
    A[142] ,
    A[141] ,
    A[140] ,
    A[139] ,
    A[138] ,
    A[137] ,
    A[136] ,
    A[135] ,
    A[134] ,
    A[133] ,
    A[132] ,
    A[131] ,
    A[130] ,
    A[129] ,
    A[128] ,
    A[127] ,
    A[126] ,
    A[125] ,
    A[124] ,
    A[123] ,
    A[122] ,
    A[121] ,
    A[120] ,
    A[119] ,
    A[118] ,
    A[117] ,
    A[116] ,
    A[115] ,
    A[114] ,
    A[113] ,
    A[112] ,
    A[111] ,
    A[110] ,
    A[109] ,
    A[108] ,
    A[107] ,
    A[106] ,
    A[105] ,
    A[104] ,
    A[103] ,
    A[102] ,
    A[101] ,
    A[100] ,
    A[99] ,
    A[98] ,
    A[97] ,
    A[96] ,
    A[95] ,
    A[94] ,
    A[93] ,
    A[92] ,
    A[91] ,
    A[90] ,
    A[89] ,
    A[88] ,
    A[87] ,
    A[86] ,
    A[85] ,
    A[84] ,
    A[83] ,
    A[82] ,
    A[81] ,
    A[80] ,
    A[79] ,
    A[78] ,
    A[77] ,
    A[76] ,
    A[75] ,
    A[74] ,
    A[73] ,
    A[72] ,
    A[71] ,
    A[70] ,
    A[69] ,
    A[68] ,
    A[67] ,
    A[66] ,
    A[65] ,
    A[64] ,
    A[63] ,
    A[62] ,
    A[61] ,
    A[60] ,
    A[59] ,
    A[58] ,
    A[57] ,
    A[56] ,
    A[55] ,
    A[54] ,
    A[53] ,
    A[52] ,
    A[51] ,
    A[50] ,
    A[49] ,
    A[48] ,
    A[47] ,
    A[46] ,
    A[45] ,
    A[44] ,
    A[43] ,
    A[42] ,
    A[41] ,
    A[40] ,
    A[39] ,
    A[38] ,
    A[37] ,
    A[36] ,
    A[35] ,
    A[34] ,
    A[33] ,
    A[32] ,
    A[31] ,
    A[30] ,
    A[29] ,
    A[28] ,
    A[27] ,
    A[26] ,
    A[25] ,
    A[24] ,
    A[23] ,
    A[22] ,
    A[21] ,
    A[20] ,
    A[19] ,
    A[18] ,
    A[17] ,
    A[16] ,
    A[15] ,
    A[14] ,
    A[13] ,
    A[12] ,
    A[11] ,
    A[10] ,
    A[9] ,
    A[8] ,
    A[7] ,
    A[6] ,
    A[5] ,
    A[4] ,
    A[3] ,
    A[2] ,
    A[1] ,
    A[0] ,
    B[143] ,
    B[142] ,
    B[141] ,
    B[140] ,
    B[139] ,
    B[138] ,
    B[137] ,
    B[136] ,
    B[135] ,
    B[134] ,
    B[133] ,
    B[132] ,
    B[131] ,
    B[130] ,
    B[129] ,
    B[128] ,
    B[127] ,
    B[126] ,
    B[125] ,
    B[124] ,
    B[123] ,
    B[122] ,
    B[121] ,
    B[120] ,
    B[119] ,
    B[118] ,
    B[117] ,
    B[116] ,
    B[115] ,
    B[114] ,
    B[113] ,
    B[112] ,
    B[111] ,
    B[110] ,
    B[109] ,
    B[108] ,
    B[107] ,
    B[106] ,
    B[105] ,
    B[104] ,
    B[103] ,
    B[102] ,
    B[101] ,
    B[100] ,
    B[99] ,
    B[98] ,
    B[97] ,
    B[96] ,
    B[95] ,
    B[94] ,
    B[93] ,
    B[92] ,
    B[91] ,
    B[90] ,
    B[89] ,
    B[88] ,
    B[87] ,
    B[86] ,
    B[85] ,
    B[84] ,
    B[83] ,
    B[82] ,
    B[81] ,
    B[80] ,
    B[79] ,
    B[78] ,
    B[77] ,
    B[76] ,
    B[75] ,
    B[74] ,
    B[73] ,
    B[72] ,
    B[71] ,
    B[70] ,
    B[69] ,
    B[68] ,
    B[67] ,
    B[66] ,
    B[65] ,
    B[64] ,
    B[63] ,
    B[62] ,
    B[61] ,
    B[60] ,
    B[59] ,
    B[58] ,
    B[57] ,
    B[56] ,
    B[55] ,
    B[54] ,
    B[53] ,
    B[52] ,
    B[51] ,
    B[50] ,
    B[49] ,
    B[48] ,
    B[47] ,
    B[46] ,
    B[45] ,
    B[44] ,
    B[43] ,
    B[42] ,
    B[41] ,
    B[40] ,
    B[39] ,
    B[38] ,
    B[37] ,
    B[36] ,
    B[35] ,
    B[34] ,
    B[33] ,
    B[32] ,
    B[31] ,
    B[30] ,
    B[29] ,
    B[28] ,
    B[27] ,
    B[26] ,
    B[25] ,
    B[24] ,
    B[23] ,
    B[22] ,
    B[21] ,
    B[20] ,
    B[19] ,
    B[18] ,
    B[17] ,
    B[16] ,
    B[15] ,
    B[14] ,
    B[13] ,
    B[12] ,
    B[11] ,
    B[10] ,
    B[9] ,
    B[8] ,
    B[7] ,
    B[6] ,
    B[5] ,
    B[4] ,
    B[3] ,
    B[2] ,
    B[1] ,
    B[0] ,
    Result[29] ,
    Result[136] ,
    Result[72] ,
    Result[7] ,
    Result[107] ,
    Result[27] ,
    Result[89] ,
    Result[88] ,
    Result[95] ,
    Result[94] ,
    Result[92] ,
    Result[40] ,
    Result[135] ,
    Result[71] ,
    Result[124] ,
    Result[134] ,
    Result[109] ,
    Result[70] ,
    Result[38] ,
    Result[30] ,
    Result[142] ,
    Result[126] ,
    Result[78] ,
    Result[46] ,
    Result[11] ,
    Result[90] ,
    Result[110] ,
    Result[24] ,
    Result[141] ,
    Result[125] ,
    Result[77] ,
    Result[45] ,
    Result[9] ,
    Result[111] ,
    Result[108] ,
    Result[55] ,
    Result[31] ,
    Result[143] ,
    Result[127] ,
    Result[79] ,
    Result[47] ,
    Result[15] ,
    Result[14] ,
    Result[93] ,
    Result[91] ,
    Result[59] ,
    Result[54] ,
    Result[120] ,
    Result[104] ,
    Result[56] ,
    Result[123] ,
    Result[122] ,
    Result[137] ,
    Result[73] ,
    Result[41] ,
    Result[106] ,
    Result[28] ,
    Result[139] ,
    Result[75] ,
    Result[43] ,
    Result[119] ,
    Result[118] ,
    Result[61] ,
    Result[103] ,
    Result[140] ,
    Result[76] ,
    Result[44] ,
    Result[62] ,
    Result[13] ,
    Result[12] ,
    Result[6] ,
    Result[121] ,
    Result[105] ,
    Result[63] ,
    Result[60] ,
    Result[57] ,
    Result[138] ,
    Result[74] ,
    Result[42] ,
    Result[39] ,
    Result[58] ,
    Result[26] ,
    Result[102] ,
    Result[86] ,
    Result[101] ,
    Result[25] ,
    Result[22] ,
    Result[87] ,
    Result[10] ,
    Result[8] ,
    Result[5] ,
    Result[133] ,
    Result[69] ,
    Result[37] ,
    Result[85] ,
    Result[117] ,
    Result[53] ,
    Result[21] ,
    Result[23] ,
    Result[100] ,
    Result[84] ,
    Result[4] ,
    Result[132] ,
    Result[116] ,
    Result[68] ,
    Result[52] ,
    Result[36] ,
    Result[20] ,
    Result[131] ,
    Result[99] ,
    Result[83] ,
    Result[67] ,
    Result[35] ,
    Result[19] ,
    Result[98] ,
    Result[82] ,
    Result[2] ,
    Result[3] ,
    Result[130] ,
    Result[115] ,
    Result[114] ,
    Result[66] ,
    Result[51] ,
    Result[50] ,
    Result[34] ,
    Result[18] ,
    Result[129] ,
    Result[113] ,
    Result[97] ,
    Result[81] ,
    Result[65] ,
    Result[49] ,
    Result[33] ,
    Result[17] ,
    Result[1] ,
    Result[128] ,
    Result[112] ,
    Result[96] ,
    Result[80] ,
    Result[64] ,
    Result[48] ,
    Result[32] ,
    Result[16] ,
    Result[0]  );
`else
   	matrix_mult_3x3_iverilog inst(.*);
`endif
initial begin
	A=0;
	B=0;
	$display ("\n\n*** Random Functionality Tests for multiplier with signed inputs are applied***\n\n");
	repeat (1000) begin
		A = $urandom;
		B = $urandom;
		#10;
		display_stimulus;
		display_output;
		#10;
	end
	$display ("\n\n***Random Functionality Tests for multiplier with signed inputs are ended***\n\n");

	A=0;
	B=0;

	$display ("\n\n***Directed Functionality Test for multiplier is applied***\n\n");
	A = 20'hfffff;
	B = 18'h3ffff;
	#10;
	display_stimulus;
	display_output;
	$display ("\n\n***Directed Functionality Test for multiplier is ended***\n\n");
	#100;
	if(mismatch == 0)
        $display("\n**** All Comparison Matched ***\nSimulation Passed");
    else
        $display("%0d comparison(s) mismatched\nERROR: SIM: Simulation Failed", mismatch);
	$finish;
	end
	

task display_stimulus;
	$display ($time,," Test stimulus is: A=%0d, B=%0d", A, B);
endtask
task display_output;
	$display ($time,," Output is: %0d" ,Result);
endtask


initial begin
    $dumpfile("tb.vcd");
    $dumpvars;
end
endmodule