// `include "register_vhd.v"
// `include "alu_top_vhd.v"
// `include "decoder_top_vhd.v"
// `include "mux_top_vhd.v"
// `include "shift_reg_top_vhd.v"
// `include "rom_top_vhd.v"

module design394_36_37_top #(parameter WIDTH=32,CHANNEL=36) (clk, rst, in, out);

	localparam OUT_BUS=CHANNEL*WIDTH;
	input clk,rst;
	input [WIDTH-1:0] in;
	output [WIDTH-1:0] out;

	reg [WIDTH-1:0] d_in0;
	reg [WIDTH-1:0] d_in1;
	reg [WIDTH-1:0] d_in2;
	reg [WIDTH-1:0] d_in3;
	reg [WIDTH-1:0] d_in4;
	reg [WIDTH-1:0] d_in5;
	reg [WIDTH-1:0] d_in6;
	reg [WIDTH-1:0] d_in7;
	reg [WIDTH-1:0] d_in8;
	reg [WIDTH-1:0] d_in9;
	reg [WIDTH-1:0] d_in10;
	reg [WIDTH-1:0] d_in11;
	reg [WIDTH-1:0] d_in12;
	reg [WIDTH-1:0] d_in13;
	reg [WIDTH-1:0] d_in14;
	reg [WIDTH-1:0] d_in15;
	reg [WIDTH-1:0] d_in16;
	reg [WIDTH-1:0] d_in17;
	reg [WIDTH-1:0] d_in18;
	reg [WIDTH-1:0] d_in19;
	reg [WIDTH-1:0] d_in20;
	reg [WIDTH-1:0] d_in21;
	reg [WIDTH-1:0] d_in22;
	reg [WIDTH-1:0] d_in23;
	reg [WIDTH-1:0] d_in24;
	reg [WIDTH-1:0] d_in25;
	reg [WIDTH-1:0] d_in26;
	reg [WIDTH-1:0] d_in27;
	reg [WIDTH-1:0] d_in28;
	reg [WIDTH-1:0] d_in29;
	reg [WIDTH-1:0] d_in30;
	reg [WIDTH-1:0] d_in31;
	reg [WIDTH-1:0] d_in32;
	reg [WIDTH-1:0] d_in33;
	reg [WIDTH-1:0] d_in34;
	reg [WIDTH-1:0] d_in35;
	wire [WIDTH-1:0] d_out0;
	wire [WIDTH-1:0] d_out1;
	wire [WIDTH-1:0] d_out2;
	wire [WIDTH-1:0] d_out3;
	wire [WIDTH-1:0] d_out4;
	wire [WIDTH-1:0] d_out5;
	wire [WIDTH-1:0] d_out6;
	wire [WIDTH-1:0] d_out7;
	wire [WIDTH-1:0] d_out8;
	wire [WIDTH-1:0] d_out9;
	wire [WIDTH-1:0] d_out10;
	wire [WIDTH-1:0] d_out11;
	wire [WIDTH-1:0] d_out12;
	wire [WIDTH-1:0] d_out13;
	wire [WIDTH-1:0] d_out14;
	wire [WIDTH-1:0] d_out15;
	wire [WIDTH-1:0] d_out16;
	wire [WIDTH-1:0] d_out17;
	wire [WIDTH-1:0] d_out18;
	wire [WIDTH-1:0] d_out19;
	wire [WIDTH-1:0] d_out20;
	wire [WIDTH-1:0] d_out21;
	wire [WIDTH-1:0] d_out22;
	wire [WIDTH-1:0] d_out23;
	wire [WIDTH-1:0] d_out24;
	wire [WIDTH-1:0] d_out25;
	wire [WIDTH-1:0] d_out26;
	wire [WIDTH-1:0] d_out27;
	wire [WIDTH-1:0] d_out28;
	wire [WIDTH-1:0] d_out29;
	wire [WIDTH-1:0] d_out30;
	wire [WIDTH-1:0] d_out31;
	wire [WIDTH-1:0] d_out32;
	wire [WIDTH-1:0] d_out33;
	wire [WIDTH-1:0] d_out34;
	wire [WIDTH-1:0] d_out35;

	reg [OUT_BUS-1:0] tmp;

	always @ (posedge clk or posedge rst) begin
		if (rst)
			tmp <= 0;
		else
			tmp <= {tmp[OUT_BUS-(WIDTH-1):0],in};
	end

	always @ (posedge clk) begin
		d_in0 <= tmp[WIDTH-1:0];
		d_in1 <= tmp[(WIDTH*2)-1:WIDTH*1];
		d_in2 <= tmp[(WIDTH*3)-1:WIDTH*2];
		d_in3 <= tmp[(WIDTH*4)-1:WIDTH*3];
		d_in4 <= tmp[(WIDTH*5)-1:WIDTH*4];
		d_in5 <= tmp[(WIDTH*6)-1:WIDTH*5];
		d_in6 <= tmp[(WIDTH*7)-1:WIDTH*6];
		d_in7 <= tmp[(WIDTH*8)-1:WIDTH*7];
		d_in8 <= tmp[(WIDTH*9)-1:WIDTH*8];
		d_in9 <= tmp[(WIDTH*10)-1:WIDTH*9];
		d_in10 <= tmp[(WIDTH*11)-1:WIDTH*10];
		d_in11 <= tmp[(WIDTH*12)-1:WIDTH*11];
		d_in12 <= tmp[(WIDTH*13)-1:WIDTH*12];
		d_in13 <= tmp[(WIDTH*14)-1:WIDTH*13];
		d_in14 <= tmp[(WIDTH*15)-1:WIDTH*14];
		d_in15 <= tmp[(WIDTH*16)-1:WIDTH*15];
		d_in16 <= tmp[(WIDTH*17)-1:WIDTH*16];
		d_in17 <= tmp[(WIDTH*18)-1:WIDTH*17];
		d_in18 <= tmp[(WIDTH*19)-1:WIDTH*18];
		d_in19 <= tmp[(WIDTH*20)-1:WIDTH*19];
		d_in20 <= tmp[(WIDTH*21)-1:WIDTH*20];
		d_in21 <= tmp[(WIDTH*22)-1:WIDTH*21];
		d_in22 <= tmp[(WIDTH*23)-1:WIDTH*22];
		d_in23 <= tmp[(WIDTH*24)-1:WIDTH*23];
		d_in24 <= tmp[(WIDTH*25)-1:WIDTH*24];
		d_in25 <= tmp[(WIDTH*26)-1:WIDTH*25];
		d_in26 <= tmp[(WIDTH*27)-1:WIDTH*26];
		d_in27 <= tmp[(WIDTH*28)-1:WIDTH*27];
		d_in28 <= tmp[(WIDTH*29)-1:WIDTH*28];
		d_in29 <= tmp[(WIDTH*30)-1:WIDTH*29];
		d_in30 <= tmp[(WIDTH*31)-1:WIDTH*30];
		d_in31 <= tmp[(WIDTH*32)-1:WIDTH*31];
		d_in32 <= tmp[(WIDTH*33)-1:WIDTH*32];
		d_in33 <= tmp[(WIDTH*34)-1:WIDTH*33];
		d_in34 <= tmp[(WIDTH*35)-1:WIDTH*34];
		d_in35 <= tmp[(WIDTH*36)-1:WIDTH*35];
	end

	design394_36_37 #(.WIDTH(WIDTH)) design394_36_37_inst(.d_in0(d_in0),.d_in1(d_in1),.d_in2(d_in2),.d_in3(d_in3),.d_in4(d_in4),.d_in5(d_in5),.d_in6(d_in6),.d_in7(d_in7),.d_in8(d_in8),.d_in9(d_in9),.d_in10(d_in10),.d_in11(d_in11),.d_in12(d_in12),.d_in13(d_in13),.d_in14(d_in14),.d_in15(d_in15),.d_in16(d_in16),.d_in17(d_in17),.d_in18(d_in18),.d_in19(d_in19),.d_in20(d_in20),.d_in21(d_in21),.d_in22(d_in22),.d_in23(d_in23),.d_in24(d_in24),.d_in25(d_in25),.d_in26(d_in26),.d_in27(d_in27),.d_in28(d_in28),.d_in29(d_in29),.d_in30(d_in30),.d_in31(d_in31),.d_in32(d_in32),.d_in33(d_in33),.d_in34(d_in34),.d_in35(d_in35),.d_out0(d_out0),.d_out1(d_out1),.d_out2(d_out2),.d_out3(d_out3),.d_out4(d_out4),.d_out5(d_out5),.d_out6(d_out6),.d_out7(d_out7),.d_out8(d_out8),.d_out9(d_out9),.d_out10(d_out10),.d_out11(d_out11),.d_out12(d_out12),.d_out13(d_out13),.d_out14(d_out14),.d_out15(d_out15),.d_out16(d_out16),.d_out17(d_out17),.d_out18(d_out18),.d_out19(d_out19),.d_out20(d_out20),.d_out21(d_out21),.d_out22(d_out22),.d_out23(d_out23),.d_out24(d_out24),.d_out25(d_out25),.d_out26(d_out26),.d_out27(d_out27),.d_out28(d_out28),.d_out29(d_out29),.d_out30(d_out30),.d_out31(d_out31),.d_out32(d_out32),.d_out33(d_out33),.d_out34(d_out34),.d_out35(d_out35),.clk(clk),.rst(rst));

	assign out = d_out0^d_out1^d_out2^d_out3^d_out4^d_out5^d_out6^d_out7^d_out8^d_out9^d_out10^d_out11^d_out12^d_out13^d_out14^d_out15^d_out16^d_out17^d_out18^d_out19^d_out20^d_out21^d_out22^d_out23^d_out24^d_out25^d_out26^d_out27^d_out28^d_out29^d_out30^d_out31^d_out32^d_out33^d_out34^d_out35;

endmodule

module design394_36_37 #(parameter WIDTH=32) (d_in0, d_in1, d_in2, d_in3, d_in4, d_in5, d_in6, d_in7, d_in8, d_in9, d_in10, d_in11, d_in12, d_in13, d_in14, d_in15, d_in16, d_in17, d_in18, d_in19, d_in20, d_in21, d_in22, d_in23, d_in24, d_in25, d_in26, d_in27, d_in28, d_in29, d_in30, d_in31, d_in32, d_in33, d_in34, d_in35, d_out0, d_out1, d_out2, d_out3, d_out4, d_out5, d_out6, d_out7, d_out8, d_out9, d_out10, d_out11, d_out12, d_out13, d_out14, d_out15, d_out16, d_out17, d_out18, d_out19, d_out20, d_out21, d_out22, d_out23, d_out24, d_out25, d_out26, d_out27, d_out28, d_out29, d_out30, d_out31, d_out32, d_out33, d_out34, d_out35, clk, rst);
	input clk;
	input rst;
	input [WIDTH-1:0] d_in0; 
	input [WIDTH-1:0] d_in1; 
	input [WIDTH-1:0] d_in2; 
	input [WIDTH-1:0] d_in3; 
	input [WIDTH-1:0] d_in4; 
	input [WIDTH-1:0] d_in5; 
	input [WIDTH-1:0] d_in6; 
	input [WIDTH-1:0] d_in7; 
	input [WIDTH-1:0] d_in8; 
	input [WIDTH-1:0] d_in9; 
	input [WIDTH-1:0] d_in10; 
	input [WIDTH-1:0] d_in11; 
	input [WIDTH-1:0] d_in12; 
	input [WIDTH-1:0] d_in13; 
	input [WIDTH-1:0] d_in14; 
	input [WIDTH-1:0] d_in15; 
	input [WIDTH-1:0] d_in16; 
	input [WIDTH-1:0] d_in17; 
	input [WIDTH-1:0] d_in18; 
	input [WIDTH-1:0] d_in19; 
	input [WIDTH-1:0] d_in20; 
	input [WIDTH-1:0] d_in21; 
	input [WIDTH-1:0] d_in22; 
	input [WIDTH-1:0] d_in23; 
	input [WIDTH-1:0] d_in24; 
	input [WIDTH-1:0] d_in25; 
	input [WIDTH-1:0] d_in26; 
	input [WIDTH-1:0] d_in27; 
	input [WIDTH-1:0] d_in28; 
	input [WIDTH-1:0] d_in29; 
	input [WIDTH-1:0] d_in30; 
	input [WIDTH-1:0] d_in31; 
	input [WIDTH-1:0] d_in32; 
	input [WIDTH-1:0] d_in33; 
	input [WIDTH-1:0] d_in34; 
	input [WIDTH-1:0] d_in35; 
	output [WIDTH-1:0] d_out0; 
	output [WIDTH-1:0] d_out1; 
	output [WIDTH-1:0] d_out2; 
	output [WIDTH-1:0] d_out3; 
	output [WIDTH-1:0] d_out4; 
	output [WIDTH-1:0] d_out5; 
	output [WIDTH-1:0] d_out6; 
	output [WIDTH-1:0] d_out7; 
	output [WIDTH-1:0] d_out8; 
	output [WIDTH-1:0] d_out9; 
	output [WIDTH-1:0] d_out10; 
	output [WIDTH-1:0] d_out11; 
	output [WIDTH-1:0] d_out12; 
	output [WIDTH-1:0] d_out13; 
	output [WIDTH-1:0] d_out14; 
	output [WIDTH-1:0] d_out15; 
	output [WIDTH-1:0] d_out16; 
	output [WIDTH-1:0] d_out17; 
	output [WIDTH-1:0] d_out18; 
	output [WIDTH-1:0] d_out19; 
	output [WIDTH-1:0] d_out20; 
	output [WIDTH-1:0] d_out21; 
	output [WIDTH-1:0] d_out22; 
	output [WIDTH-1:0] d_out23; 
	output [WIDTH-1:0] d_out24; 
	output [WIDTH-1:0] d_out25; 
	output [WIDTH-1:0] d_out26; 
	output [WIDTH-1:0] d_out27; 
	output [WIDTH-1:0] d_out28; 
	output [WIDTH-1:0] d_out29; 
	output [WIDTH-1:0] d_out30; 
	output [WIDTH-1:0] d_out31; 
	output [WIDTH-1:0] d_out32; 
	output [WIDTH-1:0] d_out33; 
	output [WIDTH-1:0] d_out34; 
	output [WIDTH-1:0] d_out35; 

	wire [WIDTH-1:0] wire_d0_0;
	wire [WIDTH-1:0] wire_d0_1;
	wire [WIDTH-1:0] wire_d0_2;
	wire [WIDTH-1:0] wire_d0_3;
	wire [WIDTH-1:0] wire_d0_4;
	wire [WIDTH-1:0] wire_d0_5;
	wire [WIDTH-1:0] wire_d0_6;
	wire [WIDTH-1:0] wire_d0_7;
	wire [WIDTH-1:0] wire_d0_8;
	wire [WIDTH-1:0] wire_d0_9;
	wire [WIDTH-1:0] wire_d0_10;
	wire [WIDTH-1:0] wire_d0_11;
	wire [WIDTH-1:0] wire_d0_12;
	wire [WIDTH-1:0] wire_d0_13;
	wire [WIDTH-1:0] wire_d0_14;
	wire [WIDTH-1:0] wire_d0_15;
	wire [WIDTH-1:0] wire_d0_16;
	wire [WIDTH-1:0] wire_d0_17;
	wire [WIDTH-1:0] wire_d0_18;
	wire [WIDTH-1:0] wire_d0_19;
	wire [WIDTH-1:0] wire_d0_20;
	wire [WIDTH-1:0] wire_d0_21;
	wire [WIDTH-1:0] wire_d0_22;
	wire [WIDTH-1:0] wire_d0_23;
	wire [WIDTH-1:0] wire_d0_24;
	wire [WIDTH-1:0] wire_d0_25;
	wire [WIDTH-1:0] wire_d0_26;
	wire [WIDTH-1:0] wire_d0_27;
	wire [WIDTH-1:0] wire_d0_28;
	wire [WIDTH-1:0] wire_d0_29;
	wire [WIDTH-1:0] wire_d0_30;
	wire [WIDTH-1:0] wire_d0_31;
	wire [WIDTH-1:0] wire_d0_32;
	wire [WIDTH-1:0] wire_d0_33;
	wire [WIDTH-1:0] wire_d0_34;
	wire [WIDTH-1:0] wire_d0_35;
	wire [WIDTH-1:0] wire_d1_0;
	wire [WIDTH-1:0] wire_d1_1;
	wire [WIDTH-1:0] wire_d1_2;
	wire [WIDTH-1:0] wire_d1_3;
	wire [WIDTH-1:0] wire_d1_4;
	wire [WIDTH-1:0] wire_d1_5;
	wire [WIDTH-1:0] wire_d1_6;
	wire [WIDTH-1:0] wire_d1_7;
	wire [WIDTH-1:0] wire_d1_8;
	wire [WIDTH-1:0] wire_d1_9;
	wire [WIDTH-1:0] wire_d1_10;
	wire [WIDTH-1:0] wire_d1_11;
	wire [WIDTH-1:0] wire_d1_12;
	wire [WIDTH-1:0] wire_d1_13;
	wire [WIDTH-1:0] wire_d1_14;
	wire [WIDTH-1:0] wire_d1_15;
	wire [WIDTH-1:0] wire_d1_16;
	wire [WIDTH-1:0] wire_d1_17;
	wire [WIDTH-1:0] wire_d1_18;
	wire [WIDTH-1:0] wire_d1_19;
	wire [WIDTH-1:0] wire_d1_20;
	wire [WIDTH-1:0] wire_d1_21;
	wire [WIDTH-1:0] wire_d1_22;
	wire [WIDTH-1:0] wire_d1_23;
	wire [WIDTH-1:0] wire_d1_24;
	wire [WIDTH-1:0] wire_d1_25;
	wire [WIDTH-1:0] wire_d1_26;
	wire [WIDTH-1:0] wire_d1_27;
	wire [WIDTH-1:0] wire_d1_28;
	wire [WIDTH-1:0] wire_d1_29;
	wire [WIDTH-1:0] wire_d1_30;
	wire [WIDTH-1:0] wire_d1_31;
	wire [WIDTH-1:0] wire_d1_32;
	wire [WIDTH-1:0] wire_d1_33;
	wire [WIDTH-1:0] wire_d1_34;
	wire [WIDTH-1:0] wire_d1_35;
	wire [WIDTH-1:0] wire_d2_0;
	wire [WIDTH-1:0] wire_d2_1;
	wire [WIDTH-1:0] wire_d2_2;
	wire [WIDTH-1:0] wire_d2_3;
	wire [WIDTH-1:0] wire_d2_4;
	wire [WIDTH-1:0] wire_d2_5;
	wire [WIDTH-1:0] wire_d2_6;
	wire [WIDTH-1:0] wire_d2_7;
	wire [WIDTH-1:0] wire_d2_8;
	wire [WIDTH-1:0] wire_d2_9;
	wire [WIDTH-1:0] wire_d2_10;
	wire [WIDTH-1:0] wire_d2_11;
	wire [WIDTH-1:0] wire_d2_12;
	wire [WIDTH-1:0] wire_d2_13;
	wire [WIDTH-1:0] wire_d2_14;
	wire [WIDTH-1:0] wire_d2_15;
	wire [WIDTH-1:0] wire_d2_16;
	wire [WIDTH-1:0] wire_d2_17;
	wire [WIDTH-1:0] wire_d2_18;
	wire [WIDTH-1:0] wire_d2_19;
	wire [WIDTH-1:0] wire_d2_20;
	wire [WIDTH-1:0] wire_d2_21;
	wire [WIDTH-1:0] wire_d2_22;
	wire [WIDTH-1:0] wire_d2_23;
	wire [WIDTH-1:0] wire_d2_24;
	wire [WIDTH-1:0] wire_d2_25;
	wire [WIDTH-1:0] wire_d2_26;
	wire [WIDTH-1:0] wire_d2_27;
	wire [WIDTH-1:0] wire_d2_28;
	wire [WIDTH-1:0] wire_d2_29;
	wire [WIDTH-1:0] wire_d2_30;
	wire [WIDTH-1:0] wire_d2_31;
	wire [WIDTH-1:0] wire_d2_32;
	wire [WIDTH-1:0] wire_d2_33;
	wire [WIDTH-1:0] wire_d2_34;
	wire [WIDTH-1:0] wire_d2_35;
	wire [WIDTH-1:0] wire_d3_0;
	wire [WIDTH-1:0] wire_d3_1;
	wire [WIDTH-1:0] wire_d3_2;
	wire [WIDTH-1:0] wire_d3_3;
	wire [WIDTH-1:0] wire_d3_4;
	wire [WIDTH-1:0] wire_d3_5;
	wire [WIDTH-1:0] wire_d3_6;
	wire [WIDTH-1:0] wire_d3_7;
	wire [WIDTH-1:0] wire_d3_8;
	wire [WIDTH-1:0] wire_d3_9;
	wire [WIDTH-1:0] wire_d3_10;
	wire [WIDTH-1:0] wire_d3_11;
	wire [WIDTH-1:0] wire_d3_12;
	wire [WIDTH-1:0] wire_d3_13;
	wire [WIDTH-1:0] wire_d3_14;
	wire [WIDTH-1:0] wire_d3_15;
	wire [WIDTH-1:0] wire_d3_16;
	wire [WIDTH-1:0] wire_d3_17;
	wire [WIDTH-1:0] wire_d3_18;
	wire [WIDTH-1:0] wire_d3_19;
	wire [WIDTH-1:0] wire_d3_20;
	wire [WIDTH-1:0] wire_d3_21;
	wire [WIDTH-1:0] wire_d3_22;
	wire [WIDTH-1:0] wire_d3_23;
	wire [WIDTH-1:0] wire_d3_24;
	wire [WIDTH-1:0] wire_d3_25;
	wire [WIDTH-1:0] wire_d3_26;
	wire [WIDTH-1:0] wire_d3_27;
	wire [WIDTH-1:0] wire_d3_28;
	wire [WIDTH-1:0] wire_d3_29;
	wire [WIDTH-1:0] wire_d3_30;
	wire [WIDTH-1:0] wire_d3_31;
	wire [WIDTH-1:0] wire_d3_32;
	wire [WIDTH-1:0] wire_d3_33;
	wire [WIDTH-1:0] wire_d3_34;
	wire [WIDTH-1:0] wire_d3_35;
	wire [WIDTH-1:0] wire_d4_0;
	wire [WIDTH-1:0] wire_d4_1;
	wire [WIDTH-1:0] wire_d4_2;
	wire [WIDTH-1:0] wire_d4_3;
	wire [WIDTH-1:0] wire_d4_4;
	wire [WIDTH-1:0] wire_d4_5;
	wire [WIDTH-1:0] wire_d4_6;
	wire [WIDTH-1:0] wire_d4_7;
	wire [WIDTH-1:0] wire_d4_8;
	wire [WIDTH-1:0] wire_d4_9;
	wire [WIDTH-1:0] wire_d4_10;
	wire [WIDTH-1:0] wire_d4_11;
	wire [WIDTH-1:0] wire_d4_12;
	wire [WIDTH-1:0] wire_d4_13;
	wire [WIDTH-1:0] wire_d4_14;
	wire [WIDTH-1:0] wire_d4_15;
	wire [WIDTH-1:0] wire_d4_16;
	wire [WIDTH-1:0] wire_d4_17;
	wire [WIDTH-1:0] wire_d4_18;
	wire [WIDTH-1:0] wire_d4_19;
	wire [WIDTH-1:0] wire_d4_20;
	wire [WIDTH-1:0] wire_d4_21;
	wire [WIDTH-1:0] wire_d4_22;
	wire [WIDTH-1:0] wire_d4_23;
	wire [WIDTH-1:0] wire_d4_24;
	wire [WIDTH-1:0] wire_d4_25;
	wire [WIDTH-1:0] wire_d4_26;
	wire [WIDTH-1:0] wire_d4_27;
	wire [WIDTH-1:0] wire_d4_28;
	wire [WIDTH-1:0] wire_d4_29;
	wire [WIDTH-1:0] wire_d4_30;
	wire [WIDTH-1:0] wire_d4_31;
	wire [WIDTH-1:0] wire_d4_32;
	wire [WIDTH-1:0] wire_d4_33;
	wire [WIDTH-1:0] wire_d4_34;
	wire [WIDTH-1:0] wire_d4_35;
	wire [WIDTH-1:0] wire_d5_0;
	wire [WIDTH-1:0] wire_d5_1;
	wire [WIDTH-1:0] wire_d5_2;
	wire [WIDTH-1:0] wire_d5_3;
	wire [WIDTH-1:0] wire_d5_4;
	wire [WIDTH-1:0] wire_d5_5;
	wire [WIDTH-1:0] wire_d5_6;
	wire [WIDTH-1:0] wire_d5_7;
	wire [WIDTH-1:0] wire_d5_8;
	wire [WIDTH-1:0] wire_d5_9;
	wire [WIDTH-1:0] wire_d5_10;
	wire [WIDTH-1:0] wire_d5_11;
	wire [WIDTH-1:0] wire_d5_12;
	wire [WIDTH-1:0] wire_d5_13;
	wire [WIDTH-1:0] wire_d5_14;
	wire [WIDTH-1:0] wire_d5_15;
	wire [WIDTH-1:0] wire_d5_16;
	wire [WIDTH-1:0] wire_d5_17;
	wire [WIDTH-1:0] wire_d5_18;
	wire [WIDTH-1:0] wire_d5_19;
	wire [WIDTH-1:0] wire_d5_20;
	wire [WIDTH-1:0] wire_d5_21;
	wire [WIDTH-1:0] wire_d5_22;
	wire [WIDTH-1:0] wire_d5_23;
	wire [WIDTH-1:0] wire_d5_24;
	wire [WIDTH-1:0] wire_d5_25;
	wire [WIDTH-1:0] wire_d5_26;
	wire [WIDTH-1:0] wire_d5_27;
	wire [WIDTH-1:0] wire_d5_28;
	wire [WIDTH-1:0] wire_d5_29;
	wire [WIDTH-1:0] wire_d5_30;
	wire [WIDTH-1:0] wire_d5_31;
	wire [WIDTH-1:0] wire_d5_32;
	wire [WIDTH-1:0] wire_d5_33;
	wire [WIDTH-1:0] wire_d5_34;
	wire [WIDTH-1:0] wire_d5_35;
	wire [WIDTH-1:0] wire_d6_0;
	wire [WIDTH-1:0] wire_d6_1;
	wire [WIDTH-1:0] wire_d6_2;
	wire [WIDTH-1:0] wire_d6_3;
	wire [WIDTH-1:0] wire_d6_4;
	wire [WIDTH-1:0] wire_d6_5;
	wire [WIDTH-1:0] wire_d6_6;
	wire [WIDTH-1:0] wire_d6_7;
	wire [WIDTH-1:0] wire_d6_8;
	wire [WIDTH-1:0] wire_d6_9;
	wire [WIDTH-1:0] wire_d6_10;
	wire [WIDTH-1:0] wire_d6_11;
	wire [WIDTH-1:0] wire_d6_12;
	wire [WIDTH-1:0] wire_d6_13;
	wire [WIDTH-1:0] wire_d6_14;
	wire [WIDTH-1:0] wire_d6_15;
	wire [WIDTH-1:0] wire_d6_16;
	wire [WIDTH-1:0] wire_d6_17;
	wire [WIDTH-1:0] wire_d6_18;
	wire [WIDTH-1:0] wire_d6_19;
	wire [WIDTH-1:0] wire_d6_20;
	wire [WIDTH-1:0] wire_d6_21;
	wire [WIDTH-1:0] wire_d6_22;
	wire [WIDTH-1:0] wire_d6_23;
	wire [WIDTH-1:0] wire_d6_24;
	wire [WIDTH-1:0] wire_d6_25;
	wire [WIDTH-1:0] wire_d6_26;
	wire [WIDTH-1:0] wire_d6_27;
	wire [WIDTH-1:0] wire_d6_28;
	wire [WIDTH-1:0] wire_d6_29;
	wire [WIDTH-1:0] wire_d6_30;
	wire [WIDTH-1:0] wire_d6_31;
	wire [WIDTH-1:0] wire_d6_32;
	wire [WIDTH-1:0] wire_d6_33;
	wire [WIDTH-1:0] wire_d6_34;
	wire [WIDTH-1:0] wire_d6_35;
	wire [WIDTH-1:0] wire_d7_0;
	wire [WIDTH-1:0] wire_d7_1;
	wire [WIDTH-1:0] wire_d7_2;
	wire [WIDTH-1:0] wire_d7_3;
	wire [WIDTH-1:0] wire_d7_4;
	wire [WIDTH-1:0] wire_d7_5;
	wire [WIDTH-1:0] wire_d7_6;
	wire [WIDTH-1:0] wire_d7_7;
	wire [WIDTH-1:0] wire_d7_8;
	wire [WIDTH-1:0] wire_d7_9;
	wire [WIDTH-1:0] wire_d7_10;
	wire [WIDTH-1:0] wire_d7_11;
	wire [WIDTH-1:0] wire_d7_12;
	wire [WIDTH-1:0] wire_d7_13;
	wire [WIDTH-1:0] wire_d7_14;
	wire [WIDTH-1:0] wire_d7_15;
	wire [WIDTH-1:0] wire_d7_16;
	wire [WIDTH-1:0] wire_d7_17;
	wire [WIDTH-1:0] wire_d7_18;
	wire [WIDTH-1:0] wire_d7_19;
	wire [WIDTH-1:0] wire_d7_20;
	wire [WIDTH-1:0] wire_d7_21;
	wire [WIDTH-1:0] wire_d7_22;
	wire [WIDTH-1:0] wire_d7_23;
	wire [WIDTH-1:0] wire_d7_24;
	wire [WIDTH-1:0] wire_d7_25;
	wire [WIDTH-1:0] wire_d7_26;
	wire [WIDTH-1:0] wire_d7_27;
	wire [WIDTH-1:0] wire_d7_28;
	wire [WIDTH-1:0] wire_d7_29;
	wire [WIDTH-1:0] wire_d7_30;
	wire [WIDTH-1:0] wire_d7_31;
	wire [WIDTH-1:0] wire_d7_32;
	wire [WIDTH-1:0] wire_d7_33;
	wire [WIDTH-1:0] wire_d7_34;
	wire [WIDTH-1:0] wire_d7_35;
	wire [WIDTH-1:0] wire_d8_0;
	wire [WIDTH-1:0] wire_d8_1;
	wire [WIDTH-1:0] wire_d8_2;
	wire [WIDTH-1:0] wire_d8_3;
	wire [WIDTH-1:0] wire_d8_4;
	wire [WIDTH-1:0] wire_d8_5;
	wire [WIDTH-1:0] wire_d8_6;
	wire [WIDTH-1:0] wire_d8_7;
	wire [WIDTH-1:0] wire_d8_8;
	wire [WIDTH-1:0] wire_d8_9;
	wire [WIDTH-1:0] wire_d8_10;
	wire [WIDTH-1:0] wire_d8_11;
	wire [WIDTH-1:0] wire_d8_12;
	wire [WIDTH-1:0] wire_d8_13;
	wire [WIDTH-1:0] wire_d8_14;
	wire [WIDTH-1:0] wire_d8_15;
	wire [WIDTH-1:0] wire_d8_16;
	wire [WIDTH-1:0] wire_d8_17;
	wire [WIDTH-1:0] wire_d8_18;
	wire [WIDTH-1:0] wire_d8_19;
	wire [WIDTH-1:0] wire_d8_20;
	wire [WIDTH-1:0] wire_d8_21;
	wire [WIDTH-1:0] wire_d8_22;
	wire [WIDTH-1:0] wire_d8_23;
	wire [WIDTH-1:0] wire_d8_24;
	wire [WIDTH-1:0] wire_d8_25;
	wire [WIDTH-1:0] wire_d8_26;
	wire [WIDTH-1:0] wire_d8_27;
	wire [WIDTH-1:0] wire_d8_28;
	wire [WIDTH-1:0] wire_d8_29;
	wire [WIDTH-1:0] wire_d8_30;
	wire [WIDTH-1:0] wire_d8_31;
	wire [WIDTH-1:0] wire_d8_32;
	wire [WIDTH-1:0] wire_d8_33;
	wire [WIDTH-1:0] wire_d8_34;
	wire [WIDTH-1:0] wire_d8_35;
	wire [WIDTH-1:0] wire_d9_0;
	wire [WIDTH-1:0] wire_d9_1;
	wire [WIDTH-1:0] wire_d9_2;
	wire [WIDTH-1:0] wire_d9_3;
	wire [WIDTH-1:0] wire_d9_4;
	wire [WIDTH-1:0] wire_d9_5;
	wire [WIDTH-1:0] wire_d9_6;
	wire [WIDTH-1:0] wire_d9_7;
	wire [WIDTH-1:0] wire_d9_8;
	wire [WIDTH-1:0] wire_d9_9;
	wire [WIDTH-1:0] wire_d9_10;
	wire [WIDTH-1:0] wire_d9_11;
	wire [WIDTH-1:0] wire_d9_12;
	wire [WIDTH-1:0] wire_d9_13;
	wire [WIDTH-1:0] wire_d9_14;
	wire [WIDTH-1:0] wire_d9_15;
	wire [WIDTH-1:0] wire_d9_16;
	wire [WIDTH-1:0] wire_d9_17;
	wire [WIDTH-1:0] wire_d9_18;
	wire [WIDTH-1:0] wire_d9_19;
	wire [WIDTH-1:0] wire_d9_20;
	wire [WIDTH-1:0] wire_d9_21;
	wire [WIDTH-1:0] wire_d9_22;
	wire [WIDTH-1:0] wire_d9_23;
	wire [WIDTH-1:0] wire_d9_24;
	wire [WIDTH-1:0] wire_d9_25;
	wire [WIDTH-1:0] wire_d9_26;
	wire [WIDTH-1:0] wire_d9_27;
	wire [WIDTH-1:0] wire_d9_28;
	wire [WIDTH-1:0] wire_d9_29;
	wire [WIDTH-1:0] wire_d9_30;
	wire [WIDTH-1:0] wire_d9_31;
	wire [WIDTH-1:0] wire_d9_32;
	wire [WIDTH-1:0] wire_d9_33;
	wire [WIDTH-1:0] wire_d9_34;
	wire [WIDTH-1:0] wire_d9_35;
	wire [WIDTH-1:0] wire_d10_0;
	wire [WIDTH-1:0] wire_d10_1;
	wire [WIDTH-1:0] wire_d10_2;
	wire [WIDTH-1:0] wire_d10_3;
	wire [WIDTH-1:0] wire_d10_4;
	wire [WIDTH-1:0] wire_d10_5;
	wire [WIDTH-1:0] wire_d10_6;
	wire [WIDTH-1:0] wire_d10_7;
	wire [WIDTH-1:0] wire_d10_8;
	wire [WIDTH-1:0] wire_d10_9;
	wire [WIDTH-1:0] wire_d10_10;
	wire [WIDTH-1:0] wire_d10_11;
	wire [WIDTH-1:0] wire_d10_12;
	wire [WIDTH-1:0] wire_d10_13;
	wire [WIDTH-1:0] wire_d10_14;
	wire [WIDTH-1:0] wire_d10_15;
	wire [WIDTH-1:0] wire_d10_16;
	wire [WIDTH-1:0] wire_d10_17;
	wire [WIDTH-1:0] wire_d10_18;
	wire [WIDTH-1:0] wire_d10_19;
	wire [WIDTH-1:0] wire_d10_20;
	wire [WIDTH-1:0] wire_d10_21;
	wire [WIDTH-1:0] wire_d10_22;
	wire [WIDTH-1:0] wire_d10_23;
	wire [WIDTH-1:0] wire_d10_24;
	wire [WIDTH-1:0] wire_d10_25;
	wire [WIDTH-1:0] wire_d10_26;
	wire [WIDTH-1:0] wire_d10_27;
	wire [WIDTH-1:0] wire_d10_28;
	wire [WIDTH-1:0] wire_d10_29;
	wire [WIDTH-1:0] wire_d10_30;
	wire [WIDTH-1:0] wire_d10_31;
	wire [WIDTH-1:0] wire_d10_32;
	wire [WIDTH-1:0] wire_d10_33;
	wire [WIDTH-1:0] wire_d10_34;
	wire [WIDTH-1:0] wire_d10_35;
	wire [WIDTH-1:0] wire_d11_0;
	wire [WIDTH-1:0] wire_d11_1;
	wire [WIDTH-1:0] wire_d11_2;
	wire [WIDTH-1:0] wire_d11_3;
	wire [WIDTH-1:0] wire_d11_4;
	wire [WIDTH-1:0] wire_d11_5;
	wire [WIDTH-1:0] wire_d11_6;
	wire [WIDTH-1:0] wire_d11_7;
	wire [WIDTH-1:0] wire_d11_8;
	wire [WIDTH-1:0] wire_d11_9;
	wire [WIDTH-1:0] wire_d11_10;
	wire [WIDTH-1:0] wire_d11_11;
	wire [WIDTH-1:0] wire_d11_12;
	wire [WIDTH-1:0] wire_d11_13;
	wire [WIDTH-1:0] wire_d11_14;
	wire [WIDTH-1:0] wire_d11_15;
	wire [WIDTH-1:0] wire_d11_16;
	wire [WIDTH-1:0] wire_d11_17;
	wire [WIDTH-1:0] wire_d11_18;
	wire [WIDTH-1:0] wire_d11_19;
	wire [WIDTH-1:0] wire_d11_20;
	wire [WIDTH-1:0] wire_d11_21;
	wire [WIDTH-1:0] wire_d11_22;
	wire [WIDTH-1:0] wire_d11_23;
	wire [WIDTH-1:0] wire_d11_24;
	wire [WIDTH-1:0] wire_d11_25;
	wire [WIDTH-1:0] wire_d11_26;
	wire [WIDTH-1:0] wire_d11_27;
	wire [WIDTH-1:0] wire_d11_28;
	wire [WIDTH-1:0] wire_d11_29;
	wire [WIDTH-1:0] wire_d11_30;
	wire [WIDTH-1:0] wire_d11_31;
	wire [WIDTH-1:0] wire_d11_32;
	wire [WIDTH-1:0] wire_d11_33;
	wire [WIDTH-1:0] wire_d11_34;
	wire [WIDTH-1:0] wire_d11_35;
	wire [WIDTH-1:0] wire_d12_0;
	wire [WIDTH-1:0] wire_d12_1;
	wire [WIDTH-1:0] wire_d12_2;
	wire [WIDTH-1:0] wire_d12_3;
	wire [WIDTH-1:0] wire_d12_4;
	wire [WIDTH-1:0] wire_d12_5;
	wire [WIDTH-1:0] wire_d12_6;
	wire [WIDTH-1:0] wire_d12_7;
	wire [WIDTH-1:0] wire_d12_8;
	wire [WIDTH-1:0] wire_d12_9;
	wire [WIDTH-1:0] wire_d12_10;
	wire [WIDTH-1:0] wire_d12_11;
	wire [WIDTH-1:0] wire_d12_12;
	wire [WIDTH-1:0] wire_d12_13;
	wire [WIDTH-1:0] wire_d12_14;
	wire [WIDTH-1:0] wire_d12_15;
	wire [WIDTH-1:0] wire_d12_16;
	wire [WIDTH-1:0] wire_d12_17;
	wire [WIDTH-1:0] wire_d12_18;
	wire [WIDTH-1:0] wire_d12_19;
	wire [WIDTH-1:0] wire_d12_20;
	wire [WIDTH-1:0] wire_d12_21;
	wire [WIDTH-1:0] wire_d12_22;
	wire [WIDTH-1:0] wire_d12_23;
	wire [WIDTH-1:0] wire_d12_24;
	wire [WIDTH-1:0] wire_d12_25;
	wire [WIDTH-1:0] wire_d12_26;
	wire [WIDTH-1:0] wire_d12_27;
	wire [WIDTH-1:0] wire_d12_28;
	wire [WIDTH-1:0] wire_d12_29;
	wire [WIDTH-1:0] wire_d12_30;
	wire [WIDTH-1:0] wire_d12_31;
	wire [WIDTH-1:0] wire_d12_32;
	wire [WIDTH-1:0] wire_d12_33;
	wire [WIDTH-1:0] wire_d12_34;
	wire [WIDTH-1:0] wire_d12_35;
	wire [WIDTH-1:0] wire_d13_0;
	wire [WIDTH-1:0] wire_d13_1;
	wire [WIDTH-1:0] wire_d13_2;
	wire [WIDTH-1:0] wire_d13_3;
	wire [WIDTH-1:0] wire_d13_4;
	wire [WIDTH-1:0] wire_d13_5;
	wire [WIDTH-1:0] wire_d13_6;
	wire [WIDTH-1:0] wire_d13_7;
	wire [WIDTH-1:0] wire_d13_8;
	wire [WIDTH-1:0] wire_d13_9;
	wire [WIDTH-1:0] wire_d13_10;
	wire [WIDTH-1:0] wire_d13_11;
	wire [WIDTH-1:0] wire_d13_12;
	wire [WIDTH-1:0] wire_d13_13;
	wire [WIDTH-1:0] wire_d13_14;
	wire [WIDTH-1:0] wire_d13_15;
	wire [WIDTH-1:0] wire_d13_16;
	wire [WIDTH-1:0] wire_d13_17;
	wire [WIDTH-1:0] wire_d13_18;
	wire [WIDTH-1:0] wire_d13_19;
	wire [WIDTH-1:0] wire_d13_20;
	wire [WIDTH-1:0] wire_d13_21;
	wire [WIDTH-1:0] wire_d13_22;
	wire [WIDTH-1:0] wire_d13_23;
	wire [WIDTH-1:0] wire_d13_24;
	wire [WIDTH-1:0] wire_d13_25;
	wire [WIDTH-1:0] wire_d13_26;
	wire [WIDTH-1:0] wire_d13_27;
	wire [WIDTH-1:0] wire_d13_28;
	wire [WIDTH-1:0] wire_d13_29;
	wire [WIDTH-1:0] wire_d13_30;
	wire [WIDTH-1:0] wire_d13_31;
	wire [WIDTH-1:0] wire_d13_32;
	wire [WIDTH-1:0] wire_d13_33;
	wire [WIDTH-1:0] wire_d13_34;
	wire [WIDTH-1:0] wire_d13_35;
	wire [WIDTH-1:0] wire_d14_0;
	wire [WIDTH-1:0] wire_d14_1;
	wire [WIDTH-1:0] wire_d14_2;
	wire [WIDTH-1:0] wire_d14_3;
	wire [WIDTH-1:0] wire_d14_4;
	wire [WIDTH-1:0] wire_d14_5;
	wire [WIDTH-1:0] wire_d14_6;
	wire [WIDTH-1:0] wire_d14_7;
	wire [WIDTH-1:0] wire_d14_8;
	wire [WIDTH-1:0] wire_d14_9;
	wire [WIDTH-1:0] wire_d14_10;
	wire [WIDTH-1:0] wire_d14_11;
	wire [WIDTH-1:0] wire_d14_12;
	wire [WIDTH-1:0] wire_d14_13;
	wire [WIDTH-1:0] wire_d14_14;
	wire [WIDTH-1:0] wire_d14_15;
	wire [WIDTH-1:0] wire_d14_16;
	wire [WIDTH-1:0] wire_d14_17;
	wire [WIDTH-1:0] wire_d14_18;
	wire [WIDTH-1:0] wire_d14_19;
	wire [WIDTH-1:0] wire_d14_20;
	wire [WIDTH-1:0] wire_d14_21;
	wire [WIDTH-1:0] wire_d14_22;
	wire [WIDTH-1:0] wire_d14_23;
	wire [WIDTH-1:0] wire_d14_24;
	wire [WIDTH-1:0] wire_d14_25;
	wire [WIDTH-1:0] wire_d14_26;
	wire [WIDTH-1:0] wire_d14_27;
	wire [WIDTH-1:0] wire_d14_28;
	wire [WIDTH-1:0] wire_d14_29;
	wire [WIDTH-1:0] wire_d14_30;
	wire [WIDTH-1:0] wire_d14_31;
	wire [WIDTH-1:0] wire_d14_32;
	wire [WIDTH-1:0] wire_d14_33;
	wire [WIDTH-1:0] wire_d14_34;
	wire [WIDTH-1:0] wire_d14_35;
	wire [WIDTH-1:0] wire_d15_0;
	wire [WIDTH-1:0] wire_d15_1;
	wire [WIDTH-1:0] wire_d15_2;
	wire [WIDTH-1:0] wire_d15_3;
	wire [WIDTH-1:0] wire_d15_4;
	wire [WIDTH-1:0] wire_d15_5;
	wire [WIDTH-1:0] wire_d15_6;
	wire [WIDTH-1:0] wire_d15_7;
	wire [WIDTH-1:0] wire_d15_8;
	wire [WIDTH-1:0] wire_d15_9;
	wire [WIDTH-1:0] wire_d15_10;
	wire [WIDTH-1:0] wire_d15_11;
	wire [WIDTH-1:0] wire_d15_12;
	wire [WIDTH-1:0] wire_d15_13;
	wire [WIDTH-1:0] wire_d15_14;
	wire [WIDTH-1:0] wire_d15_15;
	wire [WIDTH-1:0] wire_d15_16;
	wire [WIDTH-1:0] wire_d15_17;
	wire [WIDTH-1:0] wire_d15_18;
	wire [WIDTH-1:0] wire_d15_19;
	wire [WIDTH-1:0] wire_d15_20;
	wire [WIDTH-1:0] wire_d15_21;
	wire [WIDTH-1:0] wire_d15_22;
	wire [WIDTH-1:0] wire_d15_23;
	wire [WIDTH-1:0] wire_d15_24;
	wire [WIDTH-1:0] wire_d15_25;
	wire [WIDTH-1:0] wire_d15_26;
	wire [WIDTH-1:0] wire_d15_27;
	wire [WIDTH-1:0] wire_d15_28;
	wire [WIDTH-1:0] wire_d15_29;
	wire [WIDTH-1:0] wire_d15_30;
	wire [WIDTH-1:0] wire_d15_31;
	wire [WIDTH-1:0] wire_d15_32;
	wire [WIDTH-1:0] wire_d15_33;
	wire [WIDTH-1:0] wire_d15_34;
	wire [WIDTH-1:0] wire_d15_35;
	wire [WIDTH-1:0] wire_d16_0;
	wire [WIDTH-1:0] wire_d16_1;
	wire [WIDTH-1:0] wire_d16_2;
	wire [WIDTH-1:0] wire_d16_3;
	wire [WIDTH-1:0] wire_d16_4;
	wire [WIDTH-1:0] wire_d16_5;
	wire [WIDTH-1:0] wire_d16_6;
	wire [WIDTH-1:0] wire_d16_7;
	wire [WIDTH-1:0] wire_d16_8;
	wire [WIDTH-1:0] wire_d16_9;
	wire [WIDTH-1:0] wire_d16_10;
	wire [WIDTH-1:0] wire_d16_11;
	wire [WIDTH-1:0] wire_d16_12;
	wire [WIDTH-1:0] wire_d16_13;
	wire [WIDTH-1:0] wire_d16_14;
	wire [WIDTH-1:0] wire_d16_15;
	wire [WIDTH-1:0] wire_d16_16;
	wire [WIDTH-1:0] wire_d16_17;
	wire [WIDTH-1:0] wire_d16_18;
	wire [WIDTH-1:0] wire_d16_19;
	wire [WIDTH-1:0] wire_d16_20;
	wire [WIDTH-1:0] wire_d16_21;
	wire [WIDTH-1:0] wire_d16_22;
	wire [WIDTH-1:0] wire_d16_23;
	wire [WIDTH-1:0] wire_d16_24;
	wire [WIDTH-1:0] wire_d16_25;
	wire [WIDTH-1:0] wire_d16_26;
	wire [WIDTH-1:0] wire_d16_27;
	wire [WIDTH-1:0] wire_d16_28;
	wire [WIDTH-1:0] wire_d16_29;
	wire [WIDTH-1:0] wire_d16_30;
	wire [WIDTH-1:0] wire_d16_31;
	wire [WIDTH-1:0] wire_d16_32;
	wire [WIDTH-1:0] wire_d16_33;
	wire [WIDTH-1:0] wire_d16_34;
	wire [WIDTH-1:0] wire_d16_35;
	wire [WIDTH-1:0] wire_d17_0;
	wire [WIDTH-1:0] wire_d17_1;
	wire [WIDTH-1:0] wire_d17_2;
	wire [WIDTH-1:0] wire_d17_3;
	wire [WIDTH-1:0] wire_d17_4;
	wire [WIDTH-1:0] wire_d17_5;
	wire [WIDTH-1:0] wire_d17_6;
	wire [WIDTH-1:0] wire_d17_7;
	wire [WIDTH-1:0] wire_d17_8;
	wire [WIDTH-1:0] wire_d17_9;
	wire [WIDTH-1:0] wire_d17_10;
	wire [WIDTH-1:0] wire_d17_11;
	wire [WIDTH-1:0] wire_d17_12;
	wire [WIDTH-1:0] wire_d17_13;
	wire [WIDTH-1:0] wire_d17_14;
	wire [WIDTH-1:0] wire_d17_15;
	wire [WIDTH-1:0] wire_d17_16;
	wire [WIDTH-1:0] wire_d17_17;
	wire [WIDTH-1:0] wire_d17_18;
	wire [WIDTH-1:0] wire_d17_19;
	wire [WIDTH-1:0] wire_d17_20;
	wire [WIDTH-1:0] wire_d17_21;
	wire [WIDTH-1:0] wire_d17_22;
	wire [WIDTH-1:0] wire_d17_23;
	wire [WIDTH-1:0] wire_d17_24;
	wire [WIDTH-1:0] wire_d17_25;
	wire [WIDTH-1:0] wire_d17_26;
	wire [WIDTH-1:0] wire_d17_27;
	wire [WIDTH-1:0] wire_d17_28;
	wire [WIDTH-1:0] wire_d17_29;
	wire [WIDTH-1:0] wire_d17_30;
	wire [WIDTH-1:0] wire_d17_31;
	wire [WIDTH-1:0] wire_d17_32;
	wire [WIDTH-1:0] wire_d17_33;
	wire [WIDTH-1:0] wire_d17_34;
	wire [WIDTH-1:0] wire_d17_35;
	wire [WIDTH-1:0] wire_d18_0;
	wire [WIDTH-1:0] wire_d18_1;
	wire [WIDTH-1:0] wire_d18_2;
	wire [WIDTH-1:0] wire_d18_3;
	wire [WIDTH-1:0] wire_d18_4;
	wire [WIDTH-1:0] wire_d18_5;
	wire [WIDTH-1:0] wire_d18_6;
	wire [WIDTH-1:0] wire_d18_7;
	wire [WIDTH-1:0] wire_d18_8;
	wire [WIDTH-1:0] wire_d18_9;
	wire [WIDTH-1:0] wire_d18_10;
	wire [WIDTH-1:0] wire_d18_11;
	wire [WIDTH-1:0] wire_d18_12;
	wire [WIDTH-1:0] wire_d18_13;
	wire [WIDTH-1:0] wire_d18_14;
	wire [WIDTH-1:0] wire_d18_15;
	wire [WIDTH-1:0] wire_d18_16;
	wire [WIDTH-1:0] wire_d18_17;
	wire [WIDTH-1:0] wire_d18_18;
	wire [WIDTH-1:0] wire_d18_19;
	wire [WIDTH-1:0] wire_d18_20;
	wire [WIDTH-1:0] wire_d18_21;
	wire [WIDTH-1:0] wire_d18_22;
	wire [WIDTH-1:0] wire_d18_23;
	wire [WIDTH-1:0] wire_d18_24;
	wire [WIDTH-1:0] wire_d18_25;
	wire [WIDTH-1:0] wire_d18_26;
	wire [WIDTH-1:0] wire_d18_27;
	wire [WIDTH-1:0] wire_d18_28;
	wire [WIDTH-1:0] wire_d18_29;
	wire [WIDTH-1:0] wire_d18_30;
	wire [WIDTH-1:0] wire_d18_31;
	wire [WIDTH-1:0] wire_d18_32;
	wire [WIDTH-1:0] wire_d18_33;
	wire [WIDTH-1:0] wire_d18_34;
	wire [WIDTH-1:0] wire_d18_35;
	wire [WIDTH-1:0] wire_d19_0;
	wire [WIDTH-1:0] wire_d19_1;
	wire [WIDTH-1:0] wire_d19_2;
	wire [WIDTH-1:0] wire_d19_3;
	wire [WIDTH-1:0] wire_d19_4;
	wire [WIDTH-1:0] wire_d19_5;
	wire [WIDTH-1:0] wire_d19_6;
	wire [WIDTH-1:0] wire_d19_7;
	wire [WIDTH-1:0] wire_d19_8;
	wire [WIDTH-1:0] wire_d19_9;
	wire [WIDTH-1:0] wire_d19_10;
	wire [WIDTH-1:0] wire_d19_11;
	wire [WIDTH-1:0] wire_d19_12;
	wire [WIDTH-1:0] wire_d19_13;
	wire [WIDTH-1:0] wire_d19_14;
	wire [WIDTH-1:0] wire_d19_15;
	wire [WIDTH-1:0] wire_d19_16;
	wire [WIDTH-1:0] wire_d19_17;
	wire [WIDTH-1:0] wire_d19_18;
	wire [WIDTH-1:0] wire_d19_19;
	wire [WIDTH-1:0] wire_d19_20;
	wire [WIDTH-1:0] wire_d19_21;
	wire [WIDTH-1:0] wire_d19_22;
	wire [WIDTH-1:0] wire_d19_23;
	wire [WIDTH-1:0] wire_d19_24;
	wire [WIDTH-1:0] wire_d19_25;
	wire [WIDTH-1:0] wire_d19_26;
	wire [WIDTH-1:0] wire_d19_27;
	wire [WIDTH-1:0] wire_d19_28;
	wire [WIDTH-1:0] wire_d19_29;
	wire [WIDTH-1:0] wire_d19_30;
	wire [WIDTH-1:0] wire_d19_31;
	wire [WIDTH-1:0] wire_d19_32;
	wire [WIDTH-1:0] wire_d19_33;
	wire [WIDTH-1:0] wire_d19_34;
	wire [WIDTH-1:0] wire_d19_35;
	wire [WIDTH-1:0] wire_d20_0;
	wire [WIDTH-1:0] wire_d20_1;
	wire [WIDTH-1:0] wire_d20_2;
	wire [WIDTH-1:0] wire_d20_3;
	wire [WIDTH-1:0] wire_d20_4;
	wire [WIDTH-1:0] wire_d20_5;
	wire [WIDTH-1:0] wire_d20_6;
	wire [WIDTH-1:0] wire_d20_7;
	wire [WIDTH-1:0] wire_d20_8;
	wire [WIDTH-1:0] wire_d20_9;
	wire [WIDTH-1:0] wire_d20_10;
	wire [WIDTH-1:0] wire_d20_11;
	wire [WIDTH-1:0] wire_d20_12;
	wire [WIDTH-1:0] wire_d20_13;
	wire [WIDTH-1:0] wire_d20_14;
	wire [WIDTH-1:0] wire_d20_15;
	wire [WIDTH-1:0] wire_d20_16;
	wire [WIDTH-1:0] wire_d20_17;
	wire [WIDTH-1:0] wire_d20_18;
	wire [WIDTH-1:0] wire_d20_19;
	wire [WIDTH-1:0] wire_d20_20;
	wire [WIDTH-1:0] wire_d20_21;
	wire [WIDTH-1:0] wire_d20_22;
	wire [WIDTH-1:0] wire_d20_23;
	wire [WIDTH-1:0] wire_d20_24;
	wire [WIDTH-1:0] wire_d20_25;
	wire [WIDTH-1:0] wire_d20_26;
	wire [WIDTH-1:0] wire_d20_27;
	wire [WIDTH-1:0] wire_d20_28;
	wire [WIDTH-1:0] wire_d20_29;
	wire [WIDTH-1:0] wire_d20_30;
	wire [WIDTH-1:0] wire_d20_31;
	wire [WIDTH-1:0] wire_d20_32;
	wire [WIDTH-1:0] wire_d20_33;
	wire [WIDTH-1:0] wire_d20_34;
	wire [WIDTH-1:0] wire_d20_35;
	wire [WIDTH-1:0] wire_d21_0;
	wire [WIDTH-1:0] wire_d21_1;
	wire [WIDTH-1:0] wire_d21_2;
	wire [WIDTH-1:0] wire_d21_3;
	wire [WIDTH-1:0] wire_d21_4;
	wire [WIDTH-1:0] wire_d21_5;
	wire [WIDTH-1:0] wire_d21_6;
	wire [WIDTH-1:0] wire_d21_7;
	wire [WIDTH-1:0] wire_d21_8;
	wire [WIDTH-1:0] wire_d21_9;
	wire [WIDTH-1:0] wire_d21_10;
	wire [WIDTH-1:0] wire_d21_11;
	wire [WIDTH-1:0] wire_d21_12;
	wire [WIDTH-1:0] wire_d21_13;
	wire [WIDTH-1:0] wire_d21_14;
	wire [WIDTH-1:0] wire_d21_15;
	wire [WIDTH-1:0] wire_d21_16;
	wire [WIDTH-1:0] wire_d21_17;
	wire [WIDTH-1:0] wire_d21_18;
	wire [WIDTH-1:0] wire_d21_19;
	wire [WIDTH-1:0] wire_d21_20;
	wire [WIDTH-1:0] wire_d21_21;
	wire [WIDTH-1:0] wire_d21_22;
	wire [WIDTH-1:0] wire_d21_23;
	wire [WIDTH-1:0] wire_d21_24;
	wire [WIDTH-1:0] wire_d21_25;
	wire [WIDTH-1:0] wire_d21_26;
	wire [WIDTH-1:0] wire_d21_27;
	wire [WIDTH-1:0] wire_d21_28;
	wire [WIDTH-1:0] wire_d21_29;
	wire [WIDTH-1:0] wire_d21_30;
	wire [WIDTH-1:0] wire_d21_31;
	wire [WIDTH-1:0] wire_d21_32;
	wire [WIDTH-1:0] wire_d21_33;
	wire [WIDTH-1:0] wire_d21_34;
	wire [WIDTH-1:0] wire_d21_35;
	wire [WIDTH-1:0] wire_d22_0;
	wire [WIDTH-1:0] wire_d22_1;
	wire [WIDTH-1:0] wire_d22_2;
	wire [WIDTH-1:0] wire_d22_3;
	wire [WIDTH-1:0] wire_d22_4;
	wire [WIDTH-1:0] wire_d22_5;
	wire [WIDTH-1:0] wire_d22_6;
	wire [WIDTH-1:0] wire_d22_7;
	wire [WIDTH-1:0] wire_d22_8;
	wire [WIDTH-1:0] wire_d22_9;
	wire [WIDTH-1:0] wire_d22_10;
	wire [WIDTH-1:0] wire_d22_11;
	wire [WIDTH-1:0] wire_d22_12;
	wire [WIDTH-1:0] wire_d22_13;
	wire [WIDTH-1:0] wire_d22_14;
	wire [WIDTH-1:0] wire_d22_15;
	wire [WIDTH-1:0] wire_d22_16;
	wire [WIDTH-1:0] wire_d22_17;
	wire [WIDTH-1:0] wire_d22_18;
	wire [WIDTH-1:0] wire_d22_19;
	wire [WIDTH-1:0] wire_d22_20;
	wire [WIDTH-1:0] wire_d22_21;
	wire [WIDTH-1:0] wire_d22_22;
	wire [WIDTH-1:0] wire_d22_23;
	wire [WIDTH-1:0] wire_d22_24;
	wire [WIDTH-1:0] wire_d22_25;
	wire [WIDTH-1:0] wire_d22_26;
	wire [WIDTH-1:0] wire_d22_27;
	wire [WIDTH-1:0] wire_d22_28;
	wire [WIDTH-1:0] wire_d22_29;
	wire [WIDTH-1:0] wire_d22_30;
	wire [WIDTH-1:0] wire_d22_31;
	wire [WIDTH-1:0] wire_d22_32;
	wire [WIDTH-1:0] wire_d22_33;
	wire [WIDTH-1:0] wire_d22_34;
	wire [WIDTH-1:0] wire_d22_35;
	wire [WIDTH-1:0] wire_d23_0;
	wire [WIDTH-1:0] wire_d23_1;
	wire [WIDTH-1:0] wire_d23_2;
	wire [WIDTH-1:0] wire_d23_3;
	wire [WIDTH-1:0] wire_d23_4;
	wire [WIDTH-1:0] wire_d23_5;
	wire [WIDTH-1:0] wire_d23_6;
	wire [WIDTH-1:0] wire_d23_7;
	wire [WIDTH-1:0] wire_d23_8;
	wire [WIDTH-1:0] wire_d23_9;
	wire [WIDTH-1:0] wire_d23_10;
	wire [WIDTH-1:0] wire_d23_11;
	wire [WIDTH-1:0] wire_d23_12;
	wire [WIDTH-1:0] wire_d23_13;
	wire [WIDTH-1:0] wire_d23_14;
	wire [WIDTH-1:0] wire_d23_15;
	wire [WIDTH-1:0] wire_d23_16;
	wire [WIDTH-1:0] wire_d23_17;
	wire [WIDTH-1:0] wire_d23_18;
	wire [WIDTH-1:0] wire_d23_19;
	wire [WIDTH-1:0] wire_d23_20;
	wire [WIDTH-1:0] wire_d23_21;
	wire [WIDTH-1:0] wire_d23_22;
	wire [WIDTH-1:0] wire_d23_23;
	wire [WIDTH-1:0] wire_d23_24;
	wire [WIDTH-1:0] wire_d23_25;
	wire [WIDTH-1:0] wire_d23_26;
	wire [WIDTH-1:0] wire_d23_27;
	wire [WIDTH-1:0] wire_d23_28;
	wire [WIDTH-1:0] wire_d23_29;
	wire [WIDTH-1:0] wire_d23_30;
	wire [WIDTH-1:0] wire_d23_31;
	wire [WIDTH-1:0] wire_d23_32;
	wire [WIDTH-1:0] wire_d23_33;
	wire [WIDTH-1:0] wire_d23_34;
	wire [WIDTH-1:0] wire_d23_35;
	wire [WIDTH-1:0] wire_d24_0;
	wire [WIDTH-1:0] wire_d24_1;
	wire [WIDTH-1:0] wire_d24_2;
	wire [WIDTH-1:0] wire_d24_3;
	wire [WIDTH-1:0] wire_d24_4;
	wire [WIDTH-1:0] wire_d24_5;
	wire [WIDTH-1:0] wire_d24_6;
	wire [WIDTH-1:0] wire_d24_7;
	wire [WIDTH-1:0] wire_d24_8;
	wire [WIDTH-1:0] wire_d24_9;
	wire [WIDTH-1:0] wire_d24_10;
	wire [WIDTH-1:0] wire_d24_11;
	wire [WIDTH-1:0] wire_d24_12;
	wire [WIDTH-1:0] wire_d24_13;
	wire [WIDTH-1:0] wire_d24_14;
	wire [WIDTH-1:0] wire_d24_15;
	wire [WIDTH-1:0] wire_d24_16;
	wire [WIDTH-1:0] wire_d24_17;
	wire [WIDTH-1:0] wire_d24_18;
	wire [WIDTH-1:0] wire_d24_19;
	wire [WIDTH-1:0] wire_d24_20;
	wire [WIDTH-1:0] wire_d24_21;
	wire [WIDTH-1:0] wire_d24_22;
	wire [WIDTH-1:0] wire_d24_23;
	wire [WIDTH-1:0] wire_d24_24;
	wire [WIDTH-1:0] wire_d24_25;
	wire [WIDTH-1:0] wire_d24_26;
	wire [WIDTH-1:0] wire_d24_27;
	wire [WIDTH-1:0] wire_d24_28;
	wire [WIDTH-1:0] wire_d24_29;
	wire [WIDTH-1:0] wire_d24_30;
	wire [WIDTH-1:0] wire_d24_31;
	wire [WIDTH-1:0] wire_d24_32;
	wire [WIDTH-1:0] wire_d24_33;
	wire [WIDTH-1:0] wire_d24_34;
	wire [WIDTH-1:0] wire_d24_35;
	wire [WIDTH-1:0] wire_d25_0;
	wire [WIDTH-1:0] wire_d25_1;
	wire [WIDTH-1:0] wire_d25_2;
	wire [WIDTH-1:0] wire_d25_3;
	wire [WIDTH-1:0] wire_d25_4;
	wire [WIDTH-1:0] wire_d25_5;
	wire [WIDTH-1:0] wire_d25_6;
	wire [WIDTH-1:0] wire_d25_7;
	wire [WIDTH-1:0] wire_d25_8;
	wire [WIDTH-1:0] wire_d25_9;
	wire [WIDTH-1:0] wire_d25_10;
	wire [WIDTH-1:0] wire_d25_11;
	wire [WIDTH-1:0] wire_d25_12;
	wire [WIDTH-1:0] wire_d25_13;
	wire [WIDTH-1:0] wire_d25_14;
	wire [WIDTH-1:0] wire_d25_15;
	wire [WIDTH-1:0] wire_d25_16;
	wire [WIDTH-1:0] wire_d25_17;
	wire [WIDTH-1:0] wire_d25_18;
	wire [WIDTH-1:0] wire_d25_19;
	wire [WIDTH-1:0] wire_d25_20;
	wire [WIDTH-1:0] wire_d25_21;
	wire [WIDTH-1:0] wire_d25_22;
	wire [WIDTH-1:0] wire_d25_23;
	wire [WIDTH-1:0] wire_d25_24;
	wire [WIDTH-1:0] wire_d25_25;
	wire [WIDTH-1:0] wire_d25_26;
	wire [WIDTH-1:0] wire_d25_27;
	wire [WIDTH-1:0] wire_d25_28;
	wire [WIDTH-1:0] wire_d25_29;
	wire [WIDTH-1:0] wire_d25_30;
	wire [WIDTH-1:0] wire_d25_31;
	wire [WIDTH-1:0] wire_d25_32;
	wire [WIDTH-1:0] wire_d25_33;
	wire [WIDTH-1:0] wire_d25_34;
	wire [WIDTH-1:0] wire_d25_35;
	wire [WIDTH-1:0] wire_d26_0;
	wire [WIDTH-1:0] wire_d26_1;
	wire [WIDTH-1:0] wire_d26_2;
	wire [WIDTH-1:0] wire_d26_3;
	wire [WIDTH-1:0] wire_d26_4;
	wire [WIDTH-1:0] wire_d26_5;
	wire [WIDTH-1:0] wire_d26_6;
	wire [WIDTH-1:0] wire_d26_7;
	wire [WIDTH-1:0] wire_d26_8;
	wire [WIDTH-1:0] wire_d26_9;
	wire [WIDTH-1:0] wire_d26_10;
	wire [WIDTH-1:0] wire_d26_11;
	wire [WIDTH-1:0] wire_d26_12;
	wire [WIDTH-1:0] wire_d26_13;
	wire [WIDTH-1:0] wire_d26_14;
	wire [WIDTH-1:0] wire_d26_15;
	wire [WIDTH-1:0] wire_d26_16;
	wire [WIDTH-1:0] wire_d26_17;
	wire [WIDTH-1:0] wire_d26_18;
	wire [WIDTH-1:0] wire_d26_19;
	wire [WIDTH-1:0] wire_d26_20;
	wire [WIDTH-1:0] wire_d26_21;
	wire [WIDTH-1:0] wire_d26_22;
	wire [WIDTH-1:0] wire_d26_23;
	wire [WIDTH-1:0] wire_d26_24;
	wire [WIDTH-1:0] wire_d26_25;
	wire [WIDTH-1:0] wire_d26_26;
	wire [WIDTH-1:0] wire_d26_27;
	wire [WIDTH-1:0] wire_d26_28;
	wire [WIDTH-1:0] wire_d26_29;
	wire [WIDTH-1:0] wire_d26_30;
	wire [WIDTH-1:0] wire_d26_31;
	wire [WIDTH-1:0] wire_d26_32;
	wire [WIDTH-1:0] wire_d26_33;
	wire [WIDTH-1:0] wire_d26_34;
	wire [WIDTH-1:0] wire_d26_35;
	wire [WIDTH-1:0] wire_d27_0;
	wire [WIDTH-1:0] wire_d27_1;
	wire [WIDTH-1:0] wire_d27_2;
	wire [WIDTH-1:0] wire_d27_3;
	wire [WIDTH-1:0] wire_d27_4;
	wire [WIDTH-1:0] wire_d27_5;
	wire [WIDTH-1:0] wire_d27_6;
	wire [WIDTH-1:0] wire_d27_7;
	wire [WIDTH-1:0] wire_d27_8;
	wire [WIDTH-1:0] wire_d27_9;
	wire [WIDTH-1:0] wire_d27_10;
	wire [WIDTH-1:0] wire_d27_11;
	wire [WIDTH-1:0] wire_d27_12;
	wire [WIDTH-1:0] wire_d27_13;
	wire [WIDTH-1:0] wire_d27_14;
	wire [WIDTH-1:0] wire_d27_15;
	wire [WIDTH-1:0] wire_d27_16;
	wire [WIDTH-1:0] wire_d27_17;
	wire [WIDTH-1:0] wire_d27_18;
	wire [WIDTH-1:0] wire_d27_19;
	wire [WIDTH-1:0] wire_d27_20;
	wire [WIDTH-1:0] wire_d27_21;
	wire [WIDTH-1:0] wire_d27_22;
	wire [WIDTH-1:0] wire_d27_23;
	wire [WIDTH-1:0] wire_d27_24;
	wire [WIDTH-1:0] wire_d27_25;
	wire [WIDTH-1:0] wire_d27_26;
	wire [WIDTH-1:0] wire_d27_27;
	wire [WIDTH-1:0] wire_d27_28;
	wire [WIDTH-1:0] wire_d27_29;
	wire [WIDTH-1:0] wire_d27_30;
	wire [WIDTH-1:0] wire_d27_31;
	wire [WIDTH-1:0] wire_d27_32;
	wire [WIDTH-1:0] wire_d27_33;
	wire [WIDTH-1:0] wire_d27_34;
	wire [WIDTH-1:0] wire_d27_35;
	wire [WIDTH-1:0] wire_d28_0;
	wire [WIDTH-1:0] wire_d28_1;
	wire [WIDTH-1:0] wire_d28_2;
	wire [WIDTH-1:0] wire_d28_3;
	wire [WIDTH-1:0] wire_d28_4;
	wire [WIDTH-1:0] wire_d28_5;
	wire [WIDTH-1:0] wire_d28_6;
	wire [WIDTH-1:0] wire_d28_7;
	wire [WIDTH-1:0] wire_d28_8;
	wire [WIDTH-1:0] wire_d28_9;
	wire [WIDTH-1:0] wire_d28_10;
	wire [WIDTH-1:0] wire_d28_11;
	wire [WIDTH-1:0] wire_d28_12;
	wire [WIDTH-1:0] wire_d28_13;
	wire [WIDTH-1:0] wire_d28_14;
	wire [WIDTH-1:0] wire_d28_15;
	wire [WIDTH-1:0] wire_d28_16;
	wire [WIDTH-1:0] wire_d28_17;
	wire [WIDTH-1:0] wire_d28_18;
	wire [WIDTH-1:0] wire_d28_19;
	wire [WIDTH-1:0] wire_d28_20;
	wire [WIDTH-1:0] wire_d28_21;
	wire [WIDTH-1:0] wire_d28_22;
	wire [WIDTH-1:0] wire_d28_23;
	wire [WIDTH-1:0] wire_d28_24;
	wire [WIDTH-1:0] wire_d28_25;
	wire [WIDTH-1:0] wire_d28_26;
	wire [WIDTH-1:0] wire_d28_27;
	wire [WIDTH-1:0] wire_d28_28;
	wire [WIDTH-1:0] wire_d28_29;
	wire [WIDTH-1:0] wire_d28_30;
	wire [WIDTH-1:0] wire_d28_31;
	wire [WIDTH-1:0] wire_d28_32;
	wire [WIDTH-1:0] wire_d28_33;
	wire [WIDTH-1:0] wire_d28_34;
	wire [WIDTH-1:0] wire_d28_35;
	wire [WIDTH-1:0] wire_d29_0;
	wire [WIDTH-1:0] wire_d29_1;
	wire [WIDTH-1:0] wire_d29_2;
	wire [WIDTH-1:0] wire_d29_3;
	wire [WIDTH-1:0] wire_d29_4;
	wire [WIDTH-1:0] wire_d29_5;
	wire [WIDTH-1:0] wire_d29_6;
	wire [WIDTH-1:0] wire_d29_7;
	wire [WIDTH-1:0] wire_d29_8;
	wire [WIDTH-1:0] wire_d29_9;
	wire [WIDTH-1:0] wire_d29_10;
	wire [WIDTH-1:0] wire_d29_11;
	wire [WIDTH-1:0] wire_d29_12;
	wire [WIDTH-1:0] wire_d29_13;
	wire [WIDTH-1:0] wire_d29_14;
	wire [WIDTH-1:0] wire_d29_15;
	wire [WIDTH-1:0] wire_d29_16;
	wire [WIDTH-1:0] wire_d29_17;
	wire [WIDTH-1:0] wire_d29_18;
	wire [WIDTH-1:0] wire_d29_19;
	wire [WIDTH-1:0] wire_d29_20;
	wire [WIDTH-1:0] wire_d29_21;
	wire [WIDTH-1:0] wire_d29_22;
	wire [WIDTH-1:0] wire_d29_23;
	wire [WIDTH-1:0] wire_d29_24;
	wire [WIDTH-1:0] wire_d29_25;
	wire [WIDTH-1:0] wire_d29_26;
	wire [WIDTH-1:0] wire_d29_27;
	wire [WIDTH-1:0] wire_d29_28;
	wire [WIDTH-1:0] wire_d29_29;
	wire [WIDTH-1:0] wire_d29_30;
	wire [WIDTH-1:0] wire_d29_31;
	wire [WIDTH-1:0] wire_d29_32;
	wire [WIDTH-1:0] wire_d29_33;
	wire [WIDTH-1:0] wire_d29_34;
	wire [WIDTH-1:0] wire_d29_35;
	wire [WIDTH-1:0] wire_d30_0;
	wire [WIDTH-1:0] wire_d30_1;
	wire [WIDTH-1:0] wire_d30_2;
	wire [WIDTH-1:0] wire_d30_3;
	wire [WIDTH-1:0] wire_d30_4;
	wire [WIDTH-1:0] wire_d30_5;
	wire [WIDTH-1:0] wire_d30_6;
	wire [WIDTH-1:0] wire_d30_7;
	wire [WIDTH-1:0] wire_d30_8;
	wire [WIDTH-1:0] wire_d30_9;
	wire [WIDTH-1:0] wire_d30_10;
	wire [WIDTH-1:0] wire_d30_11;
	wire [WIDTH-1:0] wire_d30_12;
	wire [WIDTH-1:0] wire_d30_13;
	wire [WIDTH-1:0] wire_d30_14;
	wire [WIDTH-1:0] wire_d30_15;
	wire [WIDTH-1:0] wire_d30_16;
	wire [WIDTH-1:0] wire_d30_17;
	wire [WIDTH-1:0] wire_d30_18;
	wire [WIDTH-1:0] wire_d30_19;
	wire [WIDTH-1:0] wire_d30_20;
	wire [WIDTH-1:0] wire_d30_21;
	wire [WIDTH-1:0] wire_d30_22;
	wire [WIDTH-1:0] wire_d30_23;
	wire [WIDTH-1:0] wire_d30_24;
	wire [WIDTH-1:0] wire_d30_25;
	wire [WIDTH-1:0] wire_d30_26;
	wire [WIDTH-1:0] wire_d30_27;
	wire [WIDTH-1:0] wire_d30_28;
	wire [WIDTH-1:0] wire_d30_29;
	wire [WIDTH-1:0] wire_d30_30;
	wire [WIDTH-1:0] wire_d30_31;
	wire [WIDTH-1:0] wire_d30_32;
	wire [WIDTH-1:0] wire_d30_33;
	wire [WIDTH-1:0] wire_d30_34;
	wire [WIDTH-1:0] wire_d30_35;
	wire [WIDTH-1:0] wire_d31_0;
	wire [WIDTH-1:0] wire_d31_1;
	wire [WIDTH-1:0] wire_d31_2;
	wire [WIDTH-1:0] wire_d31_3;
	wire [WIDTH-1:0] wire_d31_4;
	wire [WIDTH-1:0] wire_d31_5;
	wire [WIDTH-1:0] wire_d31_6;
	wire [WIDTH-1:0] wire_d31_7;
	wire [WIDTH-1:0] wire_d31_8;
	wire [WIDTH-1:0] wire_d31_9;
	wire [WIDTH-1:0] wire_d31_10;
	wire [WIDTH-1:0] wire_d31_11;
	wire [WIDTH-1:0] wire_d31_12;
	wire [WIDTH-1:0] wire_d31_13;
	wire [WIDTH-1:0] wire_d31_14;
	wire [WIDTH-1:0] wire_d31_15;
	wire [WIDTH-1:0] wire_d31_16;
	wire [WIDTH-1:0] wire_d31_17;
	wire [WIDTH-1:0] wire_d31_18;
	wire [WIDTH-1:0] wire_d31_19;
	wire [WIDTH-1:0] wire_d31_20;
	wire [WIDTH-1:0] wire_d31_21;
	wire [WIDTH-1:0] wire_d31_22;
	wire [WIDTH-1:0] wire_d31_23;
	wire [WIDTH-1:0] wire_d31_24;
	wire [WIDTH-1:0] wire_d31_25;
	wire [WIDTH-1:0] wire_d31_26;
	wire [WIDTH-1:0] wire_d31_27;
	wire [WIDTH-1:0] wire_d31_28;
	wire [WIDTH-1:0] wire_d31_29;
	wire [WIDTH-1:0] wire_d31_30;
	wire [WIDTH-1:0] wire_d31_31;
	wire [WIDTH-1:0] wire_d31_32;
	wire [WIDTH-1:0] wire_d31_33;
	wire [WIDTH-1:0] wire_d31_34;
	wire [WIDTH-1:0] wire_d31_35;
	wire [WIDTH-1:0] wire_d32_0;
	wire [WIDTH-1:0] wire_d32_1;
	wire [WIDTH-1:0] wire_d32_2;
	wire [WIDTH-1:0] wire_d32_3;
	wire [WIDTH-1:0] wire_d32_4;
	wire [WIDTH-1:0] wire_d32_5;
	wire [WIDTH-1:0] wire_d32_6;
	wire [WIDTH-1:0] wire_d32_7;
	wire [WIDTH-1:0] wire_d32_8;
	wire [WIDTH-1:0] wire_d32_9;
	wire [WIDTH-1:0] wire_d32_10;
	wire [WIDTH-1:0] wire_d32_11;
	wire [WIDTH-1:0] wire_d32_12;
	wire [WIDTH-1:0] wire_d32_13;
	wire [WIDTH-1:0] wire_d32_14;
	wire [WIDTH-1:0] wire_d32_15;
	wire [WIDTH-1:0] wire_d32_16;
	wire [WIDTH-1:0] wire_d32_17;
	wire [WIDTH-1:0] wire_d32_18;
	wire [WIDTH-1:0] wire_d32_19;
	wire [WIDTH-1:0] wire_d32_20;
	wire [WIDTH-1:0] wire_d32_21;
	wire [WIDTH-1:0] wire_d32_22;
	wire [WIDTH-1:0] wire_d32_23;
	wire [WIDTH-1:0] wire_d32_24;
	wire [WIDTH-1:0] wire_d32_25;
	wire [WIDTH-1:0] wire_d32_26;
	wire [WIDTH-1:0] wire_d32_27;
	wire [WIDTH-1:0] wire_d32_28;
	wire [WIDTH-1:0] wire_d32_29;
	wire [WIDTH-1:0] wire_d32_30;
	wire [WIDTH-1:0] wire_d32_31;
	wire [WIDTH-1:0] wire_d32_32;
	wire [WIDTH-1:0] wire_d32_33;
	wire [WIDTH-1:0] wire_d32_34;
	wire [WIDTH-1:0] wire_d32_35;
	wire [WIDTH-1:0] wire_d33_0;
	wire [WIDTH-1:0] wire_d33_1;
	wire [WIDTH-1:0] wire_d33_2;
	wire [WIDTH-1:0] wire_d33_3;
	wire [WIDTH-1:0] wire_d33_4;
	wire [WIDTH-1:0] wire_d33_5;
	wire [WIDTH-1:0] wire_d33_6;
	wire [WIDTH-1:0] wire_d33_7;
	wire [WIDTH-1:0] wire_d33_8;
	wire [WIDTH-1:0] wire_d33_9;
	wire [WIDTH-1:0] wire_d33_10;
	wire [WIDTH-1:0] wire_d33_11;
	wire [WIDTH-1:0] wire_d33_12;
	wire [WIDTH-1:0] wire_d33_13;
	wire [WIDTH-1:0] wire_d33_14;
	wire [WIDTH-1:0] wire_d33_15;
	wire [WIDTH-1:0] wire_d33_16;
	wire [WIDTH-1:0] wire_d33_17;
	wire [WIDTH-1:0] wire_d33_18;
	wire [WIDTH-1:0] wire_d33_19;
	wire [WIDTH-1:0] wire_d33_20;
	wire [WIDTH-1:0] wire_d33_21;
	wire [WIDTH-1:0] wire_d33_22;
	wire [WIDTH-1:0] wire_d33_23;
	wire [WIDTH-1:0] wire_d33_24;
	wire [WIDTH-1:0] wire_d33_25;
	wire [WIDTH-1:0] wire_d33_26;
	wire [WIDTH-1:0] wire_d33_27;
	wire [WIDTH-1:0] wire_d33_28;
	wire [WIDTH-1:0] wire_d33_29;
	wire [WIDTH-1:0] wire_d33_30;
	wire [WIDTH-1:0] wire_d33_31;
	wire [WIDTH-1:0] wire_d33_32;
	wire [WIDTH-1:0] wire_d33_33;
	wire [WIDTH-1:0] wire_d33_34;
	wire [WIDTH-1:0] wire_d33_35;
	wire [WIDTH-1:0] wire_d34_0;
	wire [WIDTH-1:0] wire_d34_1;
	wire [WIDTH-1:0] wire_d34_2;
	wire [WIDTH-1:0] wire_d34_3;
	wire [WIDTH-1:0] wire_d34_4;
	wire [WIDTH-1:0] wire_d34_5;
	wire [WIDTH-1:0] wire_d34_6;
	wire [WIDTH-1:0] wire_d34_7;
	wire [WIDTH-1:0] wire_d34_8;
	wire [WIDTH-1:0] wire_d34_9;
	wire [WIDTH-1:0] wire_d34_10;
	wire [WIDTH-1:0] wire_d34_11;
	wire [WIDTH-1:0] wire_d34_12;
	wire [WIDTH-1:0] wire_d34_13;
	wire [WIDTH-1:0] wire_d34_14;
	wire [WIDTH-1:0] wire_d34_15;
	wire [WIDTH-1:0] wire_d34_16;
	wire [WIDTH-1:0] wire_d34_17;
	wire [WIDTH-1:0] wire_d34_18;
	wire [WIDTH-1:0] wire_d34_19;
	wire [WIDTH-1:0] wire_d34_20;
	wire [WIDTH-1:0] wire_d34_21;
	wire [WIDTH-1:0] wire_d34_22;
	wire [WIDTH-1:0] wire_d34_23;
	wire [WIDTH-1:0] wire_d34_24;
	wire [WIDTH-1:0] wire_d34_25;
	wire [WIDTH-1:0] wire_d34_26;
	wire [WIDTH-1:0] wire_d34_27;
	wire [WIDTH-1:0] wire_d34_28;
	wire [WIDTH-1:0] wire_d34_29;
	wire [WIDTH-1:0] wire_d34_30;
	wire [WIDTH-1:0] wire_d34_31;
	wire [WIDTH-1:0] wire_d34_32;
	wire [WIDTH-1:0] wire_d34_33;
	wire [WIDTH-1:0] wire_d34_34;
	wire [WIDTH-1:0] wire_d34_35;
	wire [WIDTH-1:0] wire_d35_0;
	wire [WIDTH-1:0] wire_d35_1;
	wire [WIDTH-1:0] wire_d35_2;
	wire [WIDTH-1:0] wire_d35_3;
	wire [WIDTH-1:0] wire_d35_4;
	wire [WIDTH-1:0] wire_d35_5;
	wire [WIDTH-1:0] wire_d35_6;
	wire [WIDTH-1:0] wire_d35_7;
	wire [WIDTH-1:0] wire_d35_8;
	wire [WIDTH-1:0] wire_d35_9;
	wire [WIDTH-1:0] wire_d35_10;
	wire [WIDTH-1:0] wire_d35_11;
	wire [WIDTH-1:0] wire_d35_12;
	wire [WIDTH-1:0] wire_d35_13;
	wire [WIDTH-1:0] wire_d35_14;
	wire [WIDTH-1:0] wire_d35_15;
	wire [WIDTH-1:0] wire_d35_16;
	wire [WIDTH-1:0] wire_d35_17;
	wire [WIDTH-1:0] wire_d35_18;
	wire [WIDTH-1:0] wire_d35_19;
	wire [WIDTH-1:0] wire_d35_20;
	wire [WIDTH-1:0] wire_d35_21;
	wire [WIDTH-1:0] wire_d35_22;
	wire [WIDTH-1:0] wire_d35_23;
	wire [WIDTH-1:0] wire_d35_24;
	wire [WIDTH-1:0] wire_d35_25;
	wire [WIDTH-1:0] wire_d35_26;
	wire [WIDTH-1:0] wire_d35_27;
	wire [WIDTH-1:0] wire_d35_28;
	wire [WIDTH-1:0] wire_d35_29;
	wire [WIDTH-1:0] wire_d35_30;
	wire [WIDTH-1:0] wire_d35_31;
	wire [WIDTH-1:0] wire_d35_32;
	wire [WIDTH-1:0] wire_d35_33;
	wire [WIDTH-1:0] wire_d35_34;
	wire [WIDTH-1:0] wire_d35_35;

	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance100(.data_in(d_in0),.data_out(wire_d0_0),.clk(clk),.rst(rst));            //channel 1
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance101(.data_in(wire_d0_0),.data_out(wire_d0_1),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance102(.data_in(wire_d0_1),.data_out(wire_d0_2),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance103(.data_in(wire_d0_2),.data_out(wire_d0_3),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance104(.data_in(wire_d0_3),.data_out(wire_d0_4),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance105(.data_in(wire_d0_4),.data_out(wire_d0_5),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance106(.data_in(wire_d0_5),.data_out(wire_d0_6),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance107(.data_in(wire_d0_6),.data_out(wire_d0_7),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance108(.data_in(wire_d0_7),.data_out(wire_d0_8),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance109(.data_in(wire_d0_8),.data_out(wire_d0_9),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1010(.data_in(wire_d0_9),.data_out(wire_d0_10),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1011(.data_in(wire_d0_10),.data_out(wire_d0_11),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1012(.data_in(wire_d0_11),.data_out(wire_d0_12),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1013(.data_in(wire_d0_12),.data_out(wire_d0_13),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1014(.data_in(wire_d0_13),.data_out(wire_d0_14),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1015(.data_in(wire_d0_14),.data_out(wire_d0_15),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1016(.data_in(wire_d0_15),.data_out(wire_d0_16),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1017(.data_in(wire_d0_16),.data_out(wire_d0_17),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1018(.data_in(wire_d0_17),.data_out(wire_d0_18),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1019(.data_in(wire_d0_18),.data_out(wire_d0_19),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1020(.data_in(wire_d0_19),.data_out(wire_d0_20),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1021(.data_in(wire_d0_20),.data_out(wire_d0_21),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1022(.data_in(wire_d0_21),.data_out(wire_d0_22),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1023(.data_in(wire_d0_22),.data_out(wire_d0_23),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1024(.data_in(wire_d0_23),.data_out(wire_d0_24),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1025(.data_in(wire_d0_24),.data_out(wire_d0_25),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1026(.data_in(wire_d0_25),.data_out(wire_d0_26),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1027(.data_in(wire_d0_26),.data_out(wire_d0_27),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1028(.data_in(wire_d0_27),.data_out(wire_d0_28),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1029(.data_in(wire_d0_28),.data_out(wire_d0_29),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1030(.data_in(wire_d0_29),.data_out(wire_d0_30),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1031(.data_in(wire_d0_30),.data_out(wire_d0_31),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1032(.data_in(wire_d0_31),.data_out(wire_d0_32),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1033(.data_in(wire_d0_32),.data_out(wire_d0_33),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1034(.data_in(wire_d0_33),.data_out(wire_d0_34),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1035(.data_in(wire_d0_34),.data_out(wire_d0_35),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1036(.data_in(wire_d0_35),.data_out(d_out0),.clk(clk),.rst(rst));

	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance210(.data_in(d_in1),.data_out(wire_d1_0),.clk(clk),.rst(rst));            //channel 2
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance211(.data_in(wire_d1_0),.data_out(wire_d1_1),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance212(.data_in(wire_d1_1),.data_out(wire_d1_2),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance213(.data_in(wire_d1_2),.data_out(wire_d1_3),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance214(.data_in(wire_d1_3),.data_out(wire_d1_4),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance215(.data_in(wire_d1_4),.data_out(wire_d1_5),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance216(.data_in(wire_d1_5),.data_out(wire_d1_6),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance217(.data_in(wire_d1_6),.data_out(wire_d1_7),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance218(.data_in(wire_d1_7),.data_out(wire_d1_8),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance219(.data_in(wire_d1_8),.data_out(wire_d1_9),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2110(.data_in(wire_d1_9),.data_out(wire_d1_10),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2111(.data_in(wire_d1_10),.data_out(wire_d1_11),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2112(.data_in(wire_d1_11),.data_out(wire_d1_12),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2113(.data_in(wire_d1_12),.data_out(wire_d1_13),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2114(.data_in(wire_d1_13),.data_out(wire_d1_14),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2115(.data_in(wire_d1_14),.data_out(wire_d1_15),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2116(.data_in(wire_d1_15),.data_out(wire_d1_16),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2117(.data_in(wire_d1_16),.data_out(wire_d1_17),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2118(.data_in(wire_d1_17),.data_out(wire_d1_18),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2119(.data_in(wire_d1_18),.data_out(wire_d1_19),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2120(.data_in(wire_d1_19),.data_out(wire_d1_20),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2121(.data_in(wire_d1_20),.data_out(wire_d1_21),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2122(.data_in(wire_d1_21),.data_out(wire_d1_22),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2123(.data_in(wire_d1_22),.data_out(wire_d1_23),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2124(.data_in(wire_d1_23),.data_out(wire_d1_24),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2125(.data_in(wire_d1_24),.data_out(wire_d1_25),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2126(.data_in(wire_d1_25),.data_out(wire_d1_26),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2127(.data_in(wire_d1_26),.data_out(wire_d1_27),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2128(.data_in(wire_d1_27),.data_out(wire_d1_28),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2129(.data_in(wire_d1_28),.data_out(wire_d1_29),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2130(.data_in(wire_d1_29),.data_out(wire_d1_30),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2131(.data_in(wire_d1_30),.data_out(wire_d1_31),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2132(.data_in(wire_d1_31),.data_out(wire_d1_32),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2133(.data_in(wire_d1_32),.data_out(wire_d1_33),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2134(.data_in(wire_d1_33),.data_out(wire_d1_34),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2135(.data_in(wire_d1_34),.data_out(wire_d1_35),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2136(.data_in(wire_d1_35),.data_out(d_out1),.clk(clk),.rst(rst));

	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance320(.data_in(d_in2),.data_out(wire_d2_0),.clk(clk),.rst(rst));            //channel 3
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance321(.data_in(wire_d2_0),.data_out(wire_d2_1),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance322(.data_in(wire_d2_1),.data_out(wire_d2_2),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance323(.data_in(wire_d2_2),.data_out(wire_d2_3),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance324(.data_in(wire_d2_3),.data_out(wire_d2_4),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance325(.data_in(wire_d2_4),.data_out(wire_d2_5),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance326(.data_in(wire_d2_5),.data_out(wire_d2_6),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance327(.data_in(wire_d2_6),.data_out(wire_d2_7),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance328(.data_in(wire_d2_7),.data_out(wire_d2_8),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance329(.data_in(wire_d2_8),.data_out(wire_d2_9),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3210(.data_in(wire_d2_9),.data_out(wire_d2_10),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3211(.data_in(wire_d2_10),.data_out(wire_d2_11),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3212(.data_in(wire_d2_11),.data_out(wire_d2_12),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3213(.data_in(wire_d2_12),.data_out(wire_d2_13),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3214(.data_in(wire_d2_13),.data_out(wire_d2_14),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3215(.data_in(wire_d2_14),.data_out(wire_d2_15),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3216(.data_in(wire_d2_15),.data_out(wire_d2_16),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3217(.data_in(wire_d2_16),.data_out(wire_d2_17),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3218(.data_in(wire_d2_17),.data_out(wire_d2_18),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3219(.data_in(wire_d2_18),.data_out(wire_d2_19),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3220(.data_in(wire_d2_19),.data_out(wire_d2_20),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3221(.data_in(wire_d2_20),.data_out(wire_d2_21),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3222(.data_in(wire_d2_21),.data_out(wire_d2_22),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3223(.data_in(wire_d2_22),.data_out(wire_d2_23),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3224(.data_in(wire_d2_23),.data_out(wire_d2_24),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3225(.data_in(wire_d2_24),.data_out(wire_d2_25),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3226(.data_in(wire_d2_25),.data_out(wire_d2_26),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3227(.data_in(wire_d2_26),.data_out(wire_d2_27),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3228(.data_in(wire_d2_27),.data_out(wire_d2_28),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3229(.data_in(wire_d2_28),.data_out(wire_d2_29),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3230(.data_in(wire_d2_29),.data_out(wire_d2_30),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3231(.data_in(wire_d2_30),.data_out(wire_d2_31),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3232(.data_in(wire_d2_31),.data_out(wire_d2_32),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3233(.data_in(wire_d2_32),.data_out(wire_d2_33),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3234(.data_in(wire_d2_33),.data_out(wire_d2_34),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3235(.data_in(wire_d2_34),.data_out(wire_d2_35),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3236(.data_in(wire_d2_35),.data_out(d_out2),.clk(clk),.rst(rst));

	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance430(.data_in(d_in3),.data_out(wire_d3_0),.clk(clk),.rst(rst));            //channel 4
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance431(.data_in(wire_d3_0),.data_out(wire_d3_1),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance432(.data_in(wire_d3_1),.data_out(wire_d3_2),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance433(.data_in(wire_d3_2),.data_out(wire_d3_3),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance434(.data_in(wire_d3_3),.data_out(wire_d3_4),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance435(.data_in(wire_d3_4),.data_out(wire_d3_5),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance436(.data_in(wire_d3_5),.data_out(wire_d3_6),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance437(.data_in(wire_d3_6),.data_out(wire_d3_7),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance438(.data_in(wire_d3_7),.data_out(wire_d3_8),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance439(.data_in(wire_d3_8),.data_out(wire_d3_9),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance4310(.data_in(wire_d3_9),.data_out(wire_d3_10),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance4311(.data_in(wire_d3_10),.data_out(wire_d3_11),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance4312(.data_in(wire_d3_11),.data_out(wire_d3_12),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance4313(.data_in(wire_d3_12),.data_out(wire_d3_13),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance4314(.data_in(wire_d3_13),.data_out(wire_d3_14),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance4315(.data_in(wire_d3_14),.data_out(wire_d3_15),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance4316(.data_in(wire_d3_15),.data_out(wire_d3_16),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance4317(.data_in(wire_d3_16),.data_out(wire_d3_17),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance4318(.data_in(wire_d3_17),.data_out(wire_d3_18),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance4319(.data_in(wire_d3_18),.data_out(wire_d3_19),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance4320(.data_in(wire_d3_19),.data_out(wire_d3_20),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance4321(.data_in(wire_d3_20),.data_out(wire_d3_21),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance4322(.data_in(wire_d3_21),.data_out(wire_d3_22),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance4323(.data_in(wire_d3_22),.data_out(wire_d3_23),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance4324(.data_in(wire_d3_23),.data_out(wire_d3_24),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance4325(.data_in(wire_d3_24),.data_out(wire_d3_25),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance4326(.data_in(wire_d3_25),.data_out(wire_d3_26),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance4327(.data_in(wire_d3_26),.data_out(wire_d3_27),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance4328(.data_in(wire_d3_27),.data_out(wire_d3_28),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance4329(.data_in(wire_d3_28),.data_out(wire_d3_29),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance4330(.data_in(wire_d3_29),.data_out(wire_d3_30),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance4331(.data_in(wire_d3_30),.data_out(wire_d3_31),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance4332(.data_in(wire_d3_31),.data_out(wire_d3_32),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance4333(.data_in(wire_d3_32),.data_out(wire_d3_33),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance4334(.data_in(wire_d3_33),.data_out(wire_d3_34),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance4335(.data_in(wire_d3_34),.data_out(wire_d3_35),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance4336(.data_in(wire_d3_35),.data_out(d_out3),.clk(clk),.rst(rst));

	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance540(.data_in(d_in4),.data_out(wire_d4_0),.clk(clk),.rst(rst));            //channel 5
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance541(.data_in(wire_d4_0),.data_out(wire_d4_1),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance542(.data_in(wire_d4_1),.data_out(wire_d4_2),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance543(.data_in(wire_d4_2),.data_out(wire_d4_3),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance544(.data_in(wire_d4_3),.data_out(wire_d4_4),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance545(.data_in(wire_d4_4),.data_out(wire_d4_5),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance546(.data_in(wire_d4_5),.data_out(wire_d4_6),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance547(.data_in(wire_d4_6),.data_out(wire_d4_7),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance548(.data_in(wire_d4_7),.data_out(wire_d4_8),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance549(.data_in(wire_d4_8),.data_out(wire_d4_9),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance5410(.data_in(wire_d4_9),.data_out(wire_d4_10),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance5411(.data_in(wire_d4_10),.data_out(wire_d4_11),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance5412(.data_in(wire_d4_11),.data_out(wire_d4_12),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance5413(.data_in(wire_d4_12),.data_out(wire_d4_13),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance5414(.data_in(wire_d4_13),.data_out(wire_d4_14),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance5415(.data_in(wire_d4_14),.data_out(wire_d4_15),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance5416(.data_in(wire_d4_15),.data_out(wire_d4_16),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance5417(.data_in(wire_d4_16),.data_out(wire_d4_17),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance5418(.data_in(wire_d4_17),.data_out(wire_d4_18),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance5419(.data_in(wire_d4_18),.data_out(wire_d4_19),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance5420(.data_in(wire_d4_19),.data_out(wire_d4_20),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance5421(.data_in(wire_d4_20),.data_out(wire_d4_21),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance5422(.data_in(wire_d4_21),.data_out(wire_d4_22),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance5423(.data_in(wire_d4_22),.data_out(wire_d4_23),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance5424(.data_in(wire_d4_23),.data_out(wire_d4_24),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance5425(.data_in(wire_d4_24),.data_out(wire_d4_25),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance5426(.data_in(wire_d4_25),.data_out(wire_d4_26),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance5427(.data_in(wire_d4_26),.data_out(wire_d4_27),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance5428(.data_in(wire_d4_27),.data_out(wire_d4_28),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance5429(.data_in(wire_d4_28),.data_out(wire_d4_29),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance5430(.data_in(wire_d4_29),.data_out(wire_d4_30),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance5431(.data_in(wire_d4_30),.data_out(wire_d4_31),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance5432(.data_in(wire_d4_31),.data_out(wire_d4_32),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance5433(.data_in(wire_d4_32),.data_out(wire_d4_33),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance5434(.data_in(wire_d4_33),.data_out(wire_d4_34),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance5435(.data_in(wire_d4_34),.data_out(wire_d4_35),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance5436(.data_in(wire_d4_35),.data_out(d_out4),.clk(clk),.rst(rst));

	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance650(.data_in(d_in5),.data_out(wire_d5_0),.clk(clk),.rst(rst));            //channel 6
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance651(.data_in(wire_d5_0),.data_out(wire_d5_1),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance652(.data_in(wire_d5_1),.data_out(wire_d5_2),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance653(.data_in(wire_d5_2),.data_out(wire_d5_3),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance654(.data_in(wire_d5_3),.data_out(wire_d5_4),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance655(.data_in(wire_d5_4),.data_out(wire_d5_5),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance656(.data_in(wire_d5_5),.data_out(wire_d5_6),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance657(.data_in(wire_d5_6),.data_out(wire_d5_7),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance658(.data_in(wire_d5_7),.data_out(wire_d5_8),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance659(.data_in(wire_d5_8),.data_out(wire_d5_9),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance6510(.data_in(wire_d5_9),.data_out(wire_d5_10),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance6511(.data_in(wire_d5_10),.data_out(wire_d5_11),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance6512(.data_in(wire_d5_11),.data_out(wire_d5_12),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance6513(.data_in(wire_d5_12),.data_out(wire_d5_13),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance6514(.data_in(wire_d5_13),.data_out(wire_d5_14),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance6515(.data_in(wire_d5_14),.data_out(wire_d5_15),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance6516(.data_in(wire_d5_15),.data_out(wire_d5_16),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance6517(.data_in(wire_d5_16),.data_out(wire_d5_17),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance6518(.data_in(wire_d5_17),.data_out(wire_d5_18),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance6519(.data_in(wire_d5_18),.data_out(wire_d5_19),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance6520(.data_in(wire_d5_19),.data_out(wire_d5_20),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance6521(.data_in(wire_d5_20),.data_out(wire_d5_21),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance6522(.data_in(wire_d5_21),.data_out(wire_d5_22),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance6523(.data_in(wire_d5_22),.data_out(wire_d5_23),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance6524(.data_in(wire_d5_23),.data_out(wire_d5_24),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance6525(.data_in(wire_d5_24),.data_out(wire_d5_25),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance6526(.data_in(wire_d5_25),.data_out(wire_d5_26),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance6527(.data_in(wire_d5_26),.data_out(wire_d5_27),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance6528(.data_in(wire_d5_27),.data_out(wire_d5_28),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance6529(.data_in(wire_d5_28),.data_out(wire_d5_29),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance6530(.data_in(wire_d5_29),.data_out(wire_d5_30),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance6531(.data_in(wire_d5_30),.data_out(wire_d5_31),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance6532(.data_in(wire_d5_31),.data_out(wire_d5_32),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance6533(.data_in(wire_d5_32),.data_out(wire_d5_33),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance6534(.data_in(wire_d5_33),.data_out(wire_d5_34),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance6535(.data_in(wire_d5_34),.data_out(wire_d5_35),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance6536(.data_in(wire_d5_35),.data_out(d_out5),.clk(clk),.rst(rst));

	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance760(.data_in(d_in6),.data_out(wire_d6_0),.clk(clk),.rst(rst));            //channel 7
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance761(.data_in(wire_d6_0),.data_out(wire_d6_1),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance762(.data_in(wire_d6_1),.data_out(wire_d6_2),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance763(.data_in(wire_d6_2),.data_out(wire_d6_3),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance764(.data_in(wire_d6_3),.data_out(wire_d6_4),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance765(.data_in(wire_d6_4),.data_out(wire_d6_5),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance766(.data_in(wire_d6_5),.data_out(wire_d6_6),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance767(.data_in(wire_d6_6),.data_out(wire_d6_7),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance768(.data_in(wire_d6_7),.data_out(wire_d6_8),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance769(.data_in(wire_d6_8),.data_out(wire_d6_9),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance7610(.data_in(wire_d6_9),.data_out(wire_d6_10),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance7611(.data_in(wire_d6_10),.data_out(wire_d6_11),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance7612(.data_in(wire_d6_11),.data_out(wire_d6_12),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance7613(.data_in(wire_d6_12),.data_out(wire_d6_13),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance7614(.data_in(wire_d6_13),.data_out(wire_d6_14),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance7615(.data_in(wire_d6_14),.data_out(wire_d6_15),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance7616(.data_in(wire_d6_15),.data_out(wire_d6_16),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance7617(.data_in(wire_d6_16),.data_out(wire_d6_17),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance7618(.data_in(wire_d6_17),.data_out(wire_d6_18),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance7619(.data_in(wire_d6_18),.data_out(wire_d6_19),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance7620(.data_in(wire_d6_19),.data_out(wire_d6_20),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance7621(.data_in(wire_d6_20),.data_out(wire_d6_21),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance7622(.data_in(wire_d6_21),.data_out(wire_d6_22),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance7623(.data_in(wire_d6_22),.data_out(wire_d6_23),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance7624(.data_in(wire_d6_23),.data_out(wire_d6_24),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance7625(.data_in(wire_d6_24),.data_out(wire_d6_25),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance7626(.data_in(wire_d6_25),.data_out(wire_d6_26),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance7627(.data_in(wire_d6_26),.data_out(wire_d6_27),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance7628(.data_in(wire_d6_27),.data_out(wire_d6_28),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance7629(.data_in(wire_d6_28),.data_out(wire_d6_29),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance7630(.data_in(wire_d6_29),.data_out(wire_d6_30),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance7631(.data_in(wire_d6_30),.data_out(wire_d6_31),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance7632(.data_in(wire_d6_31),.data_out(wire_d6_32),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance7633(.data_in(wire_d6_32),.data_out(wire_d6_33),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance7634(.data_in(wire_d6_33),.data_out(wire_d6_34),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance7635(.data_in(wire_d6_34),.data_out(wire_d6_35),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance7636(.data_in(wire_d6_35),.data_out(d_out6),.clk(clk),.rst(rst));

	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance870(.data_in(d_in7),.data_out(wire_d7_0),.clk(clk),.rst(rst));            //channel 8
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance871(.data_in(wire_d7_0),.data_out(wire_d7_1),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance872(.data_in(wire_d7_1),.data_out(wire_d7_2),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance873(.data_in(wire_d7_2),.data_out(wire_d7_3),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance874(.data_in(wire_d7_3),.data_out(wire_d7_4),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance875(.data_in(wire_d7_4),.data_out(wire_d7_5),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance876(.data_in(wire_d7_5),.data_out(wire_d7_6),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance877(.data_in(wire_d7_6),.data_out(wire_d7_7),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance878(.data_in(wire_d7_7),.data_out(wire_d7_8),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance879(.data_in(wire_d7_8),.data_out(wire_d7_9),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance8710(.data_in(wire_d7_9),.data_out(wire_d7_10),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance8711(.data_in(wire_d7_10),.data_out(wire_d7_11),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance8712(.data_in(wire_d7_11),.data_out(wire_d7_12),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance8713(.data_in(wire_d7_12),.data_out(wire_d7_13),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance8714(.data_in(wire_d7_13),.data_out(wire_d7_14),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance8715(.data_in(wire_d7_14),.data_out(wire_d7_15),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance8716(.data_in(wire_d7_15),.data_out(wire_d7_16),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance8717(.data_in(wire_d7_16),.data_out(wire_d7_17),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance8718(.data_in(wire_d7_17),.data_out(wire_d7_18),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance8719(.data_in(wire_d7_18),.data_out(wire_d7_19),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance8720(.data_in(wire_d7_19),.data_out(wire_d7_20),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance8721(.data_in(wire_d7_20),.data_out(wire_d7_21),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance8722(.data_in(wire_d7_21),.data_out(wire_d7_22),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance8723(.data_in(wire_d7_22),.data_out(wire_d7_23),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance8724(.data_in(wire_d7_23),.data_out(wire_d7_24),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance8725(.data_in(wire_d7_24),.data_out(wire_d7_25),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance8726(.data_in(wire_d7_25),.data_out(wire_d7_26),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance8727(.data_in(wire_d7_26),.data_out(wire_d7_27),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance8728(.data_in(wire_d7_27),.data_out(wire_d7_28),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance8729(.data_in(wire_d7_28),.data_out(wire_d7_29),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance8730(.data_in(wire_d7_29),.data_out(wire_d7_30),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance8731(.data_in(wire_d7_30),.data_out(wire_d7_31),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance8732(.data_in(wire_d7_31),.data_out(wire_d7_32),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance8733(.data_in(wire_d7_32),.data_out(wire_d7_33),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance8734(.data_in(wire_d7_33),.data_out(wire_d7_34),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance8735(.data_in(wire_d7_34),.data_out(wire_d7_35),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance8736(.data_in(wire_d7_35),.data_out(d_out7),.clk(clk),.rst(rst));

	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance980(.data_in(d_in8),.data_out(wire_d8_0),.clk(clk),.rst(rst));            //channel 9
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance981(.data_in(wire_d8_0),.data_out(wire_d8_1),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance982(.data_in(wire_d8_1),.data_out(wire_d8_2),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance983(.data_in(wire_d8_2),.data_out(wire_d8_3),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance984(.data_in(wire_d8_3),.data_out(wire_d8_4),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance985(.data_in(wire_d8_4),.data_out(wire_d8_5),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance986(.data_in(wire_d8_5),.data_out(wire_d8_6),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance987(.data_in(wire_d8_6),.data_out(wire_d8_7),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance988(.data_in(wire_d8_7),.data_out(wire_d8_8),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance989(.data_in(wire_d8_8),.data_out(wire_d8_9),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance9810(.data_in(wire_d8_9),.data_out(wire_d8_10),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance9811(.data_in(wire_d8_10),.data_out(wire_d8_11),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance9812(.data_in(wire_d8_11),.data_out(wire_d8_12),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance9813(.data_in(wire_d8_12),.data_out(wire_d8_13),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance9814(.data_in(wire_d8_13),.data_out(wire_d8_14),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance9815(.data_in(wire_d8_14),.data_out(wire_d8_15),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance9816(.data_in(wire_d8_15),.data_out(wire_d8_16),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance9817(.data_in(wire_d8_16),.data_out(wire_d8_17),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance9818(.data_in(wire_d8_17),.data_out(wire_d8_18),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance9819(.data_in(wire_d8_18),.data_out(wire_d8_19),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance9820(.data_in(wire_d8_19),.data_out(wire_d8_20),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance9821(.data_in(wire_d8_20),.data_out(wire_d8_21),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance9822(.data_in(wire_d8_21),.data_out(wire_d8_22),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance9823(.data_in(wire_d8_22),.data_out(wire_d8_23),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance9824(.data_in(wire_d8_23),.data_out(wire_d8_24),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance9825(.data_in(wire_d8_24),.data_out(wire_d8_25),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance9826(.data_in(wire_d8_25),.data_out(wire_d8_26),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance9827(.data_in(wire_d8_26),.data_out(wire_d8_27),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance9828(.data_in(wire_d8_27),.data_out(wire_d8_28),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance9829(.data_in(wire_d8_28),.data_out(wire_d8_29),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance9830(.data_in(wire_d8_29),.data_out(wire_d8_30),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance9831(.data_in(wire_d8_30),.data_out(wire_d8_31),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance9832(.data_in(wire_d8_31),.data_out(wire_d8_32),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance9833(.data_in(wire_d8_32),.data_out(wire_d8_33),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance9834(.data_in(wire_d8_33),.data_out(wire_d8_34),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance9835(.data_in(wire_d8_34),.data_out(wire_d8_35),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance9836(.data_in(wire_d8_35),.data_out(d_out8),.clk(clk),.rst(rst));

	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance10090(.data_in(d_in9),.data_out(wire_d9_0),.clk(clk),.rst(rst));            //channel 10
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance10091(.data_in(wire_d9_0),.data_out(wire_d9_1),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance10092(.data_in(wire_d9_1),.data_out(wire_d9_2),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance10093(.data_in(wire_d9_2),.data_out(wire_d9_3),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance10094(.data_in(wire_d9_3),.data_out(wire_d9_4),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance10095(.data_in(wire_d9_4),.data_out(wire_d9_5),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance10096(.data_in(wire_d9_5),.data_out(wire_d9_6),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance10097(.data_in(wire_d9_6),.data_out(wire_d9_7),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance10098(.data_in(wire_d9_7),.data_out(wire_d9_8),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance10099(.data_in(wire_d9_8),.data_out(wire_d9_9),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance100910(.data_in(wire_d9_9),.data_out(wire_d9_10),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance100911(.data_in(wire_d9_10),.data_out(wire_d9_11),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance100912(.data_in(wire_d9_11),.data_out(wire_d9_12),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance100913(.data_in(wire_d9_12),.data_out(wire_d9_13),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance100914(.data_in(wire_d9_13),.data_out(wire_d9_14),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance100915(.data_in(wire_d9_14),.data_out(wire_d9_15),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance100916(.data_in(wire_d9_15),.data_out(wire_d9_16),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance100917(.data_in(wire_d9_16),.data_out(wire_d9_17),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance100918(.data_in(wire_d9_17),.data_out(wire_d9_18),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance100919(.data_in(wire_d9_18),.data_out(wire_d9_19),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance100920(.data_in(wire_d9_19),.data_out(wire_d9_20),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance100921(.data_in(wire_d9_20),.data_out(wire_d9_21),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance100922(.data_in(wire_d9_21),.data_out(wire_d9_22),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance100923(.data_in(wire_d9_22),.data_out(wire_d9_23),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance100924(.data_in(wire_d9_23),.data_out(wire_d9_24),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance100925(.data_in(wire_d9_24),.data_out(wire_d9_25),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance100926(.data_in(wire_d9_25),.data_out(wire_d9_26),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance100927(.data_in(wire_d9_26),.data_out(wire_d9_27),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance100928(.data_in(wire_d9_27),.data_out(wire_d9_28),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance100929(.data_in(wire_d9_28),.data_out(wire_d9_29),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance100930(.data_in(wire_d9_29),.data_out(wire_d9_30),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance100931(.data_in(wire_d9_30),.data_out(wire_d9_31),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance100932(.data_in(wire_d9_31),.data_out(wire_d9_32),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance100933(.data_in(wire_d9_32),.data_out(wire_d9_33),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance100934(.data_in(wire_d9_33),.data_out(wire_d9_34),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance100935(.data_in(wire_d9_34),.data_out(wire_d9_35),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance100936(.data_in(wire_d9_35),.data_out(d_out9),.clk(clk),.rst(rst));

	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance110100(.data_in(d_in10),.data_out(wire_d10_0),.clk(clk),.rst(rst));            //channel 11
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance110101(.data_in(wire_d10_0),.data_out(wire_d10_1),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance110102(.data_in(wire_d10_1),.data_out(wire_d10_2),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance110103(.data_in(wire_d10_2),.data_out(wire_d10_3),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance110104(.data_in(wire_d10_3),.data_out(wire_d10_4),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance110105(.data_in(wire_d10_4),.data_out(wire_d10_5),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance110106(.data_in(wire_d10_5),.data_out(wire_d10_6),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance110107(.data_in(wire_d10_6),.data_out(wire_d10_7),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance110108(.data_in(wire_d10_7),.data_out(wire_d10_8),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance110109(.data_in(wire_d10_8),.data_out(wire_d10_9),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1101010(.data_in(wire_d10_9),.data_out(wire_d10_10),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1101011(.data_in(wire_d10_10),.data_out(wire_d10_11),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1101012(.data_in(wire_d10_11),.data_out(wire_d10_12),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1101013(.data_in(wire_d10_12),.data_out(wire_d10_13),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1101014(.data_in(wire_d10_13),.data_out(wire_d10_14),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1101015(.data_in(wire_d10_14),.data_out(wire_d10_15),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1101016(.data_in(wire_d10_15),.data_out(wire_d10_16),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1101017(.data_in(wire_d10_16),.data_out(wire_d10_17),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1101018(.data_in(wire_d10_17),.data_out(wire_d10_18),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1101019(.data_in(wire_d10_18),.data_out(wire_d10_19),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1101020(.data_in(wire_d10_19),.data_out(wire_d10_20),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1101021(.data_in(wire_d10_20),.data_out(wire_d10_21),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1101022(.data_in(wire_d10_21),.data_out(wire_d10_22),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1101023(.data_in(wire_d10_22),.data_out(wire_d10_23),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1101024(.data_in(wire_d10_23),.data_out(wire_d10_24),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1101025(.data_in(wire_d10_24),.data_out(wire_d10_25),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1101026(.data_in(wire_d10_25),.data_out(wire_d10_26),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1101027(.data_in(wire_d10_26),.data_out(wire_d10_27),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1101028(.data_in(wire_d10_27),.data_out(wire_d10_28),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1101029(.data_in(wire_d10_28),.data_out(wire_d10_29),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1101030(.data_in(wire_d10_29),.data_out(wire_d10_30),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1101031(.data_in(wire_d10_30),.data_out(wire_d10_31),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1101032(.data_in(wire_d10_31),.data_out(wire_d10_32),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1101033(.data_in(wire_d10_32),.data_out(wire_d10_33),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1101034(.data_in(wire_d10_33),.data_out(wire_d10_34),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1101035(.data_in(wire_d10_34),.data_out(wire_d10_35),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1101036(.data_in(wire_d10_35),.data_out(d_out10),.clk(clk),.rst(rst));

	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance120110(.data_in(d_in11),.data_out(wire_d11_0),.clk(clk),.rst(rst));            //channel 12
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance120111(.data_in(wire_d11_0),.data_out(wire_d11_1),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance120112(.data_in(wire_d11_1),.data_out(wire_d11_2),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance120113(.data_in(wire_d11_2),.data_out(wire_d11_3),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance120114(.data_in(wire_d11_3),.data_out(wire_d11_4),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance120115(.data_in(wire_d11_4),.data_out(wire_d11_5),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance120116(.data_in(wire_d11_5),.data_out(wire_d11_6),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance120117(.data_in(wire_d11_6),.data_out(wire_d11_7),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance120118(.data_in(wire_d11_7),.data_out(wire_d11_8),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance120119(.data_in(wire_d11_8),.data_out(wire_d11_9),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1201110(.data_in(wire_d11_9),.data_out(wire_d11_10),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1201111(.data_in(wire_d11_10),.data_out(wire_d11_11),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1201112(.data_in(wire_d11_11),.data_out(wire_d11_12),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1201113(.data_in(wire_d11_12),.data_out(wire_d11_13),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1201114(.data_in(wire_d11_13),.data_out(wire_d11_14),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1201115(.data_in(wire_d11_14),.data_out(wire_d11_15),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1201116(.data_in(wire_d11_15),.data_out(wire_d11_16),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1201117(.data_in(wire_d11_16),.data_out(wire_d11_17),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1201118(.data_in(wire_d11_17),.data_out(wire_d11_18),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1201119(.data_in(wire_d11_18),.data_out(wire_d11_19),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1201120(.data_in(wire_d11_19),.data_out(wire_d11_20),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1201121(.data_in(wire_d11_20),.data_out(wire_d11_21),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1201122(.data_in(wire_d11_21),.data_out(wire_d11_22),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1201123(.data_in(wire_d11_22),.data_out(wire_d11_23),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1201124(.data_in(wire_d11_23),.data_out(wire_d11_24),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1201125(.data_in(wire_d11_24),.data_out(wire_d11_25),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1201126(.data_in(wire_d11_25),.data_out(wire_d11_26),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1201127(.data_in(wire_d11_26),.data_out(wire_d11_27),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1201128(.data_in(wire_d11_27),.data_out(wire_d11_28),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1201129(.data_in(wire_d11_28),.data_out(wire_d11_29),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1201130(.data_in(wire_d11_29),.data_out(wire_d11_30),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1201131(.data_in(wire_d11_30),.data_out(wire_d11_31),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1201132(.data_in(wire_d11_31),.data_out(wire_d11_32),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1201133(.data_in(wire_d11_32),.data_out(wire_d11_33),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1201134(.data_in(wire_d11_33),.data_out(wire_d11_34),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1201135(.data_in(wire_d11_34),.data_out(wire_d11_35),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1201136(.data_in(wire_d11_35),.data_out(d_out11),.clk(clk),.rst(rst));

	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance130120(.data_in(d_in12),.data_out(wire_d12_0),.clk(clk),.rst(rst));            //channel 13
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance130121(.data_in(wire_d12_0),.data_out(wire_d12_1),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance130122(.data_in(wire_d12_1),.data_out(wire_d12_2),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance130123(.data_in(wire_d12_2),.data_out(wire_d12_3),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance130124(.data_in(wire_d12_3),.data_out(wire_d12_4),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance130125(.data_in(wire_d12_4),.data_out(wire_d12_5),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance130126(.data_in(wire_d12_5),.data_out(wire_d12_6),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance130127(.data_in(wire_d12_6),.data_out(wire_d12_7),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance130128(.data_in(wire_d12_7),.data_out(wire_d12_8),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance130129(.data_in(wire_d12_8),.data_out(wire_d12_9),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1301210(.data_in(wire_d12_9),.data_out(wire_d12_10),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1301211(.data_in(wire_d12_10),.data_out(wire_d12_11),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1301212(.data_in(wire_d12_11),.data_out(wire_d12_12),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1301213(.data_in(wire_d12_12),.data_out(wire_d12_13),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1301214(.data_in(wire_d12_13),.data_out(wire_d12_14),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1301215(.data_in(wire_d12_14),.data_out(wire_d12_15),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1301216(.data_in(wire_d12_15),.data_out(wire_d12_16),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1301217(.data_in(wire_d12_16),.data_out(wire_d12_17),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1301218(.data_in(wire_d12_17),.data_out(wire_d12_18),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1301219(.data_in(wire_d12_18),.data_out(wire_d12_19),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1301220(.data_in(wire_d12_19),.data_out(wire_d12_20),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1301221(.data_in(wire_d12_20),.data_out(wire_d12_21),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1301222(.data_in(wire_d12_21),.data_out(wire_d12_22),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1301223(.data_in(wire_d12_22),.data_out(wire_d12_23),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1301224(.data_in(wire_d12_23),.data_out(wire_d12_24),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1301225(.data_in(wire_d12_24),.data_out(wire_d12_25),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1301226(.data_in(wire_d12_25),.data_out(wire_d12_26),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1301227(.data_in(wire_d12_26),.data_out(wire_d12_27),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1301228(.data_in(wire_d12_27),.data_out(wire_d12_28),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1301229(.data_in(wire_d12_28),.data_out(wire_d12_29),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1301230(.data_in(wire_d12_29),.data_out(wire_d12_30),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1301231(.data_in(wire_d12_30),.data_out(wire_d12_31),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1301232(.data_in(wire_d12_31),.data_out(wire_d12_32),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1301233(.data_in(wire_d12_32),.data_out(wire_d12_33),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1301234(.data_in(wire_d12_33),.data_out(wire_d12_34),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1301235(.data_in(wire_d12_34),.data_out(wire_d12_35),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1301236(.data_in(wire_d12_35),.data_out(d_out12),.clk(clk),.rst(rst));

	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance140130(.data_in(d_in13),.data_out(wire_d13_0),.clk(clk),.rst(rst));            //channel 14
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance140131(.data_in(wire_d13_0),.data_out(wire_d13_1),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance140132(.data_in(wire_d13_1),.data_out(wire_d13_2),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance140133(.data_in(wire_d13_2),.data_out(wire_d13_3),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance140134(.data_in(wire_d13_3),.data_out(wire_d13_4),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance140135(.data_in(wire_d13_4),.data_out(wire_d13_5),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance140136(.data_in(wire_d13_5),.data_out(wire_d13_6),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance140137(.data_in(wire_d13_6),.data_out(wire_d13_7),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance140138(.data_in(wire_d13_7),.data_out(wire_d13_8),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance140139(.data_in(wire_d13_8),.data_out(wire_d13_9),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1401310(.data_in(wire_d13_9),.data_out(wire_d13_10),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1401311(.data_in(wire_d13_10),.data_out(wire_d13_11),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1401312(.data_in(wire_d13_11),.data_out(wire_d13_12),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1401313(.data_in(wire_d13_12),.data_out(wire_d13_13),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1401314(.data_in(wire_d13_13),.data_out(wire_d13_14),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1401315(.data_in(wire_d13_14),.data_out(wire_d13_15),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1401316(.data_in(wire_d13_15),.data_out(wire_d13_16),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1401317(.data_in(wire_d13_16),.data_out(wire_d13_17),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1401318(.data_in(wire_d13_17),.data_out(wire_d13_18),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1401319(.data_in(wire_d13_18),.data_out(wire_d13_19),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1401320(.data_in(wire_d13_19),.data_out(wire_d13_20),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1401321(.data_in(wire_d13_20),.data_out(wire_d13_21),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1401322(.data_in(wire_d13_21),.data_out(wire_d13_22),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1401323(.data_in(wire_d13_22),.data_out(wire_d13_23),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1401324(.data_in(wire_d13_23),.data_out(wire_d13_24),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1401325(.data_in(wire_d13_24),.data_out(wire_d13_25),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1401326(.data_in(wire_d13_25),.data_out(wire_d13_26),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1401327(.data_in(wire_d13_26),.data_out(wire_d13_27),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1401328(.data_in(wire_d13_27),.data_out(wire_d13_28),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1401329(.data_in(wire_d13_28),.data_out(wire_d13_29),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1401330(.data_in(wire_d13_29),.data_out(wire_d13_30),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1401331(.data_in(wire_d13_30),.data_out(wire_d13_31),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1401332(.data_in(wire_d13_31),.data_out(wire_d13_32),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1401333(.data_in(wire_d13_32),.data_out(wire_d13_33),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1401334(.data_in(wire_d13_33),.data_out(wire_d13_34),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1401335(.data_in(wire_d13_34),.data_out(wire_d13_35),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1401336(.data_in(wire_d13_35),.data_out(d_out13),.clk(clk),.rst(rst));

	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance150140(.data_in(d_in14),.data_out(wire_d14_0),.clk(clk),.rst(rst));            //channel 15
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance150141(.data_in(wire_d14_0),.data_out(wire_d14_1),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance150142(.data_in(wire_d14_1),.data_out(wire_d14_2),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance150143(.data_in(wire_d14_2),.data_out(wire_d14_3),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance150144(.data_in(wire_d14_3),.data_out(wire_d14_4),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance150145(.data_in(wire_d14_4),.data_out(wire_d14_5),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance150146(.data_in(wire_d14_5),.data_out(wire_d14_6),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance150147(.data_in(wire_d14_6),.data_out(wire_d14_7),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance150148(.data_in(wire_d14_7),.data_out(wire_d14_8),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance150149(.data_in(wire_d14_8),.data_out(wire_d14_9),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1501410(.data_in(wire_d14_9),.data_out(wire_d14_10),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1501411(.data_in(wire_d14_10),.data_out(wire_d14_11),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1501412(.data_in(wire_d14_11),.data_out(wire_d14_12),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1501413(.data_in(wire_d14_12),.data_out(wire_d14_13),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1501414(.data_in(wire_d14_13),.data_out(wire_d14_14),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1501415(.data_in(wire_d14_14),.data_out(wire_d14_15),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1501416(.data_in(wire_d14_15),.data_out(wire_d14_16),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1501417(.data_in(wire_d14_16),.data_out(wire_d14_17),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1501418(.data_in(wire_d14_17),.data_out(wire_d14_18),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1501419(.data_in(wire_d14_18),.data_out(wire_d14_19),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1501420(.data_in(wire_d14_19),.data_out(wire_d14_20),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1501421(.data_in(wire_d14_20),.data_out(wire_d14_21),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1501422(.data_in(wire_d14_21),.data_out(wire_d14_22),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1501423(.data_in(wire_d14_22),.data_out(wire_d14_23),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1501424(.data_in(wire_d14_23),.data_out(wire_d14_24),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1501425(.data_in(wire_d14_24),.data_out(wire_d14_25),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1501426(.data_in(wire_d14_25),.data_out(wire_d14_26),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1501427(.data_in(wire_d14_26),.data_out(wire_d14_27),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1501428(.data_in(wire_d14_27),.data_out(wire_d14_28),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1501429(.data_in(wire_d14_28),.data_out(wire_d14_29),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1501430(.data_in(wire_d14_29),.data_out(wire_d14_30),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1501431(.data_in(wire_d14_30),.data_out(wire_d14_31),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1501432(.data_in(wire_d14_31),.data_out(wire_d14_32),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1501433(.data_in(wire_d14_32),.data_out(wire_d14_33),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1501434(.data_in(wire_d14_33),.data_out(wire_d14_34),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1501435(.data_in(wire_d14_34),.data_out(wire_d14_35),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1501436(.data_in(wire_d14_35),.data_out(d_out14),.clk(clk),.rst(rst));

	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance160150(.data_in(d_in15),.data_out(wire_d15_0),.clk(clk),.rst(rst));            //channel 16
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance160151(.data_in(wire_d15_0),.data_out(wire_d15_1),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance160152(.data_in(wire_d15_1),.data_out(wire_d15_2),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance160153(.data_in(wire_d15_2),.data_out(wire_d15_3),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance160154(.data_in(wire_d15_3),.data_out(wire_d15_4),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance160155(.data_in(wire_d15_4),.data_out(wire_d15_5),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance160156(.data_in(wire_d15_5),.data_out(wire_d15_6),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance160157(.data_in(wire_d15_6),.data_out(wire_d15_7),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance160158(.data_in(wire_d15_7),.data_out(wire_d15_8),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance160159(.data_in(wire_d15_8),.data_out(wire_d15_9),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1601510(.data_in(wire_d15_9),.data_out(wire_d15_10),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1601511(.data_in(wire_d15_10),.data_out(wire_d15_11),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1601512(.data_in(wire_d15_11),.data_out(wire_d15_12),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1601513(.data_in(wire_d15_12),.data_out(wire_d15_13),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1601514(.data_in(wire_d15_13),.data_out(wire_d15_14),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1601515(.data_in(wire_d15_14),.data_out(wire_d15_15),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1601516(.data_in(wire_d15_15),.data_out(wire_d15_16),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1601517(.data_in(wire_d15_16),.data_out(wire_d15_17),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1601518(.data_in(wire_d15_17),.data_out(wire_d15_18),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1601519(.data_in(wire_d15_18),.data_out(wire_d15_19),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1601520(.data_in(wire_d15_19),.data_out(wire_d15_20),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1601521(.data_in(wire_d15_20),.data_out(wire_d15_21),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1601522(.data_in(wire_d15_21),.data_out(wire_d15_22),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1601523(.data_in(wire_d15_22),.data_out(wire_d15_23),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1601524(.data_in(wire_d15_23),.data_out(wire_d15_24),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1601525(.data_in(wire_d15_24),.data_out(wire_d15_25),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1601526(.data_in(wire_d15_25),.data_out(wire_d15_26),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1601527(.data_in(wire_d15_26),.data_out(wire_d15_27),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1601528(.data_in(wire_d15_27),.data_out(wire_d15_28),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1601529(.data_in(wire_d15_28),.data_out(wire_d15_29),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1601530(.data_in(wire_d15_29),.data_out(wire_d15_30),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1601531(.data_in(wire_d15_30),.data_out(wire_d15_31),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1601532(.data_in(wire_d15_31),.data_out(wire_d15_32),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1601533(.data_in(wire_d15_32),.data_out(wire_d15_33),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1601534(.data_in(wire_d15_33),.data_out(wire_d15_34),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1601535(.data_in(wire_d15_34),.data_out(wire_d15_35),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1601536(.data_in(wire_d15_35),.data_out(d_out15),.clk(clk),.rst(rst));

	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance170160(.data_in(d_in16),.data_out(wire_d16_0),.clk(clk),.rst(rst));            //channel 17
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance170161(.data_in(wire_d16_0),.data_out(wire_d16_1),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance170162(.data_in(wire_d16_1),.data_out(wire_d16_2),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance170163(.data_in(wire_d16_2),.data_out(wire_d16_3),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance170164(.data_in(wire_d16_3),.data_out(wire_d16_4),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance170165(.data_in(wire_d16_4),.data_out(wire_d16_5),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance170166(.data_in(wire_d16_5),.data_out(wire_d16_6),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance170167(.data_in(wire_d16_6),.data_out(wire_d16_7),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance170168(.data_in(wire_d16_7),.data_out(wire_d16_8),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance170169(.data_in(wire_d16_8),.data_out(wire_d16_9),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1701610(.data_in(wire_d16_9),.data_out(wire_d16_10),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1701611(.data_in(wire_d16_10),.data_out(wire_d16_11),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1701612(.data_in(wire_d16_11),.data_out(wire_d16_12),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1701613(.data_in(wire_d16_12),.data_out(wire_d16_13),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1701614(.data_in(wire_d16_13),.data_out(wire_d16_14),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1701615(.data_in(wire_d16_14),.data_out(wire_d16_15),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1701616(.data_in(wire_d16_15),.data_out(wire_d16_16),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1701617(.data_in(wire_d16_16),.data_out(wire_d16_17),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1701618(.data_in(wire_d16_17),.data_out(wire_d16_18),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1701619(.data_in(wire_d16_18),.data_out(wire_d16_19),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1701620(.data_in(wire_d16_19),.data_out(wire_d16_20),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1701621(.data_in(wire_d16_20),.data_out(wire_d16_21),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1701622(.data_in(wire_d16_21),.data_out(wire_d16_22),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1701623(.data_in(wire_d16_22),.data_out(wire_d16_23),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1701624(.data_in(wire_d16_23),.data_out(wire_d16_24),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1701625(.data_in(wire_d16_24),.data_out(wire_d16_25),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1701626(.data_in(wire_d16_25),.data_out(wire_d16_26),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1701627(.data_in(wire_d16_26),.data_out(wire_d16_27),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1701628(.data_in(wire_d16_27),.data_out(wire_d16_28),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1701629(.data_in(wire_d16_28),.data_out(wire_d16_29),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1701630(.data_in(wire_d16_29),.data_out(wire_d16_30),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1701631(.data_in(wire_d16_30),.data_out(wire_d16_31),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1701632(.data_in(wire_d16_31),.data_out(wire_d16_32),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1701633(.data_in(wire_d16_32),.data_out(wire_d16_33),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1701634(.data_in(wire_d16_33),.data_out(wire_d16_34),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1701635(.data_in(wire_d16_34),.data_out(wire_d16_35),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1701636(.data_in(wire_d16_35),.data_out(d_out16),.clk(clk),.rst(rst));

	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance180170(.data_in(d_in17),.data_out(wire_d17_0),.clk(clk),.rst(rst));            //channel 18
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance180171(.data_in(wire_d17_0),.data_out(wire_d17_1),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance180172(.data_in(wire_d17_1),.data_out(wire_d17_2),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance180173(.data_in(wire_d17_2),.data_out(wire_d17_3),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance180174(.data_in(wire_d17_3),.data_out(wire_d17_4),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance180175(.data_in(wire_d17_4),.data_out(wire_d17_5),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance180176(.data_in(wire_d17_5),.data_out(wire_d17_6),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance180177(.data_in(wire_d17_6),.data_out(wire_d17_7),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance180178(.data_in(wire_d17_7),.data_out(wire_d17_8),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance180179(.data_in(wire_d17_8),.data_out(wire_d17_9),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1801710(.data_in(wire_d17_9),.data_out(wire_d17_10),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1801711(.data_in(wire_d17_10),.data_out(wire_d17_11),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1801712(.data_in(wire_d17_11),.data_out(wire_d17_12),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1801713(.data_in(wire_d17_12),.data_out(wire_d17_13),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1801714(.data_in(wire_d17_13),.data_out(wire_d17_14),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1801715(.data_in(wire_d17_14),.data_out(wire_d17_15),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1801716(.data_in(wire_d17_15),.data_out(wire_d17_16),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1801717(.data_in(wire_d17_16),.data_out(wire_d17_17),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1801718(.data_in(wire_d17_17),.data_out(wire_d17_18),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1801719(.data_in(wire_d17_18),.data_out(wire_d17_19),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1801720(.data_in(wire_d17_19),.data_out(wire_d17_20),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1801721(.data_in(wire_d17_20),.data_out(wire_d17_21),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1801722(.data_in(wire_d17_21),.data_out(wire_d17_22),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1801723(.data_in(wire_d17_22),.data_out(wire_d17_23),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1801724(.data_in(wire_d17_23),.data_out(wire_d17_24),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1801725(.data_in(wire_d17_24),.data_out(wire_d17_25),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1801726(.data_in(wire_d17_25),.data_out(wire_d17_26),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1801727(.data_in(wire_d17_26),.data_out(wire_d17_27),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1801728(.data_in(wire_d17_27),.data_out(wire_d17_28),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1801729(.data_in(wire_d17_28),.data_out(wire_d17_29),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1801730(.data_in(wire_d17_29),.data_out(wire_d17_30),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1801731(.data_in(wire_d17_30),.data_out(wire_d17_31),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1801732(.data_in(wire_d17_31),.data_out(wire_d17_32),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1801733(.data_in(wire_d17_32),.data_out(wire_d17_33),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1801734(.data_in(wire_d17_33),.data_out(wire_d17_34),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1801735(.data_in(wire_d17_34),.data_out(wire_d17_35),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1801736(.data_in(wire_d17_35),.data_out(d_out17),.clk(clk),.rst(rst));

	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance190180(.data_in(d_in18),.data_out(wire_d18_0),.clk(clk),.rst(rst));            //channel 19
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance190181(.data_in(wire_d18_0),.data_out(wire_d18_1),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance190182(.data_in(wire_d18_1),.data_out(wire_d18_2),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance190183(.data_in(wire_d18_2),.data_out(wire_d18_3),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance190184(.data_in(wire_d18_3),.data_out(wire_d18_4),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance190185(.data_in(wire_d18_4),.data_out(wire_d18_5),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance190186(.data_in(wire_d18_5),.data_out(wire_d18_6),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance190187(.data_in(wire_d18_6),.data_out(wire_d18_7),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance190188(.data_in(wire_d18_7),.data_out(wire_d18_8),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance190189(.data_in(wire_d18_8),.data_out(wire_d18_9),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1901810(.data_in(wire_d18_9),.data_out(wire_d18_10),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1901811(.data_in(wire_d18_10),.data_out(wire_d18_11),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1901812(.data_in(wire_d18_11),.data_out(wire_d18_12),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1901813(.data_in(wire_d18_12),.data_out(wire_d18_13),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1901814(.data_in(wire_d18_13),.data_out(wire_d18_14),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1901815(.data_in(wire_d18_14),.data_out(wire_d18_15),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1901816(.data_in(wire_d18_15),.data_out(wire_d18_16),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1901817(.data_in(wire_d18_16),.data_out(wire_d18_17),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1901818(.data_in(wire_d18_17),.data_out(wire_d18_18),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1901819(.data_in(wire_d18_18),.data_out(wire_d18_19),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1901820(.data_in(wire_d18_19),.data_out(wire_d18_20),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1901821(.data_in(wire_d18_20),.data_out(wire_d18_21),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1901822(.data_in(wire_d18_21),.data_out(wire_d18_22),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance1901823(.data_in(wire_d18_22),.data_out(wire_d18_23),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1901824(.data_in(wire_d18_23),.data_out(wire_d18_24),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1901825(.data_in(wire_d18_24),.data_out(wire_d18_25),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1901826(.data_in(wire_d18_25),.data_out(wire_d18_26),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1901827(.data_in(wire_d18_26),.data_out(wire_d18_27),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1901828(.data_in(wire_d18_27),.data_out(wire_d18_28),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1901829(.data_in(wire_d18_28),.data_out(wire_d18_29),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1901830(.data_in(wire_d18_29),.data_out(wire_d18_30),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance1901831(.data_in(wire_d18_30),.data_out(wire_d18_31),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance1901832(.data_in(wire_d18_31),.data_out(wire_d18_32),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1901833(.data_in(wire_d18_32),.data_out(wire_d18_33),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance1901834(.data_in(wire_d18_33),.data_out(wire_d18_34),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance1901835(.data_in(wire_d18_34),.data_out(wire_d18_35),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance1901836(.data_in(wire_d18_35),.data_out(d_out18),.clk(clk),.rst(rst));

	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance200190(.data_in(d_in19),.data_out(wire_d19_0),.clk(clk),.rst(rst));            //channel 20
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance200191(.data_in(wire_d19_0),.data_out(wire_d19_1),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance200192(.data_in(wire_d19_1),.data_out(wire_d19_2),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance200193(.data_in(wire_d19_2),.data_out(wire_d19_3),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance200194(.data_in(wire_d19_3),.data_out(wire_d19_4),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance200195(.data_in(wire_d19_4),.data_out(wire_d19_5),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance200196(.data_in(wire_d19_5),.data_out(wire_d19_6),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance200197(.data_in(wire_d19_6),.data_out(wire_d19_7),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance200198(.data_in(wire_d19_7),.data_out(wire_d19_8),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance200199(.data_in(wire_d19_8),.data_out(wire_d19_9),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2001910(.data_in(wire_d19_9),.data_out(wire_d19_10),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2001911(.data_in(wire_d19_10),.data_out(wire_d19_11),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2001912(.data_in(wire_d19_11),.data_out(wire_d19_12),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2001913(.data_in(wire_d19_12),.data_out(wire_d19_13),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2001914(.data_in(wire_d19_13),.data_out(wire_d19_14),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2001915(.data_in(wire_d19_14),.data_out(wire_d19_15),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2001916(.data_in(wire_d19_15),.data_out(wire_d19_16),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2001917(.data_in(wire_d19_16),.data_out(wire_d19_17),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2001918(.data_in(wire_d19_17),.data_out(wire_d19_18),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2001919(.data_in(wire_d19_18),.data_out(wire_d19_19),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2001920(.data_in(wire_d19_19),.data_out(wire_d19_20),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2001921(.data_in(wire_d19_20),.data_out(wire_d19_21),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2001922(.data_in(wire_d19_21),.data_out(wire_d19_22),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2001923(.data_in(wire_d19_22),.data_out(wire_d19_23),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2001924(.data_in(wire_d19_23),.data_out(wire_d19_24),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2001925(.data_in(wire_d19_24),.data_out(wire_d19_25),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2001926(.data_in(wire_d19_25),.data_out(wire_d19_26),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2001927(.data_in(wire_d19_26),.data_out(wire_d19_27),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2001928(.data_in(wire_d19_27),.data_out(wire_d19_28),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2001929(.data_in(wire_d19_28),.data_out(wire_d19_29),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2001930(.data_in(wire_d19_29),.data_out(wire_d19_30),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2001931(.data_in(wire_d19_30),.data_out(wire_d19_31),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2001932(.data_in(wire_d19_31),.data_out(wire_d19_32),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2001933(.data_in(wire_d19_32),.data_out(wire_d19_33),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2001934(.data_in(wire_d19_33),.data_out(wire_d19_34),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2001935(.data_in(wire_d19_34),.data_out(wire_d19_35),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2001936(.data_in(wire_d19_35),.data_out(d_out19),.clk(clk),.rst(rst));

	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance210200(.data_in(d_in20),.data_out(wire_d20_0),.clk(clk),.rst(rst));            //channel 21
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance210201(.data_in(wire_d20_0),.data_out(wire_d20_1),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance210202(.data_in(wire_d20_1),.data_out(wire_d20_2),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance210203(.data_in(wire_d20_2),.data_out(wire_d20_3),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance210204(.data_in(wire_d20_3),.data_out(wire_d20_4),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance210205(.data_in(wire_d20_4),.data_out(wire_d20_5),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance210206(.data_in(wire_d20_5),.data_out(wire_d20_6),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance210207(.data_in(wire_d20_6),.data_out(wire_d20_7),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance210208(.data_in(wire_d20_7),.data_out(wire_d20_8),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance210209(.data_in(wire_d20_8),.data_out(wire_d20_9),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2102010(.data_in(wire_d20_9),.data_out(wire_d20_10),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2102011(.data_in(wire_d20_10),.data_out(wire_d20_11),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2102012(.data_in(wire_d20_11),.data_out(wire_d20_12),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2102013(.data_in(wire_d20_12),.data_out(wire_d20_13),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2102014(.data_in(wire_d20_13),.data_out(wire_d20_14),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2102015(.data_in(wire_d20_14),.data_out(wire_d20_15),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2102016(.data_in(wire_d20_15),.data_out(wire_d20_16),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2102017(.data_in(wire_d20_16),.data_out(wire_d20_17),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2102018(.data_in(wire_d20_17),.data_out(wire_d20_18),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2102019(.data_in(wire_d20_18),.data_out(wire_d20_19),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2102020(.data_in(wire_d20_19),.data_out(wire_d20_20),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2102021(.data_in(wire_d20_20),.data_out(wire_d20_21),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2102022(.data_in(wire_d20_21),.data_out(wire_d20_22),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2102023(.data_in(wire_d20_22),.data_out(wire_d20_23),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2102024(.data_in(wire_d20_23),.data_out(wire_d20_24),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2102025(.data_in(wire_d20_24),.data_out(wire_d20_25),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2102026(.data_in(wire_d20_25),.data_out(wire_d20_26),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2102027(.data_in(wire_d20_26),.data_out(wire_d20_27),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2102028(.data_in(wire_d20_27),.data_out(wire_d20_28),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2102029(.data_in(wire_d20_28),.data_out(wire_d20_29),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2102030(.data_in(wire_d20_29),.data_out(wire_d20_30),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2102031(.data_in(wire_d20_30),.data_out(wire_d20_31),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2102032(.data_in(wire_d20_31),.data_out(wire_d20_32),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2102033(.data_in(wire_d20_32),.data_out(wire_d20_33),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2102034(.data_in(wire_d20_33),.data_out(wire_d20_34),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2102035(.data_in(wire_d20_34),.data_out(wire_d20_35),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2102036(.data_in(wire_d20_35),.data_out(d_out20),.clk(clk),.rst(rst));

	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance220210(.data_in(d_in21),.data_out(wire_d21_0),.clk(clk),.rst(rst));            //channel 22
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance220211(.data_in(wire_d21_0),.data_out(wire_d21_1),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance220212(.data_in(wire_d21_1),.data_out(wire_d21_2),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance220213(.data_in(wire_d21_2),.data_out(wire_d21_3),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance220214(.data_in(wire_d21_3),.data_out(wire_d21_4),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance220215(.data_in(wire_d21_4),.data_out(wire_d21_5),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance220216(.data_in(wire_d21_5),.data_out(wire_d21_6),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance220217(.data_in(wire_d21_6),.data_out(wire_d21_7),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance220218(.data_in(wire_d21_7),.data_out(wire_d21_8),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance220219(.data_in(wire_d21_8),.data_out(wire_d21_9),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2202110(.data_in(wire_d21_9),.data_out(wire_d21_10),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2202111(.data_in(wire_d21_10),.data_out(wire_d21_11),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2202112(.data_in(wire_d21_11),.data_out(wire_d21_12),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2202113(.data_in(wire_d21_12),.data_out(wire_d21_13),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2202114(.data_in(wire_d21_13),.data_out(wire_d21_14),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2202115(.data_in(wire_d21_14),.data_out(wire_d21_15),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2202116(.data_in(wire_d21_15),.data_out(wire_d21_16),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2202117(.data_in(wire_d21_16),.data_out(wire_d21_17),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2202118(.data_in(wire_d21_17),.data_out(wire_d21_18),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2202119(.data_in(wire_d21_18),.data_out(wire_d21_19),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2202120(.data_in(wire_d21_19),.data_out(wire_d21_20),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2202121(.data_in(wire_d21_20),.data_out(wire_d21_21),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2202122(.data_in(wire_d21_21),.data_out(wire_d21_22),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2202123(.data_in(wire_d21_22),.data_out(wire_d21_23),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2202124(.data_in(wire_d21_23),.data_out(wire_d21_24),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2202125(.data_in(wire_d21_24),.data_out(wire_d21_25),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2202126(.data_in(wire_d21_25),.data_out(wire_d21_26),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2202127(.data_in(wire_d21_26),.data_out(wire_d21_27),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2202128(.data_in(wire_d21_27),.data_out(wire_d21_28),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2202129(.data_in(wire_d21_28),.data_out(wire_d21_29),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2202130(.data_in(wire_d21_29),.data_out(wire_d21_30),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2202131(.data_in(wire_d21_30),.data_out(wire_d21_31),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2202132(.data_in(wire_d21_31),.data_out(wire_d21_32),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2202133(.data_in(wire_d21_32),.data_out(wire_d21_33),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2202134(.data_in(wire_d21_33),.data_out(wire_d21_34),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2202135(.data_in(wire_d21_34),.data_out(wire_d21_35),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2202136(.data_in(wire_d21_35),.data_out(d_out21),.clk(clk),.rst(rst));

	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance230220(.data_in(d_in22),.data_out(wire_d22_0),.clk(clk),.rst(rst));            //channel 23
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance230221(.data_in(wire_d22_0),.data_out(wire_d22_1),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance230222(.data_in(wire_d22_1),.data_out(wire_d22_2),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance230223(.data_in(wire_d22_2),.data_out(wire_d22_3),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance230224(.data_in(wire_d22_3),.data_out(wire_d22_4),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance230225(.data_in(wire_d22_4),.data_out(wire_d22_5),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance230226(.data_in(wire_d22_5),.data_out(wire_d22_6),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance230227(.data_in(wire_d22_6),.data_out(wire_d22_7),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance230228(.data_in(wire_d22_7),.data_out(wire_d22_8),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance230229(.data_in(wire_d22_8),.data_out(wire_d22_9),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2302210(.data_in(wire_d22_9),.data_out(wire_d22_10),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2302211(.data_in(wire_d22_10),.data_out(wire_d22_11),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2302212(.data_in(wire_d22_11),.data_out(wire_d22_12),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2302213(.data_in(wire_d22_12),.data_out(wire_d22_13),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2302214(.data_in(wire_d22_13),.data_out(wire_d22_14),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2302215(.data_in(wire_d22_14),.data_out(wire_d22_15),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2302216(.data_in(wire_d22_15),.data_out(wire_d22_16),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2302217(.data_in(wire_d22_16),.data_out(wire_d22_17),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2302218(.data_in(wire_d22_17),.data_out(wire_d22_18),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2302219(.data_in(wire_d22_18),.data_out(wire_d22_19),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2302220(.data_in(wire_d22_19),.data_out(wire_d22_20),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2302221(.data_in(wire_d22_20),.data_out(wire_d22_21),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2302222(.data_in(wire_d22_21),.data_out(wire_d22_22),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2302223(.data_in(wire_d22_22),.data_out(wire_d22_23),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2302224(.data_in(wire_d22_23),.data_out(wire_d22_24),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2302225(.data_in(wire_d22_24),.data_out(wire_d22_25),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2302226(.data_in(wire_d22_25),.data_out(wire_d22_26),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2302227(.data_in(wire_d22_26),.data_out(wire_d22_27),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2302228(.data_in(wire_d22_27),.data_out(wire_d22_28),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2302229(.data_in(wire_d22_28),.data_out(wire_d22_29),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2302230(.data_in(wire_d22_29),.data_out(wire_d22_30),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2302231(.data_in(wire_d22_30),.data_out(wire_d22_31),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2302232(.data_in(wire_d22_31),.data_out(wire_d22_32),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2302233(.data_in(wire_d22_32),.data_out(wire_d22_33),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2302234(.data_in(wire_d22_33),.data_out(wire_d22_34),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2302235(.data_in(wire_d22_34),.data_out(wire_d22_35),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2302236(.data_in(wire_d22_35),.data_out(d_out22),.clk(clk),.rst(rst));

	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance240230(.data_in(d_in23),.data_out(wire_d23_0),.clk(clk),.rst(rst));            //channel 24
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance240231(.data_in(wire_d23_0),.data_out(wire_d23_1),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance240232(.data_in(wire_d23_1),.data_out(wire_d23_2),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance240233(.data_in(wire_d23_2),.data_out(wire_d23_3),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance240234(.data_in(wire_d23_3),.data_out(wire_d23_4),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance240235(.data_in(wire_d23_4),.data_out(wire_d23_5),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance240236(.data_in(wire_d23_5),.data_out(wire_d23_6),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance240237(.data_in(wire_d23_6),.data_out(wire_d23_7),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance240238(.data_in(wire_d23_7),.data_out(wire_d23_8),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance240239(.data_in(wire_d23_8),.data_out(wire_d23_9),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2402310(.data_in(wire_d23_9),.data_out(wire_d23_10),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2402311(.data_in(wire_d23_10),.data_out(wire_d23_11),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2402312(.data_in(wire_d23_11),.data_out(wire_d23_12),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2402313(.data_in(wire_d23_12),.data_out(wire_d23_13),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2402314(.data_in(wire_d23_13),.data_out(wire_d23_14),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2402315(.data_in(wire_d23_14),.data_out(wire_d23_15),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2402316(.data_in(wire_d23_15),.data_out(wire_d23_16),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2402317(.data_in(wire_d23_16),.data_out(wire_d23_17),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2402318(.data_in(wire_d23_17),.data_out(wire_d23_18),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2402319(.data_in(wire_d23_18),.data_out(wire_d23_19),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2402320(.data_in(wire_d23_19),.data_out(wire_d23_20),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2402321(.data_in(wire_d23_20),.data_out(wire_d23_21),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2402322(.data_in(wire_d23_21),.data_out(wire_d23_22),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2402323(.data_in(wire_d23_22),.data_out(wire_d23_23),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2402324(.data_in(wire_d23_23),.data_out(wire_d23_24),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2402325(.data_in(wire_d23_24),.data_out(wire_d23_25),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2402326(.data_in(wire_d23_25),.data_out(wire_d23_26),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2402327(.data_in(wire_d23_26),.data_out(wire_d23_27),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2402328(.data_in(wire_d23_27),.data_out(wire_d23_28),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2402329(.data_in(wire_d23_28),.data_out(wire_d23_29),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2402330(.data_in(wire_d23_29),.data_out(wire_d23_30),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2402331(.data_in(wire_d23_30),.data_out(wire_d23_31),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2402332(.data_in(wire_d23_31),.data_out(wire_d23_32),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2402333(.data_in(wire_d23_32),.data_out(wire_d23_33),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2402334(.data_in(wire_d23_33),.data_out(wire_d23_34),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2402335(.data_in(wire_d23_34),.data_out(wire_d23_35),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2402336(.data_in(wire_d23_35),.data_out(d_out23),.clk(clk),.rst(rst));

	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance250240(.data_in(d_in24),.data_out(wire_d24_0),.clk(clk),.rst(rst));            //channel 25
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance250241(.data_in(wire_d24_0),.data_out(wire_d24_1),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance250242(.data_in(wire_d24_1),.data_out(wire_d24_2),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance250243(.data_in(wire_d24_2),.data_out(wire_d24_3),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance250244(.data_in(wire_d24_3),.data_out(wire_d24_4),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance250245(.data_in(wire_d24_4),.data_out(wire_d24_5),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance250246(.data_in(wire_d24_5),.data_out(wire_d24_6),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance250247(.data_in(wire_d24_6),.data_out(wire_d24_7),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance250248(.data_in(wire_d24_7),.data_out(wire_d24_8),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance250249(.data_in(wire_d24_8),.data_out(wire_d24_9),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2502410(.data_in(wire_d24_9),.data_out(wire_d24_10),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2502411(.data_in(wire_d24_10),.data_out(wire_d24_11),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2502412(.data_in(wire_d24_11),.data_out(wire_d24_12),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2502413(.data_in(wire_d24_12),.data_out(wire_d24_13),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2502414(.data_in(wire_d24_13),.data_out(wire_d24_14),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2502415(.data_in(wire_d24_14),.data_out(wire_d24_15),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2502416(.data_in(wire_d24_15),.data_out(wire_d24_16),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2502417(.data_in(wire_d24_16),.data_out(wire_d24_17),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2502418(.data_in(wire_d24_17),.data_out(wire_d24_18),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2502419(.data_in(wire_d24_18),.data_out(wire_d24_19),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2502420(.data_in(wire_d24_19),.data_out(wire_d24_20),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2502421(.data_in(wire_d24_20),.data_out(wire_d24_21),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2502422(.data_in(wire_d24_21),.data_out(wire_d24_22),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2502423(.data_in(wire_d24_22),.data_out(wire_d24_23),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2502424(.data_in(wire_d24_23),.data_out(wire_d24_24),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2502425(.data_in(wire_d24_24),.data_out(wire_d24_25),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2502426(.data_in(wire_d24_25),.data_out(wire_d24_26),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2502427(.data_in(wire_d24_26),.data_out(wire_d24_27),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2502428(.data_in(wire_d24_27),.data_out(wire_d24_28),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2502429(.data_in(wire_d24_28),.data_out(wire_d24_29),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2502430(.data_in(wire_d24_29),.data_out(wire_d24_30),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2502431(.data_in(wire_d24_30),.data_out(wire_d24_31),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2502432(.data_in(wire_d24_31),.data_out(wire_d24_32),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2502433(.data_in(wire_d24_32),.data_out(wire_d24_33),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2502434(.data_in(wire_d24_33),.data_out(wire_d24_34),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2502435(.data_in(wire_d24_34),.data_out(wire_d24_35),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2502436(.data_in(wire_d24_35),.data_out(d_out24),.clk(clk),.rst(rst));

	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance260250(.data_in(d_in25),.data_out(wire_d25_0),.clk(clk),.rst(rst));            //channel 26
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance260251(.data_in(wire_d25_0),.data_out(wire_d25_1),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance260252(.data_in(wire_d25_1),.data_out(wire_d25_2),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance260253(.data_in(wire_d25_2),.data_out(wire_d25_3),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance260254(.data_in(wire_d25_3),.data_out(wire_d25_4),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance260255(.data_in(wire_d25_4),.data_out(wire_d25_5),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance260256(.data_in(wire_d25_5),.data_out(wire_d25_6),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance260257(.data_in(wire_d25_6),.data_out(wire_d25_7),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance260258(.data_in(wire_d25_7),.data_out(wire_d25_8),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance260259(.data_in(wire_d25_8),.data_out(wire_d25_9),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2602510(.data_in(wire_d25_9),.data_out(wire_d25_10),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2602511(.data_in(wire_d25_10),.data_out(wire_d25_11),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2602512(.data_in(wire_d25_11),.data_out(wire_d25_12),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2602513(.data_in(wire_d25_12),.data_out(wire_d25_13),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2602514(.data_in(wire_d25_13),.data_out(wire_d25_14),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2602515(.data_in(wire_d25_14),.data_out(wire_d25_15),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2602516(.data_in(wire_d25_15),.data_out(wire_d25_16),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2602517(.data_in(wire_d25_16),.data_out(wire_d25_17),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2602518(.data_in(wire_d25_17),.data_out(wire_d25_18),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2602519(.data_in(wire_d25_18),.data_out(wire_d25_19),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2602520(.data_in(wire_d25_19),.data_out(wire_d25_20),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2602521(.data_in(wire_d25_20),.data_out(wire_d25_21),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2602522(.data_in(wire_d25_21),.data_out(wire_d25_22),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2602523(.data_in(wire_d25_22),.data_out(wire_d25_23),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2602524(.data_in(wire_d25_23),.data_out(wire_d25_24),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2602525(.data_in(wire_d25_24),.data_out(wire_d25_25),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2602526(.data_in(wire_d25_25),.data_out(wire_d25_26),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2602527(.data_in(wire_d25_26),.data_out(wire_d25_27),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2602528(.data_in(wire_d25_27),.data_out(wire_d25_28),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2602529(.data_in(wire_d25_28),.data_out(wire_d25_29),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2602530(.data_in(wire_d25_29),.data_out(wire_d25_30),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2602531(.data_in(wire_d25_30),.data_out(wire_d25_31),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2602532(.data_in(wire_d25_31),.data_out(wire_d25_32),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2602533(.data_in(wire_d25_32),.data_out(wire_d25_33),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2602534(.data_in(wire_d25_33),.data_out(wire_d25_34),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2602535(.data_in(wire_d25_34),.data_out(wire_d25_35),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2602536(.data_in(wire_d25_35),.data_out(d_out25),.clk(clk),.rst(rst));

	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance270260(.data_in(d_in26),.data_out(wire_d26_0),.clk(clk),.rst(rst));            //channel 27
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance270261(.data_in(wire_d26_0),.data_out(wire_d26_1),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance270262(.data_in(wire_d26_1),.data_out(wire_d26_2),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance270263(.data_in(wire_d26_2),.data_out(wire_d26_3),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance270264(.data_in(wire_d26_3),.data_out(wire_d26_4),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance270265(.data_in(wire_d26_4),.data_out(wire_d26_5),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance270266(.data_in(wire_d26_5),.data_out(wire_d26_6),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance270267(.data_in(wire_d26_6),.data_out(wire_d26_7),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance270268(.data_in(wire_d26_7),.data_out(wire_d26_8),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance270269(.data_in(wire_d26_8),.data_out(wire_d26_9),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2702610(.data_in(wire_d26_9),.data_out(wire_d26_10),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2702611(.data_in(wire_d26_10),.data_out(wire_d26_11),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2702612(.data_in(wire_d26_11),.data_out(wire_d26_12),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2702613(.data_in(wire_d26_12),.data_out(wire_d26_13),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2702614(.data_in(wire_d26_13),.data_out(wire_d26_14),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2702615(.data_in(wire_d26_14),.data_out(wire_d26_15),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2702616(.data_in(wire_d26_15),.data_out(wire_d26_16),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2702617(.data_in(wire_d26_16),.data_out(wire_d26_17),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2702618(.data_in(wire_d26_17),.data_out(wire_d26_18),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2702619(.data_in(wire_d26_18),.data_out(wire_d26_19),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2702620(.data_in(wire_d26_19),.data_out(wire_d26_20),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2702621(.data_in(wire_d26_20),.data_out(wire_d26_21),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2702622(.data_in(wire_d26_21),.data_out(wire_d26_22),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2702623(.data_in(wire_d26_22),.data_out(wire_d26_23),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2702624(.data_in(wire_d26_23),.data_out(wire_d26_24),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2702625(.data_in(wire_d26_24),.data_out(wire_d26_25),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2702626(.data_in(wire_d26_25),.data_out(wire_d26_26),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2702627(.data_in(wire_d26_26),.data_out(wire_d26_27),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2702628(.data_in(wire_d26_27),.data_out(wire_d26_28),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2702629(.data_in(wire_d26_28),.data_out(wire_d26_29),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2702630(.data_in(wire_d26_29),.data_out(wire_d26_30),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2702631(.data_in(wire_d26_30),.data_out(wire_d26_31),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2702632(.data_in(wire_d26_31),.data_out(wire_d26_32),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2702633(.data_in(wire_d26_32),.data_out(wire_d26_33),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2702634(.data_in(wire_d26_33),.data_out(wire_d26_34),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2702635(.data_in(wire_d26_34),.data_out(wire_d26_35),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2702636(.data_in(wire_d26_35),.data_out(d_out26),.clk(clk),.rst(rst));

	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance280270(.data_in(d_in27),.data_out(wire_d27_0),.clk(clk),.rst(rst));            //channel 28
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance280271(.data_in(wire_d27_0),.data_out(wire_d27_1),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance280272(.data_in(wire_d27_1),.data_out(wire_d27_2),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance280273(.data_in(wire_d27_2),.data_out(wire_d27_3),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance280274(.data_in(wire_d27_3),.data_out(wire_d27_4),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance280275(.data_in(wire_d27_4),.data_out(wire_d27_5),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance280276(.data_in(wire_d27_5),.data_out(wire_d27_6),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance280277(.data_in(wire_d27_6),.data_out(wire_d27_7),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance280278(.data_in(wire_d27_7),.data_out(wire_d27_8),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance280279(.data_in(wire_d27_8),.data_out(wire_d27_9),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2802710(.data_in(wire_d27_9),.data_out(wire_d27_10),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2802711(.data_in(wire_d27_10),.data_out(wire_d27_11),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2802712(.data_in(wire_d27_11),.data_out(wire_d27_12),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2802713(.data_in(wire_d27_12),.data_out(wire_d27_13),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2802714(.data_in(wire_d27_13),.data_out(wire_d27_14),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2802715(.data_in(wire_d27_14),.data_out(wire_d27_15),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2802716(.data_in(wire_d27_15),.data_out(wire_d27_16),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2802717(.data_in(wire_d27_16),.data_out(wire_d27_17),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2802718(.data_in(wire_d27_17),.data_out(wire_d27_18),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2802719(.data_in(wire_d27_18),.data_out(wire_d27_19),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2802720(.data_in(wire_d27_19),.data_out(wire_d27_20),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2802721(.data_in(wire_d27_20),.data_out(wire_d27_21),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2802722(.data_in(wire_d27_21),.data_out(wire_d27_22),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2802723(.data_in(wire_d27_22),.data_out(wire_d27_23),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2802724(.data_in(wire_d27_23),.data_out(wire_d27_24),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2802725(.data_in(wire_d27_24),.data_out(wire_d27_25),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2802726(.data_in(wire_d27_25),.data_out(wire_d27_26),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2802727(.data_in(wire_d27_26),.data_out(wire_d27_27),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2802728(.data_in(wire_d27_27),.data_out(wire_d27_28),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2802729(.data_in(wire_d27_28),.data_out(wire_d27_29),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2802730(.data_in(wire_d27_29),.data_out(wire_d27_30),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2802731(.data_in(wire_d27_30),.data_out(wire_d27_31),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2802732(.data_in(wire_d27_31),.data_out(wire_d27_32),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2802733(.data_in(wire_d27_32),.data_out(wire_d27_33),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2802734(.data_in(wire_d27_33),.data_out(wire_d27_34),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2802735(.data_in(wire_d27_34),.data_out(wire_d27_35),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2802736(.data_in(wire_d27_35),.data_out(d_out27),.clk(clk),.rst(rst));

	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance290280(.data_in(d_in28),.data_out(wire_d28_0),.clk(clk),.rst(rst));            //channel 29
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance290281(.data_in(wire_d28_0),.data_out(wire_d28_1),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance290282(.data_in(wire_d28_1),.data_out(wire_d28_2),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance290283(.data_in(wire_d28_2),.data_out(wire_d28_3),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance290284(.data_in(wire_d28_3),.data_out(wire_d28_4),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance290285(.data_in(wire_d28_4),.data_out(wire_d28_5),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance290286(.data_in(wire_d28_5),.data_out(wire_d28_6),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance290287(.data_in(wire_d28_6),.data_out(wire_d28_7),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance290288(.data_in(wire_d28_7),.data_out(wire_d28_8),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance290289(.data_in(wire_d28_8),.data_out(wire_d28_9),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2902810(.data_in(wire_d28_9),.data_out(wire_d28_10),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2902811(.data_in(wire_d28_10),.data_out(wire_d28_11),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2902812(.data_in(wire_d28_11),.data_out(wire_d28_12),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2902813(.data_in(wire_d28_12),.data_out(wire_d28_13),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2902814(.data_in(wire_d28_13),.data_out(wire_d28_14),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2902815(.data_in(wire_d28_14),.data_out(wire_d28_15),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2902816(.data_in(wire_d28_15),.data_out(wire_d28_16),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2902817(.data_in(wire_d28_16),.data_out(wire_d28_17),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2902818(.data_in(wire_d28_17),.data_out(wire_d28_18),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2902819(.data_in(wire_d28_18),.data_out(wire_d28_19),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2902820(.data_in(wire_d28_19),.data_out(wire_d28_20),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2902821(.data_in(wire_d28_20),.data_out(wire_d28_21),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance2902822(.data_in(wire_d28_21),.data_out(wire_d28_22),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2902823(.data_in(wire_d28_22),.data_out(wire_d28_23),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2902824(.data_in(wire_d28_23),.data_out(wire_d28_24),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2902825(.data_in(wire_d28_24),.data_out(wire_d28_25),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2902826(.data_in(wire_d28_25),.data_out(wire_d28_26),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2902827(.data_in(wire_d28_26),.data_out(wire_d28_27),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2902828(.data_in(wire_d28_27),.data_out(wire_d28_28),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance2902829(.data_in(wire_d28_28),.data_out(wire_d28_29),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance2902830(.data_in(wire_d28_29),.data_out(wire_d28_30),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2902831(.data_in(wire_d28_30),.data_out(wire_d28_31),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance2902832(.data_in(wire_d28_31),.data_out(wire_d28_32),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2902833(.data_in(wire_d28_32),.data_out(wire_d28_33),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2902834(.data_in(wire_d28_33),.data_out(wire_d28_34),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance2902835(.data_in(wire_d28_34),.data_out(wire_d28_35),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance2902836(.data_in(wire_d28_35),.data_out(d_out28),.clk(clk),.rst(rst));

	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance300290(.data_in(d_in29),.data_out(wire_d29_0),.clk(clk),.rst(rst));            //channel 30
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance300291(.data_in(wire_d29_0),.data_out(wire_d29_1),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance300292(.data_in(wire_d29_1),.data_out(wire_d29_2),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance300293(.data_in(wire_d29_2),.data_out(wire_d29_3),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance300294(.data_in(wire_d29_3),.data_out(wire_d29_4),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance300295(.data_in(wire_d29_4),.data_out(wire_d29_5),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance300296(.data_in(wire_d29_5),.data_out(wire_d29_6),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance300297(.data_in(wire_d29_6),.data_out(wire_d29_7),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance300298(.data_in(wire_d29_7),.data_out(wire_d29_8),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance300299(.data_in(wire_d29_8),.data_out(wire_d29_9),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3002910(.data_in(wire_d29_9),.data_out(wire_d29_10),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3002911(.data_in(wire_d29_10),.data_out(wire_d29_11),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3002912(.data_in(wire_d29_11),.data_out(wire_d29_12),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3002913(.data_in(wire_d29_12),.data_out(wire_d29_13),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3002914(.data_in(wire_d29_13),.data_out(wire_d29_14),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3002915(.data_in(wire_d29_14),.data_out(wire_d29_15),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3002916(.data_in(wire_d29_15),.data_out(wire_d29_16),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3002917(.data_in(wire_d29_16),.data_out(wire_d29_17),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3002918(.data_in(wire_d29_17),.data_out(wire_d29_18),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3002919(.data_in(wire_d29_18),.data_out(wire_d29_19),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3002920(.data_in(wire_d29_19),.data_out(wire_d29_20),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3002921(.data_in(wire_d29_20),.data_out(wire_d29_21),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3002922(.data_in(wire_d29_21),.data_out(wire_d29_22),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3002923(.data_in(wire_d29_22),.data_out(wire_d29_23),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3002924(.data_in(wire_d29_23),.data_out(wire_d29_24),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3002925(.data_in(wire_d29_24),.data_out(wire_d29_25),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3002926(.data_in(wire_d29_25),.data_out(wire_d29_26),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3002927(.data_in(wire_d29_26),.data_out(wire_d29_27),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3002928(.data_in(wire_d29_27),.data_out(wire_d29_28),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3002929(.data_in(wire_d29_28),.data_out(wire_d29_29),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3002930(.data_in(wire_d29_29),.data_out(wire_d29_30),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3002931(.data_in(wire_d29_30),.data_out(wire_d29_31),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3002932(.data_in(wire_d29_31),.data_out(wire_d29_32),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3002933(.data_in(wire_d29_32),.data_out(wire_d29_33),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3002934(.data_in(wire_d29_33),.data_out(wire_d29_34),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3002935(.data_in(wire_d29_34),.data_out(wire_d29_35),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3002936(.data_in(wire_d29_35),.data_out(d_out29),.clk(clk),.rst(rst));

	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance310300(.data_in(d_in30),.data_out(wire_d30_0),.clk(clk),.rst(rst));            //channel 31
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance310301(.data_in(wire_d30_0),.data_out(wire_d30_1),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance310302(.data_in(wire_d30_1),.data_out(wire_d30_2),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance310303(.data_in(wire_d30_2),.data_out(wire_d30_3),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance310304(.data_in(wire_d30_3),.data_out(wire_d30_4),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance310305(.data_in(wire_d30_4),.data_out(wire_d30_5),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance310306(.data_in(wire_d30_5),.data_out(wire_d30_6),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance310307(.data_in(wire_d30_6),.data_out(wire_d30_7),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance310308(.data_in(wire_d30_7),.data_out(wire_d30_8),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance310309(.data_in(wire_d30_8),.data_out(wire_d30_9),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3103010(.data_in(wire_d30_9),.data_out(wire_d30_10),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3103011(.data_in(wire_d30_10),.data_out(wire_d30_11),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3103012(.data_in(wire_d30_11),.data_out(wire_d30_12),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3103013(.data_in(wire_d30_12),.data_out(wire_d30_13),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3103014(.data_in(wire_d30_13),.data_out(wire_d30_14),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3103015(.data_in(wire_d30_14),.data_out(wire_d30_15),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3103016(.data_in(wire_d30_15),.data_out(wire_d30_16),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3103017(.data_in(wire_d30_16),.data_out(wire_d30_17),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3103018(.data_in(wire_d30_17),.data_out(wire_d30_18),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3103019(.data_in(wire_d30_18),.data_out(wire_d30_19),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3103020(.data_in(wire_d30_19),.data_out(wire_d30_20),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3103021(.data_in(wire_d30_20),.data_out(wire_d30_21),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3103022(.data_in(wire_d30_21),.data_out(wire_d30_22),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3103023(.data_in(wire_d30_22),.data_out(wire_d30_23),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3103024(.data_in(wire_d30_23),.data_out(wire_d30_24),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3103025(.data_in(wire_d30_24),.data_out(wire_d30_25),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3103026(.data_in(wire_d30_25),.data_out(wire_d30_26),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3103027(.data_in(wire_d30_26),.data_out(wire_d30_27),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3103028(.data_in(wire_d30_27),.data_out(wire_d30_28),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3103029(.data_in(wire_d30_28),.data_out(wire_d30_29),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3103030(.data_in(wire_d30_29),.data_out(wire_d30_30),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3103031(.data_in(wire_d30_30),.data_out(wire_d30_31),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3103032(.data_in(wire_d30_31),.data_out(wire_d30_32),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3103033(.data_in(wire_d30_32),.data_out(wire_d30_33),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3103034(.data_in(wire_d30_33),.data_out(wire_d30_34),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3103035(.data_in(wire_d30_34),.data_out(wire_d30_35),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3103036(.data_in(wire_d30_35),.data_out(d_out30),.clk(clk),.rst(rst));

	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance320310(.data_in(d_in31),.data_out(wire_d31_0),.clk(clk),.rst(rst));            //channel 32
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance320311(.data_in(wire_d31_0),.data_out(wire_d31_1),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance320312(.data_in(wire_d31_1),.data_out(wire_d31_2),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance320313(.data_in(wire_d31_2),.data_out(wire_d31_3),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance320314(.data_in(wire_d31_3),.data_out(wire_d31_4),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance320315(.data_in(wire_d31_4),.data_out(wire_d31_5),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance320316(.data_in(wire_d31_5),.data_out(wire_d31_6),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance320317(.data_in(wire_d31_6),.data_out(wire_d31_7),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance320318(.data_in(wire_d31_7),.data_out(wire_d31_8),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance320319(.data_in(wire_d31_8),.data_out(wire_d31_9),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3203110(.data_in(wire_d31_9),.data_out(wire_d31_10),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3203111(.data_in(wire_d31_10),.data_out(wire_d31_11),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3203112(.data_in(wire_d31_11),.data_out(wire_d31_12),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3203113(.data_in(wire_d31_12),.data_out(wire_d31_13),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3203114(.data_in(wire_d31_13),.data_out(wire_d31_14),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3203115(.data_in(wire_d31_14),.data_out(wire_d31_15),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3203116(.data_in(wire_d31_15),.data_out(wire_d31_16),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3203117(.data_in(wire_d31_16),.data_out(wire_d31_17),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3203118(.data_in(wire_d31_17),.data_out(wire_d31_18),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3203119(.data_in(wire_d31_18),.data_out(wire_d31_19),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3203120(.data_in(wire_d31_19),.data_out(wire_d31_20),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3203121(.data_in(wire_d31_20),.data_out(wire_d31_21),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3203122(.data_in(wire_d31_21),.data_out(wire_d31_22),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3203123(.data_in(wire_d31_22),.data_out(wire_d31_23),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3203124(.data_in(wire_d31_23),.data_out(wire_d31_24),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3203125(.data_in(wire_d31_24),.data_out(wire_d31_25),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3203126(.data_in(wire_d31_25),.data_out(wire_d31_26),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3203127(.data_in(wire_d31_26),.data_out(wire_d31_27),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3203128(.data_in(wire_d31_27),.data_out(wire_d31_28),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3203129(.data_in(wire_d31_28),.data_out(wire_d31_29),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3203130(.data_in(wire_d31_29),.data_out(wire_d31_30),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3203131(.data_in(wire_d31_30),.data_out(wire_d31_31),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3203132(.data_in(wire_d31_31),.data_out(wire_d31_32),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3203133(.data_in(wire_d31_32),.data_out(wire_d31_33),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3203134(.data_in(wire_d31_33),.data_out(wire_d31_34),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3203135(.data_in(wire_d31_34),.data_out(wire_d31_35),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3203136(.data_in(wire_d31_35),.data_out(d_out31),.clk(clk),.rst(rst));

	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance330320(.data_in(d_in32),.data_out(wire_d32_0),.clk(clk),.rst(rst));            //channel 33
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance330321(.data_in(wire_d32_0),.data_out(wire_d32_1),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance330322(.data_in(wire_d32_1),.data_out(wire_d32_2),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance330323(.data_in(wire_d32_2),.data_out(wire_d32_3),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance330324(.data_in(wire_d32_3),.data_out(wire_d32_4),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance330325(.data_in(wire_d32_4),.data_out(wire_d32_5),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance330326(.data_in(wire_d32_5),.data_out(wire_d32_6),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance330327(.data_in(wire_d32_6),.data_out(wire_d32_7),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance330328(.data_in(wire_d32_7),.data_out(wire_d32_8),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance330329(.data_in(wire_d32_8),.data_out(wire_d32_9),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3303210(.data_in(wire_d32_9),.data_out(wire_d32_10),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3303211(.data_in(wire_d32_10),.data_out(wire_d32_11),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3303212(.data_in(wire_d32_11),.data_out(wire_d32_12),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3303213(.data_in(wire_d32_12),.data_out(wire_d32_13),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3303214(.data_in(wire_d32_13),.data_out(wire_d32_14),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3303215(.data_in(wire_d32_14),.data_out(wire_d32_15),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3303216(.data_in(wire_d32_15),.data_out(wire_d32_16),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3303217(.data_in(wire_d32_16),.data_out(wire_d32_17),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3303218(.data_in(wire_d32_17),.data_out(wire_d32_18),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3303219(.data_in(wire_d32_18),.data_out(wire_d32_19),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3303220(.data_in(wire_d32_19),.data_out(wire_d32_20),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3303221(.data_in(wire_d32_20),.data_out(wire_d32_21),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3303222(.data_in(wire_d32_21),.data_out(wire_d32_22),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3303223(.data_in(wire_d32_22),.data_out(wire_d32_23),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3303224(.data_in(wire_d32_23),.data_out(wire_d32_24),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3303225(.data_in(wire_d32_24),.data_out(wire_d32_25),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3303226(.data_in(wire_d32_25),.data_out(wire_d32_26),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3303227(.data_in(wire_d32_26),.data_out(wire_d32_27),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3303228(.data_in(wire_d32_27),.data_out(wire_d32_28),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3303229(.data_in(wire_d32_28),.data_out(wire_d32_29),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3303230(.data_in(wire_d32_29),.data_out(wire_d32_30),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3303231(.data_in(wire_d32_30),.data_out(wire_d32_31),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3303232(.data_in(wire_d32_31),.data_out(wire_d32_32),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3303233(.data_in(wire_d32_32),.data_out(wire_d32_33),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3303234(.data_in(wire_d32_33),.data_out(wire_d32_34),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3303235(.data_in(wire_d32_34),.data_out(wire_d32_35),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3303236(.data_in(wire_d32_35),.data_out(d_out32),.clk(clk),.rst(rst));

	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance340330(.data_in(d_in33),.data_out(wire_d33_0),.clk(clk),.rst(rst));            //channel 34
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance340331(.data_in(wire_d33_0),.data_out(wire_d33_1),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance340332(.data_in(wire_d33_1),.data_out(wire_d33_2),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance340333(.data_in(wire_d33_2),.data_out(wire_d33_3),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance340334(.data_in(wire_d33_3),.data_out(wire_d33_4),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance340335(.data_in(wire_d33_4),.data_out(wire_d33_5),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance340336(.data_in(wire_d33_5),.data_out(wire_d33_6),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance340337(.data_in(wire_d33_6),.data_out(wire_d33_7),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance340338(.data_in(wire_d33_7),.data_out(wire_d33_8),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance340339(.data_in(wire_d33_8),.data_out(wire_d33_9),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3403310(.data_in(wire_d33_9),.data_out(wire_d33_10),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3403311(.data_in(wire_d33_10),.data_out(wire_d33_11),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3403312(.data_in(wire_d33_11),.data_out(wire_d33_12),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3403313(.data_in(wire_d33_12),.data_out(wire_d33_13),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3403314(.data_in(wire_d33_13),.data_out(wire_d33_14),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3403315(.data_in(wire_d33_14),.data_out(wire_d33_15),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3403316(.data_in(wire_d33_15),.data_out(wire_d33_16),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3403317(.data_in(wire_d33_16),.data_out(wire_d33_17),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3403318(.data_in(wire_d33_17),.data_out(wire_d33_18),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3403319(.data_in(wire_d33_18),.data_out(wire_d33_19),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3403320(.data_in(wire_d33_19),.data_out(wire_d33_20),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3403321(.data_in(wire_d33_20),.data_out(wire_d33_21),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3403322(.data_in(wire_d33_21),.data_out(wire_d33_22),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3403323(.data_in(wire_d33_22),.data_out(wire_d33_23),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3403324(.data_in(wire_d33_23),.data_out(wire_d33_24),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3403325(.data_in(wire_d33_24),.data_out(wire_d33_25),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3403326(.data_in(wire_d33_25),.data_out(wire_d33_26),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3403327(.data_in(wire_d33_26),.data_out(wire_d33_27),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3403328(.data_in(wire_d33_27),.data_out(wire_d33_28),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3403329(.data_in(wire_d33_28),.data_out(wire_d33_29),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3403330(.data_in(wire_d33_29),.data_out(wire_d33_30),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3403331(.data_in(wire_d33_30),.data_out(wire_d33_31),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3403332(.data_in(wire_d33_31),.data_out(wire_d33_32),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3403333(.data_in(wire_d33_32),.data_out(wire_d33_33),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3403334(.data_in(wire_d33_33),.data_out(wire_d33_34),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3403335(.data_in(wire_d33_34),.data_out(wire_d33_35),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3403336(.data_in(wire_d33_35),.data_out(d_out33),.clk(clk),.rst(rst));

	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance350340(.data_in(d_in34),.data_out(wire_d34_0),.clk(clk),.rst(rst));            //channel 35
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance350341(.data_in(wire_d34_0),.data_out(wire_d34_1),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance350342(.data_in(wire_d34_1),.data_out(wire_d34_2),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance350343(.data_in(wire_d34_2),.data_out(wire_d34_3),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance350344(.data_in(wire_d34_3),.data_out(wire_d34_4),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance350345(.data_in(wire_d34_4),.data_out(wire_d34_5),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance350346(.data_in(wire_d34_5),.data_out(wire_d34_6),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance350347(.data_in(wire_d34_6),.data_out(wire_d34_7),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance350348(.data_in(wire_d34_7),.data_out(wire_d34_8),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance350349(.data_in(wire_d34_8),.data_out(wire_d34_9),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3503410(.data_in(wire_d34_9),.data_out(wire_d34_10),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3503411(.data_in(wire_d34_10),.data_out(wire_d34_11),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3503412(.data_in(wire_d34_11),.data_out(wire_d34_12),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3503413(.data_in(wire_d34_12),.data_out(wire_d34_13),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3503414(.data_in(wire_d34_13),.data_out(wire_d34_14),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3503415(.data_in(wire_d34_14),.data_out(wire_d34_15),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3503416(.data_in(wire_d34_15),.data_out(wire_d34_16),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3503417(.data_in(wire_d34_16),.data_out(wire_d34_17),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3503418(.data_in(wire_d34_17),.data_out(wire_d34_18),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3503419(.data_in(wire_d34_18),.data_out(wire_d34_19),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3503420(.data_in(wire_d34_19),.data_out(wire_d34_20),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3503421(.data_in(wire_d34_20),.data_out(wire_d34_21),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3503422(.data_in(wire_d34_21),.data_out(wire_d34_22),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3503423(.data_in(wire_d34_22),.data_out(wire_d34_23),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3503424(.data_in(wire_d34_23),.data_out(wire_d34_24),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3503425(.data_in(wire_d34_24),.data_out(wire_d34_25),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3503426(.data_in(wire_d34_25),.data_out(wire_d34_26),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3503427(.data_in(wire_d34_26),.data_out(wire_d34_27),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3503428(.data_in(wire_d34_27),.data_out(wire_d34_28),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3503429(.data_in(wire_d34_28),.data_out(wire_d34_29),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3503430(.data_in(wire_d34_29),.data_out(wire_d34_30),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3503431(.data_in(wire_d34_30),.data_out(wire_d34_31),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3503432(.data_in(wire_d34_31),.data_out(wire_d34_32),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3503433(.data_in(wire_d34_32),.data_out(wire_d34_33),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3503434(.data_in(wire_d34_33),.data_out(wire_d34_34),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3503435(.data_in(wire_d34_34),.data_out(wire_d34_35),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3503436(.data_in(wire_d34_35),.data_out(d_out34),.clk(clk),.rst(rst));

	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance360350(.data_in(d_in35),.data_out(wire_d35_0),.clk(clk),.rst(rst));            //channel 36
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance360351(.data_in(wire_d35_0),.data_out(wire_d35_1),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance360352(.data_in(wire_d35_1),.data_out(wire_d35_2),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance360353(.data_in(wire_d35_2),.data_out(wire_d35_3),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance360354(.data_in(wire_d35_3),.data_out(wire_d35_4),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance360355(.data_in(wire_d35_4),.data_out(wire_d35_5),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance360356(.data_in(wire_d35_5),.data_out(wire_d35_6),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance360357(.data_in(wire_d35_6),.data_out(wire_d35_7),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance360358(.data_in(wire_d35_7),.data_out(wire_d35_8),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance360359(.data_in(wire_d35_8),.data_out(wire_d35_9),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3603510(.data_in(wire_d35_9),.data_out(wire_d35_10),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3603511(.data_in(wire_d35_10),.data_out(wire_d35_11),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3603512(.data_in(wire_d35_11),.data_out(wire_d35_12),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3603513(.data_in(wire_d35_12),.data_out(wire_d35_13),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3603514(.data_in(wire_d35_13),.data_out(wire_d35_14),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3603515(.data_in(wire_d35_14),.data_out(wire_d35_15),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3603516(.data_in(wire_d35_15),.data_out(wire_d35_16),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3603517(.data_in(wire_d35_16),.data_out(wire_d35_17),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3603518(.data_in(wire_d35_17),.data_out(wire_d35_18),.clk(clk),.rst(rst));
	mux_top_vhd #(.WIDTH(WIDTH)) mux_top_vhd_instance3603519(.data_in(wire_d35_18),.data_out(wire_d35_19),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3603520(.data_in(wire_d35_19),.data_out(wire_d35_20),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3603521(.data_in(wire_d35_20),.data_out(wire_d35_21),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3603522(.data_in(wire_d35_21),.data_out(wire_d35_22),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3603523(.data_in(wire_d35_22),.data_out(wire_d35_23),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3603524(.data_in(wire_d35_23),.data_out(wire_d35_24),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3603525(.data_in(wire_d35_24),.data_out(wire_d35_25),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3603526(.data_in(wire_d35_25),.data_out(wire_d35_26),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3603527(.data_in(wire_d35_26),.data_out(wire_d35_27),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3603528(.data_in(wire_d35_27),.data_out(wire_d35_28),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3603529(.data_in(wire_d35_28),.data_out(wire_d35_29),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3603530(.data_in(wire_d35_29),.data_out(wire_d35_30),.clk(clk),.rst(rst));
	register_vhd #(.WIDTH(WIDTH)) register_vhd_instance3603531(.data_in(wire_d35_30),.data_out(wire_d35_31),.clk(clk),.rst(rst));
	shift_reg_top_vhd #(.WIDTH(WIDTH)) shift_reg_top_vhd_instance3603532(.data_in(wire_d35_31),.data_out(wire_d35_32),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3603533(.data_in(wire_d35_32),.data_out(wire_d35_33),.clk(clk),.rst(rst));
	rom_top_vhd #(.WIDTH(WIDTH)) rom_top_vhd_instance3603534(.data_in(wire_d35_33),.data_out(wire_d35_34),.clk(clk),.rst(rst));
	alu_top_vhd #(.WIDTH(WIDTH)) alu_top_vhd_instance3603535(.data_in(wire_d35_34),.data_out(wire_d35_35),.clk(clk),.rst(rst));
	decoder_top_vhd #(.WIDTH(WIDTH)) decoder_top_vhd_instance3603536(.data_in(wire_d35_35),.data_out(d_out35),.clk(clk),.rst(rst));


endmodule