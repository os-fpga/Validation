-- (C) 2010 Altera Corporation. All rights reserved.
-- Your use of Altera Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions, and any output
-- files any of the foregoing (including device programming or simulation
-- files), and any associated documentation or information are expressly subject
-- to the terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other applicable
-- license agreement, including, without limitation, that your use is for the
-- sole purpose of programming logic devices manufactured by Altera and sold by
-- Altera or its authorized distributors.  Please refer to the applicable
-- agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   DOUBLE PRECISION CORE LIBRARY             ***
--***                                             ***
--***   DP_ADDB.VHD                               ***
--***                                             ***
--***   Function: Behavioral Fixed Point Adder    ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_addb IS 
GENERIC (
         width : positive := 64;
         pipes : positive := 1
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      carryin : IN STD_LOGIC;
      
      cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
     );
END dp_addb;

ARCHITECTURE rtl OF dp_addb IS

  type pipefftype IS ARRAY (pipes DOWNTO 1) OF STD_LOGIC_VECTOR (width DOWNTO 1);
  
  signal delff : STD_LOGIC_VECTOR (width DOWNTO 1);
  signal pipeff : pipefftype;
  signal ccnode : STD_LOGIC_VECTOR (width DOWNTO 1);
  signal zerovec : STD_LOGIC_VECTOR (width-1 DOWNTO 1);
    
BEGIN
  
  gza: FOR k IN 1 TO width-1 GENERATE
    zerovec(k) <= '0';
  END GENERATE;

  ccnode <= aa + bb + (zerovec & carryin);
  
  gda: IF (pipes = 1) GENERATE
  
    pda: PROCESS (sysclk,reset)
    BEGIN

      IF (reset = '1') THEN
    
        FOR k IN 1 TO width LOOP
          delff(k) <= '0';
        END LOOP;
     
      ELSIF (rising_edge(sysclk)) THEN

        IF (enable = '1') THEN   
          delff <= ccnode;
        END IF;

      END IF;

    END PROCESS;
    
    cc <= delff;
    
  END GENERATE;
  
  gpa: IF (pipes > 1) GENERATE
  
    ppa: PROCESS (sysclk,reset)
    BEGIN

      IF (reset = '1') THEN
        
        FOR k IN 1 TO pipes LOOP 
          FOR j IN 1 TO width LOOP
            pipeff(k)(j) <= '0';
          END LOOP;
        END LOOP;
   
      ELSIF (rising_edge(sysclk)) THEN

        IF (enable = '1') THEN   
          pipeff(1)(width DOWNTO 1) <= ccnode;
          FOR k IN 2 TO pipes LOOP
            pipeff(k)(width DOWNTO 1) <= pipeff(k-1)(width DOWNTO 1);
          END LOOP;
        END IF;

      END IF;

    END PROCESS;

    cc <= pipeff(pipes)(width DOWNTO 1);
          
  END GENERATE;
       
END rtl;


LIBRARY ieee;
LIBRARY work;
LIBRARY lpm;
USE lpm.all;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CONVERSION - CORE LEVEL    ***
--***                                             ***
--***   DP_ADDPIPE.VHD                            ***
--***                                             ***
--***   Function: Adder                           ***
--***                                             ***
--***   14/07/07 ML                               ***
--***                                             ***
--***   (c) 2007 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_addpipe IS
GENERIC (
         width : positive := 64;
         pipes : positive := 1
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      carryin : IN STD_LOGIC;
      
      cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
     );
END dp_addpipe;

ARCHITECTURE syn of dp_addpipe IS

  component lpm_add_sub
  GENERIC (
		     lpm_direction		: STRING;
		     lpm_hint		: STRING;
		     lpm_pipeline		: NATURAL;
		     lpm_type		: STRING;
		     lpm_width		: NATURAL
	       );
	PORT (
			dataa	: IN STD_LOGIC_VECTOR (lpm_width-1 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (lpm_width-1 DOWNTO 0);
			cin	: IN STD_LOGIC ;
			clken	: IN STD_LOGIC ;
			aclr	: IN STD_LOGIC ;
			clock	: IN STD_LOGIC ;
			result	: OUT STD_LOGIC_VECTOR (lpm_width-1 DOWNTO 0)
	     );
  end component;

BEGIN
  
  addtwo: lpm_add_sub
  GENERIC MAP (
		       lpm_direction => "ADD",
		       lpm_hint => "ONE_INPUT_IS_CONSTANT=NO,CIN_USED=YES",
		       lpm_pipeline => pipes,
		       lpm_type => "LPM_ADD_SUB",
		       lpm_width => width
	           )
  PORT MAP (
  		    dataa => aa,
		    datab => bb,
		    cin => carryin,
		    clken => enable,
		    aclr => reset,
		    clock => sysclk,
		    result => cc
	       );  
  
END syn;


LIBRARY ieee;
LIBRARY work;
LIBRARY lpm;
USE lpm.all;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   DOUBLE PRECISION CORE LIBRARY             ***
--***                                             ***
--***   DP_ADDS.VHD                               ***
--***                                             ***
--***   Function: Synthesizable Fixed Point Adder ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_adds IS
GENERIC (
         width : positive := 64;
         pipes : positive := 1
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      carryin : IN STD_LOGIC;
      
      cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
     );
END dp_adds;

ARCHITECTURE syn of dp_adds IS

  component lpm_add_sub
  GENERIC (
		     lpm_direction		: STRING;
		     lpm_hint		: STRING;
		     lpm_pipeline		: NATURAL;
		     lpm_type		: STRING;
		     lpm_width		: NATURAL
	       );
	PORT (
			dataa	: IN STD_LOGIC_VECTOR (lpm_width-1 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (lpm_width-1 DOWNTO 0);
			cin	: IN STD_LOGIC ;
			clken	: IN STD_LOGIC ;
			aclr	: IN STD_LOGIC ;
			clock	: IN STD_LOGIC ;
			result	: OUT STD_LOGIC_VECTOR (lpm_width-1 DOWNTO 0)
	     );
  end component;

BEGIN
  
  addtwo: lpm_add_sub
  GENERIC MAP (
		       lpm_direction => "ADD",
		       lpm_hint => "ONE_INPUT_IS_CONSTANT=NO,CIN_USED=YES",
		       lpm_pipeline => pipes,
		       lpm_type => "LPM_ADD_SUB",
		       lpm_width => width
	           )
  PORT MAP (
  		    dataa => aa,
		    datab => bb,
		    cin => carryin,
		    clken => enable,
		    aclr => reset,
		    clock => sysclk,
		    result => cc
	       );  
  
END syn;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOAT CONVERT - CORE LEVEL                ***
--***                                             ***
--***   DP_CLZ64.VHD                              ***
--***                                             ***
--***   Function: Combinatorial Count Leading     ***
--***             Zeroes (64 bits)                ***
--***                                             ***
--***   01/12/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_clz64 IS
PORT (
      mantissa : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
      
      leading : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
     );
END dp_clz64;

ARCHITECTURE rtl of dp_clz64 IS

  type positiontype IS ARRAY (11 DOWNTO 1) OF STD_LOGIC_VECTOR (6 DOWNTO 1);
  
  signal position, positionmux : positiontype;
  signal zerogroup, firstzero : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal lastman : STD_LOGIC_VECTOR (6 DOWNTO 1);
  
  component dp_pos
  GENERIC (start: integer := 0);
  PORT 
       (
        ingroup : IN STD_LOGIC_VECTOR (6 DOWNTO 1); 
        
        position : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
       );
  end component;
  
BEGIN
     
  zerogroup(1) <= mantissa(64) OR mantissa(63) OR mantissa(62) OR mantissa(61) OR mantissa(60) OR mantissa(59);
  zerogroup(2) <= mantissa(58) OR mantissa(57) OR mantissa(56) OR mantissa(55) OR mantissa(54) OR mantissa(53);
  zerogroup(3) <= mantissa(52) OR mantissa(51) OR mantissa(50) OR mantissa(49) OR mantissa(48) OR mantissa(47);
  zerogroup(4) <= mantissa(46) OR mantissa(45) OR mantissa(44) OR mantissa(43) OR mantissa(42) OR mantissa(41);
  zerogroup(5) <= mantissa(40) OR mantissa(39) OR mantissa(38) OR mantissa(37) OR mantissa(36) OR mantissa(35);
  zerogroup(6) <= mantissa(34) OR mantissa(33) OR mantissa(32) OR mantissa(31) OR mantissa(30) OR mantissa(29);
  zerogroup(7) <= mantissa(28) OR mantissa(27) OR mantissa(26) OR mantissa(25) OR mantissa(24) OR mantissa(23);
  zerogroup(8) <= mantissa(22) OR mantissa(21) OR mantissa(20) OR mantissa(19) OR mantissa(18) OR mantissa(17);
  zerogroup(9) <= mantissa(16) OR mantissa(15) OR mantissa(14) OR mantissa(13) OR mantissa(12) OR mantissa(11); 
  zerogroup(10) <= mantissa(10) OR mantissa(9) OR mantissa(8) OR mantissa(7) OR mantissa(6) OR mantissa(5); 
  zerogroup(11) <= mantissa(4) OR mantissa(3) OR mantissa(2) OR mantissa(1); 

  lastman <= mantissa(4 DOWNTO 1) & "00";
  
  pone: dp_pos 
  GENERIC MAP (start=>60) 
  PORT MAP (ingroup=>lastman,position=>position(11)(6 DOWNTO 1));
  ptwo: dp_pos 
  GENERIC MAP (start=>54) 
  PORT MAP (ingroup=>mantissa(10 DOWNTO 5),position=>position(10)(6 DOWNTO 1));
  pthr: dp_pos 
  GENERIC MAP (start=>48) 
  PORT MAP (ingroup=>mantissa(16 DOWNTO 11),position=>position(9)(6 DOWNTO 1));
  pfor: dp_pos 
  GENERIC MAP (start=>42) 
  PORT MAP (ingroup=>mantissa(22 DOWNTO 17),position=>position(8)(6 DOWNTO 1));
  pfiv: dp_pos
  GENERIC MAP (start=>36) 
  PORT MAP (ingroup=>mantissa(28 DOWNTO 23),position=>position(7)(6 DOWNTO 1));
  psix: dp_pos 
  GENERIC MAP (start=>30) 
  PORT MAP (ingroup=>mantissa(34 DOWNTO 29),position=>position(6)(6 DOWNTO 1));
  psev: dp_pos 
  GENERIC MAP (start=>24) 
  PORT MAP (ingroup=>mantissa(40 DOWNTO 35),position=>position(5)(6 DOWNTO 1));
  pegt: dp_pos 
  GENERIC MAP (start=>18) 
  PORT MAP (ingroup=>mantissa(46 DOWNTO 41),position=>position(4)(6 DOWNTO 1));  
  pnin: dp_pos 
  GENERIC MAP (start=>12) 
  PORT MAP (ingroup=>mantissa(52 DOWNTO 47),position=>position(3)(6 DOWNTO 1));
  pten: dp_pos 
  GENERIC MAP (start=>6) 
  PORT MAP (ingroup=>mantissa(58 DOWNTO 53),position=>position(2)(6 DOWNTO 1));
  pelv: dp_pos 
  GENERIC MAP (start=>0) 
  PORT MAP (ingroup=>mantissa(64 DOWNTO 59),position=>position(1)(6 DOWNTO 1));

  firstzero(1) <= zerogroup(1);
  firstzero(2) <= NOT(zerogroup(1)) AND zerogroup(2);
  firstzero(3) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND zerogroup(3);
  firstzero(4) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND zerogroup(4);
  firstzero(5) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND NOT(zerogroup(4)) 
                  AND zerogroup(5);
  firstzero(6) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND NOT(zerogroup(4)) 
                  AND NOT(zerogroup(5)) AND zerogroup(6);                
  firstzero(7) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND NOT(zerogroup(4)) 
                  AND NOT(zerogroup(5)) AND NOT(zerogroup(6)) AND zerogroup(7); 
  firstzero(8) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND NOT(zerogroup(4)) 
                  AND NOT(zerogroup(5)) AND NOT(zerogroup(6)) AND NOT(zerogroup(7)) AND zerogroup(8); 
  firstzero(9) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND NOT(zerogroup(4)) 
                  AND NOT(zerogroup(5)) AND NOT(zerogroup(6)) AND NOT(zerogroup(7)) AND NOT(zerogroup(8)) 
                  AND zerogroup(9);
  firstzero(10) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND NOT(zerogroup(4)) 
                   AND NOT(zerogroup(5)) AND NOT(zerogroup(6)) AND NOT(zerogroup(7)) AND NOT(zerogroup(8)) 
                   AND NOT(zerogroup(9)) AND zerogroup(10);
  firstzero(11) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND NOT(zerogroup(4)) 
                   AND NOT(zerogroup(5)) AND NOT(zerogroup(6)) AND NOT(zerogroup(7)) AND NOT(zerogroup(8)) 
                   AND NOT(zerogroup(9)) AND NOT(zerogroup(10)) AND zerogroup(11); 
                
gma: FOR k IN 1 TO 6 GENERATE
  positionmux(1)(k) <= position(1)(k) AND firstzero(1);
  gmb: FOR j IN 2 TO 11 GENERATE
    positionmux(j)(k) <= positionmux(j-1)(k) OR (position(j)(k) AND firstzero(j));
  END GENERATE;
END GENERATE;
  
leading <= positionmux(11)(6 DOWNTO 1);
                                               
END rtl;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOAT CONVERT - CORE LEVEL                ***
--***                                             ***
--***   DP_CLZPIPE64.VHD                          ***
--***                                             ***
--***   Function: Pipelined, Count Leading Zeroes ***
--***                                             ***
--***   01/12/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_clzpipe64 IS
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      mantissa : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
      
      leading : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
     );
END dp_clzpipe64;

ARCHITECTURE rtl of dp_clzpipe64 IS

  type positiontype IS ARRAY (11 DOWNTO 1) OF STD_LOGIC_VECTOR (6 DOWNTO 1);
  
  signal position, positionff, positionmux : positiontype;
  signal zerogroupff, firstzero : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal lastman : STD_LOGIC_VECTOR (6 DOWNTO 1);
  
  component dp_pos
  GENERIC (start: integer := 0);
  PORT 
       (
        ingroup : IN STD_LOGIC_VECTOR (6 DOWNTO 1); 
        
        position : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
       );
  end component;
  
BEGIN

  pp: PROCESS (sysclk,reset)
  BEGIN
    
    IF (reset = '1') THEN
      
      FOR k IN 1 TO 11 LOOP
        zerogroupff(k) <= '0';
        FOR j IN 1 TO 6 LOOP
          positionff(k)(j) <= '0';
        END LOOP;
      END LOOP;
  
    ELSIF (rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN
     
        zerogroupff(1) <= mantissa(64) OR mantissa(63) OR mantissa(62) OR mantissa(61) OR mantissa(60) OR mantissa(59);
        zerogroupff(2) <= mantissa(58) OR mantissa(57) OR mantissa(56) OR mantissa(55) OR mantissa(54) OR mantissa(53);
        zerogroupff(3) <= mantissa(52) OR mantissa(51) OR mantissa(50) OR mantissa(49) OR mantissa(48) OR mantissa(47);
        zerogroupff(4) <= mantissa(46) OR mantissa(45) OR mantissa(44) OR mantissa(43) OR mantissa(42) OR mantissa(41);
        zerogroupff(5) <= mantissa(40) OR mantissa(39) OR mantissa(38) OR mantissa(37) OR mantissa(36) OR mantissa(35);
        zerogroupff(6) <= mantissa(34) OR mantissa(33) OR mantissa(32) OR mantissa(31) OR mantissa(30) OR mantissa(29);
        zerogroupff(7) <= mantissa(28) OR mantissa(27) OR mantissa(26) OR mantissa(25) OR mantissa(24) OR mantissa(23);
        zerogroupff(8) <= mantissa(22) OR mantissa(21) OR mantissa(20) OR mantissa(19) OR mantissa(18) OR mantissa(17);
        zerogroupff(9) <= mantissa(16) OR mantissa(15) OR mantissa(14) OR mantissa(13) OR mantissa(12) OR mantissa(11); 
        zerogroupff(10) <= mantissa(10) OR mantissa(9) OR mantissa(8) OR mantissa(7) OR mantissa(6) OR mantissa(5); 
        zerogroupff(11) <= mantissa(4) OR mantissa(3) OR mantissa(2) OR mantissa(1);  
        FOR k IN 1 TO 11 LOOP
          positionff(k)(6 DOWNTO 1) <= position(k)(6 DOWNTO 1);
        END LOOP;
     
      END IF;
    
    END IF;
  
  END PROCESS;

  lastman <= mantissa(4 DOWNTO 1) & "00";
  
  pone: dp_pos 
  GENERIC MAP (start=>60) 
  PORT MAP (ingroup=>lastman,position=>position(11)(6 DOWNTO 1));
  ptwo: dp_pos 
  GENERIC MAP (start=>54) 
  PORT MAP (ingroup=>mantissa(10 DOWNTO 5),position=>position(10)(6 DOWNTO 1));
  pthr: dp_pos 
  GENERIC MAP (start=>48) 
  PORT MAP (ingroup=>mantissa(16 DOWNTO 11),position=>position(9)(6 DOWNTO 1));
  pfor: dp_pos 
  GENERIC MAP (start=>42) 
  PORT MAP (ingroup=>mantissa(22 DOWNTO 17),position=>position(8)(6 DOWNTO 1));
  pfiv: dp_pos
  GENERIC MAP (start=>36) 
  PORT MAP (ingroup=>mantissa(28 DOWNTO 23),position=>position(7)(6 DOWNTO 1));
  psix: dp_pos 
  GENERIC MAP (start=>30) 
  PORT MAP (ingroup=>mantissa(34 DOWNTO 29),position=>position(6)(6 DOWNTO 1));
  psev: dp_pos 
  GENERIC MAP (start=>24) 
  PORT MAP (ingroup=>mantissa(40 DOWNTO 35),position=>position(5)(6 DOWNTO 1));
  pegt: dp_pos 
  GENERIC MAP (start=>18) 
  PORT MAP (ingroup=>mantissa(46 DOWNTO 41),position=>position(4)(6 DOWNTO 1));  
  pnin: dp_pos 
  GENERIC MAP (start=>12) 
  PORT MAP (ingroup=>mantissa(52 DOWNTO 47),position=>position(3)(6 DOWNTO 1));
  pten: dp_pos 
  GENERIC MAP (start=>6) 
  PORT MAP (ingroup=>mantissa(58 DOWNTO 53),position=>position(2)(6 DOWNTO 1));
  pelv: dp_pos 
  GENERIC MAP (start=>0) 
  PORT MAP (ingroup=>mantissa(64 DOWNTO 59),position=>position(1)(6 DOWNTO 1));

  firstzero(1) <= zerogroupff(1);
  firstzero(2) <= NOT(zerogroupff(1)) AND zerogroupff(2);
  firstzero(3) <= NOT(zerogroupff(1)) AND NOT(zerogroupff(2)) AND zerogroupff(3);
  firstzero(4) <= NOT(zerogroupff(1)) AND NOT(zerogroupff(2)) AND NOT(zerogroupff(3)) AND zerogroupff(4);
  firstzero(5) <= NOT(zerogroupff(1)) AND NOT(zerogroupff(2)) AND NOT(zerogroupff(3)) AND NOT(zerogroupff(4)) 
                  AND zerogroupff(5);
  firstzero(6) <= NOT(zerogroupff(1)) AND NOT(zerogroupff(2)) AND NOT(zerogroupff(3)) AND NOT(zerogroupff(4)) 
                  AND NOT(zerogroupff(5)) AND zerogroupff(6);                
  firstzero(7) <= NOT(zerogroupff(1)) AND NOT(zerogroupff(2)) AND NOT(zerogroupff(3)) AND NOT(zerogroupff(4)) 
                  AND NOT(zerogroupff(5)) AND NOT(zerogroupff(6)) AND zerogroupff(7); 
  firstzero(8) <= NOT(zerogroupff(1)) AND NOT(zerogroupff(2)) AND NOT(zerogroupff(3)) AND NOT(zerogroupff(4)) 
                  AND NOT(zerogroupff(5)) AND NOT(zerogroupff(6)) AND NOT(zerogroupff(7)) AND zerogroupff(8); 
  firstzero(9) <= NOT(zerogroupff(1)) AND NOT(zerogroupff(2)) AND NOT(zerogroupff(3)) AND NOT(zerogroupff(4)) 
                  AND NOT(zerogroupff(5)) AND NOT(zerogroupff(6)) AND NOT(zerogroupff(7)) AND NOT(zerogroupff(8)) 
                  AND zerogroupff(9); 
  firstzero(10) <= NOT(zerogroupff(1)) AND NOT(zerogroupff(2)) AND NOT(zerogroupff(3)) AND NOT(zerogroupff(4)) 
                   AND NOT(zerogroupff(5)) AND NOT(zerogroupff(6)) AND NOT(zerogroupff(7)) AND NOT(zerogroupff(8)) 
                   AND NOT(zerogroupff(9)) AND zerogroupff(10);
  firstzero(11) <= NOT(zerogroupff(1)) AND NOT(zerogroupff(2)) AND NOT(zerogroupff(3)) AND NOT(zerogroupff(4)) 
                   AND NOT(zerogroupff(5)) AND NOT(zerogroupff(6)) AND NOT(zerogroupff(7)) AND NOT(zerogroupff(8)) 
                   AND NOT(zerogroupff(9)) AND NOT(zerogroupff(10)) AND zerogroupff(11);
                                   
gma: FOR k IN 1 TO 6 GENERATE
  positionmux(1)(k) <= positionff(1)(k) AND firstzero(1);
  gmb: FOR j IN 2 TO 11 GENERATE
    positionmux(j)(k) <= positionmux(j-1)(k) OR (positionff(j)(k) AND firstzero(j));
  END GENERATE;
END GENERATE;
  
leading <= positionmux(11)(6 DOWNTO 1);
                                               
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   DOUBLE PRECISION DIVIDER - CORE           ***
--***                                             ***
--***   DP_DIV_CORE.VHD                           ***
--***                                             ***
--***   Function: Fixed Point 54 Bit Divider      ***
--***                                             ***
--***   Multiplier Convergence Algorithm          ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***   24/04/09 - SIII/SIV multiplier support    ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** SII Latency = 19 + 4*doublespeed            ***
--*** SIII/IV Latency = 18 + 2*doublespeed        ***
--***************************************************

ENTITY dp_div_core IS 
GENERIC (
         doublespeed : integer := 0; -- 0/1
         doubleaccuracy : integer := 0;  -- 0 = pruned multiplier, 1 = normal multiplier
         device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
         synthesize : integer := 1      -- 0/1      
        ); 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      dividend : IN STD_LOGIC_VECTOR (54 DOWNTO 1);
      divisor : IN STD_LOGIC_VECTOR (54 DOWNTO 1);

		quotient : OUT STD_LOGIC_VECTOR (55 DOWNTO 1)
		);
END dp_div_core;

ARCHITECTURE rtl OF dp_div_core IS

  --SII mullatency = doublespeed+5, SIII/IV mullatency = 4
  constant mullatency : positive := doublespeed+5 - device*(1+doublespeed);
  --SII addlatency = 2*doublespeed+1, SIII/IV addlatency = doublespeed+1
  constant addlatency : positive := 2*doublespeed+1 - device*doublespeed;
 
  signal zerovec : STD_LOGIC_VECTOR (54 DOWNTO 1);
  
  -- estimate
  signal invdivisor : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal dividenddel, divisordel : STD_LOGIC_VECTOR (54 DOWNTO 1);
  -- scale
  signal scaleden, scalenum : STD_LOGIC_VECTOR (54 DOWNTO 1);
  -- iteration
  signal twonode, subscaleden : STD_LOGIC_VECTOR (55 DOWNTO 1);
  signal guessone : STD_LOGIC_VECTOR (55 DOWNTO 1);
  signal guessonevec : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal absoluteval : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal absolutevalff, absoluteff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal abscarryff : STD_LOGIC;
  signal delscalenum : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal iteratenumnode : STD_LOGIC_VECTOR (72 DOWNTO 1);
  signal iteratenum : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal absoluteerror : STD_LOGIC_VECTOR (72 DOWNTO 1);
  signal mulabsguesslower : STD_LOGIC_VECTOR (19 DOWNTO 1);
  signal mulabsguessnode : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal mulabsguess : STD_LOGIC_VECTOR (54 DOWNTO 1);

  signal quotientnode : STD_LOGIC_VECTOR (72 DOWNTO 1);
  
  component fp_div_est IS 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        divisor : IN STD_LOGIC_VECTOR (19 DOWNTO 1);

		  invdivisor : OUT STD_LOGIC_VECTOR (18 DOWNTO 1)
		  );
  end component;
  
  component fp_fxmul  
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36;
           pipes : positive := 1;
           accuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1); 
      
        result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
       );
  end component;
  
  component dp_fxadd 
  GENERIC (
           width : positive := 64;
           pipes : positive := 1;
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
        carryin : IN STD_LOGIC;
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
  end component;
   
  component fp_del
  GENERIC (
           width : positive := 64;
           pipes : positive := 2
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
       
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
   end component;  
       
BEGIN
  
  gza: FOR k IN 1 TO 54 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  invcore: fp_div_est 
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            divisor=>divisor(54 DOWNTO 36),invdivisor=>invdivisor);
  
  delinone: fp_del
  GENERIC MAP (width=>54,pipes=>5)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>dividend,cc=>dividenddel);
            
  delintwo: fp_del
  GENERIC MAP (width=>54,pipes=>5)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>divisor,cc=>divisordel);
            
  --**********************************
  --*** ITERATION 0 - SCALE INPUTS ***
  --**********************************
  
  -- in level 5, out level 8+doublespeed
  mulscaleone: fp_fxmul
  GENERIC MAP (widthaa=>54,widthbb=>18,widthcc=>54,
               pipes=>3+doublespeed,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>divisordel,databb=>invdivisor,
            result=>scaleden);
  
  mulscaletwo: fp_fxmul
  GENERIC MAP (widthaa=>54,widthbb=>18,widthcc=>54,
               pipes=>3+doublespeed,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>dividenddel,databb=>invdivisor,
            result=>scalenum);
  
  --********************
  --*** ITERATION 1  ***
  --********************
  
  twonode <= '1' & zerovec(54 DOWNTO 1);
  
  gta: FOR k IN 1 TO 54 GENERATE
    subscaleden(k) <= NOT(scaleden(k));
  END GENERATE;
  subscaleden(55) <= '1';

  -- in level 8+speed, outlevel 9+2*speed
  addtwoone: dp_fxadd 
  GENERIC MAP (width=>55,pipes=>doublespeed+1,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>twonode,bb=>subscaleden,carryin=>'1',
            cc=>guessone);  
  
  guessonevec <= guessone(54 DOWNTO 1);
  
  -- absolute value of guess lower 36 bits
  -- this is still correct, because (for positive), value will be 1.(17 zeros)error
  -- can also be calculated from guessonevec (code below)
  -- gabs: FOR k IN 1 TO 36 GENERATE
  --   absoluteval(k) <= guessonevec(k) XOR NOT(guessonevec(54));
  -- END GENERATE;
  gabs: FOR k IN 1 TO 36 GENERATE
    absoluteval(k) <= scaleden(k) XOR NOT(scaleden(54));
  END GENERATE;
  
  pta: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN

      FOR k IN 1 TO 36 LOOP
        absolutevalff(k) <= '0';
        absoluteff(k) <= '0';
      END LOOP;
      abscarryff <= '0';
      
    ELSIF (rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN
          
        absolutevalff <= absoluteval; -- out level 9+speed
        abscarryff <= NOT(scaleden(54)); 
        absoluteff <= absolutevalff + 
                     (zerovec(35 DOWNTO 1) & abscarryff); -- out level 10+speed
        
      END IF;
    
    END IF;
    
  END PROCESS;

  deloneone: fp_del
  GENERIC MAP (width=>54,pipes=>doublespeed+1)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>scalenum,
            cc=>delscalenum);
    
  -- in level 9+2*doublespeed
  -- SII out level 14+3*doublespeed
  -- SIII/IV out level 13+2*doublespeed
  muloneone: fp_fxmul
  GENERIC MAP (widthaa=>54,widthbb=>54,widthcc=>72,pipes=>mullatency,
               accuracy=>doubleaccuracy,device=>device,
               synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>delscalenum,databb=>guessonevec,
            result=>iteratenumnode);
         
  gia: IF (device = 0) GENERATE     
    iteratenum <= iteratenumnode(71 DOWNTO 18);
  END GENERATE;

  gib: IF (device = 1) GENERATE 
    -- SIII/IV out level 14+2*doublespeed
    delit: fp_del
    GENERIC MAP (width=>54,pipes=>1)   
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>iteratenumnode(71 DOWNTO 18),
              cc=>iteratenum);
  END GENERATE;
  
  -- in level 10+doublespeed, out level 13+doublespeed
  mulonetwo: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>36,widthcc=>72,pipes=>3,
               synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>absoluteff,databb=>absoluteff,
            result=>absoluteerror);

  -- if speed = 0, delay absoluteerror 1 clock, else 2
  -- this guess always positive (check??)
  -- change here, error can be [19:1], not [18:1] - this is because (1.[17 zeros].error)^2
  -- gives 1.[34 zeros].error
  
  -- in level 13+speed
  -- SII out level 14+3*speed
  -- SIII/IV out level 14+2*speed
  addtwotwo: dp_fxadd 
  GENERIC MAP (width=>19,pipes=>addlatency,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>absoluteerror(72 DOWNTO 54),
            bb=>zerovec(19 DOWNTO 1),
            carryin=>absoluteerror(53),
            cc=>mulabsguesslower);  
            
  mulabsguessnode(19 DOWNTO 1) <= mulabsguesslower;
  gmga: FOR k IN 20 TO 53 GENERATE
    mulabsguessnode(k) <= '0';
  END GENERATE;
  mulabsguessnode(54) <= '1';

  mulabsguess <= mulabsguessnode;
  
  --*********************
  --*** OUTPUT SCALE  ***
  --*********************
  
  -- SII: in level 14+3*doublespeed, out level 19+4*doublespeed
  -- SIII/IV: in level 14+2*doublespeed, out level 18+2*doublespeed
  mulout: fp_fxmul
  GENERIC MAP (widthaa=>54,widthbb=>54,widthcc=>72,pipes=>mullatency,
               accuracy=>doubleaccuracy,device=>device,
               synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>iteratenum,databb=>mulabsguess,
            result=>quotientnode);
            
  quotient <= quotientnode(71 DOWNTO 17);
                  
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   DOUBLE PRECISION DIVIDER - OUTPUT STAGE   ***
--***                                             ***
--***   DP_DIVNORND.VHD                           ***
--***                                             ***
--***   Function: Output Stage, No Rounding       ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes: Latency = 1                          ***
--***************************************************

ENTITY dp_divnornd IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentdiv : IN STD_LOGIC_VECTOR (13 DOWNTO 1);
      mantissadiv : IN STD_LOGIC_VECTOR (53 DOWNTO 1); -- includes roundbit
      nanin : IN STD_LOGIC;
      dividebyzeroin : IN STD_LOGIC;

		signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
      --------------------------------------------------
      nanout : OUT STD_LOGIC;
      invalidout : OUT STD_LOGIC;
      dividebyzeroout : OUT STD_LOGIC
		);
END dp_divnornd;

ARCHITECTURE rtl OF dp_divnornd IS

  constant expwidth : positive := 11;
  constant manwidth : positive := 52;
  
  type exponentfftype IS ARRAY (2 DOWNTO 1) OF STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  
  signal zerovec : STD_LOGIC_VECTOR (manwidth-1 DOWNTO 1);
  signal signff : STD_LOGIC;
  signal nanff : STD_LOGIC;
  signal dividebyzeroff : STD_LOGIC;  
  signal mantissaff : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal exponentff : STD_LOGIC_VECTOR (expwidth+2 DOWNTO 1);
  
  signal infinitygen : STD_LOGIC_VECTOR (expwidth+1 DOWNTO 1);
  signal zerogen : STD_LOGIC_VECTOR (expwidth+1 DOWNTO 1);  
  signal setmanzero, setmanmax : STD_LOGIC;
  signal setexpzero, setexpmax : STD_LOGIC;

BEGIN
    
  gzv: FOR k IN 1 TO manwidth-1 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  pra: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN
        
      signff <= '0';
      nanff <= '0';
      dividebyzeroff <= '0';
      FOR k IN 1 TO manwidth LOOP
        mantissaff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        exponentff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF(enable = '1') THEN 
      
        signff <= signin;
        nanff <= nanin;
        dividebyzeroff <= dividebyzeroin;

        -- nan takes precedence (set max)
        -- nan takes precedence (set max)  
        FOR k IN 1 TO manwidth LOOP
          mantissaff(k) <= (mantissadiv(k+1) AND setmanzero) OR setmanmax;
        END LOOP;
               
        FOR k IN 1 TO expwidth LOOP
          exponentff(k) <= (exponentdiv(k) AND setexpzero) OR setexpmax;
        END LOOP;
      
      END IF;
             
    END IF;
      
  END PROCESS;
                                                  
--**********************************
--*** CHECK GENERATED CONDITIONS ***   
--**********************************

  -- infinity if exponent >= 255
  infinitygen(1) <= exponentdiv(1);
  gia: FOR k IN 2 TO expwidth GENERATE
    infinitygen(k) <= infinitygen(k-1) AND exponentdiv(k);
  END GENERATE;
  infinitygen(expwidth+1) <= infinitygen(expwidth) OR 
                            (exponentdiv(expwidth+1) AND 
                             NOT(exponentdiv(expwidth+2))); -- ;1' if infinity
                         
  -- zero if exponent <= 0
  zerogen(1) <= exponentdiv(1);
  gza: FOR k IN 2 TO expwidth GENERATE
    zerogen(k) <= zerogen(k-1) OR exponentdiv(k);
  END GENERATE;
  zerogen(expwidth+1) <= zerogen(expwidth) AND 
                         NOT(exponentdiv(expwidth+2)); -- '0' if zero
                    
  -- set mantissa to 0 when infinity or zero condition
  setmanzero <= NOT(infinitygen(expwidth+1)) AND zerogen(expwidth+1) AND NOT(dividebyzeroin);
  -- setmantissa to "11..11" when nan
  setmanmax <= nanin;
  -- set exponent to 0 when zero condition 
  setexpzero <= zerogen(expwidth+1);
  -- set exponent to "11..11" when nan, infinity, or divide by 0
  setexpmax <= nanin OR infinitygen(expwidth+1) OR dividebyzeroin;
                             
--***************
--*** OUTPUTS ***
--***************

  signout <= signff;   
  mantissaout <= mantissaff;
  exponentout <= exponentff(expwidth DOWNTO 1); 
  -----------------------------------------------
  nanout <= nanff;
  invalidout <= nanff;
  dividebyzeroout <= dividebyzeroff;

END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   DOUBLE PRECISION EXPONENT(e) - TOP LEVEL  ***
--***                                             ***
--***   DP_EXP.VHD                                ***
--***                                             ***
--***   Function: IEEE754 DP EXP()                ***
--***                                             ***
--***   12/08/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** Stratix II                                  ***
--*** Latency = 20 + 2*DoubleSpeed +              ***
--***           Roundconvert*(1+DoubleSpeed)      ***
--*** DoubleSpeed = 0, Roundconvert = 0 : 20      ***
--*** DoubleSpeed = 1, Roundconvert = 0 : 22      ***
--*** DoubleSpeed = 0, Roundconvert = 1 : 21      ***
--*** DoubleSpeed = 1, Roundconvert = 1 : 24      ***
--***                                             ***
--*** Stratix III                                 ***
--*** Latency = 18 +                              ***
--***           Roundconvert*(1+DoubleSpeed)      ***
--*** DoubleSpeed = 0, Roundconvert = 0 : 18      ***
--*** DoubleSpeed = 1, Roundconvert = 0 : 18      ***
--*** DoubleSpeed = 0, Roundconvert = 1 : 19      ***
--*** DoubleSpeed = 1, Roundconvert = 1 : 20      ***
--***                                             ***
--***************************************************

ENTITY dp_exp IS 
GENERIC (
         roundconvert : integer := 0; -- 0 = no round, 1 = round
         doubleaccuracy : integer := 0;  -- 0 = pruned multiplier, 1 = normal multiplier
         doublespeed : integer := 0;   -- 0/1
         device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
         synthesize : integer := 1      -- 0/1    
        );          
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (52 DOWNTO 1);

		  signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
      --------------------------------------------------
      nanout : OUT STD_LOGIC;
      overflowout : OUT STD_LOGIC;
      underflowout : OUT STD_LOGIC
		);
END dp_exp;

ARCHITECTURE rtl OF dp_exp IS
  
  constant expwidth : positive := 11;
  constant manwidth : positive := 52;
  
  constant coredepth : positive := 19 + 2*doublespeed - device*(4 + 2*doublespeed);

  signal signinff : STD_LOGIC;
  signal maninff : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal expinff : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal signff : STD_LOGIC_VECTOR (coredepth-1 DOWNTO 1);    
  signal mantissanode : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal exponentnode : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal rangeerror : STD_LOGIC;
      
  -- conditions
  signal zeroman : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal zeroexp : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal maxexp : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal zeromaninff : STD_LOGIC;
  signal maxexpinff : STD_LOGIC;
  signal naninff : STD_LOGIC;
  signal nanff : STD_LOGIC_VECTOR (coredepth-3 DOWNTO 1);
  
  --*** SII Latency = 19 + 2*doublespeed            ***
  --*** SIII/IV Latency = 14                        ***    
  component dp_exp_core
  GENERIC (
           doublespeed : integer := 0;   -- 0/1
           doubleaccuracy : integer := 0;  -- 0 = pruned multiplier, 1 = normal multiplier
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 1      -- 0/1       
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aasgn : IN STD_LOGIC;
        aaman : IN STD_LOGIC_VECTOR (52 DOWNTO 1);
        aaexp : IN STD_LOGIC_VECTOR (11 DOWNTO 1);

        ccman : OUT STD_LOGIC_VECTOR (54 DOWNTO 1);
        ccexp : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
        rangeerror : OUT STD_LOGIC
      );
  end component;

  component dp_expnornd
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        signin : IN STD_LOGIC;
        exponentexp : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
        mantissaexp : IN STD_LOGIC_VECTOR (53 DOWNTO 1);
        nanin : IN STD_LOGIC;
        rangeerror : IN STD_LOGIC;

        exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
        mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
        --------------------------------------------------
        nanout : OUT STD_LOGIC;
        overflowout : OUT STD_LOGIC;
        underflowout : OUT STD_LOGIC
		  );
  end component;
       	
  component dp_exprnd
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        signin : IN STD_LOGIC;
        exponentexp : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
        mantissaexp : IN STD_LOGIC_VECTOR (53 DOWNTO 1);
        nanin : IN STD_LOGIC;
        rangeerror : IN STD_LOGIC;

        exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
        mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
        --------------------------------------------------
        nanout : OUT STD_LOGIC;
        overflowout : OUT STD_LOGIC;
        underflowout : OUT STD_LOGIC
		  );
  end component;

  component dp_exprndpipe
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        signin : IN STD_LOGIC;
        exponentexp : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
        mantissaexp : IN STD_LOGIC_VECTOR (53 DOWNTO 1);
        nanin : IN STD_LOGIC;
        rangeerror : IN STD_LOGIC;

        exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
        mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
        --------------------------------------------------
        nanout : OUT STD_LOGIC;
        overflowout : OUT STD_LOGIC;
        underflowout : OUT STD_LOGIC
		  );
  end component;
  
BEGIN

  pma: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
  
      signinff <= '0';
      FOR k IN 1 TO manwidth LOOP
        maninff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        expinff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO coredepth-1 LOOP
        signff(k) <= '0';
      END LOOP;
    
    ELSIF (rising_edge(sysclk)) THEN

      IF (enable = '1') THEN
        
        signinff <= signin;
        maninff <= mantissain;
        expinff <= exponentin;

        signff(1) <= signinff;
        FOR k IN 2 TO coredepth-1 LOOP
          signff(k) <= signff(k-1);
        END LOOP;
                                                  
      END IF;
  
    END IF;
  
  END PROCESS;

--********************
--*** CHECK INPUTS ***
--********************

  zeroman(1) <= maninff(1);
  gca: FOR k IN 2 TO manwidth GENERATE
    zeroman(k) <= zeroman(k-1) OR maninff(k);
  END GENERATE; 
  zeroexp(1) <= expinff(1);
  gcb: FOR k IN 2 TO expwidth GENERATE
    zeroexp(k) <= zeroexp(k-1) OR expinff(k);
  END GENERATE;
  maxexp(1) <= expinff(1);
  gcc: FOR k IN 2 TO expwidth GENERATE
    maxexp(k) <= maxexp(k-1) AND expinff(k);
  END GENERATE;

  pcc: PROCESS (sysclk,reset)
  BEGIN
    
    IF (reset = '1') THEN
      
      zeromaninff <= '0';
      maxexpinff <= '0';  
      naninff <= '0';
      FOR k IN 1 TO coredepth-3 LOOP
        nanff(k) <= '0';
      END LOOP;
     
    ELSIF (rising_edge(sysclk)) THEN
            
      IF (enable = '1') THEN
     
        zeromaninff <= zeroman(manwidth);
        maxexpinff <= maxexp(expwidth);
    
        -- zero when man = 0, exp = 0
        -- infinity when man = 0, exp = max
        -- nan when man != 0, exp = max
    
        -- all ffs '1' when condition true
        naninff <= zeromaninff AND maxexpinff;

        -- nan output when nan input
        nanff(1) <= naninff;
        FOR k IN 2 TO coredepth-3 LOOP
          nanff(k) <= nanff(k-1);
        END LOOP;
      
      END IF;
   
    END IF;

  END PROCESS;


--****************
--*** EXP CORE ***
--****************

  expcore: dp_exp_core
  GENERIC MAP (doublespeed=>doublespeed,doubleaccuracy=>doubleaccuracy,
               device=>device,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aasgn=>signin,aaman=>mantissain,aaexp=>exponentin,
            ccman=>mantissanode,ccexp=>exponentnode,
            rangeerror=>rangeerror);
           
--************************
--*** ROUND AND OUTPUT ***
--************************

  gra: IF (roundconvert = 0) GENERATE

    norndout: dp_expnornd
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              signin=>signff(coredepth-1),
              exponentexp=>exponentnode,
              mantissaexp=>mantissanode(53 DOWNTO 1),
              nanin=>nanff(coredepth-3),
              rangeerror=>rangeerror,

              exponentout=>exponentout,mantissaout=>mantissaout,
              nanout=>nanout,overflowout=>overflowout,underflowout=>underflowout);
            
  END GENERATE;
  
  grb: IF (roundconvert = 1 AND doublespeed = 0) GENERATE

    rndout: dp_exprnd
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              signin=>signff(coredepth-1),
              exponentexp=>exponentnode,
              mantissaexp=>mantissanode(53 DOWNTO 1),
              nanin=>nanff(coredepth-3),
              rangeerror=>rangeerror,

              exponentout=>exponentout,mantissaout=>mantissaout,
              nanout=>nanout,overflowout=>overflowout,underflowout=>underflowout);
            
  END GENERATE;

  grc: IF (roundconvert = 1 AND doublespeed = 1) GENERATE
    
    rndoutpipe: dp_exprndpipe
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              signin=>signff(coredepth-1),
              exponentexp=>exponentnode,
              mantissaexp=>mantissanode(53 DOWNTO 1),
              nanin=>nanff(coredepth-3),
              rangeerror=>rangeerror,

              exponentout=>exponentout,mantissaout=>mantissaout,
              nanout=>nanout,overflowout=>overflowout,underflowout=>underflowout);
            
  END GENERATE;
  
  signout <= '0';
  
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   DOUBLE PRECISION EXPONENT(e) - CORE       ***
--***                                             ***
--***   DP_EXP_CORE.VHD                           ***
--***                                             ***
--***   Function: Double Precision Exponent Core  ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***   24/04/09 - SIII/SIV multiplier support    ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** SII Latency = 19 + 2*doublespeed            ***
--*** SIII/IV Latency = 17                        ***
--***************************************************

ENTITY dp_exp_core IS
GENERIC (
         doublespeed : integer := 0;   -- 0/1
         doubleaccuracy : integer := 0;  -- 0 = pruned multiplier, 1 = normal multiplier
         device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
         synthesize : integer := 1      -- 0/1       
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      aasgn : IN STD_LOGIC;
      aaman : IN STD_LOGIC_VECTOR (52 DOWNTO 1);
      aaexp : IN STD_LOGIC_VECTOR (11 DOWNTO 1);

      ccman : OUT STD_LOGIC_VECTOR (54 DOWNTO 1);
      ccexp : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
      rangeerror : OUT STD_LOGIC
     );
END dp_exp_core;

ARCHITECTURE rtl OF dp_exp_core IS

  --SII mullatency = doublespeed+5, SIII/IV mullatency = 4
  constant mullatency : positive := doublespeed+5 - device*(1+doublespeed);
  constant ranlatency : positive := 15+2*doublespeed-device*(2+2*doublespeed);
  
  type expcalcfftype IS ARRAY ((ranlatency-4) DOWNTO 1) OF 
       STD_LOGIC_VECTOR (11 DOWNTO 1);
  
  signal zerovec : STD_LOGIC_VECTOR (54 DOWNTO 1);
  -- INPUT BLOCK & SHIFTER
  signal signff : STD_LOGIC_VECTOR (ranlatency+3 DOWNTO 1);
  signal aamanff, aamandelff : STD_LOGIC_VECTOR (52 DOWNTO 1);
  signal aaexpff : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal leftshift, rightshift : STD_LOGIC_VECTOR (12 DOWNTO 1);
  signal leftshiftff, rightshiftff : STD_LOGIC_VECTOR (10 DOWNTO 1);
  signal cmpexp : STD_LOGIC_VECTOR(11 DOWNTO 1);
  signal bigexpff : STD_LOGIC_VECTOR(2 DOWNTO 1);
  signal smallrightshift : STD_LOGIC;
  signal selshiftff : STD_LOGIC_VECTOR (2 DOWNTO 1);
  signal powerbus : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal leftone, lefttwo : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal rightone, righttwo, rightthree : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal leftff, rightff : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal powerff : STD_LOGIC_VECTOR (65 DOWNTO 1);
  signal decimalleft : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal decimalright : STD_LOGIC_VECTOR (10 DOWNTO 1);
  signal fractionalleft, fractionalright : STD_LOGIC_VECTOR (54 DOWNTO 1);
  -- TABLES
  signal addlutposff, addlutnegff : STD_LOGIC_VECTOR (10 DOWNTO 1);
  signal addluttwoff, addlutthrff : STD_LOGIC_VECTOR (10 DOWNTO 1);
  signal lutposmanff, lutnegmanff : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal luttwomanff, lutthrmanff : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal lutposexpff, lutnegexpff : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal luttwoexpff : STD_LOGIC;
  signal manpos, manneg, mantwo, manthr : STD_LOGIC_VECTOR (52 DOWNTO 1);
  signal exppos, expneg : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal exptwo : STD_LOGIC;
  signal lutonemanff, luttwomandelff : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal lutoneexpff : STD_LOGIC_VECTOR (11 DOWNTO 1); 
  signal luttwoexpdelff : STD_LOGIC;
  signal expcalcff : expcalcfftype;  
  -- OVER & UNDERFLOW
  signal powercheck : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal rangeff : STD_LOGIC_VECTOR (ranlatency DOWNTO 1);
  -- TAYLOR SERIES
  signal fraction : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal xterm : STD_LOGIC_VECTOR (33 DOWNTO 1);
  signal xsquareterm : STD_LOGIC_VECTOR (12 DOWNTO 1);
  signal approxff : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal lutthrmandel : STD_LOGIC_VECTOR (54 DOWNTO 1);
  -- MULTIPLY
  signal resultone : STD_LOGIC_VECTOR (72 DOWNTO 1);
  signal resultonedel : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal resulttwo, resultthr : STD_LOGIC_VECTOR (72 DOWNTO 1);
  -- NORMALIZE
  signal normshift : STD_LOGIC_VECTOR (2 DOWNTO 1);
  signal manoutff : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal expout, expoutff : STD_LOGIC_VECTOR (11 DOWNTO 1);
    
  component dp_explutpos
  PORT (
        add : IN STD_LOGIC_VECTOR (10 DOWNTO 1);
        manhi : OUT STD_LOGIC_VECTOR (24 DOWNTO 1);
        manlo : OUT STD_LOGIC_VECTOR (28 DOWNTO 1);
        exponent : OUT STD_LOGIC_VECTOR (11 DOWNTO 1)
       );
  end component;

  component dp_explutneg 
  PORT (
        add : IN STD_LOGIC_VECTOR (10 DOWNTO 1);
        manhi : OUT STD_LOGIC_VECTOR (24 DOWNTO 1);
        manlo : OUT STD_LOGIC_VECTOR (28 DOWNTO 1);
        exponent : OUT STD_LOGIC_VECTOR (11 DOWNTO 1)
       );
  end component;
    
  component dp_explut10 
  PORT (
        add : IN STD_LOGIC_VECTOR (10 DOWNTO 1);
        manhi : OUT STD_LOGIC_VECTOR (24 DOWNTO 1);
        manlo : OUT STD_LOGIC_VECTOR (28 DOWNTO 1);
        exponent : OUT STD_LOGIC
       );
  end component;
  
  component dp_explut20 
  PORT (
        add : IN STD_LOGIC_VECTOR (10 DOWNTO 1);
        manhi : OUT STD_LOGIC_VECTOR (24 DOWNTO 1);
        manlo : OUT STD_LOGIC_VECTOR (28 DOWNTO 1)
       );
  end component;

  component fp_fxmul
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36;
           pipes : positive := 1;
           accuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1); 
      
        result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
       );
  end component;

  component fp_del
  GENERIC (
           width : positive := 64;
           pipes : positive := 2
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
       
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
   end component;  
     
BEGIN
    
  gza: FOR k IN 1 TO 54 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  --*******************
  --*** INPUT BLOCK ***
  --*******************
  
  psa: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN
    
      FOR k IN 1 TO (ranlatency+3) LOOP
        signff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 52 LOOP
        aamanff(k) <= '0';
        aamandelff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 11 LOOP
        aaexpff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 10 LOOP
        leftshiftff(k) <= '0';
        rightshiftff(k) <= '0';
	  END LOOP;
      selshiftff <= "00";
      FOR k IN 1 TO 64 LOOP
        leftff(k) <= '0';
        rightff(k) <= '0';
        powerff(k) <= '0';
      END LOOP;
	  powerff(65) <= '0';
	  bigexpff <= "00";
          
    ELSIF (rising_edge(sysclk)) THEN
    
      IF (enable = '1') THEN
          
        signff(1) <= aasgn;
        FOR k IN 2 TO (ranlatency+3) LOOP
          signff(k) <= signff(k-1);
        END LOOP;
        aamanff <= aaman;
        aamandelff <= aamanff;
        aaexpff <= aaexp;
            
        leftshiftff <= leftshift(10 DOWNTO 1);
        rightshiftff <= rightshift(10 DOWNTO 1);
        
        selshiftff(1) <= leftshift(12);
        selshiftff(2) <= selshiftff(1);
          
        -- level 3
        leftff <= lefttwo;
		-- mask out right barrel shifter output when shifting by 64 or more positions
		FOR k IN 1 TO 64 LOOP
		  rightff(k) <= rightthree(k) AND smallrightshift;
		END LOOP;
		-- overflow of left shifter matters only when the left shifted mantissa result is to be used
		bigexpff(2) <= bigexpff(1) AND NOT(selshiftff(2));
		bigexpff(1) <= NOT(cmpexp(11));
        
        -- level 4
        FOR k IN 1 TO 54 LOOP
          powerff(k) <= (fractionalleft(k) AND NOT(selshiftff(2))) OR 
                        (fractionalright(k) AND selshiftff(2));
        END LOOP;
        FOR k IN 1 TO 10 LOOP
          powerff(k+54) <= (decimalleft(k) AND NOT(selshiftff(2))) OR 
                           (decimalright(k) AND selshiftff(2));
        END LOOP;
		powerff(65) <= (decimalleft(11) AND NOT(selshiftff(2)));
		-- overflow bit required to catch exp(-1023.frac) case
     
      END IF;
 
    END IF;    
      
      
  END PROCESS;
 
  leftshift <= ('0' & aaexpff) - "001111111111";
  rightshift <= "001111111111" - ('0' & aaexpff);
          
  powerbus <= "0000000001" & aamandelff & "00";
  
  decimalleft <= ('0' & leftff(64 DOWNTO 55)) + ("0000000000" & signff(3));
  -- decimalleft may overflow to bit 11 when exp(x), -1024 < x <= -1023
  decimalright <= rightff(64 DOWNTO 55) + ("000000000" & signff(3));
  gfa: FOR k IN 1 TO 54 GENERATE
    fractionalleft(k) <= leftff(k) XOR signff(3);
    fractionalright(k) <= rightff(k) XOR signff(3);
  END GENERATE;
  
  --**********************    
  --*** BARREL SHIFTER ***
  --**********************
  
  leftone(1) <=  powerbus(1)     AND NOT(leftshiftff(2)) AND NOT(leftshiftff(1));
  leftone(2) <= (powerbus(2)     AND NOT(leftshiftff(2)) AND NOT(leftshiftff(1))) OR
                (powerbus(1)     AND NOT(leftshiftff(2)) AND     leftshiftff(1)); 
  leftone(3) <= (powerbus(3)     AND NOT(leftshiftff(2)) AND NOT(leftshiftff(1))) OR
                (powerbus(2)     AND NOT(leftshiftff(2)) AND     leftshiftff(1)) OR
                (powerbus(1)     AND     leftshiftff(2)  AND NOT(leftshiftff(1))); 
  gla: FOR k IN 4 TO 64 GENERATE
    leftone(k) <= (powerbus(k)   AND NOT(leftshiftff(2)) AND NOT(leftshiftff(1))) OR
                  (powerbus(k-1) AND NOT(leftshiftff(2)) AND     leftshiftff(1)) OR
                  (powerbus(k-2) AND     leftshiftff(2)  AND NOT(leftshiftff(1))) OR
                  (powerbus(k-3) AND     leftshiftff(2)  AND     leftshiftff(1));
  END GENERATE;
             
  glb: FOR k IN 1 TO 4 GENERATE
    lefttwo(k) <=  leftone(k)    AND NOT(leftshiftff(4)) AND NOT(leftshiftff(3));
  END GENERATE;
  glc: FOR k IN 5 TO 8 GENERATE
    lefttwo(k) <= (leftone(k)    AND NOT(leftshiftff(4)) AND NOT(leftshiftff(3))) OR
                  (leftone(k-4)  AND NOT(leftshiftff(4)) AND     leftshiftff(3)); 
  END GENERATE;
  gld: FOR k IN 9 TO 12 GENERATE
    lefttwo(k) <= (leftone(k)    AND NOT(leftshiftff(4)) AND NOT(leftshiftff(3))) OR
                  (leftone(k-4)  AND NOT(leftshiftff(4)) AND     leftshiftff(3)) OR
                  (leftone(k-8)  AND     leftshiftff(4)  AND NOT(leftshiftff(3))); 
  END GENERATE;
  gle: FOR k IN 13 TO 64 GENERATE
    lefttwo(k) <= (leftone(k)    AND NOT(leftshiftff(4)) AND NOT(leftshiftff(3))) OR
                  (leftone(k-4)  AND NOT(leftshiftff(4)) AND     leftshiftff(3)) OR
                  (leftone(k-8)  AND     leftshiftff(4)  AND NOT(leftshiftff(3)))  OR
                  (leftone(k-12) AND     leftshiftff(4)  AND     leftshiftff(3)); 
  END GENERATE;
  cmpexp <=  ('0' & leftshiftff) - "00000001010";
  -- detect when left barrel shifter overflows (i.e. leftshiftff > 9)
  
  gra: FOR k IN 1 TO 61 GENERATE
    rightone(k) <= (powerbus(k)   AND NOT(rightshiftff(2)) AND NOT(rightshiftff(1))) OR
                   (powerbus(k+1) AND NOT(rightshiftff(2)) AND     rightshiftff(1)) OR
                   (powerbus(k+2) AND     rightshiftff(2)  AND NOT(rightshiftff(1))) OR
                   (powerbus(k+3) AND     rightshiftff(2)  AND     rightshiftff(1));
  END GENERATE;
  rightone(62) <= (powerbus(62) AND NOT(rightshiftff(2)) AND NOT(rightshiftff(1))) OR
                  (powerbus(63) AND NOT(rightshiftff(2)) AND     rightshiftff(1)) OR
                  (powerbus(64) AND     rightshiftff(2)  AND NOT(rightshiftff(1))); 
  rightone(63) <= (powerbus(63) AND NOT(rightshiftff(2)) AND NOT(rightshiftff(1))) OR
                  (powerbus(64) AND NOT(rightshiftff(2)) AND     rightshiftff(1));
  rightone(64) <=  powerbus(64) AND NOT(rightshiftff(2)) AND NOT(rightshiftff(1));
  
  grb: FOR k IN 1 TO 52 GENERATE
    righttwo(k) <= (rightone(k)    AND NOT(rightshiftff(4)) AND NOT(rightshiftff(3))) OR
                   (rightone(k+4)  AND NOT(rightshiftff(4)) AND     rightshiftff(3)) OR
                   (rightone(k+8)  AND     rightshiftff(4)  AND NOT(rightshiftff(3))) OR
                   (rightone(k+12) AND     rightshiftff(4)  AND     rightshiftff(3)); 
  END GENERATE;
  grc: FOR k IN 53 TO 56 GENERATE
    righttwo(k) <= (rightone(k)   AND NOT(rightshiftff(4)) AND NOT(rightshiftff(3))) OR
                   (rightone(k+4) AND NOT(rightshiftff(4)) AND     rightshiftff(3)) OR
                   (rightone(k+8) AND     rightshiftff(4)  AND NOT(rightshiftff(3))); 
  END GENERATE; 
  grd: FOR k IN 57 TO 60 GENERATE
    righttwo(k) <= (rightone(k)   AND NOT(rightshiftff(4)) AND NOT(rightshiftff(3))) OR
                   (rightone(k+4) AND NOT(rightshiftff(4)) AND     rightshiftff(3));
  END GENERATE; 
  gre: FOR k IN 61 TO 64 GENERATE
    righttwo(k) <= (rightone(k)   AND NOT(rightshiftff(4)) AND NOT(rightshiftff(3)));
  END GENERATE; 

  grf: FOR k IN 1 TO 16 GENERATE
    rightthree(k) <= (righttwo(k)    AND NOT(rightshiftff(6)) AND NOT(rightshiftff(5))) OR
                     (righttwo(k+16) AND NOT(rightshiftff(6)) AND     rightshiftff(5)) OR
                     (righttwo(k+32) AND     rightshiftff(6)  AND NOT(rightshiftff(5))) OR
                     (righttwo(k+48) AND     rightshiftff(6)  AND     rightshiftff(5)); 
  END GENERATE;
  grg: FOR k IN 17 TO 32 GENERATE
    rightthree(k) <= (righttwo(k)    AND NOT(rightshiftff(6)) AND NOT(rightshiftff(5))) OR
                     (righttwo(k+16) AND NOT(rightshiftff(6)) AND     rightshiftff(5)) OR
                     (righttwo(k+32) AND     rightshiftff(6)  AND NOT(rightshiftff(5)));
  END GENERATE;
  grh: FOR k IN 33 TO 48 GENERATE
    rightthree(k) <= (righttwo(k)    AND NOT(rightshiftff(6)) AND NOT(rightshiftff(5))) OR
                     (righttwo(k+16) AND NOT(rightshiftff(6)) AND     rightshiftff(5));
  END GENERATE;
  gri: FOR k IN 49 TO 64 GENERATE
    rightthree(k) <= (righttwo(k)    AND NOT(rightshiftff(6)) AND NOT(rightshiftff(5)));
  END GENERATE;
  -- is rightshiftff < 64, otherwise right barrel shifter output will be masked out
  smallrightshift <= NOT(rightshiftff(7) OR rightshiftff(8) OR rightshiftff(9) OR rightshiftff(10));
  
  --******************************************
  --*** TABLES - NO RESET, FORCE TO MEMORY ***
  --******************************************
  
  -- level: 4 in, 6 out
  pla: PROCESS (sysclk)
  BEGIN
  
    IF (rising_edge(sysclk)) THEN
        
      IF (enable = '1') THEN
          
        addlutposff <= powerff(64 DOWNTO 55);
        addlutnegff <= powerff(64 DOWNTO 55);
        addluttwoff <= powerff(54 DOWNTO 45);
        addlutthrff <= powerff(44 DOWNTO 35);
        
        lutposmanff <= '1' & manpos & '0';
        lutposexpff <= exppos;
        lutnegmanff <= '1' & manneg & '0';
        lutnegexpff <= expneg;
        luttwomanff <= '1' & mantwo & '0';
        luttwoexpff <= exptwo;
        lutthrmanff <= '1' & manthr & '0';
            
      END IF;
      
    END IF;
  
  END PROCESS;
  
  declut: dp_explutpos
  PORT MAP (add=>addlutposff,
            manhi=>manpos(52 DOWNTO 29),manlo=>manpos(28 DOWNTO 1),exponent=>exppos);
            
  neglut: dp_explutneg
  PORT MAP (add=>addlutnegff,
            manhi=>manneg(52 DOWNTO 29),manlo=>manneg(28 DOWNTO 1),exponent=>expneg);
                     
  frachilut: dp_explut10
  PORT MAP (add=>addluttwoff,
            manhi=>mantwo(52 DOWNTO 29),manlo=>mantwo(28 DOWNTO 1),exponent=>exptwo);
            
  fraclolut: dp_explut20
  PORT MAP (add=>addlutthrff,
            manhi=>manthr(52 DOWNTO 29),manlo=>manthr(28 DOWNTO 1));

  -- level: 6 in, 7 out
  pma: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
    
      FOR k IN 1 TO 54 LOOP
        lutonemanff(k) <= '0';
        luttwomandelff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 11 LOOP
        lutoneexpff(k) <= '0';
      END LOOP;
      luttwoexpdelff <= '0';
      FOR k IN 1 TO (ranlatency-4) LOOP
        expcalcff(k)(11 DOWNTO 1) <= "00000000000";
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
        
      IF (enable = '1') THEN
          
        FOR k IN 1 TO 54 LOOP
          lutonemanff(k) <= (lutposmanff(k) AND NOT(signff(6))) OR (lutnegmanff(k) AND signff(6));
        END LOOP;
        luttwomandelff <= luttwomanff;
        FOR k IN 1 TO 11 LOOP
          lutoneexpff(k) <= (lutposexpff(k) AND NOT(signff(6))) OR (lutnegexpff(k) AND signff(6));
        END LOOP;
        luttwoexpdelff <= luttwoexpff;
        
        -- level: 8 in
        -- SII: 19+2*doublespeed out
        -- SII: 17+2*doublespeed out
        expcalcff(1)(11 DOWNTO 1) <= lutoneexpff + ("0000000000" & luttwoexpdelff);
        FOR k IN 2 TO (ranlatency-4) LOOP
          expcalcff(k)(11 DOWNTO 1) <= expcalcff(k-1)(11 DOWNTO 1);
        END LOOP;
            
      END IF;
      
    END IF;
          
  END PROCESS;
  
  --**************************************
  --*** PREDICT OVERFLOW AND UNDERFLOW ***
  --**************************************
  
  -- overflow or underflow if power > 709
  -- overflow or underflow if power != 0 and explut = 0
  
  powercheck <= powerff(65 DOWNTO 55) - "1011000110";  -- 710
  
  -- level 4 in
  -- SII: level 19+2 out
  -- SIII/IV: level 17 out
  ppca: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
    
      FOR k IN 1 TO ranlatency LOOP
        rangeff(k) <= '0';
      END LOOP;
    
    ELSIF (rising_edge(sysclk)) THEN
        
      IF (enable = '1') THEN
       
         rangeff(1) <= bigexpff(2) OR NOT(powercheck(11));
		 -- exp(x) -> 0 or Inf, when abs(x)>=710 or has overflowed the left shifter
         FOR k IN 2 TO (ranlatency-1) LOOP
           rangeff(k) <= rangeff(k-1);
         END LOOP;
		 rangeff(ranlatency) <= rangeff(ranlatency-1) AND NOT(signff(ranlatency+3));
		 -- overflow only if input x is large and positive, exp(x) -> Inf
       
      END IF;
      
    END IF;
          
  END PROCESS;
  
  --***********************
  --*** TAYLOR's SERIES ***
  --***********************
  
  -- approximation : sequence = 1 + x + x^2/2 + x^3/6 + x^4/24
  -- but x^3/6 term is about 62 bits down, so just try 1 + x + x^2/2
  -- ('1' & zero) + (zero(21:1) & x(34:2)) + (zero(42:1) & square(72:61))
  
  fraction <= powerff(34 DOWNTO 1) & "00";
  
  -- level: 4 in, 7 out
  mulsqr: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>36,widthcc=>12,
               pipes=>3,device=>device,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>fraction,databb=>fraction,
            result=>xsquareterm);
 
  delfrac: fp_del
  GENERIC MAP (width=>33,pipes=>3)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>powerff(34 DOWNTO 2),
            cc=>xterm); 
            
  delthr: fp_del
  GENERIC MAP (width=>54,pipes=>2)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>lutthrmanff,
            cc=>lutthrmandel); 
           
  -- level 8
  pta: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
    
      FOR k IN 1 TO 54 LOOP
        approxff(k) <= '0';
      END LOOP;
     
    ELSIF (rising_edge(sysclk)) THEN
        
      IF (enable = '1') THEN
          
        approxff <= ('1' & zerovec(20 DOWNTO 1) & xterm) + (zerovec(42 DOWNTO 1) & xsquareterm);
            
      END IF;
      
    END IF;
          
  END PROCESS;          

  --*************************************
  --*** MULTIPLY ALL EXP(X) SUBRANGES ***
  --*************************************
  
  -- SII level in 7, level out 12+speed
  -- SIII/IV level in 7, level out 11
  mulone: fp_fxmul
  GENERIC MAP (widthaa=>54,widthbb=>54,widthcc=>72,
               pipes=>mullatency,accuracy=>doubleaccuracy,
               device=>device,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>lutonemanff,databb=>luttwomandelff,
            result=>resultone);
  
  -- SII level in 12+speed, level out 13+speed
  -- SIII/IV level in 11, level out 12        
  delone: fp_del
  GENERIC MAP (width=>54,pipes=>1)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>resultone(72 DOWNTO 19),
            cc=>resultonedel); 
  
  -- SII level in 8, level out 13+speed
  -- SIII/IV level in 8, level out 12 
  multwo: fp_fxmul
  GENERIC MAP (widthaa=>54,widthbb=>54,widthcc=>72,
               pipes=>mullatency,accuracy=>doubleaccuracy,
               device=>device,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>lutthrmandel,databb=>approxff,
            result=>resulttwo);
  
  -- SII level in 13+speed, level out 18+2*speed
  -- SIII/IV level in 12, level out 16   
  multhr: fp_fxmul
  GENERIC MAP (widthaa=>54,widthbb=>54,widthcc=>72,
               pipes=>mullatency,accuracy=>doubleaccuracy,
               device=>device,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>resultonedel,databb=>resulttwo(72 DOWNTO 19),
            result=>resultthr);

  --************************
  --*** NORMALIZE OUTPUT ***
  --************************
              
  pns: PROCESS (resultthr)
  BEGIN
      
    CASE resultthr(72 DOWNTO 69) IS
      WHEN "0000" => normshift <= "11";
      WHEN "0001" => normshift <= "11";
      WHEN "0010" => normshift <= "10";
      WHEN "0011" => normshift <= "10";
      WHEN "0100" => normshift <= "01";
      WHEN "0101" => normshift <= "01";
      WHEN "0110" => normshift <= "01";
      WHEN "0111" => normshift <= "01";
      WHEN "1000" => normshift <= "00";
      WHEN "1001" => normshift <= "00";
      WHEN "1010" => normshift <= "00";
      WHEN "1011" => normshift <= "00";
      WHEN "1100" => normshift <= "00";
      WHEN "1101" => normshift <= "00";
      WHEN "1110" => normshift <= "00";
      WHEN "1111" => normshift <= "00";   
      WHEN others => normshift <= "00";
    END CASE;
        
  END PROCESS;
  
  pna: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
    
      FOR k IN 1 TO 54 LOOP
        manoutff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 11 LOOP
        expoutff(k) <= '0';
      END LOOP;
     
    ELSIF (rising_edge(sysclk)) THEN
        
      IF (enable = '1') THEN
         
        -- SII level in 18+2*doublespeed, level out 19+2*doublespeed
        -- SIII/IV level in 16, level out 17 
        FOR k IN 1 TO 54 LOOP
          manoutff(k) <= (resultthr(k+18) AND NOT(normshift(2)) AND NOT(normshift(1))) OR
                         (resultthr(k+17) AND NOT(normshift(2)) AND     normshift(1)) OR
                         (resultthr(k+16) AND     normshift(2)  AND NOT(normshift(1))) OR
                         (resultthr(k+15) AND     normshift(2)  AND     normshift(1));
        END LOOP;
		FOR k IN 1 TO 11 LOOP
          expoutff(k) <= expout(k) AND NOT(rangeff(ranlatency-1) AND signff(ranlatency+3));
		END LOOP;
        -- IEEE exponent field is set to zero when x = large negative, exp(x) -> 0
      END IF;
      
    END IF;
          
  END PROCESS; 
  expout <= expcalcff(ranlatency-4)(11 DOWNTO 1) - ("000000000" & normshift) + "00000000011";

  --***************
  --*** OUTPUTS ***
  --***************
  
  ccman <= manoutff;
  ccexp <= expoutff;
  rangeerror <= rangeff(ranlatency);
        
END rtl;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   DP_EXPLUT10.VHD                           ***
--***                                             ***
--***   Function: Look Up Table - EXP()           ***
--***                                             ***
--***   Generated by MATLAB Utility               ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_explut10 IS
PORT (
      add : IN STD_LOGIC_VECTOR (10 DOWNTO 1);
      manhi : OUT STD_LOGIC_VECTOR (24 DOWNTO 1);
      manlo : OUT STD_LOGIC_VECTOR (28 DOWNTO 1);
      exponent : OUT STD_LOGIC
     );
END dp_explut10;

ARCHITECTURE rtl OF dp_explut10 IS

BEGIN

  pca: PROCESS (add)
  BEGIN
    CASE add IS
      WHEN "0000000000" =>
            manhi <= conv_std_logic_vector(0,24);
            manlo <= conv_std_logic_vector(0,28);
           exponent <= '0';
      WHEN "0000000001" =>
            manhi <= conv_std_logic_vector(16392,24);
            manlo <= conv_std_logic_vector(699221,28);
           exponent <= '0';
      WHEN "0000000010" =>
            manhi <= conv_std_logic_vector(32800,24);
            manlo <= conv_std_logic_vector(5595137,28);
           exponent <= '0';
      WHEN "0000000011" =>
            manhi <= conv_std_logic_vector(49224,24);
            manlo <= conv_std_logic_vector(18888200,28);
           exponent <= '0';
      WHEN "0000000100" =>
            manhi <= conv_std_logic_vector(65664,24);
            manlo <= conv_std_logic_vector(44782967,28);
           exponent <= '0';
      WHEN "0000000101" =>
            manhi <= conv_std_logic_vector(82120,24);
            manlo <= conv_std_logic_vector(87488104,28);
           exponent <= '0';
      WHEN "0000000110" =>
            manhi <= conv_std_logic_vector(98592,24);
            manlo <= conv_std_logic_vector(151216387,28);
           exponent <= '0';
      WHEN "0000000111" =>
            manhi <= conv_std_logic_vector(115080,24);
            manlo <= conv_std_logic_vector(240184710,28);
           exponent <= '0';
      WHEN "0000001000" =>
            manhi <= conv_std_logic_vector(131585,24);
            manlo <= conv_std_logic_vector(90178630,28);
           exponent <= '0';
      WHEN "0000001001" =>
            manhi <= conv_std_logic_vector(148105,24);
            manlo <= conv_std_logic_vector(242294195,28);
           exponent <= '0';
      WHEN "0000001010" =>
            manhi <= conv_std_logic_vector(164642,24);
            manlo <= conv_std_logic_vector(163889760,28);
           exponent <= '0';
      WHEN "0000001011" =>
            manhi <= conv_std_logic_vector(181195,24);
            manlo <= conv_std_logic_vector(127634178,28);
           exponent <= '0';
      WHEN "0000001100" =>
            manhi <= conv_std_logic_vector(197764,24);
            manlo <= conv_std_logic_vector(137764983,28);
           exponent <= '0';
      WHEN "0000001101" =>
            manhi <= conv_std_logic_vector(214349,24);
            manlo <= conv_std_logic_vector(198523848,28);
           exponent <= '0';
      WHEN "0000001110" =>
            manhi <= conv_std_logic_vector(230951,24);
            manlo <= conv_std_logic_vector(45721136,28);
           exponent <= '0';
      WHEN "0000001111" =>
            manhi <= conv_std_logic_vector(247568,24);
            manlo <= conv_std_logic_vector(220477726,28);
           exponent <= '0';
      WHEN "0000010000" =>
            manhi <= conv_std_logic_vector(264202,24);
            manlo <= conv_std_logic_vector(190176825,28);
           exponent <= '0';
      WHEN "0000010001" =>
            manhi <= conv_std_logic_vector(280852,24);
            manlo <= conv_std_logic_vector(227512164,28);
           exponent <= '0';
      WHEN "0000010010" =>
            manhi <= conv_std_logic_vector(297519,24);
            manlo <= conv_std_logic_vector(68310723,28);
           exponent <= '0';
      WHEN "0000010011" =>
            manhi <= conv_std_logic_vector(314201,24);
            manlo <= conv_std_logic_vector(253710014,28);
           exponent <= '0';
      WHEN "0000010100" =>
            manhi <= conv_std_logic_vector(330900,24);
            manlo <= conv_std_logic_vector(251109895,28);
           exponent <= '0';
      WHEN "0000010101" =>
            manhi <= conv_std_logic_vector(347616,24);
            manlo <= conv_std_logic_vector(64785307,28);
           exponent <= '0';
      WHEN "0000010110" =>
            manhi <= conv_std_logic_vector(364347,24);
            manlo <= conv_std_logic_vector(235886282,28);
           exponent <= '0';
      WHEN "0000010111" =>
            manhi <= conv_std_logic_vector(381095,24);
            manlo <= conv_std_logic_vector(231825206,28);
           exponent <= '0';
      WHEN "0000011000" =>
            manhi <= conv_std_logic_vector(397860,24);
            manlo <= conv_std_logic_vector(56889565,28);
           exponent <= '0';
      WHEN "0000011001" =>
            manhi <= conv_std_logic_vector(414640,24);
            manlo <= conv_std_logic_vector(252241943,28);
           exponent <= '0';
      WHEN "0000011010" =>
            manhi <= conv_std_logic_vector(431438,24);
            manlo <= conv_std_logic_vector(16871840,28);
           exponent <= '0';
      WHEN "0000011011" =>
            manhi <= conv_std_logic_vector(448251,24);
            manlo <= conv_std_logic_vector(160385687,28);
           exponent <= '0';
      WHEN "0000011100" =>
            manhi <= conv_std_logic_vector(465081,24);
            manlo <= conv_std_logic_vector(150216837,28);
           exponent <= '0';
      WHEN "0000011101" =>
            manhi <= conv_std_logic_vector(481927,24);
            manlo <= conv_std_logic_vector(259109217,28);
           exponent <= '0';
      WHEN "0000011110" =>
            manhi <= conv_std_logic_vector(498790,24);
            manlo <= conv_std_logic_vector(222940052,28);
           exponent <= '0';
      WHEN "0000011111" =>
            manhi <= conv_std_logic_vector(515670,24);
            manlo <= conv_std_logic_vector(46026234,28);
           exponent <= '0';
      WHEN "0000100000" =>
            manhi <= conv_std_logic_vector(532566,24);
            manlo <= conv_std_logic_vector(1124333,28);
           exponent <= '0';
      WHEN "0000100001" =>
            manhi <= conv_std_logic_vector(549478,24);
            manlo <= conv_std_logic_vector(92559680,28);
           exponent <= '0';
      WHEN "0000100010" =>
            manhi <= conv_std_logic_vector(566407,24);
            manlo <= conv_std_logic_vector(56226380,28);
           exponent <= '0';
      WHEN "0000100011" =>
            manhi <= conv_std_logic_vector(583352,24);
            manlo <= conv_std_logic_vector(164893679,28);
           exponent <= '0';
      WHEN "0000100100" =>
            manhi <= conv_std_logic_vector(600314,24);
            manlo <= conv_std_logic_vector(154464145,28);
           exponent <= '0';
      WHEN "0000100101" =>
            manhi <= conv_std_logic_vector(617293,24);
            manlo <= conv_std_logic_vector(29280039,28);
           exponent <= '0';
      WHEN "0000100110" =>
            manhi <= conv_std_logic_vector(634288,24);
            manlo <= conv_std_logic_vector(62123323,28);
           exponent <= '0';
      WHEN "0000100111" =>
            manhi <= conv_std_logic_vector(651299,24);
            manlo <= conv_std_logic_vector(257344748,28);
           exponent <= '0';
      WHEN "0000101000" =>
            manhi <= conv_std_logic_vector(668328,24);
            manlo <= conv_std_logic_vector(82428406,28);
           exponent <= '0';
      WHEN "0000101001" =>
            manhi <= conv_std_logic_vector(685373,24);
            manlo <= conv_std_logic_vector(78604464,28);
           exponent <= '0';
      WHEN "0000101010" =>
            manhi <= conv_std_logic_vector(702434,24);
            manlo <= conv_std_logic_vector(250236442,28);
           exponent <= '0';
      WHEN "0000101011" =>
            manhi <= conv_std_logic_vector(719513,24);
            manlo <= conv_std_logic_vector(64821205,28);
           exponent <= '0';
      WHEN "0000101100" =>
            manhi <= conv_std_logic_vector(736608,24);
            manlo <= conv_std_logic_vector(63601714,28);
           exponent <= '0';
      WHEN "0000101101" =>
            manhi <= conv_std_logic_vector(753719,24);
            manlo <= conv_std_logic_vector(250954289,28);
           exponent <= '0';
      WHEN "0000101110" =>
            manhi <= conv_std_logic_vector(770848,24);
            manlo <= conv_std_logic_vector(94388611,28);
           exponent <= '0';
      WHEN "0000101111" =>
            manhi <= conv_std_logic_vector(787993,24);
            manlo <= conv_std_logic_vector(135160468,28);
           exponent <= '0';
      WHEN "0000110000" =>
            manhi <= conv_std_logic_vector(805155,24);
            manlo <= conv_std_logic_vector(109223564,28);
           exponent <= '0';
      WHEN "0000110001" =>
            manhi <= conv_std_logic_vector(822334,24);
            manlo <= conv_std_logic_vector(20971345,28);
           exponent <= '0';
      WHEN "0000110010" =>
            manhi <= conv_std_logic_vector(839529,24);
            manlo <= conv_std_logic_vector(143237009,28);
           exponent <= '0';
      WHEN "0000110011" =>
            manhi <= conv_std_logic_vector(856741,24);
            manlo <= conv_std_logic_vector(211987135,28);
           exponent <= '0';
      WHEN "0000110100" =>
            manhi <= conv_std_logic_vector(873970,24);
            manlo <= conv_std_logic_vector(231628063,28);
           exponent <= '0';
      WHEN "0000110101" =>
            manhi <= conv_std_logic_vector(891216,24);
            manlo <= conv_std_logic_vector(206570434,28);
           exponent <= '0';
      WHEN "0000110110" =>
            manhi <= conv_std_logic_vector(908479,24);
            manlo <= conv_std_logic_vector(141229202,28);
           exponent <= '0';
      WHEN "0000110111" =>
            manhi <= conv_std_logic_vector(925759,24);
            manlo <= conv_std_logic_vector(40023632,28);
           exponent <= '0';
      WHEN "0000111000" =>
            manhi <= conv_std_logic_vector(943055,24);
            manlo <= conv_std_logic_vector(175812765,28);
           exponent <= '0';
      WHEN "0000111001" =>
            manhi <= conv_std_logic_vector(960369,24);
            manlo <= conv_std_logic_vector(16153594,28);
           exponent <= '0';
      WHEN "0000111010" =>
            manhi <= conv_std_logic_vector(977699,24);
            manlo <= conv_std_logic_vector(102349263,28);
           exponent <= '0';
      WHEN "0000111011" =>
            manhi <= conv_std_logic_vector(995046,24);
            manlo <= conv_std_logic_vector(170400879,28);
           exponent <= '0';
      WHEN "0000111100" =>
            manhi <= conv_std_logic_vector(1012410,24);
            manlo <= conv_std_logic_vector(224749339,28);
           exponent <= '0';
      WHEN "0000111101" =>
            manhi <= conv_std_logic_vector(1029792,24);
            manlo <= conv_std_logic_vector(1404424,28);
           exponent <= '0';
      WHEN "0000111110" =>
            manhi <= conv_std_logic_vector(1047190,24);
            manlo <= conv_std_logic_vector(41686624,28);
           exponent <= '0';
      WHEN "0000111111" =>
            manhi <= conv_std_logic_vector(1064605,24);
            manlo <= conv_std_logic_vector(81614410,28);
           exponent <= '0';
      WHEN "0001000000" =>
            manhi <= conv_std_logic_vector(1082037,24);
            manlo <= conv_std_logic_vector(125646062,28);
           exponent <= '0';
      WHEN "0001000001" =>
            manhi <= conv_std_logic_vector(1099486,24);
            manlo <= conv_std_logic_vector(178244212,28);
           exponent <= '0';
      WHEN "0001000010" =>
            manhi <= conv_std_logic_vector(1116952,24);
            manlo <= conv_std_logic_vector(243875856,28);
           exponent <= '0';
      WHEN "0001000011" =>
            manhi <= conv_std_logic_vector(1134436,24);
            manlo <= conv_std_logic_vector(58576897,28);
           exponent <= '0';
      WHEN "0001000100" =>
            manhi <= conv_std_logic_vector(1151936,24);
            manlo <= conv_std_logic_vector(163693974,28);
           exponent <= '0';
      WHEN "0001000101" =>
            manhi <= conv_std_logic_vector(1169454,24);
            manlo <= conv_std_logic_vector(26836276,28);
           exponent <= '0';
      WHEN "0001000110" =>
            manhi <= conv_std_logic_vector(1186988,24);
            manlo <= conv_std_logic_vector(189359192,28);
           exponent <= '0';
      WHEN "0001000111" =>
            manhi <= conv_std_logic_vector(1204540,24);
            manlo <= conv_std_logic_vector(118880671,28);
           exponent <= '0';
      WHEN "0001001000" =>
            manhi <= conv_std_logic_vector(1222109,24);
            manlo <= conv_std_logic_vector(88329413,28);
           exponent <= '0';
      WHEN "0001001001" =>
            manhi <= conv_std_logic_vector(1239695,24);
            manlo <= conv_std_logic_vector(102203053,28);
           exponent <= '0';
      WHEN "0001001010" =>
            manhi <= conv_std_logic_vector(1257298,24);
            manlo <= conv_std_logic_vector(165003622,28);
           exponent <= '0';
      WHEN "0001001011" =>
            manhi <= conv_std_logic_vector(1274919,24);
            manlo <= conv_std_logic_vector(12802090,28);
           exponent <= '0';
      WHEN "0001001100" =>
            manhi <= conv_std_logic_vector(1292556,24);
            manlo <= conv_std_logic_vector(186980202,28);
           exponent <= '0';
      WHEN "0001001101" =>
            manhi <= conv_std_logic_vector(1310211,24);
            manlo <= conv_std_logic_vector(155182284,28);
           exponent <= '0';
      WHEN "0001001110" =>
            manhi <= conv_std_logic_vector(1327883,24);
            manlo <= conv_std_logic_vector(190363442,28);
           exponent <= '0';
      WHEN "0001001111" =>
            manhi <= conv_std_logic_vector(1345573,24);
            manlo <= conv_std_logic_vector(28612286,28);
           exponent <= '0';
      WHEN "0001010000" =>
            manhi <= conv_std_logic_vector(1363279,24);
            manlo <= conv_std_logic_vector(211328214,28);
           exponent <= '0';
      WHEN "0001010001" =>
            manhi <= conv_std_logic_vector(1381003,24);
            manlo <= conv_std_logic_vector(206173225,28);
           exponent <= '0';
      WHEN "0001010010" =>
            manhi <= conv_std_logic_vector(1398745,24);
            manlo <= conv_std_logic_vector(17684657,28);
           exponent <= '0';
      WHEN "0001010011" =>
            manhi <= conv_std_logic_vector(1416503,24);
            manlo <= conv_std_logic_vector(187275197,28);
           exponent <= '0';
      WHEN "0001010100" =>
            manhi <= conv_std_logic_vector(1434279,24);
            manlo <= conv_std_logic_vector(182620141,28);
           exponent <= '0';
      WHEN "0001010101" =>
            manhi <= conv_std_logic_vector(1452073,24);
            manlo <= conv_std_logic_vector(8270141,28);
           exponent <= '0';
      WHEN "0001010110" =>
            manhi <= conv_std_logic_vector(1469883,24);
            manlo <= conv_std_logic_vector(205651209,28);
           exponent <= '0';
      WHEN "0001010111" =>
            manhi <= conv_std_logic_vector(1487711,24);
            manlo <= conv_std_logic_vector(242451980,28);
           exponent <= '0';
      WHEN "0001011000" =>
            manhi <= conv_std_logic_vector(1505557,24);
            manlo <= conv_std_logic_vector(123236457,28);
           exponent <= '0';
      WHEN "0001011001" =>
            manhi <= conv_std_logic_vector(1523420,24);
            manlo <= conv_std_logic_vector(121008560,28);
           exponent <= '0';
      WHEN "0001011010" =>
            manhi <= conv_std_logic_vector(1541300,24);
            manlo <= conv_std_logic_vector(240341215,28);
           exponent <= '0';
      WHEN "0001011011" =>
            manhi <= conv_std_logic_vector(1559198,24);
            manlo <= conv_std_logic_vector(217376360,28);
           exponent <= '0';
      WHEN "0001011100" =>
            manhi <= conv_std_logic_vector(1577114,24);
            manlo <= conv_std_logic_vector(56695861,28);
           exponent <= '0';
      WHEN "0001011101" =>
            manhi <= conv_std_logic_vector(1595047,24);
            manlo <= conv_std_logic_vector(31321518,28);
           exponent <= '0';
      WHEN "0001011110" =>
            manhi <= conv_std_logic_vector(1612997,24);
            manlo <= conv_std_logic_vector(145844154,28);
           exponent <= '0';
      WHEN "0001011111" =>
            manhi <= conv_std_logic_vector(1630965,24);
            manlo <= conv_std_logic_vector(136423623,28);
           exponent <= '0';
      WHEN "0001100000" =>
            manhi <= conv_std_logic_vector(1648951,24);
            manlo <= conv_std_logic_vector(7659725,28);
           exponent <= '0';
      WHEN "0001100001" =>
            manhi <= conv_std_logic_vector(1666954,24);
            manlo <= conv_std_logic_vector(32592210,28);
           exponent <= '0';
      WHEN "0001100010" =>
            manhi <= conv_std_logic_vector(1684974,24);
            manlo <= conv_std_logic_vector(215829868,28);
           exponent <= '0';
      WHEN "0001100011" =>
            manhi <= conv_std_logic_vector(1703013,24);
            manlo <= conv_std_logic_vector(25115084,28);
           exponent <= '0';
      WHEN "0001100100" =>
            manhi <= conv_std_logic_vector(1721069,24);
            manlo <= conv_std_logic_vector(1936572,28);
           exponent <= '0';
      WHEN "0001100101" =>
            manhi <= conv_std_logic_vector(1739142,24);
            manlo <= conv_std_logic_vector(150916647,28);
           exponent <= '0';
      WHEN "0001100110" =>
            manhi <= conv_std_logic_vector(1757233,24);
            manlo <= conv_std_logic_vector(208246681,28);
           exponent <= '0';
      WHEN "0001100111" =>
            manhi <= conv_std_logic_vector(1775342,24);
            manlo <= conv_std_logic_vector(178558028,28);
           exponent <= '0';
      WHEN "0001101000" =>
            manhi <= conv_std_logic_vector(1793469,24);
            manlo <= conv_std_logic_vector(66486562,28);
           exponent <= '0';
      WHEN "0001101001" =>
            manhi <= conv_std_logic_vector(1811613,24);
            manlo <= conv_std_logic_vector(145108146,28);
           exponent <= '0';
      WHEN "0001101010" =>
            manhi <= conv_std_logic_vector(1829775,24);
            manlo <= conv_std_logic_vector(150632262,28);
           exponent <= '0';
      WHEN "0001101011" =>
            manhi <= conv_std_logic_vector(1847955,24);
            manlo <= conv_std_logic_vector(87708388,28);
           exponent <= '0';
      WHEN "0001101100" =>
            manhi <= conv_std_logic_vector(1866152,24);
            manlo <= conv_std_logic_vector(229426001,28);
           exponent <= '0';
      WHEN "0001101101" =>
            manhi <= conv_std_logic_vector(1884368,24);
            manlo <= conv_std_logic_vector(43572756,28);
           exponent <= '0';
      WHEN "0001101110" =>
            manhi <= conv_std_logic_vector(1902601,24);
            manlo <= conv_std_logic_vector(71682684,28);
           exponent <= '0';
      WHEN "0001101111" =>
            manhi <= conv_std_logic_vector(1920852,24);
            manlo <= conv_std_logic_vector(49988005,28);
           exponent <= '0';
      WHEN "0001110000" =>
            manhi <= conv_std_logic_vector(1939120,24);
            manlo <= conv_std_logic_vector(251596409,28);
           exponent <= '0';
      WHEN "0001110001" =>
            manhi <= conv_std_logic_vector(1957407,24);
            manlo <= conv_std_logic_vector(144313787,28);
           exponent <= '0';
      WHEN "0001110010" =>
            manhi <= conv_std_logic_vector(1975712,24);
            manlo <= conv_std_logic_vector(1256963,28);
           exponent <= '0';
      WHEN "0001110011" =>
            manhi <= conv_std_logic_vector(1994034,24);
            manlo <= conv_std_logic_vector(95547338,28);
           exponent <= '0';
      WHEN "0001110100" =>
            manhi <= conv_std_logic_vector(2012374,24);
            manlo <= conv_std_logic_vector(163439978,28);
           exponent <= '0';
      WHEN "0001110101" =>
            manhi <= conv_std_logic_vector(2030732,24);
            manlo <= conv_std_logic_vector(209629988,28);
           exponent <= '0';
      WHEN "0001110110" =>
            manhi <= conv_std_logic_vector(2049108,24);
            manlo <= conv_std_logic_vector(238817060,28);
           exponent <= '0';
      WHEN "0001110111" =>
            manhi <= conv_std_logic_vector(2067502,24);
            manlo <= conv_std_logic_vector(255705480,28);
           exponent <= '0';
      WHEN "0001111000" =>
            manhi <= conv_std_logic_vector(2085914,24);
            manlo <= conv_std_logic_vector(265004126,28);
           exponent <= '0';
      WHEN "0001111001" =>
            manhi <= conv_std_logic_vector(2104345,24);
            manlo <= conv_std_logic_vector(2991026,28);
           exponent <= '0';
      WHEN "0001111010" =>
            manhi <= conv_std_logic_vector(2122793,24);
            manlo <= conv_std_logic_vector(11255176,28);
           exponent <= '0';
      WHEN "0001111011" =>
            manhi <= conv_std_logic_vector(2141259,24);
            manlo <= conv_std_logic_vector(26083817,28);
           exponent <= '0';
      WHEN "0001111100" =>
            manhi <= conv_std_logic_vector(2159743,24);
            manlo <= conv_std_logic_vector(52204260,28);
           exponent <= '0';
      WHEN "0001111101" =>
            manhi <= conv_std_logic_vector(2178245,24);
            manlo <= conv_std_logic_vector(94348435,28);
           exponent <= '0';
      WHEN "0001111110" =>
            manhi <= conv_std_logic_vector(2196765,24);
            manlo <= conv_std_logic_vector(157252892,28);
           exponent <= '0';
      WHEN "0001111111" =>
            manhi <= conv_std_logic_vector(2215303,24);
            manlo <= conv_std_logic_vector(245658814,28);
           exponent <= '0';
      WHEN "0010000000" =>
            manhi <= conv_std_logic_vector(2233860,24);
            manlo <= conv_std_logic_vector(95876557,28);
           exponent <= '0';
      WHEN "0010000001" =>
            manhi <= conv_std_logic_vector(2252434,24);
            manlo <= conv_std_logic_vector(249527482,28);
           exponent <= '0';
      WHEN "0010000010" =>
            manhi <= conv_std_logic_vector(2271027,24);
            manlo <= conv_std_logic_vector(174495768,28);
           exponent <= '0';
      WHEN "0010000011" =>
            manhi <= conv_std_logic_vector(2289638,24);
            manlo <= conv_std_logic_vector(143976608,28);
           exponent <= '0';
      WHEN "0010000100" =>
            manhi <= conv_std_logic_vector(2308267,24);
            manlo <= conv_std_logic_vector(162734389,28);
           exponent <= '0';
      WHEN "0010000101" =>
            manhi <= conv_std_logic_vector(2326914,24);
            manlo <= conv_std_logic_vector(235538153,28);
           exponent <= '0';
      WHEN "0010000110" =>
            manhi <= conv_std_logic_vector(2345580,24);
            manlo <= conv_std_logic_vector(98726147,28);
           exponent <= '0';
      WHEN "0010000111" =>
            manhi <= conv_std_logic_vector(2364264,24);
            manlo <= conv_std_logic_vector(25512192,28);
           exponent <= '0';
      WHEN "0010001000" =>
            manhi <= conv_std_logic_vector(2382966,24);
            manlo <= conv_std_logic_vector(20679323,28);
           exponent <= '0';
      WHEN "0010001001" =>
            manhi <= conv_std_logic_vector(2401686,24);
            manlo <= conv_std_logic_vector(89015247,28);
           exponent <= '0';
      WHEN "0010001010" =>
            manhi <= conv_std_logic_vector(2420424,24);
            manlo <= conv_std_logic_vector(235312351,28);
           exponent <= '0';
      WHEN "0010001011" =>
            manhi <= conv_std_logic_vector(2439181,24);
            manlo <= conv_std_logic_vector(195932245,28);
           exponent <= '0';
      WHEN "0010001100" =>
            manhi <= conv_std_logic_vector(2457956,24);
            manlo <= conv_std_logic_vector(244112142,28);
           exponent <= '0';
      WHEN "0010001101" =>
            manhi <= conv_std_logic_vector(2476750,24);
            manlo <= conv_std_logic_vector(116223030,28);
           exponent <= '0';
      WHEN "0010001110" =>
            manhi <= conv_std_logic_vector(2495562,24);
            manlo <= conv_std_logic_vector(85511509,28);
           exponent <= '0';
      WHEN "0010001111" =>
            manhi <= conv_std_logic_vector(2514392,24);
            manlo <= conv_std_logic_vector(156793422,28);
           exponent <= '0';
      WHEN "0010010000" =>
            manhi <= conv_std_logic_vector(2533241,24);
            manlo <= conv_std_logic_vector(66453860,28);
           exponent <= '0';
      WHEN "0010010001" =>
            manhi <= conv_std_logic_vector(2552108,24);
            manlo <= conv_std_logic_vector(87753539,28);
           exponent <= '0';
      WHEN "0010010010" =>
            manhi <= conv_std_logic_vector(2570993,24);
            manlo <= conv_std_logic_vector(225522431,28);
           exponent <= '0';
      WHEN "0010010011" =>
            manhi <= conv_std_logic_vector(2589897,24);
            manlo <= conv_std_logic_vector(216159772,28);
           exponent <= '0';
      WHEN "0010010100" =>
            manhi <= conv_std_logic_vector(2608820,24);
            manlo <= conv_std_logic_vector(64504976,28);
           exponent <= '0';
      WHEN "0010010101" =>
            manhi <= conv_std_logic_vector(2627761,24);
            manlo <= conv_std_logic_vector(43837645,28);
           exponent <= '0';
      WHEN "0010010110" =>
            manhi <= conv_std_logic_vector(2646720,24);
            manlo <= conv_std_logic_vector(159006654,28);
           exponent <= '0';
      WHEN "0010010111" =>
            manhi <= conv_std_logic_vector(2665698,24);
            manlo <= conv_std_logic_vector(146430162,28);
           exponent <= '0';
      WHEN "0010011000" =>
            manhi <= conv_std_logic_vector(2684695,24);
            manlo <= conv_std_logic_vector(10966526,28);
           exponent <= '0';
      WHEN "0010011001" =>
            manhi <= conv_std_logic_vector(2703710,24);
            manlo <= conv_std_logic_vector(25914303,28);
           exponent <= '0';
      WHEN "0010011010" =>
            manhi <= conv_std_logic_vector(2722743,24);
            manlo <= conv_std_logic_vector(196141350,28);
           exponent <= '0';
      WHEN "0010011011" =>
            manhi <= conv_std_logic_vector(2741795,24);
            manlo <= conv_std_logic_vector(258084820,28);
           exponent <= '0';
      WHEN "0010011100" =>
            manhi <= conv_std_logic_vector(2760866,24);
            manlo <= conv_std_logic_vector(216622086,28);
           exponent <= '0';
      WHEN "0010011101" =>
            manhi <= conv_std_logic_vector(2779956,24);
            manlo <= conv_std_logic_vector(76635284,28);
           exponent <= '0';
      WHEN "0010011110" =>
            manhi <= conv_std_logic_vector(2799064,24);
            manlo <= conv_std_logic_vector(111446777,28);
           exponent <= '0';
      WHEN "0010011111" =>
            manhi <= conv_std_logic_vector(2818191,24);
            manlo <= conv_std_logic_vector(57512790,28);
           exponent <= '0';
      WHEN "0010100000" =>
            manhi <= conv_std_logic_vector(2837336,24);
            manlo <= conv_std_logic_vector(188165241,28);
           exponent <= '0';
      WHEN "0010100001" =>
            manhi <= conv_std_logic_vector(2856500,24);
            manlo <= conv_std_logic_vector(239869919,28);
           exponent <= '0';
      WHEN "0010100010" =>
            manhi <= conv_std_logic_vector(2875683,24);
            manlo <= conv_std_logic_vector(217532856,28);
           exponent <= '0';
      WHEN "0010100011" =>
            manhi <= conv_std_logic_vector(2894885,24);
            manlo <= conv_std_logic_vector(126064881,28);
           exponent <= '0';
      WHEN "0010100100" =>
            manhi <= conv_std_logic_vector(2914105,24);
            manlo <= conv_std_logic_vector(238817075,28);
           exponent <= '0';
      WHEN "0010100101" =>
            manhi <= conv_std_logic_vector(2933345,24);
            manlo <= conv_std_logic_vector(23838952,28);
           exponent <= '0';
      WHEN "0010100110" =>
            manhi <= conv_std_logic_vector(2952603,24);
            manlo <= conv_std_logic_vector(22926662,28);
           exponent <= '0';
      WHEN "0010100111" =>
            manhi <= conv_std_logic_vector(2971879,24);
            manlo <= conv_std_logic_vector(241010251,28);
           exponent <= '0';
      WHEN "0010101000" =>
            manhi <= conv_std_logic_vector(2991175,24);
            manlo <= conv_std_logic_vector(146153671,28);
           exponent <= '0';
      WHEN "0010101001" =>
            manhi <= conv_std_logic_vector(3010490,24);
            manlo <= conv_std_logic_vector(11732065,28);
           exponent <= '0';
      WHEN "0010101010" =>
            manhi <= conv_std_logic_vector(3029823,24);
            manlo <= conv_std_logic_vector(111125401,28);
           exponent <= '0';
      WHEN "0010101011" =>
            manhi <= conv_std_logic_vector(3049175,24);
            manlo <= conv_std_logic_vector(180847566,28);
           exponent <= '0';
      WHEN "0010101100" =>
            manhi <= conv_std_logic_vector(3068546,24);
            manlo <= conv_std_logic_vector(225852738,28);
           exponent <= '0';
      WHEN "0010101101" =>
            manhi <= conv_std_logic_vector(3087936,24);
            manlo <= conv_std_logic_vector(251099938,28);
           exponent <= '0';
      WHEN "0010101110" =>
            manhi <= conv_std_logic_vector(3107345,24);
            manlo <= conv_std_logic_vector(261553029,28);
           exponent <= '0';
      WHEN "0010101111" =>
            manhi <= conv_std_logic_vector(3126773,24);
            manlo <= conv_std_logic_vector(262180727,28);
           exponent <= '0';
      WHEN "0010110000" =>
            manhi <= conv_std_logic_vector(3146220,24);
            manlo <= conv_std_logic_vector(257956599,28);
           exponent <= '0';
      WHEN "0010110001" =>
            manhi <= conv_std_logic_vector(3165686,24);
            manlo <= conv_std_logic_vector(253859075,28);
           exponent <= '0';
      WHEN "0010110010" =>
            manhi <= conv_std_logic_vector(3185171,24);
            manlo <= conv_std_logic_vector(254871446,28);
           exponent <= '0';
      WHEN "0010110011" =>
            manhi <= conv_std_logic_vector(3204675,24);
            manlo <= conv_std_logic_vector(265981875,28);
           exponent <= '0';
      WHEN "0010110100" =>
            manhi <= conv_std_logic_vector(3224199,24);
            manlo <= conv_std_logic_vector(23747940,28);
           exponent <= '0';
      WHEN "0010110101" =>
            manhi <= conv_std_logic_vector(3243741,24);
            manlo <= conv_std_logic_vector(70038466,28);
           exponent <= '0';
      WHEN "0010110110" =>
            manhi <= conv_std_logic_vector(3263302,24);
            manlo <= conv_std_logic_vector(141420795,28);
           exponent <= '0';
      WHEN "0010110111" =>
            manhi <= conv_std_logic_vector(3282882,24);
            manlo <= conv_std_logic_vector(242902610,28);
           exponent <= '0';
      WHEN "0010111000" =>
            manhi <= conv_std_logic_vector(3302482,24);
            manlo <= conv_std_logic_vector(111061033,28);
           exponent <= '0';
      WHEN "0010111001" =>
            manhi <= conv_std_logic_vector(3322101,24);
            manlo <= conv_std_logic_vector(19348994,28);
           exponent <= '0';
      WHEN "0010111010" =>
            manhi <= conv_std_logic_vector(3341738,24);
            manlo <= conv_std_logic_vector(241224327,28);
           exponent <= '0';
      WHEN "0010111011" =>
            manhi <= conv_std_logic_vector(3361395,24);
            manlo <= conv_std_logic_vector(244843403,28);
           exponent <= '0';
      WHEN "0010111100" =>
            manhi <= conv_std_logic_vector(3381072,24);
            manlo <= conv_std_logic_vector(35238419,28);
           exponent <= '0';
      WHEN "0010111101" =>
            manhi <= conv_std_logic_vector(3400767,24);
            manlo <= conv_std_logic_vector(154317398,28);
           exponent <= '0';
      WHEN "0010111110" =>
            manhi <= conv_std_logic_vector(3420482,24);
            manlo <= conv_std_logic_vector(70251462,28);
           exponent <= '0';
      WHEN "0010111111" =>
            manhi <= conv_std_logic_vector(3440216,24);
            manlo <= conv_std_logic_vector(56523029,28);
           exponent <= '0';
      WHEN "0011000000" =>
            manhi <= conv_std_logic_vector(3459969,24);
            manlo <= conv_std_logic_vector(118183989,28);
           exponent <= '0';
      WHEN "0011000001" =>
            manhi <= conv_std_logic_vector(3479741,24);
            manlo <= conv_std_logic_vector(260291170,28);
           exponent <= '0';
      WHEN "0011000010" =>
            manhi <= conv_std_logic_vector(3499533,24);
            manlo <= conv_std_logic_vector(219470882,28);
           exponent <= '0';
      WHEN "0011000011" =>
            manhi <= conv_std_logic_vector(3519345,24);
            manlo <= conv_std_logic_vector(789841,28);
           exponent <= '0';
      WHEN "0011000100" =>
            manhi <= conv_std_logic_vector(3539175,24);
            manlo <= conv_std_logic_vector(146190621,28);
           exponent <= '0';
      WHEN "0011000101" =>
            manhi <= conv_std_logic_vector(3559025,24);
            manlo <= conv_std_logic_vector(123878930,28);
           exponent <= '0';
      WHEN "0011000110" =>
            manhi <= conv_std_logic_vector(3578894,24);
            manlo <= conv_std_logic_vector(207371803,28);
           exponent <= '0';
      WHEN "0011000111" =>
            manhi <= conv_std_logic_vector(3598783,24);
            manlo <= conv_std_logic_vector(133320328,28);
           exponent <= '0';
      WHEN "0011001000" =>
            manhi <= conv_std_logic_vector(3618691,24);
            manlo <= conv_std_logic_vector(175251474,28);
           exponent <= '0';
      WHEN "0011001001" =>
            manhi <= conv_std_logic_vector(3638619,24);
            manlo <= conv_std_logic_vector(69826275,28);
           exponent <= '0';
      WHEN "0011001010" =>
            manhi <= conv_std_logic_vector(3658566,24);
            manlo <= conv_std_logic_vector(90581653,28);
           exponent <= '0';
      WHEN "0011001011" =>
            manhi <= conv_std_logic_vector(3678532,24);
            manlo <= conv_std_logic_vector(242624062,28);
           exponent <= '0';
      WHEN "0011001100" =>
            manhi <= conv_std_logic_vector(3698518,24);
            manlo <= conv_std_logic_vector(262629486,28);
           exponent <= '0';
      WHEN "0011001101" =>
            manhi <= conv_std_logic_vector(3718524,24);
            manlo <= conv_std_logic_vector(155714362,28);
           exponent <= '0';
      WHEN "0011001110" =>
            manhi <= conv_std_logic_vector(3738549,24);
            manlo <= conv_std_logic_vector(195435578,28);
           exponent <= '0';
      WHEN "0011001111" =>
            manhi <= conv_std_logic_vector(3758594,24);
            manlo <= conv_std_logic_vector(118484119,28);
           exponent <= '0';
      WHEN "0011010000" =>
            manhi <= conv_std_logic_vector(3778658,24);
            manlo <= conv_std_logic_vector(198426886,28);
           exponent <= '0';
      WHEN "0011010001" =>
            manhi <= conv_std_logic_vector(3798742,24);
            manlo <= conv_std_logic_vector(171964885,28);
           exponent <= '0';
      WHEN "0011010010" =>
            manhi <= conv_std_logic_vector(3818846,24);
            manlo <= conv_std_logic_vector(44239595,28);
           exponent <= '0';
      WHEN "0011010011" =>
            manhi <= conv_std_logic_vector(3838969,24);
            manlo <= conv_std_logic_vector(88832973,28);
           exponent <= '0';
      WHEN "0011010100" =>
            manhi <= conv_std_logic_vector(3859112,24);
            manlo <= conv_std_logic_vector(42461096,28);
           exponent <= '0';
      WHEN "0011010101" =>
            manhi <= conv_std_logic_vector(3879274,24);
            manlo <= conv_std_logic_vector(178715983,28);
           exponent <= '0';
      WHEN "0011010110" =>
            manhi <= conv_std_logic_vector(3899456,24);
            manlo <= conv_std_logic_vector(234323781,28);
           exponent <= '0';
      WHEN "0011010111" =>
            manhi <= conv_std_logic_vector(3919658,24);
            manlo <= conv_std_logic_vector(214451135,28);
           exponent <= '0';
      WHEN "0011011000" =>
            manhi <= conv_std_logic_vector(3939880,24);
            manlo <= conv_std_logic_vector(124269738,28);
           exponent <= '0';
      WHEN "0011011001" =>
            manhi <= conv_std_logic_vector(3960121,24);
            manlo <= conv_std_logic_vector(237391794,28);
           exponent <= '0';
      WHEN "0011011010" =>
            manhi <= conv_std_logic_vector(3980383,24);
            manlo <= conv_std_logic_vector(22128194,28);
           exponent <= '0';
      WHEN "0011011011" =>
            manhi <= conv_std_logic_vector(4000664,24);
            manlo <= conv_std_logic_vector(20536717,28);
           exponent <= '0';
      WHEN "0011011100" =>
            manhi <= conv_std_logic_vector(4020964,24);
            manlo <= conv_std_logic_vector(237809299,28);
           exponent <= '0';
      WHEN "0011011101" =>
            manhi <= conv_std_logic_vector(4041285,24);
            manlo <= conv_std_logic_vector(142272034,28);
           exponent <= '0';
      WHEN "0011011110" =>
            manhi <= conv_std_logic_vector(4061626,24);
            manlo <= conv_std_logic_vector(7562465,28);
           exponent <= '0';
      WHEN "0011011111" =>
            manhi <= conv_std_logic_vector(4081986,24);
            manlo <= conv_std_logic_vector(107323215,28);
           exponent <= '0';
      WHEN "0011100000" =>
            manhi <= conv_std_logic_vector(4102366,24);
            manlo <= conv_std_logic_vector(178331084,28);
           exponent <= '0';
      WHEN "0011100001" =>
            manhi <= conv_std_logic_vector(4122766,24);
            manlo <= conv_std_logic_vector(225803419,28);
           exponent <= '0';
      WHEN "0011100010" =>
            manhi <= conv_std_logic_vector(4143186,24);
            manlo <= conv_std_logic_vector(254962667,28);
           exponent <= '0';
      WHEN "0011100011" =>
            manhi <= conv_std_logic_vector(4163627,24);
            manlo <= conv_std_logic_vector(2600920,28);
           exponent <= '0';
      WHEN "0011100100" =>
            manhi <= conv_std_logic_vector(4184087,24);
            manlo <= conv_std_logic_vector(10821746,28);
           exponent <= '0';
      WHEN "0011100101" =>
            manhi <= conv_std_logic_vector(4204567,24);
            manlo <= conv_std_logic_vector(16427456,28);
           exponent <= '0';
      WHEN "0011100110" =>
            manhi <= conv_std_logic_vector(4225067,24);
            manlo <= conv_std_logic_vector(24660936,28);
           exponent <= '0';
      WHEN "0011100111" =>
            manhi <= conv_std_logic_vector(4245587,24);
            manlo <= conv_std_logic_vector(40770196,28);
           exponent <= '0';
      WHEN "0011101000" =>
            manhi <= conv_std_logic_vector(4266127,24);
            manlo <= conv_std_logic_vector(70008370,28);
           exponent <= '0';
      WHEN "0011101001" =>
            manhi <= conv_std_logic_vector(4286687,24);
            manlo <= conv_std_logic_vector(117633727,28);
           exponent <= '0';
      WHEN "0011101010" =>
            manhi <= conv_std_logic_vector(4307267,24);
            manlo <= conv_std_logic_vector(188909673,28);
           exponent <= '0';
      WHEN "0011101011" =>
            manhi <= conv_std_logic_vector(4327868,24);
            manlo <= conv_std_logic_vector(20669300,28);
           exponent <= '0';
      WHEN "0011101100" =>
            manhi <= conv_std_logic_vector(4348488,24);
            manlo <= conv_std_logic_vector(155057216,28);
           exponent <= '0';
      WHEN "0011101101" =>
            manhi <= conv_std_logic_vector(4369129,24);
            manlo <= conv_std_logic_vector(60481357,28);
           exponent <= '0';
      WHEN "0011101110" =>
            manhi <= conv_std_logic_vector(4389790,24);
            manlo <= conv_std_logic_vector(10661187,28);
           exponent <= '0';
      WHEN "0011101111" =>
            manhi <= conv_std_logic_vector(4410471,24);
            manlo <= conv_std_logic_vector(10885873,28);
           exponent <= '0';
      WHEN "0011110000" =>
            manhi <= conv_std_logic_vector(4431172,24);
            manlo <= conv_std_logic_vector(66449753,28);
           exponent <= '0';
      WHEN "0011110001" =>
            manhi <= conv_std_logic_vector(4451893,24);
            manlo <= conv_std_logic_vector(182652336,28);
           exponent <= '0';
      WHEN "0011110010" =>
            manhi <= conv_std_logic_vector(4472635,24);
            manlo <= conv_std_logic_vector(96362852,28);
           exponent <= '0';
      WHEN "0011110011" =>
            manhi <= conv_std_logic_vector(4493397,24);
            manlo <= conv_std_logic_vector(81326629,28);
           exponent <= '0';
      WHEN "0011110100" =>
            manhi <= conv_std_logic_vector(4514179,24);
            manlo <= conv_std_logic_vector(142858724,28);
           exponent <= '0';
      WHEN "0011110101" =>
            manhi <= conv_std_logic_vector(4534982,24);
            manlo <= conv_std_logic_vector(17843933,28);
           exponent <= '0';
      WHEN "0011110110" =>
            manhi <= conv_std_logic_vector(4555804,24);
            manlo <= conv_std_logic_vector(248478616,28);
           exponent <= '0';
      WHEN "0011110111" =>
            manhi <= conv_std_logic_vector(4576648,24);
            manlo <= conv_std_logic_vector(34787059,28);
           exponent <= '0';
      WHEN "0011111000" =>
            manhi <= conv_std_logic_vector(4597511,24);
            manlo <= conv_std_logic_vector(187411489,28);
           exponent <= '0';
      WHEN "0011111001" =>
            manhi <= conv_std_logic_vector(4618395,24);
            manlo <= conv_std_logic_vector(174822068,28);
           exponent <= '0';
      WHEN "0011111010" =>
            manhi <= conv_std_logic_vector(4639300,24);
            manlo <= conv_std_logic_vector(2365090,28);
           exponent <= '0';
      WHEN "0011111011" =>
            manhi <= conv_std_logic_vector(4660224,24);
            manlo <= conv_std_logic_vector(212262982,28);
           exponent <= '0';
      WHEN "0011111100" =>
            manhi <= conv_std_logic_vector(4681170,24);
            manlo <= conv_std_logic_vector(4566120,28);
           exponent <= '0';
      WHEN "0011111101" =>
            manhi <= conv_std_logic_vector(4702135,24);
            manlo <= conv_std_logic_vector(189942850,28);
           exponent <= '0';
      WHEN "0011111110" =>
            manhi <= conv_std_logic_vector(4723121,24);
            manlo <= conv_std_logic_vector(236889480,28);
           exponent <= '0';
      WHEN "0011111111" =>
            manhi <= conv_std_logic_vector(4744128,24);
            manlo <= conv_std_logic_vector(150778468,28);
           exponent <= '0';
      WHEN "0100000000" =>
            manhi <= conv_std_logic_vector(4765155,24);
            manlo <= conv_std_logic_vector(205422982,28);
           exponent <= '0';
      WHEN "0100000001" =>
            manhi <= conv_std_logic_vector(4786203,24);
            manlo <= conv_std_logic_vector(137770531,28);
           exponent <= '0';
      WHEN "0100000010" =>
            manhi <= conv_std_logic_vector(4807271,24);
            manlo <= conv_std_logic_vector(221644793,28);
           exponent <= '0';
      WHEN "0100000011" =>
            manhi <= conv_std_logic_vector(4828360,24);
            manlo <= conv_std_logic_vector(194003802,28);
           exponent <= '0';
      WHEN "0100000100" =>
            manhi <= conv_std_logic_vector(4849470,24);
            manlo <= conv_std_logic_vector(60246316,28);
           exponent <= '0';
      WHEN "0100000101" =>
            manhi <= conv_std_logic_vector(4870600,24);
            manlo <= conv_std_logic_vector(94211823,28);
           exponent <= '0';
      WHEN "0100000110" =>
            manhi <= conv_std_logic_vector(4891751,24);
            manlo <= conv_std_logic_vector(32874180,28);
           exponent <= '0';
      WHEN "0100000111" =>
            manhi <= conv_std_logic_vector(4912922,24);
            manlo <= conv_std_logic_vector(150083442,28);
           exponent <= '0';
      WHEN "0100001000" =>
            manhi <= conv_std_logic_vector(4934114,24);
            manlo <= conv_std_logic_vector(182824039,28);
           exponent <= '0';
      WHEN "0100001001" =>
            manhi <= conv_std_logic_vector(4955327,24);
            manlo <= conv_std_logic_vector(136521157,28);
           exponent <= '0';
      WHEN "0100001010" =>
            manhi <= conv_std_logic_vector(4976561,24);
            manlo <= conv_std_logic_vector(16605280,28);
           exponent <= '0';
      WHEN "0100001011" =>
            manhi <= conv_std_logic_vector(4997815,24);
            manlo <= conv_std_logic_vector(96947652,28);
           exponent <= '0';
      WHEN "0100001100" =>
            manhi <= conv_std_logic_vector(5019090,24);
            manlo <= conv_std_logic_vector(114553920,28);
           exponent <= '0';
      WHEN "0100001101" =>
            manhi <= conv_std_logic_vector(5040386,24);
            manlo <= conv_std_logic_vector(74870501,28);
           exponent <= '0';
      WHEN "0100001110" =>
            manhi <= conv_std_logic_vector(5061702,24);
            manlo <= conv_std_logic_vector(251784590,28);
           exponent <= '0';
      WHEN "0100001111" =>
            manhi <= conv_std_logic_vector(5083040,24);
            manlo <= conv_std_logic_vector(113882338,28);
           exponent <= '0';
      WHEN "0100010000" =>
            manhi <= conv_std_logic_vector(5104398,24);
            manlo <= conv_std_logic_vector(203497056,28);
           exponent <= '0';
      WHEN "0100010001" =>
            manhi <= conv_std_logic_vector(5125777,24);
            manlo <= conv_std_logic_vector(257661021,28);
           exponent <= '0';
      WHEN "0100010010" =>
            manhi <= conv_std_logic_vector(5147178,24);
            manlo <= conv_std_logic_vector(13411854,28);
           exponent <= '0';
      WHEN "0100010011" =>
            manhi <= conv_std_logic_vector(5168599,24);
            manlo <= conv_std_logic_vector(13098889,28);
           exponent <= '0';
      WHEN "0100010100" =>
            manhi <= conv_std_logic_vector(5190040,24);
            manlo <= conv_std_logic_vector(262205904,28);
           exponent <= '0';
      WHEN "0100010101" =>
            manhi <= conv_std_logic_vector(5211503,24);
            manlo <= conv_std_logic_vector(229351119,28);
           exponent <= '0';
      WHEN "0100010110" =>
            manhi <= conv_std_logic_vector(5232987,24);
            manlo <= conv_std_logic_vector(188464488,28);
           exponent <= '0';
      WHEN "0100010111" =>
            manhi <= conv_std_logic_vector(5254492,24);
            manlo <= conv_std_logic_vector(145045878,28);
           exponent <= '0';
      WHEN "0100011000" =>
            manhi <= conv_std_logic_vector(5276018,24);
            manlo <= conv_std_logic_vector(104600525,28);
           exponent <= '0';
      WHEN "0100011001" =>
            manhi <= conv_std_logic_vector(5297565,24);
            manlo <= conv_std_logic_vector(72639049,28);
           exponent <= '0';
      WHEN "0100011010" =>
            manhi <= conv_std_logic_vector(5319133,24);
            manlo <= conv_std_logic_vector(54677451,28);
           exponent <= '0';
      WHEN "0100011011" =>
            manhi <= conv_std_logic_vector(5340722,24);
            manlo <= conv_std_logic_vector(56237123,28);
           exponent <= '0';
      WHEN "0100011100" =>
            manhi <= conv_std_logic_vector(5362332,24);
            manlo <= conv_std_logic_vector(82844851,28);
           exponent <= '0';
      WHEN "0100011101" =>
            manhi <= conv_std_logic_vector(5383963,24);
            manlo <= conv_std_logic_vector(140032820,28);
           exponent <= '0';
      WHEN "0100011110" =>
            manhi <= conv_std_logic_vector(5405615,24);
            manlo <= conv_std_logic_vector(233338622,28);
           exponent <= '0';
      WHEN "0100011111" =>
            manhi <= conv_std_logic_vector(5427289,24);
            manlo <= conv_std_logic_vector(99869801,28);
           exponent <= '0';
      WHEN "0100100000" =>
            manhi <= conv_std_logic_vector(5448984,24);
            manlo <= conv_std_logic_vector(13610232,28);
           exponent <= '0';
      WHEN "0100100001" =>
            manhi <= conv_std_logic_vector(5470699,24);
            manlo <= conv_std_logic_vector(248549207,28);
           exponent <= '0';
      WHEN "0100100010" =>
            manhi <= conv_std_logic_vector(5492437,24);
            manlo <= conv_std_logic_vector(4939624,28);
           exponent <= '0';
      WHEN "0100100011" =>
            manhi <= conv_std_logic_vector(5514195,24);
            manlo <= conv_std_logic_vector(93652547,28);
           exponent <= '0';
      WHEN "0100100100" =>
            manhi <= conv_std_logic_vector(5535974,24);
            manlo <= conv_std_logic_vector(251822653,28);
           exponent <= '0';
      WHEN "0100100101" =>
            manhi <= conv_std_logic_vector(5557775,24);
            manlo <= conv_std_logic_vector(216590061,28);
           exponent <= '0';
      WHEN "0100100110" =>
            manhi <= conv_std_logic_vector(5579597,24);
            manlo <= conv_std_logic_vector(261971250,28);
           exponent <= '0';
      WHEN "0100100111" =>
            manhi <= conv_std_logic_vector(5601441,24);
            manlo <= conv_std_logic_vector(125117240,28);
           exponent <= '0';
      WHEN "0100101000" =>
            manhi <= conv_std_logic_vector(5623306,24);
            manlo <= conv_std_logic_vector(80055420,28);
           exponent <= '0';
      WHEN "0100101001" =>
            manhi <= conv_std_logic_vector(5645192,24);
            manlo <= conv_std_logic_vector(132383188,28);
           exponent <= '0';
      WHEN "0100101010" =>
            manhi <= conv_std_logic_vector(5667100,24);
            manlo <= conv_std_logic_vector(19267955,28);
           exponent <= '0';
      WHEN "0100101011" =>
            manhi <= conv_std_logic_vector(5689029,24);
            manlo <= conv_std_logic_vector(14753516,28);
           exponent <= '0';
      WHEN "0100101100" =>
            manhi <= conv_std_logic_vector(5710979,24);
            manlo <= conv_std_logic_vector(124453694,28);
           exponent <= '0';
      WHEN "0100101101" =>
            manhi <= conv_std_logic_vector(5732951,24);
            manlo <= conv_std_logic_vector(85552334,28);
           exponent <= '0';
      WHEN "0100101110" =>
            manhi <= conv_std_logic_vector(5754944,24);
            manlo <= conv_std_logic_vector(172109691,28);
           exponent <= '0';
      WHEN "0100101111" =>
            manhi <= conv_std_logic_vector(5776959,24);
            manlo <= conv_std_logic_vector(121320598,28);
           exponent <= '0';
      WHEN "0100110000" =>
            manhi <= conv_std_logic_vector(5798995,24);
            manlo <= conv_std_logic_vector(207256304,28);
           exponent <= '0';
      WHEN "0100110001" =>
            manhi <= conv_std_logic_vector(5821053,24);
            manlo <= conv_std_logic_vector(167122651,28);
           exponent <= '0';
      WHEN "0100110010" =>
            manhi <= conv_std_logic_vector(5843133,24);
            manlo <= conv_std_logic_vector(6566449,28);
           exponent <= '0';
      WHEN "0100110011" =>
            manhi <= conv_std_logic_vector(5865233,24);
            manlo <= conv_std_logic_vector(268110937,28);
           exponent <= '0';
      WHEN "0100110100" =>
            manhi <= conv_std_logic_vector(5887356,24);
            manlo <= conv_std_logic_vector(152107598,28);
           exponent <= '0';
      WHEN "0100110101" =>
            manhi <= conv_std_logic_vector(5909500,24);
            manlo <= conv_std_logic_vector(201090721,28);
           exponent <= '0';
      WHEN "0100110110" =>
            manhi <= conv_std_logic_vector(5931666,24);
            manlo <= conv_std_logic_vector(152293761,28);
           exponent <= '0';
      WHEN "0100110111" =>
            manhi <= conv_std_logic_vector(5953854,24);
            manlo <= conv_std_logic_vector(11391168,28);
           exponent <= '0';
      WHEN "0100111000" =>
            manhi <= conv_std_logic_vector(5976063,24);
            manlo <= conv_std_logic_vector(52498394,28);
           exponent <= '0';
      WHEN "0100111001" =>
            manhi <= conv_std_logic_vector(5998294,24);
            manlo <= conv_std_logic_vector(12865523,28);
           exponent <= '0';
      WHEN "0100111010" =>
            manhi <= conv_std_logic_vector(6020546,24);
            manlo <= conv_std_logic_vector(166619112,28);
           exponent <= '0';
      WHEN "0100111011" =>
            manhi <= conv_std_logic_vector(6042820,24);
            manlo <= conv_std_logic_vector(251020365,28);
           exponent <= '0';
      WHEN "0100111100" =>
            manhi <= conv_std_logic_vector(6065117,24);
            manlo <= conv_std_logic_vector(3336048,28);
           exponent <= '0';
      WHEN "0100111101" =>
            manhi <= conv_std_logic_vector(6087434,24);
            manlo <= conv_std_logic_vector(234580328,28);
           exponent <= '0';
      WHEN "0100111110" =>
            manhi <= conv_std_logic_vector(6109774,24);
            manlo <= conv_std_logic_vector(145160209,28);
           exponent <= '0';
      WHEN "0100111111" =>
            manhi <= conv_std_logic_vector(6132136,24);
            manlo <= conv_std_logic_vector(9230102,28);
           exponent <= '0';
      WHEN "0101000000" =>
            manhi <= conv_std_logic_vector(6154519,24);
            manlo <= conv_std_logic_vector(100950005,28);
           exponent <= '0';
      WHEN "0101000001" =>
            manhi <= conv_std_logic_vector(6176924,24);
            manlo <= conv_std_logic_vector(157614600,28);
           exponent <= '0';
      WHEN "0101000010" =>
            manhi <= conv_std_logic_vector(6199351,24);
            manlo <= conv_std_logic_vector(184959620,28);
           exponent <= '0';
      WHEN "0101000011" =>
            manhi <= conv_std_logic_vector(6221800,24);
            manlo <= conv_std_logic_vector(188726403,28);
           exponent <= '0';
      WHEN "0101000100" =>
            manhi <= conv_std_logic_vector(6244271,24);
            manlo <= conv_std_logic_vector(174661898,28);
           exponent <= '0';
      WHEN "0101000101" =>
            manhi <= conv_std_logic_vector(6266764,24);
            manlo <= conv_std_logic_vector(148518669,28);
           exponent <= '0';
      WHEN "0101000110" =>
            manhi <= conv_std_logic_vector(6289279,24);
            manlo <= conv_std_logic_vector(116054898,28);
           exponent <= '0';
      WHEN "0101000111" =>
            manhi <= conv_std_logic_vector(6311816,24);
            manlo <= conv_std_logic_vector(83034395,28);
           exponent <= '0';
      WHEN "0101001000" =>
            manhi <= conv_std_logic_vector(6334375,24);
            manlo <= conv_std_logic_vector(55226600,28);
           exponent <= '0';
      WHEN "0101001001" =>
            manhi <= conv_std_logic_vector(6356956,24);
            manlo <= conv_std_logic_vector(38406593,28);
           exponent <= '0';
      WHEN "0101001010" =>
            manhi <= conv_std_logic_vector(6379559,24);
            manlo <= conv_std_logic_vector(38355093,28);
           exponent <= '0';
      WHEN "0101001011" =>
            manhi <= conv_std_logic_vector(6402184,24);
            manlo <= conv_std_logic_vector(60858469,28);
           exponent <= '0';
      WHEN "0101001100" =>
            manhi <= conv_std_logic_vector(6424831,24);
            manlo <= conv_std_logic_vector(111708742,28);
           exponent <= '0';
      WHEN "0101001101" =>
            manhi <= conv_std_logic_vector(6447500,24);
            manlo <= conv_std_logic_vector(196703594,28);
           exponent <= '0';
      WHEN "0101001110" =>
            manhi <= conv_std_logic_vector(6470192,24);
            manlo <= conv_std_logic_vector(53210914,28);
           exponent <= '0';
      WHEN "0101001111" =>
            manhi <= conv_std_logic_vector(6492905,24);
            manlo <= conv_std_logic_vector(223910630,28);
           exponent <= '0';
      WHEN "0101010000" =>
            manhi <= conv_std_logic_vector(6515641,24);
            manlo <= conv_std_logic_vector(177746520,28);
           exponent <= '0';
      WHEN "0101010001" =>
            manhi <= conv_std_logic_vector(6538399,24);
            manlo <= conv_std_logic_vector(188974414,28);
           exponent <= '0';
      WHEN "0101010010" =>
            manhi <= conv_std_logic_vector(6561179,24);
            manlo <= conv_std_logic_vector(263420371,28);
           exponent <= '0';
      WHEN "0101010011" =>
            manhi <= conv_std_logic_vector(6583982,24);
            manlo <= conv_std_logic_vector(138480686,28);
           exponent <= '0';
      WHEN "0101010100" =>
            manhi <= conv_std_logic_vector(6606807,24);
            manlo <= conv_std_logic_vector(88428264,28);
           exponent <= '0';
      WHEN "0101010101" =>
            manhi <= conv_std_logic_vector(6629654,24);
            manlo <= conv_std_logic_vector(119106258,28);
           exponent <= '0';
      WHEN "0101010110" =>
            manhi <= conv_std_logic_vector(6652523,24);
            manlo <= conv_std_logic_vector(236363530,28);
           exponent <= '0';
      WHEN "0101010111" =>
            manhi <= conv_std_logic_vector(6675415,24);
            manlo <= conv_std_logic_vector(177619200,28);
           exponent <= '0';
      WHEN "0101011000" =>
            manhi <= conv_std_logic_vector(6698329,24);
            manlo <= conv_std_logic_vector(217169020,28);
           exponent <= '0';
      WHEN "0101011001" =>
            manhi <= conv_std_logic_vector(6721266,24);
            manlo <= conv_std_logic_vector(92443558,28);
           exponent <= '0';
      WHEN "0101011010" =>
            manhi <= conv_std_logic_vector(6744225,24);
            manlo <= conv_std_logic_vector(77750021,28);
           exponent <= '0';
      WHEN "0101011011" =>
            manhi <= conv_std_logic_vector(6767206,24);
            manlo <= conv_std_logic_vector(178965902,28);
           exponent <= '0';
      WHEN "0101011100" =>
            manhi <= conv_std_logic_vector(6790210,24);
            manlo <= conv_std_logic_vector(133538975,28);
           exponent <= '0';
      WHEN "0101011101" =>
            manhi <= conv_std_logic_vector(6813236,24);
            manlo <= conv_std_logic_vector(215793680,28);
           exponent <= '0';
      WHEN "0101011110" =>
            manhi <= conv_std_logic_vector(6836285,24);
            manlo <= conv_std_logic_vector(163189294,28);
           exponent <= '0';
      WHEN "0101011111" =>
            manhi <= conv_std_logic_vector(6859356,24);
            manlo <= conv_std_logic_vector(250061769,28);
           exponent <= '0';
      WHEN "0101100000" =>
            manhi <= conv_std_logic_vector(6882450,24);
            manlo <= conv_std_logic_vector(213881907,28);
           exponent <= '0';
      WHEN "0101100001" =>
            manhi <= conv_std_logic_vector(6905567,24);
            manlo <= conv_std_logic_vector(60561738,28);
           exponent <= '0';
      WHEN "0101100010" =>
            manhi <= conv_std_logic_vector(6928706,24);
            manlo <= conv_std_logic_vector(64454525,28);
           exponent <= '0';
      WHEN "0101100011" =>
            manhi <= conv_std_logic_vector(6951867,24);
            manlo <= conv_std_logic_vector(231483856,28);
           exponent <= '0';
      WHEN "0101100100" =>
            manhi <= conv_std_logic_vector(6975052,24);
            manlo <= conv_std_logic_vector(30708194,28);
           exponent <= '0';
      WHEN "0101100101" =>
            manhi <= conv_std_logic_vector(6998259,24);
            manlo <= conv_std_logic_vector(4933620,28);
           exponent <= '0';
      WHEN "0101100110" =>
            manhi <= conv_std_logic_vector(7021488,24);
            manlo <= conv_std_logic_vector(160101103,28);
           exponent <= '0';
      WHEN "0101100111" =>
            manhi <= conv_std_logic_vector(7044740,24);
            manlo <= conv_std_logic_vector(233721959,28);
           exponent <= '0';
      WHEN "0101101000" =>
            manhi <= conv_std_logic_vector(7068015,24);
            manlo <= conv_std_logic_vector(231748770,28);
           exponent <= '0';
      WHEN "0101101001" =>
            manhi <= conv_std_logic_vector(7091313,24);
            manlo <= conv_std_logic_vector(160139936,28);
           exponent <= '0';
      WHEN "0101101010" =>
            manhi <= conv_std_logic_vector(7114634,24);
            manlo <= conv_std_logic_vector(24859676,28);
           exponent <= '0';
      WHEN "0101101011" =>
            manhi <= conv_std_logic_vector(7137977,24);
            manlo <= conv_std_logic_vector(100313494,28);
           exponent <= '0';
      WHEN "0101101100" =>
            manhi <= conv_std_logic_vector(7161343,24);
            manlo <= conv_std_logic_vector(124041814,28);
           exponent <= '0';
      WHEN "0101101101" =>
            manhi <= conv_std_logic_vector(7184732,24);
            manlo <= conv_std_logic_vector(102026355,28);
           exponent <= '0';
      WHEN "0101101110" =>
            manhi <= conv_std_logic_vector(7208144,24);
            manlo <= conv_std_logic_vector(40254681,28);
           exponent <= '0';
      WHEN "0101101111" =>
            manhi <= conv_std_logic_vector(7231578,24);
            manlo <= conv_std_logic_vector(213155662,28);
           exponent <= '0';
      WHEN "0101110000" =>
            manhi <= conv_std_logic_vector(7255036,24);
            manlo <= conv_std_logic_vector(89857654,28);
           exponent <= '0';
      WHEN "0101110001" =>
            manhi <= conv_std_logic_vector(7278516,24);
            manlo <= conv_std_logic_vector(213236700,28);
           exponent <= '0';
      WHEN "0101110010" =>
            manhi <= conv_std_logic_vector(7302020,24);
            manlo <= conv_std_logic_vector(52432888,28);
           exponent <= '0';
      WHEN "0101110011" =>
            manhi <= conv_std_logic_vector(7325546,24);
            manlo <= conv_std_logic_vector(150334000,28);
           exponent <= '0';
      WHEN "0101110100" =>
            manhi <= conv_std_logic_vector(7349095,24);
            manlo <= conv_std_logic_vector(244527329,28);
           exponent <= '0';
      WHEN "0101110101" =>
            manhi <= conv_std_logic_vector(7372668,24);
            manlo <= conv_std_logic_vector(72606054,28);
           exponent <= '0';
      WHEN "0101110110" =>
            manhi <= conv_std_logic_vector(7396263,24);
            manlo <= conv_std_logic_vector(177475612,28);
           exponent <= '0';
      WHEN "0101110111" =>
            manhi <= conv_std_logic_vector(7419882,24);
            manlo <= conv_std_logic_vector(28305511,28);
           exponent <= '0';
      WHEN "0101111000" =>
            manhi <= conv_std_logic_vector(7443523,24);
            manlo <= conv_std_logic_vector(168012985,28);
           exponent <= '0';
      WHEN "0101111001" =>
            manhi <= conv_std_logic_vector(7467188,24);
            manlo <= conv_std_logic_vector(65779352,28);
           exponent <= '0';
      WHEN "0101111010" =>
            manhi <= conv_std_logic_vector(7490875,24);
            manlo <= conv_std_logic_vector(264533668,28);
           exponent <= '0';
      WHEN "0101111011" =>
            manhi <= conv_std_logic_vector(7514586,24);
            manlo <= conv_std_logic_vector(233469080,28);
           exponent <= '0';
      WHEN "0101111100" =>
            manhi <= conv_std_logic_vector(7538320,24);
            manlo <= conv_std_logic_vector(247091035,28);
           exponent <= '0';
      WHEN "0101111101" =>
            manhi <= conv_std_logic_vector(7562078,24);
            manlo <= conv_std_logic_vector(43039991,28);
           exponent <= '0';
      WHEN "0101111110" =>
            manhi <= conv_std_logic_vector(7585858,24);
            manlo <= conv_std_logic_vector(164268716,28);
           exponent <= '0';
      WHEN "0101111111" =>
            manhi <= conv_std_logic_vector(7609662,24);
            manlo <= conv_std_logic_vector(79994093,28);
           exponent <= '0';
      WHEN "0110000000" =>
            manhi <= conv_std_logic_vector(7633489,24);
            manlo <= conv_std_logic_vector(64745322,28);
           exponent <= '0';
      WHEN "0110000001" =>
            manhi <= conv_std_logic_vector(7657339,24);
            manlo <= conv_std_logic_vector(124622102,28);
           exponent <= '0';
      WHEN "0110000010" =>
            manhi <= conv_std_logic_vector(7681212,24);
            manlo <= conv_std_logic_vector(265730090,28);
           exponent <= '0';
      WHEN "0110000011" =>
            manhi <= conv_std_logic_vector(7705109,24);
            manlo <= conv_std_logic_vector(225745453,28);
           exponent <= '0';
      WHEN "0110000100" =>
            manhi <= conv_std_logic_vector(7729030,24);
            manlo <= conv_std_logic_vector(10785785,28);
           exponent <= '0';
      WHEN "0110000101" =>
            manhi <= conv_std_logic_vector(7752973,24);
            manlo <= conv_std_logic_vector(163845570,28);
           exponent <= '0';
      WHEN "0110000110" =>
            manhi <= conv_std_logic_vector(7776940,24);
            manlo <= conv_std_logic_vector(154183450,28);
           exponent <= '0';
      WHEN "0110000111" =>
            manhi <= conv_std_logic_vector(7800930,24);
            manlo <= conv_std_logic_vector(256370426,28);
           exponent <= '0';
      WHEN "0110001000" =>
            manhi <= conv_std_logic_vector(7824944,24);
            manlo <= conv_std_logic_vector(208112577,28);
           exponent <= '0';
      WHEN "0110001001" =>
            manhi <= conv_std_logic_vector(7848982,24);
            manlo <= conv_std_logic_vector(15557444,28);
           exponent <= '0';
      WHEN "0110001010" =>
            manhi <= conv_std_logic_vector(7873042,24);
            manlo <= conv_std_logic_vector(221729482,28);
           exponent <= '0';
      WHEN "0110001011" =>
            manhi <= conv_std_logic_vector(7897127,24);
            manlo <= conv_std_logic_vector(27481881,28);
           exponent <= '0';
      WHEN "0110001100" =>
            manhi <= conv_std_logic_vector(7921234,24);
            manlo <= conv_std_logic_vector(244286584,28);
           exponent <= '0';
      WHEN "0110001101" =>
            manhi <= conv_std_logic_vector(7945366,24);
            manlo <= conv_std_logic_vector(73008824,28);
           exponent <= '0';
      WHEN "0110001110" =>
            manhi <= conv_std_logic_vector(7969521,24);
            manlo <= conv_std_logic_vector(56697140,28);
           exponent <= '0';
      WHEN "0110001111" =>
            manhi <= conv_std_logic_vector(7993699,24);
            manlo <= conv_std_logic_vector(201535196,28);
           exponent <= '0';
      WHEN "0110010000" =>
            manhi <= conv_std_logic_vector(8017901,24);
            manlo <= conv_std_logic_vector(245277246,28);
           exponent <= '0';
      WHEN "0110010001" =>
            manhi <= conv_std_logic_vector(8042127,24);
            manlo <= conv_std_logic_vector(194119042,28);
           exponent <= '0';
      WHEN "0110010010" =>
            manhi <= conv_std_logic_vector(8066377,24);
            manlo <= conv_std_logic_vector(54262392,28);
           exponent <= '0';
      WHEN "0110010011" =>
            manhi <= conv_std_logic_vector(8090650,24);
            manlo <= conv_std_logic_vector(100350618,28);
           exponent <= '0';
      WHEN "0110010100" =>
            manhi <= conv_std_logic_vector(8114947,24);
            manlo <= conv_std_logic_vector(70162199,28);
           exponent <= '0';
      WHEN "0110010101" =>
            manhi <= conv_std_logic_vector(8139267,24);
            manlo <= conv_std_logic_vector(238352593,28);
           exponent <= '0';
      WHEN "0110010110" =>
            manhi <= conv_std_logic_vector(8163612,24);
            manlo <= conv_std_logic_vector(74276969,28);
           exponent <= '0';
      WHEN "0110010111" =>
            manhi <= conv_std_logic_vector(8187980,24);
            manlo <= conv_std_logic_vector(121038404,28);
           exponent <= '0';
      WHEN "0110011000" =>
            manhi <= conv_std_logic_vector(8212372,24);
            manlo <= conv_std_logic_vector(116439694,28);
           exponent <= '0';
      WHEN "0110011001" =>
            manhi <= conv_std_logic_vector(8236788,24);
            manlo <= conv_std_logic_vector(66725186,28);
           exponent <= '0';
      WHEN "0110011010" =>
            manhi <= conv_std_logic_vector(8261227,24);
            manlo <= conv_std_logic_vector(246580788,28);
           exponent <= '0';
      WHEN "0110011011" =>
            manhi <= conv_std_logic_vector(8285691,24);
            manlo <= conv_std_logic_vector(125392143,28);
           exponent <= '0';
      WHEN "0110011100" =>
            manhi <= conv_std_logic_vector(8310178,24);
            manlo <= conv_std_logic_vector(246292830,28);
           exponent <= '0';
      WHEN "0110011101" =>
            manhi <= conv_std_logic_vector(8334690,24);
            manlo <= conv_std_logic_vector(78680728,28);
           exponent <= '0';
      WHEN "0110011110" =>
            manhi <= conv_std_logic_vector(8359225,24);
            manlo <= conv_std_logic_vector(165701659,28);
           exponent <= '0';
      WHEN "0110011111" =>
            manhi <= conv_std_logic_vector(8383784,24);
            manlo <= conv_std_logic_vector(245201212,28);
           exponent <= '0';
      WHEN "0110100000" =>
            manhi <= conv_std_logic_vector(8408368,24);
            manlo <= conv_std_logic_vector(55031110,28);
           exponent <= '0';
      WHEN "0110100001" =>
            manhi <= conv_std_logic_vector(8432975,24);
            manlo <= conv_std_logic_vector(138355589,28);
           exponent <= '0';
      WHEN "0110100010" =>
            manhi <= conv_std_logic_vector(8457606,24);
            manlo <= conv_std_logic_vector(233038665,28);
           exponent <= '0';
      WHEN "0110100011" =>
            manhi <= conv_std_logic_vector(8482262,24);
            manlo <= conv_std_logic_vector(76950508,28);
           exponent <= '0';
      WHEN "0110100100" =>
            manhi <= conv_std_logic_vector(8506941,24);
            manlo <= conv_std_logic_vector(213273820,28);
           exponent <= '0';
      WHEN "0110100101" =>
            manhi <= conv_std_logic_vector(8531645,24);
            manlo <= conv_std_logic_vector(111455640,28);
           exponent <= '0';
      WHEN "0110100110" =>
            manhi <= conv_std_logic_vector(8556373,24);
            manlo <= conv_std_logic_vector(46255554,28);
           exponent <= '0';
      WHEN "0110100111" =>
            manhi <= conv_std_logic_vector(8581125,24);
            manlo <= conv_std_logic_vector(24003868,28);
           exponent <= '0';
      WHEN "0110101000" =>
            manhi <= conv_std_logic_vector(8605901,24);
            manlo <= conv_std_logic_vector(51037072,28);
           exponent <= '0';
      WHEN "0110101001" =>
            manhi <= conv_std_logic_vector(8630701,24);
            manlo <= conv_std_logic_vector(133697849,28);
           exponent <= '0';
      WHEN "0110101010" =>
            manhi <= conv_std_logic_vector(8655526,24);
            manlo <= conv_std_logic_vector(9899623,28);
           exponent <= '0';
      WHEN "0110101011" =>
            manhi <= conv_std_logic_vector(8680374,24);
            manlo <= conv_std_logic_vector(222868388,28);
           exponent <= '0';
      WHEN "0110101100" =>
            manhi <= conv_std_logic_vector(8705247,24);
            manlo <= conv_std_logic_vector(242094523,28);
           exponent <= '0';
      WHEN "0110101101" =>
            manhi <= conv_std_logic_vector(8730145,24);
            manlo <= conv_std_logic_vector(73945536,28);
           exponent <= '0';
      WHEN "0110101110" =>
            manhi <= conv_std_logic_vector(8755066,24);
            manlo <= conv_std_logic_vector(261666066,28);
           exponent <= '0';
      WHEN "0110101111" =>
            manhi <= conv_std_logic_vector(8780013,24);
            manlo <= conv_std_logic_vector(6329700,28);
           exponent <= '0';
      WHEN "0110110000" =>
            manhi <= conv_std_logic_vector(8804983,24);
            manlo <= conv_std_logic_vector(119628997,28);
           exponent <= '0';
      WHEN "0110110001" =>
            manhi <= conv_std_logic_vector(8829978,24);
            manlo <= conv_std_logic_vector(71085473,28);
           exponent <= '0';
      WHEN "0110110010" =>
            manhi <= conv_std_logic_vector(8854997,24);
            manlo <= conv_std_logic_vector(135533257,28);
           exponent <= '0';
      WHEN "0110110011" =>
            manhi <= conv_std_logic_vector(8880041,24);
            manlo <= conv_std_logic_vector(50941820,28);
           exponent <= '0';
      WHEN "0110110100" =>
            manhi <= conv_std_logic_vector(8905109,24);
            manlo <= conv_std_logic_vector(92157802,28);
           exponent <= '0';
      WHEN "0110110101" =>
            manhi <= conv_std_logic_vector(8930201,24);
            manlo <= conv_std_logic_vector(265598650,28);
           exponent <= '0';
      WHEN "0110110110" =>
            manhi <= conv_std_logic_vector(8955319,24);
            manlo <= conv_std_logic_vector(40817170,28);
           exponent <= '0';
      WHEN "0110110111" =>
            manhi <= conv_std_logic_vector(8980460,24);
            manlo <= conv_std_logic_vector(229549724,28);
           exponent <= '0';
      WHEN "0110111000" =>
            manhi <= conv_std_logic_vector(9005627,24);
            manlo <= conv_std_logic_vector(32926222,28);
           exponent <= '0';
      WHEN "0110111001" =>
            manhi <= conv_std_logic_vector(9030817,24);
            manlo <= conv_std_logic_vector(262695596,28);
           exponent <= '0';
      WHEN "0110111010" =>
            manhi <= conv_std_logic_vector(9056033,24);
            manlo <= conv_std_logic_vector(120000337,28);
           exponent <= '0';
      WHEN "0110111011" =>
            manhi <= conv_std_logic_vector(9081273,24);
            manlo <= conv_std_logic_vector(148166518,28);
           exponent <= '0';
      WHEN "0110111100" =>
            manhi <= conv_std_logic_vector(9106538,24);
            manlo <= conv_std_logic_vector(85220151,28);
           exponent <= '0';
      WHEN "0110111101" =>
            manhi <= conv_std_logic_vector(9131827,24);
            manlo <= conv_std_logic_vector(206064472,28);
           exponent <= '0';
      WHEN "0110111110" =>
            manhi <= conv_std_logic_vector(9157141,24);
            manlo <= conv_std_logic_vector(248738124,28);
           exponent <= '0';
      WHEN "0110111111" =>
            manhi <= conv_std_logic_vector(9182480,24);
            manlo <= conv_std_logic_vector(219721533,28);
           exponent <= '0';
      WHEN "0111000000" =>
            manhi <= conv_std_logic_vector(9207844,24);
            manlo <= conv_std_logic_vector(125501456,28);
           exponent <= '0';
      WHEN "0111000001" =>
            manhi <= conv_std_logic_vector(9233232,24);
            manlo <= conv_std_logic_vector(241006443,28);
           exponent <= '0';
      WHEN "0111000010" =>
            manhi <= conv_std_logic_vector(9258646,24);
            manlo <= conv_std_logic_vector(35865021,28);
           exponent <= '0';
      WHEN "0111000011" =>
            manhi <= conv_std_logic_vector(9284084,24);
            manlo <= conv_std_logic_vector(53453891,28);
           exponent <= '0';
      WHEN "0111000100" =>
            manhi <= conv_std_logic_vector(9309547,24);
            manlo <= conv_std_logic_vector(31849742,28);
           exponent <= '0';
      WHEN "0111000101" =>
            manhi <= conv_std_logic_vector(9335034,24);
            manlo <= conv_std_logic_vector(246006538,28);
           exponent <= '0';
      WHEN "0111000110" =>
            manhi <= conv_std_logic_vector(9360547,24);
            manlo <= conv_std_logic_vector(165578245,28);
           exponent <= '0';
      WHEN "0111000111" =>
            manhi <= conv_std_logic_vector(9386085,24);
            manlo <= conv_std_logic_vector(65531569,28);
           exponent <= '0';
      WHEN "0111001000" =>
            manhi <= conv_std_logic_vector(9411647,24);
            manlo <= conv_std_logic_vector(220839600,28);
           exponent <= '0';
      WHEN "0111001001" =>
            manhi <= conv_std_logic_vector(9437235,24);
            manlo <= conv_std_logic_vector(101175446,28);
           exponent <= '0';
      WHEN "0111001010" =>
            manhi <= conv_std_logic_vector(9462847,24);
            manlo <= conv_std_logic_vector(249960434,28);
           exponent <= '0';
      WHEN "0111001011" =>
            manhi <= conv_std_logic_vector(9488485,24);
            manlo <= conv_std_logic_vector(136880466,28);
           exponent <= '0';
      WHEN "0111001100" =>
            manhi <= conv_std_logic_vector(9514148,24);
            manlo <= conv_std_logic_vector(36934219,28);
           exponent <= '0';
      WHEN "0111001101" =>
            manhi <= conv_std_logic_vector(9539835,24);
            manlo <= conv_std_logic_vector(225126782,28);
           exponent <= '0';
      WHEN "0111001110" =>
            manhi <= conv_std_logic_vector(9565548,24);
            manlo <= conv_std_logic_vector(171163295,28);
           exponent <= '0';
      WHEN "0111001111" =>
            manhi <= conv_std_logic_vector(9591286,24);
            manlo <= conv_std_logic_vector(150061692,28);
           exponent <= '0';
      WHEN "0111010000" =>
            manhi <= conv_std_logic_vector(9617049,24);
            manlo <= conv_std_logic_vector(168410880,28);
           exponent <= '0';
      WHEN "0111010001" =>
            manhi <= conv_std_logic_vector(9642837,24);
            manlo <= conv_std_logic_vector(232806206,28);
           exponent <= '0';
      WHEN "0111010010" =>
            manhi <= conv_std_logic_vector(9668651,24);
            manlo <= conv_std_logic_vector(81414002,28);
           exponent <= '0';
      WHEN "0111010011" =>
            manhi <= conv_std_logic_vector(9694489,24);
            manlo <= conv_std_logic_vector(257713424,28);
           exponent <= '0';
      WHEN "0111010100" =>
            manhi <= conv_std_logic_vector(9720353,24);
            manlo <= conv_std_logic_vector(231448253,28);
           exponent <= '0';
      WHEN "0111010101" =>
            manhi <= conv_std_logic_vector(9746243,24);
            manlo <= conv_std_logic_vector(9239650,28);
           exponent <= '0';
      WHEN "0111010110" =>
            manhi <= conv_std_logic_vector(9772157,24);
            manlo <= conv_std_logic_vector(134586155,28);
           exponent <= '0';
      WHEN "0111010111" =>
            manhi <= conv_std_logic_vector(9798097,24);
            manlo <= conv_std_logic_vector(77250961,28);
           exponent <= '0';
      WHEN "0111011000" =>
            manhi <= conv_std_logic_vector(9824062,24);
            manlo <= conv_std_logic_vector(112310110,28);
           exponent <= '0';
      WHEN "0111011001" =>
            manhi <= conv_std_logic_vector(9850052,24);
            manlo <= conv_std_logic_vector(246410674,28);
           exponent <= '0';
      WHEN "0111011010" =>
            manhi <= conv_std_logic_vector(9876068,24);
            manlo <= conv_std_logic_vector(217770768,28);
           exponent <= '0';
      WHEN "0111011011" =>
            manhi <= conv_std_logic_vector(9902110,24);
            manlo <= conv_std_logic_vector(33050459,28);
           exponent <= '0';
      WHEN "0111011100" =>
            manhi <= conv_std_logic_vector(9928176,24);
            manlo <= conv_std_logic_vector(235787236,28);
           exponent <= '0';
      WHEN "0111011101" =>
            manhi <= conv_std_logic_vector(9954269,24);
            manlo <= conv_std_logic_vector(27347822,28);
           exponent <= '0';
      WHEN "0111011110" =>
            manhi <= conv_std_logic_vector(9980386,24);
            manlo <= conv_std_logic_vector(219718194,28);
           exponent <= '0';
      WHEN "0111011111" =>
            manhi <= conv_std_logic_vector(10006530,24);
            manlo <= conv_std_logic_vector(14278120,28);
           exponent <= '0';
      WHEN "0111100000" =>
            manhi <= conv_std_logic_vector(10032698,24);
            manlo <= conv_std_logic_vector(223026636,28);
           exponent <= '0';
      WHEN "0111100001" =>
            manhi <= conv_std_logic_vector(10058893,24);
            manlo <= conv_std_logic_vector(47356582,28);
           exponent <= '0';
      WHEN "0111100010" =>
            manhi <= conv_std_logic_vector(10085113,24);
            manlo <= conv_std_logic_vector(30844624,28);
           exponent <= '0';
      WHEN "0111100011" =>
            manhi <= conv_std_logic_vector(10111358,24);
            manlo <= conv_std_logic_vector(180203065,28);
           exponent <= '0';
      WHEN "0111100100" =>
            manhi <= conv_std_logic_vector(10137629,24);
            manlo <= conv_std_logic_vector(233715314,28);
           exponent <= '0';
      WHEN "0111100101" =>
            manhi <= conv_std_logic_vector(10163926,24);
            manlo <= conv_std_logic_vector(198106796,28);
           exponent <= '0';
      WHEN "0111100110" =>
            manhi <= conv_std_logic_vector(10190249,24);
            manlo <= conv_std_logic_vector(80109512,28);
           exponent <= '0';
      WHEN "0111100111" =>
            manhi <= conv_std_logic_vector(10216597,24);
            manlo <= conv_std_logic_vector(154897493,28);
           exponent <= '0';
      WHEN "0111101000" =>
            manhi <= conv_std_logic_vector(10242971,24);
            manlo <= conv_std_logic_vector(160780443,28);
           exponent <= '0';
      WHEN "0111101001" =>
            manhi <= conv_std_logic_vector(10269371,24);
            manlo <= conv_std_logic_vector(104510112,28);
           exponent <= '0';
      WHEN "0111101010" =>
            manhi <= conv_std_logic_vector(10295796,24);
            manlo <= conv_std_logic_vector(261280303,28);
           exponent <= '0';
      WHEN "0111101011" =>
            manhi <= conv_std_logic_vector(10322248,24);
            manlo <= conv_std_logic_vector(100985054,28);
           exponent <= '0';
      WHEN "0111101100" =>
            manhi <= conv_std_logic_vector(10348725,24);
            manlo <= conv_std_logic_vector(167266836,28);
           exponent <= '0';
      WHEN "0111101101" =>
            manhi <= conv_std_logic_vector(10375228,24);
            manlo <= conv_std_logic_vector(198468370,28);
           exponent <= '0';
      WHEN "0111101110" =>
            manhi <= conv_std_logic_vector(10401757,24);
            manlo <= conv_std_logic_vector(201374454,28);
           exponent <= '0';
      WHEN "0111101111" =>
            manhi <= conv_std_logic_vector(10428312,24);
            manlo <= conv_std_logic_vector(182776514,28);
           exponent <= '0';
      WHEN "0111110000" =>
            manhi <= conv_std_logic_vector(10454893,24);
            manlo <= conv_std_logic_vector(149472614,28);
           exponent <= '0';
      WHEN "0111110001" =>
            manhi <= conv_std_logic_vector(10481500,24);
            manlo <= conv_std_logic_vector(108267459,28);
           exponent <= '0';
      WHEN "0111110010" =>
            manhi <= conv_std_logic_vector(10508133,24);
            manlo <= conv_std_logic_vector(65972402,28);
           exponent <= '0';
      WHEN "0111110011" =>
            manhi <= conv_std_logic_vector(10534792,24);
            manlo <= conv_std_logic_vector(29405451,28);
           exponent <= '0';
      WHEN "0111110100" =>
            manhi <= conv_std_logic_vector(10561477,24);
            manlo <= conv_std_logic_vector(5391275,28);
           exponent <= '0';
      WHEN "0111110101" =>
            manhi <= conv_std_logic_vector(10588188,24);
            manlo <= conv_std_logic_vector(761213,28);
           exponent <= '0';
      WHEN "0111110110" =>
            manhi <= conv_std_logic_vector(10614925,24);
            manlo <= conv_std_logic_vector(22353276,28);
           exponent <= '0';
      WHEN "0111110111" =>
            manhi <= conv_std_logic_vector(10641688,24);
            manlo <= conv_std_logic_vector(77012158,28);
           exponent <= '0';
      WHEN "0111111000" =>
            manhi <= conv_std_logic_vector(10668477,24);
            manlo <= conv_std_logic_vector(171589240,28);
           exponent <= '0';
      WHEN "0111111001" =>
            manhi <= conv_std_logic_vector(10695293,24);
            manlo <= conv_std_logic_vector(44507139,28);
           exponent <= '0';
      WHEN "0111111010" =>
            manhi <= conv_std_logic_vector(10722134,24);
            manlo <= conv_std_logic_vector(239501544,28);
           exponent <= '0';
      WHEN "0111111011" =>
            manhi <= conv_std_logic_vector(10749002,24);
            manlo <= conv_std_logic_vector(226573024,28);
           exponent <= '0';
      WHEN "0111111100" =>
            manhi <= conv_std_logic_vector(10775897,24);
            manlo <= conv_std_logic_vector(12599777,28);
           exponent <= '0';
      WHEN "0111111101" =>
            manhi <= conv_std_logic_vector(10802817,24);
            manlo <= conv_std_logic_vector(141337630,28);
           exponent <= '0';
      WHEN "0111111110" =>
            manhi <= conv_std_logic_vector(10829764,24);
            manlo <= conv_std_logic_vector(82807315,28);
           exponent <= '0';
      WHEN "0111111111" =>
            manhi <= conv_std_logic_vector(10856737,24);
            manlo <= conv_std_logic_vector(112342665,28);
           exponent <= '0';
      WHEN "1000000000" =>
            manhi <= conv_std_logic_vector(10883736,24);
            manlo <= conv_std_logic_vector(236848796,28);
           exponent <= '0';
      WHEN "1000000001" =>
            manhi <= conv_std_logic_vector(10910762,24);
            manlo <= conv_std_logic_vector(194802116,28);
           exponent <= '0';
      WHEN "1000000010" =>
            manhi <= conv_std_logic_vector(10937814,24);
            manlo <= conv_std_logic_vector(261556696,28);
           exponent <= '0';
      WHEN "1000000011" =>
            manhi <= conv_std_logic_vector(10964893,24);
            manlo <= conv_std_logic_vector(175602458,28);
           exponent <= '0';
      WHEN "1000000100" =>
            manhi <= conv_std_logic_vector(10991998,24);
            manlo <= conv_std_logic_vector(212307000,28);
           exponent <= '0';
      WHEN "1000000101" =>
            manhi <= conv_std_logic_vector(11019130,24);
            manlo <= conv_std_logic_vector(110173782,28);
           exponent <= '0';
      WHEN "1000000110" =>
            manhi <= conv_std_logic_vector(11046288,24);
            manlo <= conv_std_logic_vector(144583954,28);
           exponent <= '0';
      WHEN "1000000111" =>
            manhi <= conv_std_logic_vector(11073473,24);
            manlo <= conv_std_logic_vector(54054542,28);
           exponent <= '0';
      WHEN "1000001000" =>
            manhi <= conv_std_logic_vector(11100684,24);
            manlo <= conv_std_logic_vector(113980276,28);
           exponent <= '0';
      WHEN "1000001001" =>
            manhi <= conv_std_logic_vector(11127922,24);
            manlo <= conv_std_logic_vector(62891774,28);
           exponent <= '0';
      WHEN "1000001010" =>
            manhi <= conv_std_logic_vector(11155186,24);
            manlo <= conv_std_logic_vector(176197372,28);
           exponent <= '0';
      WHEN "1000001011" =>
            manhi <= conv_std_logic_vector(11182477,24);
            manlo <= conv_std_logic_vector(192441306,28);
           exponent <= '0';
      WHEN "1000001100" =>
            manhi <= conv_std_logic_vector(11209795,24);
            manlo <= conv_std_logic_vector(118610088,28);
           exponent <= '0';
      WHEN "1000001101" =>
            manhi <= conv_std_logic_vector(11237139,24);
            manlo <= conv_std_logic_vector(230132514,28);
           exponent <= '0';
      WHEN "1000001110" =>
            manhi <= conv_std_logic_vector(11264510,24);
            manlo <= conv_std_logic_vector(265573296,28);
           exponent <= '0';
      WHEN "1000001111" =>
            manhi <= conv_std_logic_vector(11291908,24);
            manlo <= conv_std_logic_vector(231939446,28);
           exponent <= '0';
      WHEN "1000010000" =>
            manhi <= conv_std_logic_vector(11319333,24);
            manlo <= conv_std_logic_vector(136244820,28);
           exponent <= '0';
      WHEN "1000010001" =>
            manhi <= conv_std_logic_vector(11346784,24);
            manlo <= conv_std_logic_vector(253945584,28);
           exponent <= '0';
      WHEN "1000010010" =>
            manhi <= conv_std_logic_vector(11374263,24);
            manlo <= conv_std_logic_vector(55198395,28);
           exponent <= '0';
      WHEN "1000010011" =>
            manhi <= conv_std_logic_vector(11401768,24);
            manlo <= conv_std_logic_vector(83908598,28);
           exponent <= '0';
      WHEN "1000010100" =>
            manhi <= conv_std_logic_vector(11429300,24);
            manlo <= conv_std_logic_vector(78682048,28);
           exponent <= '0';
      WHEN "1000010101" =>
            manhi <= conv_std_logic_vector(11456859,24);
            manlo <= conv_std_logic_vector(46566930,28);
           exponent <= '0';
      WHEN "1000010110" =>
            manhi <= conv_std_logic_vector(11484444,24);
            manlo <= conv_std_logic_vector(263053774,28);
           exponent <= '0';
      WHEN "1000010111" =>
            manhi <= conv_std_logic_vector(11512057,24);
            manlo <= conv_std_logic_vector(198333637,28);
           exponent <= '0';
      WHEN "1000011000" =>
            manhi <= conv_std_logic_vector(11539697,24);
            manlo <= conv_std_logic_vector(127910840,28);
           exponent <= '0';
      WHEN "1000011001" =>
            manhi <= conv_std_logic_vector(11567364,24);
            manlo <= conv_std_logic_vector(58861158,28);
           exponent <= '0';
      WHEN "1000011010" =>
            manhi <= conv_std_logic_vector(11595057,24);
            manlo <= conv_std_logic_vector(266702732,28);
           exponent <= '0';
      WHEN "1000011011" =>
            manhi <= conv_std_logic_vector(11622778,24);
            manlo <= conv_std_logic_vector(221654258,28);
           exponent <= '0';
      WHEN "1000011100" =>
            manhi <= conv_std_logic_vector(11650526,24);
            manlo <= conv_std_logic_vector(199247725,28);
           exponent <= '0';
      WHEN "1000011101" =>
            manhi <= conv_std_logic_vector(11678301,24);
            manlo <= conv_std_logic_vector(206586600,28);
           exponent <= '0';
      WHEN "1000011110" =>
            manhi <= conv_std_logic_vector(11706103,24);
            manlo <= conv_std_logic_vector(250781292,28);
           exponent <= '0';
      WHEN "1000011111" =>
            manhi <= conv_std_logic_vector(11733933,24);
            manlo <= conv_std_logic_vector(70513697,28);
           exponent <= '0';
      WHEN "1000100000" =>
            manhi <= conv_std_logic_vector(11761789,24);
            manlo <= conv_std_logic_vector(209779039,28);
           exponent <= '0';
      WHEN "1000100001" =>
            manhi <= conv_std_logic_vector(11789673,24);
            manlo <= conv_std_logic_vector(138837672,28);
           exponent <= '0';
      WHEN "1000100010" =>
            manhi <= conv_std_logic_vector(11817584,24);
            manlo <= conv_std_logic_vector(133263292,28);
           exponent <= '0';
      WHEN "1000100011" =>
            manhi <= conv_std_logic_vector(11845522,24);
            manlo <= conv_std_logic_vector(200201109,28);
           exponent <= '0';
      WHEN "1000100100" =>
            manhi <= conv_std_logic_vector(11873488,24);
            manlo <= conv_std_logic_vector(78367858,28);
           exponent <= '0';
      WHEN "1000100101" =>
            manhi <= conv_std_logic_vector(11901481,24);
            manlo <= conv_std_logic_vector(43358178,28);
           exponent <= '0';
      WHEN "1000100110" =>
            manhi <= conv_std_logic_vector(11929501,24);
            manlo <= conv_std_logic_vector(102338242,28);
           exponent <= '0';
      WHEN "1000100111" =>
            manhi <= conv_std_logic_vector(11957548,24);
            manlo <= conv_std_logic_vector(262481228,28);
           exponent <= '0';
      WHEN "1000101000" =>
            manhi <= conv_std_logic_vector(11985623,24);
            manlo <= conv_std_logic_vector(262531864,28);
           exponent <= '0';
      WHEN "1000101001" =>
            manhi <= conv_std_logic_vector(12013726,24);
            manlo <= conv_std_logic_vector(109677352,28);
           exponent <= '0';
      WHEN "1000101010" =>
            manhi <= conv_std_logic_vector(12041856,24);
            manlo <= conv_std_logic_vector(79547371,28);
           exponent <= '0';
      WHEN "1000101011" =>
            manhi <= conv_std_logic_vector(12070013,24);
            manlo <= conv_std_logic_vector(179343172,28);
           exponent <= '0';
      WHEN "1000101100" =>
            manhi <= conv_std_logic_vector(12098198,24);
            manlo <= conv_std_logic_vector(147837587,28);
           exponent <= '0';
      WHEN "1000101101" =>
            manhi <= conv_std_logic_vector(12126410,24);
            manlo <= conv_std_logic_vector(260681402,28);
           exponent <= '0';
      WHEN "1000101110" =>
            manhi <= conv_std_logic_vector(12154650,24);
            manlo <= conv_std_logic_vector(256661542,28);
           exponent <= '0';
      WHEN "1000101111" =>
            manhi <= conv_std_logic_vector(12182918,24);
            manlo <= conv_std_logic_vector(143007443,28);
           exponent <= '0';
      WHEN "1000110000" =>
            manhi <= conv_std_logic_vector(12211213,24);
            manlo <= conv_std_logic_vector(195391062,28);
           exponent <= '0';
      WHEN "1000110001" =>
            manhi <= conv_std_logic_vector(12239536,24);
            manlo <= conv_std_logic_vector(152620513,28);
           exponent <= '0';
      WHEN "1000110010" =>
            manhi <= conv_std_logic_vector(12267887,24);
            manlo <= conv_std_logic_vector(21946444,28);
           exponent <= '0';
      WHEN "1000110011" =>
            manhi <= conv_std_logic_vector(12296265,24);
            manlo <= conv_std_logic_vector(79062042,28);
           exponent <= '0';
      WHEN "1000110100" =>
            manhi <= conv_std_logic_vector(12324671,24);
            manlo <= conv_std_logic_vector(62796676,28);
           exponent <= '0';
      WHEN "1000110101" =>
            manhi <= conv_std_logic_vector(12353104,24);
            manlo <= conv_std_logic_vector(248857722,28);
           exponent <= '0';
      WHEN "1000110110" =>
            manhi <= conv_std_logic_vector(12381566,24);
            manlo <= conv_std_logic_vector(107653293,28);
           exponent <= '0';
      WHEN "1000110111" =>
            manhi <= conv_std_logic_vector(12410055,24);
            manlo <= conv_std_logic_vector(183340440,28);
           exponent <= '0';
      WHEN "1000111000" =>
            manhi <= conv_std_logic_vector(12438572,24);
            manlo <= conv_std_logic_vector(214776964,28);
           exponent <= '0';
      WHEN "1000111001" =>
            manhi <= conv_std_logic_vector(12467117,24);
            manlo <= conv_std_logic_vector(209263248,28);
           exponent <= '0';
      WHEN "1000111010" =>
            manhi <= conv_std_logic_vector(12495690,24);
            manlo <= conv_std_logic_vector(174106806,28);
           exponent <= '0';
      WHEN "1000111011" =>
            manhi <= conv_std_logic_vector(12524291,24);
            manlo <= conv_std_logic_vector(116622293,28);
           exponent <= '0';
      WHEN "1000111100" =>
            manhi <= conv_std_logic_vector(12552920,24);
            manlo <= conv_std_logic_vector(44131512,28);
           exponent <= '0';
      WHEN "1000111101" =>
            manhi <= conv_std_logic_vector(12581576,24);
            manlo <= conv_std_logic_vector(232398874,28);
           exponent <= '0';
      WHEN "1000111110" =>
            manhi <= conv_std_logic_vector(12610261,24);
            manlo <= conv_std_logic_vector(151889582,28);
           exponent <= '0';
      WHEN "1000111111" =>
            manhi <= conv_std_logic_vector(12638974,24);
            manlo <= conv_std_logic_vector(78382378,28);
           exponent <= '0';
      WHEN "1001000000" =>
            manhi <= conv_std_logic_vector(12667715,24);
            manlo <= conv_std_logic_vector(19227718,28);
           exponent <= '0';
      WHEN "1001000001" =>
            manhi <= conv_std_logic_vector(12696483,24);
            manlo <= conv_std_logic_vector(250218700,28);
           exponent <= '0';
      WHEN "1001000010" =>
            manhi <= conv_std_logic_vector(12725280,24);
            manlo <= conv_std_logic_vector(241849240,28);
           exponent <= '0';
      WHEN "1001000011" =>
            manhi <= conv_std_logic_vector(12754106,24);
            manlo <= conv_std_logic_vector(1491364,28);
           exponent <= '0';
      WHEN "1001000100" =>
            manhi <= conv_std_logic_vector(12782959,24);
            manlo <= conv_std_logic_vector(73395209,28);
           exponent <= '0';
      WHEN "1001000101" =>
            manhi <= conv_std_logic_vector(12811840,24);
            manlo <= conv_std_logic_vector(196511758,28);
           exponent <= '0';
      WHEN "1001000110" =>
            manhi <= conv_std_logic_vector(12840750,24);
            manlo <= conv_std_logic_vector(109799208,28);
           exponent <= '0';
      WHEN "1001000111" =>
            manhi <= conv_std_logic_vector(12869688,24);
            manlo <= conv_std_logic_vector(89093893,28);
           exponent <= '0';
      WHEN "1001001000" =>
            manhi <= conv_std_logic_vector(12898654,24);
            manlo <= conv_std_logic_vector(141803923,28);
           exponent <= '0';
      WHEN "1001001001" =>
            manhi <= conv_std_logic_vector(12927649,24);
            manlo <= conv_std_logic_vector(6909187,28);
           exponent <= '0';
      WHEN "1001001010" =>
            manhi <= conv_std_logic_vector(12956671,24);
            manlo <= conv_std_logic_vector(228703191,28);
           exponent <= '0';
      WHEN "1001001011" =>
            manhi <= conv_std_logic_vector(12985723,24);
            manlo <= conv_std_logic_vector(9309409,28);
           exponent <= '0';
      WHEN "1001001100" =>
            manhi <= conv_std_logic_vector(13014802,24);
            manlo <= conv_std_logic_vector(161471314,28);
           exponent <= '0';
      WHEN "1001001101" =>
            manhi <= conv_std_logic_vector(13043910,24);
            manlo <= conv_std_logic_vector(155762363,28);
           exponent <= '0';
      WHEN "1001001110" =>
            manhi <= conv_std_logic_vector(13073046,24);
            manlo <= conv_std_logic_vector(268069656,28);
           exponent <= '0';
      WHEN "1001001111" =>
            manhi <= conv_std_logic_vector(13102211,24);
            manlo <= conv_std_logic_vector(237416659,28);
           exponent <= '0';
      WHEN "1001010000" =>
            manhi <= conv_std_logic_vector(13131405,24);
            manlo <= conv_std_logic_vector(71269584,28);
           exponent <= '0';
      WHEN "1001010001" =>
            manhi <= conv_std_logic_vector(13160627,24);
            manlo <= conv_std_logic_vector(45537394,28);
           exponent <= '0';
      WHEN "1001010010" =>
            manhi <= conv_std_logic_vector(13189877,24);
            manlo <= conv_std_logic_vector(167700897,28);
           exponent <= '0';
      WHEN "1001010011" =>
            manhi <= conv_std_logic_vector(13219156,24);
            manlo <= conv_std_logic_vector(176812753,28);
           exponent <= '0';
      WHEN "1001010100" =>
            manhi <= conv_std_logic_vector(13248464,24);
            manlo <= conv_std_logic_vector(80368396,28);
           exponent <= '0';
      WHEN "1001010101" =>
            manhi <= conv_std_logic_vector(13277800,24);
            manlo <= conv_std_logic_vector(154306039,28);
           exponent <= '0';
      WHEN "1001010110" =>
            manhi <= conv_std_logic_vector(13307165,24);
            manlo <= conv_std_logic_vector(137700312,28);
           exponent <= '0';
      WHEN "1001010111" =>
            manhi <= conv_std_logic_vector(13336559,24);
            manlo <= conv_std_logic_vector(38068641,28);
           exponent <= '0';
      WHEN "1001011000" =>
            manhi <= conv_std_logic_vector(13365981,24);
            manlo <= conv_std_logic_vector(131371250,28);
           exponent <= '0';
      WHEN "1001011001" =>
            manhi <= conv_std_logic_vector(13395432,24);
            manlo <= conv_std_logic_vector(156704806,28);
           exponent <= '0';
      WHEN "1001011010" =>
            manhi <= conv_std_logic_vector(13424912,24);
            manlo <= conv_std_logic_vector(121608790,28);
           exponent <= '0';
      WHEN "1001011011" =>
            manhi <= conv_std_logic_vector(13454421,24);
            manlo <= conv_std_logic_vector(33630048,28);
           exponent <= '0';
      WHEN "1001011100" =>
            manhi <= conv_std_logic_vector(13483958,24);
            manlo <= conv_std_logic_vector(168758257,28);
           exponent <= '0';
      WHEN "1001011101" =>
            manhi <= conv_std_logic_vector(13513524,24);
            manlo <= conv_std_logic_vector(266119562,28);
           exponent <= '0';
      WHEN "1001011110" =>
            manhi <= conv_std_logic_vector(13543120,24);
            manlo <= conv_std_logic_vector(64847498,28);
           exponent <= '0';
      WHEN "1001011111" =>
            manhi <= conv_std_logic_vector(13572744,24);
            manlo <= conv_std_logic_vector(109389360,28);
           exponent <= '0';
      WHEN "1001100000" =>
            manhi <= conv_std_logic_vector(13602397,24);
            manlo <= conv_std_logic_vector(138893481,28);
           exponent <= '0';
      WHEN "1001100001" =>
            manhi <= conv_std_logic_vector(13632079,24);
            manlo <= conv_std_logic_vector(160951056,28);
           exponent <= '0';
      WHEN "1001100010" =>
            manhi <= conv_std_logic_vector(13661790,24);
            manlo <= conv_std_logic_vector(183160698,28);
           exponent <= '0';
      WHEN "1001100011" =>
            manhi <= conv_std_logic_vector(13691530,24);
            manlo <= conv_std_logic_vector(213128447,28);
           exponent <= '0';
      WHEN "1001100100" =>
            manhi <= conv_std_logic_vector(13721299,24);
            manlo <= conv_std_logic_vector(258467771,28);
           exponent <= '0';
      WHEN "1001100101" =>
            manhi <= conv_std_logic_vector(13751098,24);
            manlo <= conv_std_logic_vector(58364122,28);
           exponent <= '0';
      WHEN "1001100110" =>
            manhi <= conv_std_logic_vector(13780925,24);
            manlo <= conv_std_logic_vector(157316766,28);
           exponent <= '0';
      WHEN "1001100111" =>
            manhi <= conv_std_logic_vector(13810782,24);
            manlo <= conv_std_logic_vector(26090597,28);
           exponent <= '0';
      WHEN "1001101000" =>
            manhi <= conv_std_logic_vector(13840667,24);
            manlo <= conv_std_logic_vector(209199796,28);
           exponent <= '0';
      WHEN "1001101001" =>
            manhi <= conv_std_logic_vector(13870582,24);
            manlo <= conv_std_logic_vector(177424185,28);
           exponent <= '0';
      WHEN "1001101010" =>
            manhi <= conv_std_logic_vector(13900526,24);
            manlo <= conv_std_logic_vector(206857431,28);
           exponent <= '0';
      WHEN "1001101011" =>
            manhi <= conv_std_logic_vector(13930500,24);
            manlo <= conv_std_logic_vector(36729770,28);
           exponent <= '0';
      WHEN "1001101100" =>
            manhi <= conv_std_logic_vector(13960502,24);
            manlo <= conv_std_logic_vector(211585297,28);
           exponent <= '0';
      WHEN "1001101101" =>
            manhi <= conv_std_logic_vector(13990534,24);
            manlo <= conv_std_logic_vector(202233780,28);
           exponent <= '0';
      WHEN "1001101110" =>
            manhi <= conv_std_logic_vector(14020596,24);
            manlo <= conv_std_logic_vector(16363400,28);
           exponent <= '0';
      WHEN "1001101111" =>
            manhi <= conv_std_logic_vector(14050686,24);
            manlo <= conv_std_logic_vector(198540768,28);
           exponent <= '0';
      WHEN "1001110000" =>
            manhi <= conv_std_logic_vector(14080806,24);
            manlo <= conv_std_logic_vector(219598184,28);
           exponent <= '0';
      WHEN "1001110001" =>
            manhi <= conv_std_logic_vector(14110956,24);
            manlo <= conv_std_logic_vector(87246388,28);
           exponent <= '0';
      WHEN "1001110010" =>
            manhi <= conv_std_logic_vector(14141135,24);
            manlo <= conv_std_logic_vector(77639113,28);
           exponent <= '0';
      WHEN "1001110011" =>
            manhi <= conv_std_logic_vector(14171343,24);
            manlo <= conv_std_logic_vector(198502173,28);
           exponent <= '0';
      WHEN "1001110100" =>
            manhi <= conv_std_logic_vector(14201581,24);
            manlo <= conv_std_logic_vector(189133475,28);
           exponent <= '0';
      WHEN "1001110101" =>
            manhi <= conv_std_logic_vector(14231849,24);
            manlo <= conv_std_logic_vector(57273941,28);
           exponent <= '0';
      WHEN "1001110110" =>
            manhi <= conv_std_logic_vector(14262146,24);
            manlo <= conv_std_logic_vector(79107508,28);
           exponent <= '0';
      WHEN "1001110111" =>
            manhi <= conv_std_logic_vector(14292472,24);
            manlo <= conv_std_logic_vector(262390229,28);
           exponent <= '0';
      WHEN "1001111000" =>
            manhi <= conv_std_logic_vector(14322829,24);
            manlo <= conv_std_logic_vector(78014825,28);
           exponent <= '0';
      WHEN "1001111001" =>
            manhi <= conv_std_logic_vector(14353215,24);
            manlo <= conv_std_logic_vector(70623424,28);
           exponent <= '0';
      WHEN "1001111010" =>
            manhi <= conv_std_logic_vector(14383630,24);
            manlo <= conv_std_logic_vector(247994836,28);
           exponent <= '0';
      WHEN "1001111011" =>
            manhi <= conv_std_logic_vector(14414076,24);
            manlo <= conv_std_logic_vector(81044559,28);
           exponent <= '0';
      WHEN "1001111100" =>
            manhi <= conv_std_logic_vector(14444551,24);
            manlo <= conv_std_logic_vector(114437521,28);
           exponent <= '0';
      WHEN "1001111101" =>
            manhi <= conv_std_logic_vector(14475056,24);
            manlo <= conv_std_logic_vector(87539900,28);
           exponent <= '0';
      WHEN "1001111110" =>
            manhi <= conv_std_logic_vector(14505591,24);
            manlo <= conv_std_logic_vector(8160950,28);
           exponent <= '0';
      WHEN "1001111111" =>
            manhi <= conv_std_logic_vector(14536155,24);
            manlo <= conv_std_logic_vector(152553012,28);
           exponent <= '0';
      WHEN "1010000000" =>
            manhi <= conv_std_logic_vector(14566749,24);
            manlo <= conv_std_logic_vector(260105152,28);
           exponent <= '0';
      WHEN "1010000001" =>
            manhi <= conv_std_logic_vector(14597374,24);
            manlo <= conv_std_logic_vector(70214083,28);
           exponent <= '0';
      WHEN "1010000010" =>
            manhi <= conv_std_logic_vector(14628028,24);
            manlo <= conv_std_logic_vector(127590534,28);
           exponent <= '0';
      WHEN "1010000011" =>
            manhi <= conv_std_logic_vector(14658712,24);
            manlo <= conv_std_logic_vector(171646531,28);
           exponent <= '0';
      WHEN "1010000100" =>
            manhi <= conv_std_logic_vector(14689426,24);
            manlo <= conv_std_logic_vector(210237219,28);
           exponent <= '0';
      WHEN "1010000101" =>
            manhi <= conv_std_logic_vector(14720170,24);
            manlo <= conv_std_logic_vector(251225419,28);
           exponent <= '0';
      WHEN "1010000110" =>
            manhi <= conv_std_logic_vector(14750945,24);
            manlo <= conv_std_logic_vector(34046180,28);
           exponent <= '0';
      WHEN "1010000111" =>
            manhi <= conv_std_logic_vector(14781749,24);
            manlo <= conv_std_logic_vector(103448606,28);
           exponent <= '0';
      WHEN "1010001000" =>
            manhi <= conv_std_logic_vector(14812583,24);
            manlo <= conv_std_logic_vector(198883134,28);
           exponent <= '0';
      WHEN "1010001001" =>
            manhi <= conv_std_logic_vector(14843448,24);
            manlo <= conv_std_logic_vector(59807901,28);
           exponent <= '0';
      WHEN "1010001010" =>
            manhi <= conv_std_logic_vector(14874342,24);
            manlo <= conv_std_logic_vector(230995129,28);
           exponent <= '0';
      WHEN "1010001011" =>
            manhi <= conv_std_logic_vector(14905267,24);
            manlo <= conv_std_logic_vector(183482934,28);
           exponent <= '0';
      WHEN "1010001100" =>
            manhi <= conv_std_logic_vector(14936222,24);
            manlo <= conv_std_logic_vector(193623526,28);
           exponent <= '0';
      WHEN "1010001101" =>
            manhi <= conv_std_logic_vector(14967208,24);
            manlo <= conv_std_logic_vector(905939,28);
           exponent <= '0';
      WHEN "1010001110" =>
            manhi <= conv_std_logic_vector(14998223,24);
            manlo <= conv_std_logic_vector(150133320,28);
           exponent <= '0';
      WHEN "1010001111" =>
            manhi <= conv_std_logic_vector(15029269,24);
            manlo <= conv_std_logic_vector(112374738,28);
           exponent <= '0';
      WHEN "1010010000" =>
            manhi <= conv_std_logic_vector(15060345,24);
            manlo <= conv_std_logic_vector(164013390,28);
           exponent <= '0';
      WHEN "1010010001" =>
            manhi <= conv_std_logic_vector(15091452,24);
            manlo <= conv_std_logic_vector(44569327,28);
           exponent <= '0';
      WHEN "1010010010" =>
            manhi <= conv_std_logic_vector(15122589,24);
            manlo <= conv_std_logic_vector(30441282,28);
           exponent <= '0';
      WHEN "1010010011" =>
            manhi <= conv_std_logic_vector(15153756,24);
            manlo <= conv_std_logic_vector(129600316,28);
           exponent <= '0';
      WHEN "1010010100" =>
            manhi <= conv_std_logic_vector(15184954,24);
            manlo <= conv_std_logic_vector(81589818,28);
           exponent <= '0';
      WHEN "1010010101" =>
            manhi <= conv_std_logic_vector(15216182,24);
            manlo <= conv_std_logic_vector(162831889,28);
           exponent <= '0';
      WHEN "1010010110" =>
            manhi <= conv_std_logic_vector(15247441,24);
            manlo <= conv_std_logic_vector(112885518,28);
           exponent <= '0';
      WHEN "1010010111" =>
            manhi <= conv_std_logic_vector(15278730,24);
            manlo <= conv_std_logic_vector(208188418,28);
           exponent <= '0';
      WHEN "1010011000" =>
            manhi <= conv_std_logic_vector(15310050,24);
            manlo <= conv_std_logic_vector(188315209,28);
           exponent <= '0';
      WHEN "1010011001" =>
            manhi <= conv_std_logic_vector(15341401,24);
            manlo <= conv_std_logic_vector(61283792,28);
           exponent <= '0';
      WHEN "1010011010" =>
            manhi <= conv_std_logic_vector(15372782,24);
            manlo <= conv_std_logic_vector(103555359,28);
           exponent <= '0';
      WHEN "1010011011" =>
            manhi <= conv_std_logic_vector(15404194,24);
            manlo <= conv_std_logic_vector(54728032,28);
           exponent <= '0';
      WHEN "1010011100" =>
            manhi <= conv_std_logic_vector(15435636,24);
            manlo <= conv_std_logic_vector(191278690,28);
           exponent <= '0';
      WHEN "1010011101" =>
            manhi <= conv_std_logic_vector(15467109,24);
            manlo <= conv_std_logic_vector(252821163,28);
           exponent <= '0';
      WHEN "1010011110" =>
            manhi <= conv_std_logic_vector(15498613,24);
            manlo <= conv_std_logic_vector(247412597,28);
           exponent <= '0';
      WHEN "1010011111" =>
            manhi <= conv_std_logic_vector(15530148,24);
            manlo <= conv_std_logic_vector(183118012,28);
           exponent <= '0';
      WHEN "1010100000" =>
            manhi <= conv_std_logic_vector(15561714,24);
            manlo <= conv_std_logic_vector(68010306,28);
           exponent <= '0';
      WHEN "1010100001" =>
            manhi <= conv_std_logic_vector(15593310,24);
            manlo <= conv_std_logic_vector(178605723,28);
           exponent <= '0';
      WHEN "1010100010" =>
            manhi <= conv_std_logic_vector(15624937,24);
            manlo <= conv_std_logic_vector(254557489,28);
           exponent <= '0';
      WHEN "1010100011" =>
            manhi <= conv_std_logic_vector(15656596,24);
            manlo <= conv_std_logic_vector(35526733,28);
           exponent <= '0';
      WHEN "1010100100" =>
            manhi <= conv_std_logic_vector(15688285,24);
            manlo <= conv_std_logic_vector(66488863,28);
           exponent <= '0';
      WHEN "1010100101" =>
            manhi <= conv_std_logic_vector(15720005,24);
            manlo <= conv_std_logic_vector(87120837,28);
           exponent <= '0';
      WHEN "1010100110" =>
            manhi <= conv_std_logic_vector(15751756,24);
            manlo <= conv_std_logic_vector(105542995,28);
           exponent <= '0';
      WHEN "1010100111" =>
            manhi <= conv_std_logic_vector(15783538,24);
            manlo <= conv_std_logic_vector(129883612,28);
           exponent <= '0';
      WHEN "1010101000" =>
            manhi <= conv_std_logic_vector(15815351,24);
            manlo <= conv_std_logic_vector(168278902,28);
           exponent <= '0';
      WHEN "1010101001" =>
            manhi <= conv_std_logic_vector(15847195,24);
            manlo <= conv_std_logic_vector(228873033,28);
           exponent <= '0';
      WHEN "1010101010" =>
            manhi <= conv_std_logic_vector(15879071,24);
            manlo <= conv_std_logic_vector(51382669,28);
           exponent <= '0';
      WHEN "1010101011" =>
            manhi <= conv_std_logic_vector(15910977,24);
            manlo <= conv_std_logic_vector(180838811,28);
           exponent <= '0';
      WHEN "1010101100" =>
            manhi <= conv_std_logic_vector(15942915,24);
            manlo <= conv_std_logic_vector(88538606,28);
           exponent <= '0';
      WHEN "1010101101" =>
            manhi <= conv_std_logic_vector(15974884,24);
            manlo <= conv_std_logic_vector(51093552,28);
           exponent <= '0';
      WHEN "1010101110" =>
            manhi <= conv_std_logic_vector(16006884,24);
            manlo <= conv_std_logic_vector(76687676,28);
           exponent <= '0';
      WHEN "1010101111" =>
            manhi <= conv_std_logic_vector(16038915,24);
            manlo <= conv_std_logic_vector(173513005,28);
           exponent <= '0';
      WHEN "1010110000" =>
            manhi <= conv_std_logic_vector(16070978,24);
            manlo <= conv_std_logic_vector(81334110,28);
           exponent <= '0';
      WHEN "1010110001" =>
            manhi <= conv_std_logic_vector(16103072,24);
            manlo <= conv_std_logic_vector(76794490,28);
           exponent <= '0';
      WHEN "1010110010" =>
            manhi <= conv_std_logic_vector(16135197,24);
            manlo <= conv_std_logic_vector(168110204,28);
           exponent <= '0';
      WHEN "1010110011" =>
            manhi <= conv_std_logic_vector(16167354,24);
            manlo <= conv_std_logic_vector(95069884,28);
           exponent <= '0';
      WHEN "1010110100" =>
            manhi <= conv_std_logic_vector(16199542,24);
            manlo <= conv_std_logic_vector(134341108,28);
           exponent <= '0';
      WHEN "1010110101" =>
            manhi <= conv_std_logic_vector(16231762,24);
            manlo <= conv_std_logic_vector(25728588,28);
           exponent <= '0';
      WHEN "1010110110" =>
            manhi <= conv_std_logic_vector(16264013,24);
            manlo <= conv_std_logic_vector(45915996,28);
           exponent <= '0';
      WHEN "1010110111" =>
            manhi <= conv_std_logic_vector(16296295,24);
            manlo <= conv_std_logic_vector(203159607,28);
           exponent <= '0';
      WHEN "1010111000" =>
            manhi <= conv_std_logic_vector(16328609,24);
            manlo <= conv_std_logic_vector(237288310,28);
           exponent <= '0';
      WHEN "1010111001" =>
            manhi <= conv_std_logic_vector(16360955,24);
            manlo <= conv_std_logic_vector(156574520,28);
           exponent <= '0';
      WHEN "1010111010" =>
            manhi <= conv_std_logic_vector(16393332,24);
            manlo <= conv_std_logic_vector(237734194,28);
           exponent <= '0';
      WHEN "1010111011" =>
            manhi <= conv_std_logic_vector(16425741,24);
            manlo <= conv_std_logic_vector(220620465,28);
           exponent <= '0';
      WHEN "1010111100" =>
            manhi <= conv_std_logic_vector(16458182,24);
            manlo <= conv_std_logic_vector(113530022,28);
           exponent <= '0';
      WHEN "1010111101" =>
            manhi <= conv_std_logic_vector(16490654,24);
            manlo <= conv_std_logic_vector(193203116,28);
           exponent <= '0';
      WHEN "1010111110" =>
            manhi <= conv_std_logic_vector(16523158,24);
            manlo <= conv_std_logic_vector(199517199,28);
           exponent <= '0';
      WHEN "1010111111" =>
            manhi <= conv_std_logic_vector(16555694,24);
            manlo <= conv_std_logic_vector(140793302,28);
           exponent <= '0';
      WHEN "1011000000" =>
            manhi <= conv_std_logic_vector(16588262,24);
            manlo <= conv_std_logic_vector(25360585,28);
           exponent <= '0';
      WHEN "1011000001" =>
            manhi <= conv_std_logic_vector(16620861,24);
            manlo <= conv_std_logic_vector(129991803,28);
           exponent <= '0';
      WHEN "1011000010" =>
            manhi <= conv_std_logic_vector(16653492,24);
            manlo <= conv_std_logic_vector(194596944,28);
           exponent <= '0';
      WHEN "1011000011" =>
            manhi <= conv_std_logic_vector(16686155,24);
            manlo <= conv_std_logic_vector(227529607,28);
           exponent <= '0';
      WHEN "1011000100" =>
            manhi <= conv_std_logic_vector(16718850,24);
            manlo <= conv_std_logic_vector(237151552,28);
           exponent <= '0';
      WHEN "1011000101" =>
            manhi <= conv_std_logic_vector(16751577,24);
            manlo <= conv_std_logic_vector(231832709,28);
           exponent <= '0';
      WHEN "1011000110" =>
            manhi <= conv_std_logic_vector(3560,24);
            manlo <= conv_std_logic_vector(109975592,28);
           exponent <= '1';
      WHEN "1011000111" =>
            manhi <= conv_std_logic_vector(19955,24);
            manlo <= conv_std_logic_vector(239164365,28);
           exponent <= '1';
      WHEN "1011001000" =>
            manhi <= conv_std_logic_vector(36367,24);
            manlo <= conv_std_logic_vector(105026731,28);
           exponent <= '1';
      WHEN "1011001001" =>
            manhi <= conv_std_logic_vector(52794,24);
            manlo <= conv_std_logic_vector(248634947,28);
           exponent <= '1';
      WHEN "1011001010" =>
            manhi <= conv_std_logic_vector(69238,24);
            manlo <= conv_std_logic_vector(137323551,28);
           exponent <= '1';
      WHEN "1011001011" =>
            manhi <= conv_std_logic_vector(85698,24);
            manlo <= conv_std_logic_vector(43737556,28);
           exponent <= '1';
      WHEN "1011001100" =>
            manhi <= conv_std_logic_vector(102173,24);
            manlo <= conv_std_logic_vector(240526091,28);
           exponent <= '1';
      WHEN "1011001101" =>
            manhi <= conv_std_logic_vector(118665,24);
            manlo <= conv_std_logic_vector(195036030,28);
           exponent <= '1';
      WHEN "1011001110" =>
            manhi <= conv_std_logic_vector(135173,24);
            manlo <= conv_std_logic_vector(179924739,28);
           exponent <= '1';
      WHEN "1011001111" =>
            manhi <= conv_std_logic_vector(151697,24);
            manlo <= conv_std_logic_vector(199418251,28);
           exponent <= '1';
      WHEN "1011010000" =>
            manhi <= conv_std_logic_vector(168237,24);
            manlo <= conv_std_logic_vector(257746730,28);
           exponent <= '1';
      WHEN "1011010001" =>
            manhi <= conv_std_logic_vector(184794,24);
            manlo <= conv_std_logic_vector(90709016,28);
           exponent <= '1';
      WHEN "1011010010" =>
            manhi <= conv_std_logic_vector(201366,24);
            manlo <= conv_std_logic_vector(239414453,28);
           exponent <= '1';
      WHEN "1011010011" =>
            manhi <= conv_std_logic_vector(217955,24);
            manlo <= conv_std_logic_vector(171234704,28);
           exponent <= '1';
      WHEN "1011010100" =>
            manhi <= conv_std_logic_vector(234560,24);
            manlo <= conv_std_logic_vector(158851944,28);
           exponent <= '1';
      WHEN "1011010101" =>
            manhi <= conv_std_logic_vector(251181,24);
            manlo <= conv_std_logic_vector(206517042,28);
           exponent <= '1';
      WHEN "1011010110" =>
            manhi <= conv_std_logic_vector(267819,24);
            manlo <= conv_std_logic_vector(50049563,28);
           exponent <= '1';
      WHEN "1011010111" =>
            manhi <= conv_std_logic_vector(284472,24);
            manlo <= conv_std_logic_vector(230579599,28);
           exponent <= '1';
      WHEN "1011011000" =>
            manhi <= conv_std_logic_vector(301142,24);
            manlo <= conv_std_logic_vector(215499577,28);
           exponent <= '1';
      WHEN "1011011001" =>
            manhi <= conv_std_logic_vector(317829,24);
            manlo <= conv_std_logic_vector(9077005,28);
           exponent <= '1';
      WHEN "1011011010" =>
            manhi <= conv_std_logic_vector(334531,24);
            manlo <= conv_std_logic_vector(152454469,28);
           exponent <= '1';
      WHEN "1011011011" =>
            manhi <= conv_std_logic_vector(351250,24);
            manlo <= conv_std_logic_vector(113036907,28);
           exponent <= '1';
      WHEN "1011011100" =>
            manhi <= conv_std_logic_vector(367985,24);
            manlo <= conv_std_logic_vector(163539801,28);
           exponent <= '1';
      WHEN "1011011101" =>
            manhi <= conv_std_logic_vector(384737,24);
            manlo <= conv_std_logic_vector(39811903,28);
           exponent <= '1';
      WHEN "1011011110" =>
            manhi <= conv_std_logic_vector(401505,24);
            manlo <= conv_std_logic_vector(14577065,28);
           exponent <= '1';
      WHEN "1011011111" =>
            manhi <= conv_std_logic_vector(418289,24);
            manlo <= conv_std_logic_vector(92127870,28);
           exponent <= '1';
      WHEN "1011100000" =>
            manhi <= conv_std_logic_vector(435090,24);
            manlo <= conv_std_logic_vector(8325641,28);
           exponent <= '1';
      WHEN "1011100001" =>
            manhi <= conv_std_logic_vector(451907,24);
            manlo <= conv_std_logic_vector(35906810,28);
           exponent <= '1';
      WHEN "1011100010" =>
            manhi <= conv_std_logic_vector(468740,24);
            manlo <= conv_std_logic_vector(179176556,28);
           exponent <= '1';
      WHEN "1011100011" =>
            manhi <= conv_std_logic_vector(485590,24);
            manlo <= conv_std_logic_vector(174008808,28);
           exponent <= '1';
      WHEN "1011100100" =>
            manhi <= conv_std_logic_vector(502457,24);
            manlo <= conv_std_logic_vector(24717160,28);
           exponent <= '1';
      WHEN "1011100101" =>
            manhi <= conv_std_logic_vector(519340,24);
            manlo <= conv_std_logic_vector(4054880,28);
           exponent <= '1';
      WHEN "1011100110" =>
            manhi <= conv_std_logic_vector(536239,24);
            manlo <= conv_std_logic_vector(116343996,28);
           exponent <= '1';
      WHEN "1011100111" =>
            manhi <= conv_std_logic_vector(553155,24);
            manlo <= conv_std_logic_vector(97475302,28);
           exponent <= '1';
      WHEN "1011101000" =>
            manhi <= conv_std_logic_vector(570087,24);
            manlo <= conv_std_logic_vector(220214735,28);
           exponent <= '1';
      WHEN "1011101001" =>
            manhi <= conv_std_logic_vector(587036,24);
            manlo <= conv_std_logic_vector(220461546,28);
           exponent <= '1';
      WHEN "1011101010" =>
            manhi <= conv_std_logic_vector(604002,24);
            manlo <= conv_std_logic_vector(102554681,28);
           exponent <= '1';
      WHEN "1011101011" =>
            manhi <= conv_std_logic_vector(620984,24);
            manlo <= conv_std_logic_vector(139272779,28);
           exponent <= '1';
      WHEN "1011101100" =>
            manhi <= conv_std_logic_vector(637983,24);
            manlo <= conv_std_logic_vector(66527812,28);
           exponent <= '1';
      WHEN "1011101101" =>
            manhi <= conv_std_logic_vector(654998,24);
            manlo <= conv_std_logic_vector(157106911,28);
           exponent <= '1';
      WHEN "1011101110" =>
            manhi <= conv_std_logic_vector(672030,24);
            manlo <= conv_std_logic_vector(146930546,28);
           exponent <= '1';
      WHEN "1011101111" =>
            manhi <= conv_std_logic_vector(689079,24);
            manlo <= conv_std_logic_vector(40358901,28);
           exponent <= '1';
      WHEN "1011110000" =>
            manhi <= conv_std_logic_vector(706144,24);
            manlo <= conv_std_logic_vector(110191873,28);
           exponent <= '1';
      WHEN "1011110001" =>
            manhi <= conv_std_logic_vector(723226,24);
            manlo <= conv_std_logic_vector(92362714,28);
           exponent <= '1';
      WHEN "1011110010" =>
            manhi <= conv_std_logic_vector(740324,24);
            manlo <= conv_std_logic_vector(259679855,28);
           exponent <= '1';
      WHEN "1011110011" =>
            manhi <= conv_std_logic_vector(757440,24);
            manlo <= conv_std_logic_vector(79649632,28);
           exponent <= '1';
      WHEN "1011110100" =>
            manhi <= conv_std_logic_vector(774572,24);
            manlo <= conv_std_logic_vector(93524482,28);
           exponent <= '1';
      WHEN "1011110101" =>
            manhi <= conv_std_logic_vector(791721,24);
            manlo <= conv_std_logic_vector(37254754,28);
           exponent <= '1';
      WHEN "1011110110" =>
            manhi <= conv_std_logic_vector(808886,24);
            manlo <= conv_std_logic_vector(183665996,28);
           exponent <= '1';
      WHEN "1011110111" =>
            manhi <= conv_std_logic_vector(826069,24);
            manlo <= conv_std_logic_vector(281674,28);
           exponent <= '1';
      WHEN "1011111000" =>
            manhi <= conv_std_logic_vector(843268,24);
            manlo <= conv_std_logic_vector(28371374,28);
           exponent <= '1';
      WHEN "1011111001" =>
            manhi <= conv_std_logic_vector(860484,24);
            manlo <= conv_std_logic_vector(3902612,28);
           exponent <= '1';
      WHEN "1011111010" =>
            manhi <= conv_std_logic_vector(877716,24);
            manlo <= conv_std_logic_vector(199718117,28);
           exponent <= '1';
      WHEN "1011111011" =>
            manhi <= conv_std_logic_vector(894966,24);
            manlo <= conv_std_logic_vector(83358555,28);
           exponent <= '1';
      WHEN "1011111100" =>
            manhi <= conv_std_logic_vector(912232,24);
            manlo <= conv_std_logic_vector(196110728,28);
           exponent <= '1';
      WHEN "1011111101" =>
            manhi <= conv_std_logic_vector(929516,24);
            manlo <= conv_std_logic_vector(5523929,28);
           exponent <= '1';
      WHEN "1011111110" =>
            manhi <= conv_std_logic_vector(946816,24);
            manlo <= conv_std_logic_vector(52893590,28);
           exponent <= '1';
      WHEN "1011111111" =>
            manhi <= conv_std_logic_vector(964133,24);
            manlo <= conv_std_logic_vector(74213103,28);
           exponent <= '1';
      WHEN "1100000000" =>
            manhi <= conv_std_logic_vector(981467,24);
            manlo <= conv_std_logic_vector(73915640,28);
           exponent <= '1';
      WHEN "1100000001" =>
            manhi <= conv_std_logic_vector(998818,24);
            manlo <= conv_std_logic_vector(56438704,28);
           exponent <= '1';
      WHEN "1100000010" =>
            manhi <= conv_std_logic_vector(1016186,24);
            manlo <= conv_std_logic_vector(26224136,28);
           exponent <= '1';
      WHEN "1100000011" =>
            manhi <= conv_std_logic_vector(1033570,24);
            manlo <= conv_std_logic_vector(256153571,28);
           exponent <= '1';
      WHEN "1100000100" =>
            manhi <= conv_std_logic_vector(1050972,24);
            manlo <= conv_std_logic_vector(213806620,28);
           exponent <= '1';
      WHEN "1100000101" =>
            manhi <= conv_std_logic_vector(1068391,24);
            manlo <= conv_std_logic_vector(172073612,28);
           exponent <= '1';
      WHEN "1100000110" =>
            manhi <= conv_std_logic_vector(1085827,24);
            manlo <= conv_std_logic_vector(135413771,28);
           exponent <= '1';
      WHEN "1100000111" =>
            manhi <= conv_std_logic_vector(1103280,24);
            manlo <= conv_std_logic_vector(108290679,28);
           exponent <= '1';
      WHEN "1100001000" =>
            manhi <= conv_std_logic_vector(1120750,24);
            manlo <= conv_std_logic_vector(95172278,28);
           exponent <= '1';
      WHEN "1100001001" =>
            manhi <= conv_std_logic_vector(1138237,24);
            manlo <= conv_std_logic_vector(100530876,28);
           exponent <= '1';
      WHEN "1100001010" =>
            manhi <= conv_std_logic_vector(1155741,24);
            manlo <= conv_std_logic_vector(128843150,28);
           exponent <= '1';
      WHEN "1100001011" =>
            manhi <= conv_std_logic_vector(1173262,24);
            manlo <= conv_std_logic_vector(184590152,28);
           exponent <= '1';
      WHEN "1100001100" =>
            manhi <= conv_std_logic_vector(1190801,24);
            manlo <= conv_std_logic_vector(3821855,28);
           exponent <= '1';
      WHEN "1100001101" =>
            manhi <= conv_std_logic_vector(1208356,24);
            manlo <= conv_std_logic_vector(127898983,28);
           exponent <= '1';
      WHEN "1100001110" =>
            manhi <= conv_std_logic_vector(1225929,24);
            manlo <= conv_std_logic_vector(24444823,28);
           exponent <= '1';
      WHEN "1100001111" =>
            manhi <= conv_std_logic_vector(1243518,24);
            manlo <= conv_std_logic_vector(234828877,28);
           exponent <= '1';
      WHEN "1100010000" =>
            manhi <= conv_std_logic_vector(1261125,24);
            manlo <= conv_std_logic_vector(226683218,28);
           exponent <= '1';
      WHEN "1100010001" =>
            manhi <= conv_std_logic_vector(1278750,24);
            manlo <= conv_std_logic_vector(4515229,28);
           exponent <= '1';
      WHEN "1100010010" =>
            manhi <= conv_std_logic_vector(1296391,24);
            manlo <= conv_std_logic_vector(109707612,28);
           exponent <= '1';
      WHEN "1100010011" =>
            manhi <= conv_std_logic_vector(1314050,24);
            manlo <= conv_std_logic_vector(9905652,28);
           exponent <= '1';
      WHEN "1100010100" =>
            manhi <= conv_std_logic_vector(1331725,24);
            manlo <= conv_std_logic_vector(246500869,28);
           exponent <= '1';
      WHEN "1100010101" =>
            manhi <= conv_std_logic_vector(1349419,24);
            manlo <= conv_std_logic_vector(18711921,28);
           exponent <= '1';
      WHEN "1100010110" =>
            manhi <= conv_std_logic_vector(1367129,24);
            manlo <= conv_std_logic_vector(136374624,28);
           exponent <= '1';
      WHEN "1100010111" =>
            manhi <= conv_std_logic_vector(1384857,24);
            manlo <= conv_std_logic_vector(67151939,28);
           exponent <= '1';
      WHEN "1100011000" =>
            manhi <= conv_std_logic_vector(1402602,24);
            manlo <= conv_std_logic_vector(84017623,28);
           exponent <= '1';
      WHEN "1100011001" =>
            manhi <= conv_std_logic_vector(1420364,24);
            manlo <= conv_std_logic_vector(191514413,28);
           exponent <= '1';
      WHEN "1100011010" =>
            manhi <= conv_std_logic_vector(1438144,24);
            manlo <= conv_std_logic_vector(125754028,28);
           exponent <= '1';
      WHEN "1100011011" =>
            manhi <= conv_std_logic_vector(1455941,24);
            manlo <= conv_std_logic_vector(159723541,28);
           exponent <= '1';
      WHEN "1100011100" =>
            manhi <= conv_std_logic_vector(1473756,24);
            manlo <= conv_std_logic_vector(29543561,28);
           exponent <= '1';
      WHEN "1100011101" =>
            manhi <= conv_std_logic_vector(1491588,24);
            manlo <= conv_std_logic_vector(8210062,28);
           exponent <= '1';
      WHEN "1100011110" =>
            manhi <= conv_std_logic_vector(1509437,24);
            manlo <= conv_std_logic_vector(100288013,28);
           exponent <= '1';
      WHEN "1100011111" =>
            manhi <= conv_std_logic_vector(1527304,24);
            manlo <= conv_std_logic_vector(41911392,28);
           exponent <= '1';
      WHEN "1100100000" =>
            manhi <= conv_std_logic_vector(1545188,24);
            manlo <= conv_std_logic_vector(106089552,28);
           exponent <= '1';
      WHEN "1100100001" =>
            manhi <= conv_std_logic_vector(1563090,24);
            manlo <= conv_std_logic_vector(28965402,28);
           exponent <= '1';
      WHEN "1100100010" =>
            manhi <= conv_std_logic_vector(1581009,24);
            manlo <= conv_std_logic_vector(83557236,28);
           exponent <= '1';
      WHEN "1100100011" =>
            manhi <= conv_std_logic_vector(1598946,24);
            manlo <= conv_std_logic_vector(6016916,28);
           exponent <= '1';
      WHEN "1100100100" =>
            manhi <= conv_std_logic_vector(1616900,24);
            manlo <= conv_std_logic_vector(69371695,28);
           exponent <= '1';
      WHEN "1100100101" =>
            manhi <= conv_std_logic_vector(1634872,24);
            manlo <= conv_std_logic_vector(9782402,28);
           exponent <= '1';
      WHEN "1100100110" =>
            manhi <= conv_std_logic_vector(1652861,24);
            manlo <= conv_std_logic_vector(100285270,28);
           exponent <= '1';
      WHEN "1100100111" =>
            manhi <= conv_std_logic_vector(1670868,24);
            manlo <= conv_std_logic_vector(77050112,28);
           exponent <= '1';
      WHEN "1100101000" =>
            manhi <= conv_std_logic_vector(1688892,24);
            manlo <= conv_std_logic_vector(213122155,28);
           exponent <= '1';
      WHEN "1100101001" =>
            manhi <= conv_std_logic_vector(1706934,24);
            manlo <= conv_std_logic_vector(244680216,28);
           exponent <= '1';
      WHEN "1100101010" =>
            manhi <= conv_std_logic_vector(1724994,24);
            manlo <= conv_std_logic_vector(176343080,28);
           exponent <= '1';
      WHEN "1100101011" =>
            manhi <= conv_std_logic_vector(1743072,24);
            manlo <= conv_std_logic_vector(12734040,28);
           exponent <= '1';
      WHEN "1100101100" =>
            manhi <= conv_std_logic_vector(1761167,24);
            manlo <= conv_std_logic_vector(26916364,28);
           exponent <= '1';
      WHEN "1100101101" =>
            manhi <= conv_std_logic_vector(1779279,24);
            manlo <= conv_std_logic_vector(223522388,28);
           exponent <= '1';
      WHEN "1100101110" =>
            manhi <= conv_std_logic_vector(1797410,24);
            manlo <= conv_std_logic_vector(70318058,28);
           exponent <= '1';
      WHEN "1100101111" =>
            manhi <= conv_std_logic_vector(1815558,24);
            manlo <= conv_std_logic_vector(108815677,28);
           exponent <= '1';
      WHEN "1100110000" =>
            manhi <= conv_std_logic_vector(1833724,24);
            manlo <= conv_std_logic_vector(75225715,28);
           exponent <= '1';
      WHEN "1100110001" =>
            manhi <= conv_std_logic_vector(1851907,24);
            manlo <= conv_std_logic_vector(242634090,28);
           exponent <= '1';
      WHEN "1100110010" =>
            manhi <= conv_std_logic_vector(1870109,24);
            manlo <= conv_std_logic_vector(78824900,28);
           exponent <= '1';
      WHEN "1100110011" =>
            manhi <= conv_std_logic_vector(1888328,24);
            manlo <= conv_std_logic_vector(125328613,28);
           exponent <= '1';
      WHEN "1100110100" =>
            manhi <= conv_std_logic_vector(1906565,24);
            manlo <= conv_std_logic_vector(118373881,28);
           exponent <= '1';
      WHEN "1100110101" =>
            manhi <= conv_std_logic_vector(1924820,24);
            manlo <= conv_std_logic_vector(62629370,28);
           exponent <= '1';
      WHEN "1100110110" =>
            manhi <= conv_std_logic_vector(1943092,24);
            manlo <= conv_std_logic_vector(231203763,28);
           exponent <= '1';
      WHEN "1100110111" =>
            manhi <= conv_std_logic_vector(1961383,24);
            manlo <= conv_std_logic_vector(91903942,28);
           exponent <= '1';
      WHEN "1100111000" =>
            manhi <= conv_std_logic_vector(1979691,24);
            manlo <= conv_std_logic_vector(186283181,28);
           exponent <= '1';
      WHEN "1100111001" =>
            manhi <= conv_std_logic_vector(1998017,24);
            manlo <= conv_std_logic_vector(250592964,28);
           exponent <= '1';
      WHEN "1100111010" =>
            manhi <= conv_std_logic_vector(2016362,24);
            manlo <= conv_std_logic_vector(21089351,28);
           exponent <= '1';
      WHEN "1100111011" =>
            manhi <= conv_std_logic_vector(2034724,24);
            manlo <= conv_std_logic_vector(39339357,28);
           exponent <= '1';
      WHEN "1100111100" =>
            manhi <= conv_std_logic_vector(2053104,24);
            manlo <= conv_std_logic_vector(41608216,28);
           exponent <= '1';
      WHEN "1100111101" =>
            manhi <= conv_std_logic_vector(2071502,24);
            manlo <= conv_std_logic_vector(32601209,28);
           exponent <= '1';
      WHEN "1100111110" =>
            manhi <= conv_std_logic_vector(2089918,24);
            manlo <= conv_std_logic_vector(17028217,28);
           exponent <= '1';
      WHEN "1100111111" =>
            manhi <= conv_std_logic_vector(2108351,24);
            manlo <= conv_std_logic_vector(268039176,28);
           exponent <= '1';
      WHEN "1101000000" =>
            manhi <= conv_std_logic_vector(2126803,24);
            manlo <= conv_std_logic_vector(253482264,28);
           exponent <= '1';
      WHEN "1101000001" =>
            manhi <= conv_std_logic_vector(2145273,24);
            manlo <= conv_std_logic_vector(246516634,28);
           exponent <= '1';
      WHEN "1101000010" =>
            manhi <= conv_std_logic_vector(2163761,24);
            manlo <= conv_std_logic_vector(251870600,28);
           exponent <= '1';
      WHEN "1101000011" =>
            manhi <= conv_std_logic_vector(2182268,24);
            manlo <= conv_std_logic_vector(5841640,28);
           exponent <= '1';
      WHEN "1101000100" =>
            manhi <= conv_std_logic_vector(2200792,24);
            manlo <= conv_std_logic_vector(50038222,28);
           exponent <= '1';
      WHEN "1101000101" =>
            manhi <= conv_std_logic_vector(2219334,24);
            manlo <= conv_std_logic_vector(120767079,28);
           exponent <= '1';
      WHEN "1101000110" =>
            manhi <= conv_std_logic_vector(2237894,24);
            manlo <= conv_std_logic_vector(222775030,28);
           exponent <= '1';
      WHEN "1101000111" =>
            manhi <= conv_std_logic_vector(2256473,24);
            manlo <= conv_std_logic_vector(92378075,28);
           exponent <= '1';
      WHEN "1101001000" =>
            manhi <= conv_std_logic_vector(2275070,24);
            manlo <= conv_std_logic_vector(2767772,28);
           exponent <= '1';
      WHEN "1101001001" =>
            manhi <= conv_std_logic_vector(2293684,24);
            manlo <= conv_std_logic_vector(227140324,28);
           exponent <= '1';
      WHEN "1101001010" =>
            manhi <= conv_std_logic_vector(2312317,24);
            manlo <= conv_std_logic_vector(233390216,28);
           exponent <= '1';
      WHEN "1101001011" =>
            manhi <= conv_std_logic_vector(2330969,24);
            manlo <= conv_std_logic_vector(26287503,28);
           exponent <= '1';
      WHEN "1101001100" =>
            manhi <= conv_std_logic_vector(2349638,24);
            manlo <= conv_std_logic_vector(147477811,28);
           exponent <= '1';
      WHEN "1101001101" =>
            manhi <= conv_std_logic_vector(2368326,24);
            manlo <= conv_std_logic_vector(64869610,28);
           exponent <= '1';
      WHEN "1101001110" =>
            manhi <= conv_std_logic_vector(2387032,24);
            manlo <= conv_std_logic_vector(51682404,28);
           exponent <= '1';
      WHEN "1101001111" =>
            manhi <= conv_std_logic_vector(2405756,24);
            manlo <= conv_std_logic_vector(112704917,28);
           exponent <= '1';
      WHEN "1101010000" =>
            manhi <= conv_std_logic_vector(2424498,24);
            manlo <= conv_std_logic_vector(252730552,28);
           exponent <= '1';
      WHEN "1101010001" =>
            manhi <= conv_std_logic_vector(2443259,24);
            manlo <= conv_std_logic_vector(208121938,28);
           exponent <= '1';
      WHEN "1101010010" =>
            manhi <= conv_std_logic_vector(2462038,24);
            manlo <= conv_std_logic_vector(252117306,28);
           exponent <= '1';
      WHEN "1101010011" =>
            manhi <= conv_std_logic_vector(2480836,24);
            manlo <= conv_std_logic_vector(121088666,28);
           exponent <= '1';
      WHEN "1101010100" =>
            manhi <= conv_std_logic_vector(2499652,24);
            manlo <= conv_std_logic_vector(88283637,28);
           exponent <= '1';
      WHEN "1101010101" =>
            manhi <= conv_std_logic_vector(2518486,24);
            manlo <= conv_std_logic_vector(158519085,28);
           exponent <= '1';
      WHEN "1101010110" =>
            manhi <= conv_std_logic_vector(2537339,24);
            manlo <= conv_std_logic_vector(68181124,28);
           exponent <= '1';
      WHEN "1101010111" =>
            manhi <= conv_std_logic_vector(2556210,24);
            manlo <= conv_std_logic_vector(90531494,28);
           exponent <= '1';
      WHEN "1101011000" =>
            manhi <= conv_std_logic_vector(2575099,24);
            manlo <= conv_std_logic_vector(230401190,28);
           exponent <= '1';
      WHEN "1101011001" =>
            manhi <= conv_std_logic_vector(2594007,24);
            manlo <= conv_std_logic_vector(224190477,28);
           exponent <= '1';
      WHEN "1101011010" =>
            manhi <= conv_std_logic_vector(2612934,24);
            manlo <= conv_std_logic_vector(76739795,28);
           exponent <= '1';
      WHEN "1101011011" =>
            manhi <= conv_std_logic_vector(2631879,24);
            manlo <= conv_std_logic_vector(61329773,28);
           exponent <= '1';
      WHEN "1101011100" =>
            manhi <= conv_std_logic_vector(2650842,24);
            manlo <= conv_std_logic_vector(182810317,28);
           exponent <= '1';
      WHEN "1101011101" =>
            manhi <= conv_std_logic_vector(2669824,24);
            manlo <= conv_std_logic_vector(177600614,28);
           exponent <= '1';
      WHEN "1101011110" =>
            manhi <= conv_std_logic_vector(2688825,24);
            manlo <= conv_std_logic_vector(50560052,28);
           exponent <= '1';
      WHEN "1101011111" =>
            manhi <= conv_std_logic_vector(2707844,24);
            manlo <= conv_std_logic_vector(74988222,28);
           exponent <= '1';
      WHEN "1101100000" =>
            manhi <= conv_std_logic_vector(2726881,24);
            manlo <= conv_std_logic_vector(255754012,28);
           exponent <= '1';
      WHEN "1101100001" =>
            manhi <= conv_std_logic_vector(2745938,24);
            manlo <= conv_std_logic_vector(60860155,28);
           exponent <= '1';
      WHEN "1101100010" =>
            manhi <= conv_std_logic_vector(2765013,24);
            manlo <= conv_std_logic_vector(32055969,28);
           exponent <= '1';
      WHEN "1101100011" =>
            manhi <= conv_std_logic_vector(2784106,24);
            manlo <= conv_std_logic_vector(174224628,28);
           exponent <= '1';
      WHEN "1101100100" =>
            manhi <= conv_std_logic_vector(2803218,24);
            manlo <= conv_std_logic_vector(223818618,28);
           exponent <= '1';
      WHEN "1101100101" =>
            manhi <= conv_std_logic_vector(2822349,24);
            manlo <= conv_std_logic_vector(185730660,28);
           exponent <= '1';
      WHEN "1101100110" =>
            manhi <= conv_std_logic_vector(2841499,24);
            manlo <= conv_std_logic_vector(64858254,28);
           exponent <= '1';
      WHEN "1101100111" =>
            manhi <= conv_std_logic_vector(2860667,24);
            manlo <= conv_std_logic_vector(134539142,28);
           exponent <= '1';
      WHEN "1101101000" =>
            manhi <= conv_std_logic_vector(2879854,24);
            manlo <= conv_std_logic_vector(131244940,28);
           exponent <= '1';
      WHEN "1101101001" =>
            manhi <= conv_std_logic_vector(2899060,24);
            manlo <= conv_std_logic_vector(59887520,28);
           exponent <= '1';
      WHEN "1101101010" =>
            manhi <= conv_std_logic_vector(2918284,24);
            manlo <= conv_std_logic_vector(193819006,28);
           exponent <= '1';
      WHEN "1101101011" =>
            manhi <= conv_std_logic_vector(2937528,24);
            manlo <= conv_std_logic_vector(1089957,28);
           exponent <= '1';
      WHEN "1101101100" =>
            manhi <= conv_std_logic_vector(2956790,24);
            manlo <= conv_std_logic_vector(23497566,28);
           exponent <= '1';
      WHEN "1101101101" =>
            manhi <= conv_std_logic_vector(2976070,24);
            manlo <= conv_std_logic_vector(265972927,28);
           exponent <= '1';
      WHEN "1101101110" =>
            manhi <= conv_std_logic_vector(2995370,24);
            manlo <= conv_std_logic_vector(196581040,28);
           exponent <= '1';
      WHEN "1101101111" =>
            manhi <= conv_std_logic_vector(3014689,24);
            manlo <= conv_std_logic_vector(88698094,28);
           exponent <= '1';
      WHEN "1101110000" =>
            manhi <= conv_std_logic_vector(3034026,24);
            manlo <= conv_std_logic_vector(215705108,28);
           exponent <= '1';
      WHEN "1101110001" =>
            manhi <= conv_std_logic_vector(3053383,24);
            manlo <= conv_std_logic_vector(45681562,28);
           exponent <= '1';
      WHEN "1101110010" =>
            manhi <= conv_std_logic_vector(3072758,24);
            manlo <= conv_std_logic_vector(120453600,28);
           exponent <= '1';
      WHEN "1101110011" =>
            manhi <= conv_std_logic_vector(3092152,24);
            manlo <= conv_std_logic_vector(176545836,28);
           exponent <= '1';
      WHEN "1101110100" =>
            manhi <= conv_std_logic_vector(3111565,24);
            manlo <= conv_std_logic_vector(218923189,28);
           exponent <= '1';
      WHEN "1101110101" =>
            manhi <= conv_std_logic_vector(3130997,24);
            manlo <= conv_std_logic_vector(252555427,28);
           exponent <= '1';
      WHEN "1101110110" =>
            manhi <= conv_std_logic_vector(3150449,24);
            manlo <= conv_std_logic_vector(13981719,28);
           exponent <= '1';
      WHEN "1101110111" =>
            manhi <= conv_std_logic_vector(3169919,24);
            manlo <= conv_std_logic_vector(45052462,28);
           exponent <= '1';
      WHEN "1101111000" =>
            manhi <= conv_std_logic_vector(3189408,24);
            manlo <= conv_std_logic_vector(82316549,28);
           exponent <= '1';
      WHEN "1101111001" =>
            manhi <= conv_std_logic_vector(3208916,24);
            manlo <= conv_std_logic_vector(130763202,28);
           exponent <= '1';
      WHEN "1101111010" =>
            manhi <= conv_std_logic_vector(3228443,24);
            manlo <= conv_std_logic_vector(195386513,28);
           exponent <= '1';
      WHEN "1101111011" =>
            manhi <= conv_std_logic_vector(3247990,24);
            manlo <= conv_std_logic_vector(12750002,28);
           exponent <= '1';
      WHEN "1101111100" =>
            manhi <= conv_std_logic_vector(3267555,24);
            manlo <= conv_std_logic_vector(124728439,28);
           exponent <= '1';
      WHEN "1101111101" =>
            manhi <= conv_std_logic_vector(3287139,24);
            manlo <= conv_std_logic_vector(267895114,28);
           exponent <= '1';
      WHEN "1101111110" =>
            manhi <= conv_std_logic_vector(3306743,24);
            manlo <= conv_std_logic_vector(178828213,28);
           exponent <= '1';
      WHEN "1101111111" =>
            manhi <= conv_std_logic_vector(3326366,24);
            manlo <= conv_std_logic_vector(130981732,28);
           exponent <= '1';
      WHEN "1110000000" =>
            manhi <= conv_std_logic_vector(3346008,24);
            manlo <= conv_std_logic_vector(129379112,28);
           exponent <= '1';
      WHEN "1110000001" =>
            manhi <= conv_std_logic_vector(3365669,24);
            manlo <= conv_std_logic_vector(179048704,28);
           exponent <= '1';
      WHEN "1110000010" =>
            manhi <= conv_std_logic_vector(3385350,24);
            manlo <= conv_std_logic_vector(16588318,28);
           exponent <= '1';
      WHEN "1110000011" =>
            manhi <= conv_std_logic_vector(3405049,24);
            manlo <= conv_std_logic_vector(183907046,28);
           exponent <= '1';
      WHEN "1110000100" =>
            manhi <= conv_std_logic_vector(3424768,24);
            manlo <= conv_std_logic_vector(149177079,28);
           exponent <= '1';
      WHEN "1110000101" =>
            manhi <= conv_std_logic_vector(3444506,24);
            manlo <= conv_std_logic_vector(185881906,28);
           exponent <= '1';
      WHEN "1110000110" =>
            manhi <= conv_std_logic_vector(3464264,24);
            manlo <= conv_std_logic_vector(30639033,28);
           exponent <= '1';
      WHEN "1110000111" =>
            manhi <= conv_std_logic_vector(3484040,24);
            manlo <= conv_std_logic_vector(225377274,28);
           exponent <= '1';
      WHEN "1110001000" =>
            manhi <= conv_std_logic_vector(3503836,24);
            manlo <= conv_std_logic_vector(238288557,28);
           exponent <= '1';
      WHEN "1110001001" =>
            manhi <= conv_std_logic_vector(3523652,24);
            manlo <= conv_std_logic_vector(74440673,28);
           exponent <= '1';
      WHEN "1110001010" =>
            manhi <= conv_std_logic_vector(3543487,24);
            manlo <= conv_std_logic_vector(7341816,28);
           exponent <= '1';
      WHEN "1110001011" =>
            manhi <= conv_std_logic_vector(3563341,24);
            manlo <= conv_std_logic_vector(42069684,28);
           exponent <= '1';
      WHEN "1110001100" =>
            manhi <= conv_std_logic_vector(3583214,24);
            manlo <= conv_std_logic_vector(183706934,28);
           exponent <= '1';
      WHEN "1110001101" =>
            manhi <= conv_std_logic_vector(3603107,24);
            manlo <= conv_std_logic_vector(168905734,28);
           exponent <= '1';
      WHEN "1110001110" =>
            manhi <= conv_std_logic_vector(3623020,24);
            manlo <= conv_std_logic_vector(2758677,28);
           exponent <= '1';
      WHEN "1110001111" =>
            manhi <= conv_std_logic_vector(3642951,24);
            manlo <= conv_std_logic_vector(227234245,28);
           exponent <= '1';
      WHEN "1110010000" =>
            manhi <= conv_std_logic_vector(3662903,24);
            manlo <= conv_std_logic_vector(42128622,28);
           exponent <= '1';
      WHEN "1110010001" =>
            manhi <= conv_std_logic_vector(3682873,24);
            manlo <= conv_std_logic_vector(257855711,28);
           exponent <= '1';
      WHEN "1110010010" =>
            manhi <= conv_std_logic_vector(3702864,24);
            manlo <= conv_std_logic_vector(74221670,28);
           exponent <= '1';
      WHEN "1110010011" =>
            manhi <= conv_std_logic_vector(3722874,24);
            manlo <= conv_std_logic_vector(33214933,28);
           exponent <= '1';
      WHEN "1110010100" =>
            manhi <= conv_std_logic_vector(3742903,24);
            manlo <= conv_std_logic_vector(139958020,28);
           exponent <= '1';
      WHEN "1110010101" =>
            manhi <= conv_std_logic_vector(3762952,24);
            manlo <= conv_std_logic_vector(131143002,28);
           exponent <= '1';
      WHEN "1110010110" =>
            manhi <= conv_std_logic_vector(3783021,24);
            manlo <= conv_std_logic_vector(11902416,28);
           exponent <= '1';
      WHEN "1110010111" =>
            manhi <= conv_std_logic_vector(3803109,24);
            manlo <= conv_std_logic_vector(55809266,28);
           exponent <= '1';
      WHEN "1110011000" =>
            manhi <= conv_std_logic_vector(3823216,24);
            manlo <= conv_std_logic_vector(268006125,28);
           exponent <= '1';
      WHEN "1110011001" =>
            manhi <= conv_std_logic_vector(3843344,24);
            manlo <= conv_std_logic_vector(116769675,28);
           exponent <= '1';
      WHEN "1110011010" =>
            manhi <= conv_std_logic_vector(3863491,24);
            manlo <= conv_std_logic_vector(144123451,28);
           exponent <= '1';
      WHEN "1110011011" =>
            manhi <= conv_std_logic_vector(3883658,24);
            manlo <= conv_std_logic_vector(86789657,28);
           exponent <= '1';
      WHEN "1110011100" =>
            manhi <= conv_std_logic_vector(3903844,24);
            manlo <= conv_std_logic_vector(218366446,28);
           exponent <= '1';
      WHEN "1110011101" =>
            manhi <= conv_std_logic_vector(3924051,24);
            manlo <= conv_std_logic_vector(7150648,28);
           exponent <= '1';
      WHEN "1110011110" =>
            manhi <= conv_std_logic_vector(3944276,24);
            manlo <= conv_std_logic_vector(263621422,28);
           exponent <= '1';
      WHEN "1110011111" =>
            manhi <= conv_std_logic_vector(3964522,24);
            manlo <= conv_std_logic_vector(187650244,28);
           exponent <= '1';
      WHEN "1110100000" =>
            manhi <= conv_std_logic_vector(3984788,24);
            manlo <= conv_std_logic_vector(52855476,28);
           exponent <= '1';
      WHEN "1110100001" =>
            manhi <= conv_std_logic_vector(4005073,24);
            manlo <= conv_std_logic_vector(132860541,28);
           exponent <= '1';
      WHEN "1110100010" =>
            manhi <= conv_std_logic_vector(4025378,24);
            manlo <= conv_std_logic_vector(164423019,28);
           exponent <= '1';
      WHEN "1110100011" =>
            manhi <= conv_std_logic_vector(4045703,24);
            manlo <= conv_std_logic_vector(152741021,28);
           exponent <= '1';
      WHEN "1110100100" =>
            manhi <= conv_std_logic_vector(4066048,24);
            manlo <= conv_std_logic_vector(103017737,28);
           exponent <= '1';
      WHEN "1110100101" =>
            manhi <= conv_std_logic_vector(4086413,24);
            manlo <= conv_std_logic_vector(20461438,28);
           exponent <= '1';
      WHEN "1110100110" =>
            manhi <= conv_std_logic_vector(4106797,24);
            manlo <= conv_std_logic_vector(178720944,28);
           exponent <= '1';
      WHEN "1110100111" =>
            manhi <= conv_std_logic_vector(4127202,24);
            manlo <= conv_std_logic_vector(46143798,28);
           exponent <= '1';
      WHEN "1110101000" =>
            manhi <= conv_std_logic_vector(4147626,24);
            manlo <= conv_std_logic_vector(164824464,28);
           exponent <= '1';
      WHEN "1110101001" =>
            manhi <= conv_std_logic_vector(4168071,24);
            manlo <= conv_std_logic_vector(3120689,28);
           exponent <= '1';
      WHEN "1110101010" =>
            manhi <= conv_std_logic_vector(4188535,24);
            manlo <= conv_std_logic_vector(103137152,28);
           exponent <= '1';
      WHEN "1110101011" =>
            manhi <= conv_std_logic_vector(4209019,24);
            manlo <= conv_std_logic_vector(201677275,28);
           exponent <= '1';
      WHEN "1110101100" =>
            manhi <= conv_std_logic_vector(4229524,24);
            manlo <= conv_std_logic_vector(35549602,28);
           exponent <= '1';
      WHEN "1110101101" =>
            manhi <= conv_std_logic_vector(4250048,24);
            manlo <= conv_std_logic_vector(146874166,28);
           exponent <= '1';
      WHEN "1110101110" =>
            manhi <= conv_std_logic_vector(4270593,24);
            manlo <= conv_std_logic_vector(4034305,28);
           exponent <= '1';
      WHEN "1110101111" =>
            manhi <= conv_std_logic_vector(4291157,24);
            manlo <= conv_std_logic_vector(149160317,28);
           exponent <= '1';
      WHEN "1110110000" =>
            manhi <= conv_std_logic_vector(4311742,24);
            manlo <= conv_std_logic_vector(50645812,28);
           exponent <= '1';
      WHEN "1110110001" =>
            manhi <= conv_std_logic_vector(4332346,24);
            manlo <= conv_std_logic_vector(250631368,28);
           exponent <= '1';
      WHEN "1110110010" =>
            manhi <= conv_std_logic_vector(4352971,24);
            manlo <= conv_std_logic_vector(217520889,28);
           exponent <= '1';
      WHEN "1110110011" =>
            manhi <= conv_std_logic_vector(4373616,24);
            manlo <= conv_std_logic_vector(225029798,28);
           exponent <= '1';
      WHEN "1110110100" =>
            manhi <= conv_std_logic_vector(4394282,24);
            manlo <= conv_std_logic_vector(10007770,28);
           exponent <= '1';
      WHEN "1110110101" =>
            manhi <= conv_std_logic_vector(4414967,24);
            manlo <= conv_std_logic_vector(114616005,28);
           exponent <= '1';
      WHEN "1110110110" =>
            manhi <= conv_std_logic_vector(4435673,24);
            manlo <= conv_std_logic_vector(7279052,28);
           exponent <= '1';
      WHEN "1110110111" =>
            manhi <= conv_std_logic_vector(4456398,24);
            manlo <= conv_std_logic_vector(230168458,28);
           exponent <= '1';
      WHEN "1110111000" =>
            manhi <= conv_std_logic_vector(4477144,24);
            manlo <= conv_std_logic_vector(251719124,28);
           exponent <= '1';
      WHEN "1110111001" =>
            manhi <= conv_std_logic_vector(4497911,24);
            manlo <= conv_std_logic_vector(77242046,28);
           exponent <= '1';
      WHEN "1110111010" =>
            manhi <= conv_std_logic_vector(4518697,24);
            manlo <= conv_std_logic_vector(248924323,28);
           exponent <= '1';
      WHEN "1110111011" =>
            manhi <= conv_std_logic_vector(4539504,24);
            manlo <= conv_std_logic_vector(235216422,28);
           exponent <= '1';
      WHEN "1110111100" =>
            manhi <= conv_std_logic_vector(4560332,24);
            manlo <= conv_std_logic_vector(41444923,28);
           exponent <= '1';
      WHEN "1110111101" =>
            manhi <= conv_std_logic_vector(4581179,24);
            manlo <= conv_std_logic_vector(209812522,28);
           exponent <= '1';
      WHEN "1110111110" =>
            manhi <= conv_std_logic_vector(4602047,24);
            manlo <= conv_std_logic_vector(208785300,28);
           exponent <= '1';
      WHEN "1110111111" =>
            manhi <= conv_std_logic_vector(4622936,24);
            manlo <= conv_std_logic_vector(43705464,28);
           exponent <= '1';
      WHEN "1111000000" =>
            manhi <= conv_std_logic_vector(4643844,24);
            manlo <= conv_std_logic_vector(256791352,28);
           exponent <= '1';
      WHEN "1111000001" =>
            manhi <= conv_std_logic_vector(4664774,24);
            manlo <= conv_std_logic_vector(48089250,28);
           exponent <= '1';
      WHEN "1111000010" =>
            manhi <= conv_std_logic_vector(4685723,24);
            manlo <= conv_std_logic_vector(228263405,28);
           exponent <= '1';
      WHEN "1111000011" =>
            manhi <= conv_std_logic_vector(4706693,24);
            manlo <= conv_std_logic_vector(265806023,28);
           exponent <= '1';
      WHEN "1111000100" =>
            manhi <= conv_std_logic_vector(4727684,24);
            manlo <= conv_std_logic_vector(166085460,28);
           exponent <= '1';
      WHEN "1111000101" =>
            manhi <= conv_std_logic_vector(4748695,24);
            manlo <= conv_std_logic_vector(202910772,28);
           exponent <= '1';
      WHEN "1111000110" =>
            manhi <= conv_std_logic_vector(4769727,24);
            manlo <= conv_std_logic_vector(113225356,28);
           exponent <= '1';
      WHEN "1111000111" =>
            manhi <= conv_std_logic_vector(4790779,24);
            manlo <= conv_std_logic_vector(170848774,28);
           exponent <= '1';
      WHEN "1111001000" =>
            manhi <= conv_std_logic_vector(4811852,24);
            manlo <= conv_std_logic_vector(112734938,28);
           exponent <= '1';
      WHEN "1111001001" =>
            manhi <= conv_std_logic_vector(4832945,24);
            manlo <= conv_std_logic_vector(212713936,28);
           exponent <= '1';
      WHEN "1111001010" =>
            manhi <= conv_std_logic_vector(4854059,24);
            manlo <= conv_std_logic_vector(207750218,28);
           exponent <= '1';
      WHEN "1111001011" =>
            manhi <= conv_std_logic_vector(4875194,24);
            manlo <= conv_std_logic_vector(103248961,28);
           exponent <= '1';
      WHEN "1111001100" =>
            manhi <= conv_std_logic_vector(4896349,24);
            manlo <= conv_std_logic_vector(173056083,28);
           exponent <= '1';
      WHEN "1111001101" =>
            manhi <= conv_std_logic_vector(4917525,24);
            manlo <= conv_std_logic_vector(154151876,28);
           exponent <= '1';
      WHEN "1111001110" =>
            manhi <= conv_std_logic_vector(4938722,24);
            manlo <= conv_std_logic_vector(51957376,28);
           exponent <= '1';
      WHEN "1111001111" =>
            manhi <= conv_std_logic_vector(4959939,24);
            manlo <= conv_std_logic_vector(140334376,28);
           exponent <= '1';
      WHEN "1111010000" =>
            manhi <= conv_std_logic_vector(4981177,24);
            manlo <= conv_std_logic_vector(156279056,28);
           exponent <= '1';
      WHEN "1111010001" =>
            manhi <= conv_std_logic_vector(5002436,24);
            manlo <= conv_std_logic_vector(105228360,28);
           exponent <= '1';
      WHEN "1111010010" =>
            manhi <= conv_std_logic_vector(5023715,24);
            manlo <= conv_std_logic_vector(261060000,28);
           exponent <= '1';
      WHEN "1111010011" =>
            manhi <= conv_std_logic_vector(5045016,24);
            manlo <= conv_std_logic_vector(92350636,28);
           exponent <= '1';
      WHEN "1111010100" =>
            manhi <= conv_std_logic_vector(5066337,24);
            manlo <= conv_std_logic_vector(141424076,28);
           exponent <= '1';
      WHEN "1111010101" =>
            manhi <= conv_std_logic_vector(5087679,24);
            manlo <= conv_std_logic_vector(145303087,28);
           exponent <= '1';
      WHEN "1111010110" =>
            manhi <= conv_std_logic_vector(5109042,24);
            manlo <= conv_std_logic_vector(109451226,28);
           exponent <= '1';
      WHEN "1111010111" =>
            manhi <= conv_std_logic_vector(5130426,24);
            manlo <= conv_std_logic_vector(39337386,28);
           exponent <= '1';
      WHEN "1111011000" =>
            manhi <= conv_std_logic_vector(5151830,24);
            manlo <= conv_std_logic_vector(208871261,28);
           exponent <= '1';
      WHEN "1111011001" =>
            manhi <= conv_std_logic_vector(5173256,24);
            manlo <= conv_std_logic_vector(86661526,28);
           exponent <= '1';
      WHEN "1111011010" =>
            manhi <= conv_std_logic_vector(5194702,24);
            manlo <= conv_std_logic_vector(215064032,28);
           exponent <= '1';
      WHEN "1111011011" =>
            manhi <= conv_std_logic_vector(5216170,24);
            manlo <= conv_std_logic_vector(62698166,28);
           exponent <= '1';
      WHEN "1111011100" =>
            manhi <= conv_std_logic_vector(5237658,24);
            manlo <= conv_std_logic_vector(171930504,28);
           exponent <= '1';
      WHEN "1111011101" =>
            manhi <= conv_std_logic_vector(5259168,24);
            manlo <= conv_std_logic_vector(11391165,28);
           exponent <= '1';
      WHEN "1111011110" =>
            manhi <= conv_std_logic_vector(5280698,24);
            manlo <= conv_std_logic_vector(123457470,28);
           exponent <= '1';
      WHEN "1111011111" =>
            manhi <= conv_std_logic_vector(5302249,24);
            manlo <= conv_std_logic_vector(245205748,28);
           exponent <= '1';
      WHEN "1111100000" =>
            manhi <= conv_std_logic_vector(5323822,24);
            manlo <= conv_std_logic_vector(113717718,28);
           exponent <= '1';
      WHEN "1111100001" =>
            manhi <= conv_std_logic_vector(5345416,24);
            manlo <= conv_std_logic_vector(2951399,28);
           exponent <= '1';
      WHEN "1111100010" =>
            manhi <= conv_std_logic_vector(5367030,24);
            manlo <= conv_std_logic_vector(186870204,28);
           exponent <= '1';
      WHEN "1111100011" =>
            manhi <= conv_std_logic_vector(5388666,24);
            manlo <= conv_std_logic_vector(134136582,28);
           exponent <= '1';
      WHEN "1111100100" =>
            manhi <= conv_std_logic_vector(5410323,24);
            manlo <= conv_std_logic_vector(118724754,28);
           exponent <= '1';
      WHEN "1111100101" =>
            manhi <= conv_std_logic_vector(5432001,24);
            manlo <= conv_std_logic_vector(146178900,28);
           exponent <= '1';
      WHEN "1111100110" =>
            manhi <= conv_std_logic_vector(5453700,24);
            manlo <= conv_std_logic_vector(222048612,28);
           exponent <= '1';
      WHEN "1111100111" =>
            manhi <= conv_std_logic_vector(5475421,24);
            manlo <= conv_std_logic_vector(83453453,28);
           exponent <= '1';
      WHEN "1111101000" =>
            manhi <= conv_std_logic_vector(5497163,24);
            manlo <= conv_std_logic_vector(4389322,28);
           exponent <= '1';
      WHEN "1111101001" =>
            manhi <= conv_std_logic_vector(5518925,24);
            manlo <= conv_std_logic_vector(258857552,28);
           exponent <= '1';
      WHEN "1111101010" =>
            manhi <= conv_std_logic_vector(5540710,24);
            manlo <= conv_std_logic_vector(47123091,28);
           exponent <= '1';
      WHEN "1111101011" =>
            manhi <= conv_std_logic_vector(5562515,24);
            manlo <= conv_std_logic_vector(180069064,28);
           exponent <= '1';
      WHEN "1111101100" =>
            manhi <= conv_std_logic_vector(5584342,24);
            manlo <= conv_std_logic_vector(126406768,28);
           exponent <= '1';
      WHEN "1111101101" =>
            manhi <= conv_std_logic_vector(5606190,24);
            manlo <= conv_std_logic_vector(160159320,28);
           exponent <= '1';
      WHEN "1111101110" =>
            manhi <= conv_std_logic_vector(5628060,24);
            manlo <= conv_std_logic_vector(18484384,28);
           exponent <= '1';
      WHEN "1111101111" =>
            manhi <= conv_std_logic_vector(5649950,24);
            manlo <= conv_std_logic_vector(243851457,28);
           exponent <= '1';
      WHEN "1111110000" =>
            manhi <= conv_std_logic_vector(5671863,24);
            manlo <= conv_std_logic_vector(36558227,28);
           exponent <= '1';
      WHEN "1111110001" =>
            manhi <= conv_std_logic_vector(5693796,24);
            manlo <= conv_std_logic_vector(207520592,28);
           exponent <= '1';
      WHEN "1111110010" =>
            manhi <= conv_std_logic_vector(5715751,24);
            manlo <= conv_std_logic_vector(225482653,28);
           exponent <= '1';
      WHEN "1111110011" =>
            manhi <= conv_std_logic_vector(5737728,24);
            manlo <= conv_std_logic_vector(96064906,28);
           exponent <= '1';
      WHEN "1111110100" =>
            manhi <= conv_std_logic_vector(5759726,24);
            manlo <= conv_std_logic_vector(93328797,28);
           exponent <= '1';
      WHEN "1111110101" =>
            manhi <= conv_std_logic_vector(5781745,24);
            manlo <= conv_std_logic_vector(222905812,28);
           exponent <= '1';
      WHEN "1111110110" =>
            manhi <= conv_std_logic_vector(5803786,24);
            manlo <= conv_std_logic_vector(221997482,28);
           exponent <= '1';
      WHEN "1111110111" =>
            manhi <= conv_std_logic_vector(5825849,24);
            manlo <= conv_std_logic_vector(96246303,28);
           exponent <= '1';
      WHEN "1111111000" =>
            manhi <= conv_std_logic_vector(5847933,24);
            manlo <= conv_std_logic_vector(119735740,28);
           exponent <= '1';
      WHEN "1111111001" =>
            manhi <= conv_std_logic_vector(5870039,24);
            manlo <= conv_std_logic_vector(29683863,28);
           exponent <= '1';
      WHEN "1111111010" =>
            manhi <= conv_std_logic_vector(5892166,24);
            manlo <= conv_std_logic_vector(100185179,28);
           exponent <= '1';
      WHEN "1111111011" =>
            manhi <= conv_std_logic_vector(5914315,24);
            manlo <= conv_std_logic_vector(68468812,28);
           exponent <= '1';
      WHEN "1111111100" =>
            manhi <= conv_std_logic_vector(5936485,24);
            manlo <= conv_std_logic_vector(208640332,28);
           exponent <= '1';
      WHEN "1111111101" =>
            manhi <= conv_std_logic_vector(5958677,24);
            manlo <= conv_std_logic_vector(257939938,28);
           exponent <= '1';
      WHEN "1111111110" =>
            manhi <= conv_std_logic_vector(5980891,24);
            manlo <= conv_std_logic_vector(222048827,28);
           exponent <= '1';
      WHEN "1111111111" =>
            manhi <= conv_std_logic_vector(6003127,24);
            manlo <= conv_std_logic_vector(106653752,28);
           exponent <= '1';
      WHEN others =>
           manhi <= conv_std_logic_vector(0,24);
           manlo <= conv_std_logic_vector(0,28);
           exponent <= '0';
    END CASE;
  END PROCESS;

END rtl;
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   DP_EXPLUT20.VHD                           ***
--***                                             ***
--***   Function: Look Up Table - EXP()           ***
--***                                             ***
--***   Generated by MATLAB Utility               ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_explut20 IS
PORT (
      add : IN STD_LOGIC_VECTOR (10 DOWNTO 1);
      manhi : OUT STD_LOGIC_VECTOR (24 DOWNTO 1);
      manlo : OUT STD_LOGIC_VECTOR (28 DOWNTO 1)
     );
END dp_explut20;

ARCHITECTURE rtl OF dp_explut20 IS

BEGIN

  pca: PROCESS (add)
  BEGIN
    CASE add IS
      WHEN "0000000000" =>
            manhi <= conv_std_logic_vector(0,24);
            manlo <= conv_std_logic_vector(0,28);
      WHEN "0000000001" =>
            manhi <= conv_std_logic_vector(16,24);
            manlo <= conv_std_logic_vector(2048,28);
      WHEN "0000000010" =>
            manhi <= conv_std_logic_vector(32,24);
            manlo <= conv_std_logic_vector(8192,28);
      WHEN "0000000011" =>
            manhi <= conv_std_logic_vector(48,24);
            manlo <= conv_std_logic_vector(18432,28);
      WHEN "0000000100" =>
            manhi <= conv_std_logic_vector(64,24);
            manlo <= conv_std_logic_vector(32768,28);
      WHEN "0000000101" =>
            manhi <= conv_std_logic_vector(80,24);
            manlo <= conv_std_logic_vector(51200,28);
      WHEN "0000000110" =>
            manhi <= conv_std_logic_vector(96,24);
            manlo <= conv_std_logic_vector(73728,28);
      WHEN "0000000111" =>
            manhi <= conv_std_logic_vector(112,24);
            manlo <= conv_std_logic_vector(100352,28);
      WHEN "0000001000" =>
            manhi <= conv_std_logic_vector(128,24);
            manlo <= conv_std_logic_vector(131072,28);
      WHEN "0000001001" =>
            manhi <= conv_std_logic_vector(144,24);
            manlo <= conv_std_logic_vector(165888,28);
      WHEN "0000001010" =>
            manhi <= conv_std_logic_vector(160,24);
            manlo <= conv_std_logic_vector(204801,28);
      WHEN "0000001011" =>
            manhi <= conv_std_logic_vector(176,24);
            manlo <= conv_std_logic_vector(247809,28);
      WHEN "0000001100" =>
            manhi <= conv_std_logic_vector(192,24);
            manlo <= conv_std_logic_vector(294913,28);
      WHEN "0000001101" =>
            manhi <= conv_std_logic_vector(208,24);
            manlo <= conv_std_logic_vector(346113,28);
      WHEN "0000001110" =>
            manhi <= conv_std_logic_vector(224,24);
            manlo <= conv_std_logic_vector(401410,28);
      WHEN "0000001111" =>
            manhi <= conv_std_logic_vector(240,24);
            manlo <= conv_std_logic_vector(460802,28);
      WHEN "0000010000" =>
            manhi <= conv_std_logic_vector(256,24);
            manlo <= conv_std_logic_vector(524291,28);
      WHEN "0000010001" =>
            manhi <= conv_std_logic_vector(272,24);
            manlo <= conv_std_logic_vector(591875,28);
      WHEN "0000010010" =>
            manhi <= conv_std_logic_vector(288,24);
            manlo <= conv_std_logic_vector(663556,28);
      WHEN "0000010011" =>
            manhi <= conv_std_logic_vector(304,24);
            manlo <= conv_std_logic_vector(739332,28);
      WHEN "0000010100" =>
            manhi <= conv_std_logic_vector(320,24);
            manlo <= conv_std_logic_vector(819205,28);
      WHEN "0000010101" =>
            manhi <= conv_std_logic_vector(336,24);
            manlo <= conv_std_logic_vector(903174,28);
      WHEN "0000010110" =>
            manhi <= conv_std_logic_vector(352,24);
            manlo <= conv_std_logic_vector(991239,28);
      WHEN "0000010111" =>
            manhi <= conv_std_logic_vector(368,24);
            manlo <= conv_std_logic_vector(1083400,28);
      WHEN "0000011000" =>
            manhi <= conv_std_logic_vector(384,24);
            manlo <= conv_std_logic_vector(1179657,28);
      WHEN "0000011001" =>
            manhi <= conv_std_logic_vector(400,24);
            manlo <= conv_std_logic_vector(1280010,28);
      WHEN "0000011010" =>
            manhi <= conv_std_logic_vector(416,24);
            manlo <= conv_std_logic_vector(1384459,28);
      WHEN "0000011011" =>
            manhi <= conv_std_logic_vector(432,24);
            manlo <= conv_std_logic_vector(1493005,28);
      WHEN "0000011100" =>
            manhi <= conv_std_logic_vector(448,24);
            manlo <= conv_std_logic_vector(1605646,28);
      WHEN "0000011101" =>
            manhi <= conv_std_logic_vector(464,24);
            manlo <= conv_std_logic_vector(1722384,28);
      WHEN "0000011110" =>
            manhi <= conv_std_logic_vector(480,24);
            manlo <= conv_std_logic_vector(1843218,28);
      WHEN "0000011111" =>
            manhi <= conv_std_logic_vector(496,24);
            manlo <= conv_std_logic_vector(1968147,28);
      WHEN "0000100000" =>
            manhi <= conv_std_logic_vector(512,24);
            manlo <= conv_std_logic_vector(2097173,28);
      WHEN "0000100001" =>
            manhi <= conv_std_logic_vector(528,24);
            manlo <= conv_std_logic_vector(2230295,28);
      WHEN "0000100010" =>
            manhi <= conv_std_logic_vector(544,24);
            manlo <= conv_std_logic_vector(2367514,28);
      WHEN "0000100011" =>
            manhi <= conv_std_logic_vector(560,24);
            manlo <= conv_std_logic_vector(2508828,28);
      WHEN "0000100100" =>
            manhi <= conv_std_logic_vector(576,24);
            manlo <= conv_std_logic_vector(2654238,28);
      WHEN "0000100101" =>
            manhi <= conv_std_logic_vector(592,24);
            manlo <= conv_std_logic_vector(2803745,28);
      WHEN "0000100110" =>
            manhi <= conv_std_logic_vector(608,24);
            manlo <= conv_std_logic_vector(2957348,28);
      WHEN "0000100111" =>
            manhi <= conv_std_logic_vector(624,24);
            manlo <= conv_std_logic_vector(3115047,28);
      WHEN "0000101000" =>
            manhi <= conv_std_logic_vector(640,24);
            manlo <= conv_std_logic_vector(3276842,28);
      WHEN "0000101001" =>
            manhi <= conv_std_logic_vector(656,24);
            manlo <= conv_std_logic_vector(3442733,28);
      WHEN "0000101010" =>
            manhi <= conv_std_logic_vector(672,24);
            manlo <= conv_std_logic_vector(3612720,28);
      WHEN "0000101011" =>
            manhi <= conv_std_logic_vector(688,24);
            manlo <= conv_std_logic_vector(3786804,28);
      WHEN "0000101100" =>
            manhi <= conv_std_logic_vector(704,24);
            manlo <= conv_std_logic_vector(3964983,28);
      WHEN "0000101101" =>
            manhi <= conv_std_logic_vector(720,24);
            manlo <= conv_std_logic_vector(4147259,28);
      WHEN "0000101110" =>
            manhi <= conv_std_logic_vector(736,24);
            manlo <= conv_std_logic_vector(4333631,28);
      WHEN "0000101111" =>
            manhi <= conv_std_logic_vector(752,24);
            manlo <= conv_std_logic_vector(4524100,28);
      WHEN "0000110000" =>
            manhi <= conv_std_logic_vector(768,24);
            manlo <= conv_std_logic_vector(4718664,28);
      WHEN "0000110001" =>
            manhi <= conv_std_logic_vector(784,24);
            manlo <= conv_std_logic_vector(4917325,28);
      WHEN "0000110010" =>
            manhi <= conv_std_logic_vector(800,24);
            manlo <= conv_std_logic_vector(5120081,28);
      WHEN "0000110011" =>
            manhi <= conv_std_logic_vector(816,24);
            manlo <= conv_std_logic_vector(5326934,28);
      WHEN "0000110100" =>
            manhi <= conv_std_logic_vector(832,24);
            manlo <= conv_std_logic_vector(5537884,28);
      WHEN "0000110101" =>
            manhi <= conv_std_logic_vector(848,24);
            manlo <= conv_std_logic_vector(5752929,28);
      WHEN "0000110110" =>
            manhi <= conv_std_logic_vector(864,24);
            manlo <= conv_std_logic_vector(5972071,28);
      WHEN "0000110111" =>
            manhi <= conv_std_logic_vector(880,24);
            manlo <= conv_std_logic_vector(6195308,28);
      WHEN "0000111000" =>
            manhi <= conv_std_logic_vector(896,24);
            manlo <= conv_std_logic_vector(6422642,28);
      WHEN "0000111001" =>
            manhi <= conv_std_logic_vector(912,24);
            manlo <= conv_std_logic_vector(6654073,28);
      WHEN "0000111010" =>
            manhi <= conv_std_logic_vector(928,24);
            manlo <= conv_std_logic_vector(6889599,28);
      WHEN "0000111011" =>
            manhi <= conv_std_logic_vector(944,24);
            manlo <= conv_std_logic_vector(7129222,28);
      WHEN "0000111100" =>
            manhi <= conv_std_logic_vector(960,24);
            manlo <= conv_std_logic_vector(7372941,28);
      WHEN "0000111101" =>
            manhi <= conv_std_logic_vector(976,24);
            manlo <= conv_std_logic_vector(7620756,28);
      WHEN "0000111110" =>
            manhi <= conv_std_logic_vector(992,24);
            manlo <= conv_std_logic_vector(7872667,28);
      WHEN "0000111111" =>
            manhi <= conv_std_logic_vector(1008,24);
            manlo <= conv_std_logic_vector(8128675,28);
      WHEN "0001000000" =>
            manhi <= conv_std_logic_vector(1024,24);
            manlo <= conv_std_logic_vector(8388779,28);
      WHEN "0001000001" =>
            manhi <= conv_std_logic_vector(1040,24);
            manlo <= conv_std_logic_vector(8652979,28);
      WHEN "0001000010" =>
            manhi <= conv_std_logic_vector(1056,24);
            manlo <= conv_std_logic_vector(8921275,28);
      WHEN "0001000011" =>
            manhi <= conv_std_logic_vector(1072,24);
            manlo <= conv_std_logic_vector(9193668,28);
      WHEN "0001000100" =>
            manhi <= conv_std_logic_vector(1088,24);
            manlo <= conv_std_logic_vector(9470157,28);
      WHEN "0001000101" =>
            manhi <= conv_std_logic_vector(1104,24);
            manlo <= conv_std_logic_vector(9750742,28);
      WHEN "0001000110" =>
            manhi <= conv_std_logic_vector(1120,24);
            manlo <= conv_std_logic_vector(10035423,28);
      WHEN "0001000111" =>
            manhi <= conv_std_logic_vector(1136,24);
            manlo <= conv_std_logic_vector(10324201,28);
      WHEN "0001001000" =>
            manhi <= conv_std_logic_vector(1152,24);
            manlo <= conv_std_logic_vector(10617075,28);
      WHEN "0001001001" =>
            manhi <= conv_std_logic_vector(1168,24);
            manlo <= conv_std_logic_vector(10914045,28);
      WHEN "0001001010" =>
            manhi <= conv_std_logic_vector(1184,24);
            manlo <= conv_std_logic_vector(11215112,28);
      WHEN "0001001011" =>
            manhi <= conv_std_logic_vector(1200,24);
            manlo <= conv_std_logic_vector(11520275,28);
      WHEN "0001001100" =>
            manhi <= conv_std_logic_vector(1216,24);
            manlo <= conv_std_logic_vector(11829534,28);
      WHEN "0001001101" =>
            manhi <= conv_std_logic_vector(1232,24);
            manlo <= conv_std_logic_vector(12142889,28);
      WHEN "0001001110" =>
            manhi <= conv_std_logic_vector(1248,24);
            manlo <= conv_std_logic_vector(12460341,28);
      WHEN "0001001111" =>
            manhi <= conv_std_logic_vector(1264,24);
            manlo <= conv_std_logic_vector(12781889,28);
      WHEN "0001010000" =>
            manhi <= conv_std_logic_vector(1280,24);
            manlo <= conv_std_logic_vector(13107533,28);
      WHEN "0001010001" =>
            manhi <= conv_std_logic_vector(1296,24);
            manlo <= conv_std_logic_vector(13437274,28);
      WHEN "0001010010" =>
            manhi <= conv_std_logic_vector(1312,24);
            manlo <= conv_std_logic_vector(13771111,28);
      WHEN "0001010011" =>
            manhi <= conv_std_logic_vector(1328,24);
            manlo <= conv_std_logic_vector(14109044,28);
      WHEN "0001010100" =>
            manhi <= conv_std_logic_vector(1344,24);
            manlo <= conv_std_logic_vector(14451074,28);
      WHEN "0001010101" =>
            manhi <= conv_std_logic_vector(1360,24);
            manlo <= conv_std_logic_vector(14797200,28);
      WHEN "0001010110" =>
            manhi <= conv_std_logic_vector(1376,24);
            manlo <= conv_std_logic_vector(15147422,28);
      WHEN "0001010111" =>
            manhi <= conv_std_logic_vector(1392,24);
            manlo <= conv_std_logic_vector(15501741,28);
      WHEN "0001011000" =>
            manhi <= conv_std_logic_vector(1408,24);
            manlo <= conv_std_logic_vector(15860156,28);
      WHEN "0001011001" =>
            manhi <= conv_std_logic_vector(1424,24);
            manlo <= conv_std_logic_vector(16222667,28);
      WHEN "0001011010" =>
            manhi <= conv_std_logic_vector(1440,24);
            manlo <= conv_std_logic_vector(16589275,28);
      WHEN "0001011011" =>
            manhi <= conv_std_logic_vector(1456,24);
            manlo <= conv_std_logic_vector(16959979,28);
      WHEN "0001011100" =>
            manhi <= conv_std_logic_vector(1472,24);
            manlo <= conv_std_logic_vector(17334779,28);
      WHEN "0001011101" =>
            manhi <= conv_std_logic_vector(1488,24);
            manlo <= conv_std_logic_vector(17713676,28);
      WHEN "0001011110" =>
            manhi <= conv_std_logic_vector(1504,24);
            manlo <= conv_std_logic_vector(18096669,28);
      WHEN "0001011111" =>
            manhi <= conv_std_logic_vector(1520,24);
            manlo <= conv_std_logic_vector(18483758,28);
      WHEN "0001100000" =>
            manhi <= conv_std_logic_vector(1536,24);
            manlo <= conv_std_logic_vector(18874944,28);
      WHEN "0001100001" =>
            manhi <= conv_std_logic_vector(1552,24);
            manlo <= conv_std_logic_vector(19270226,28);
      WHEN "0001100010" =>
            manhi <= conv_std_logic_vector(1568,24);
            manlo <= conv_std_logic_vector(19669605,28);
      WHEN "0001100011" =>
            manhi <= conv_std_logic_vector(1584,24);
            manlo <= conv_std_logic_vector(20073080,28);
      WHEN "0001100100" =>
            manhi <= conv_std_logic_vector(1600,24);
            manlo <= conv_std_logic_vector(20480651,28);
      WHEN "0001100101" =>
            manhi <= conv_std_logic_vector(1616,24);
            manlo <= conv_std_logic_vector(20892319,28);
      WHEN "0001100110" =>
            manhi <= conv_std_logic_vector(1632,24);
            manlo <= conv_std_logic_vector(21308083,28);
      WHEN "0001100111" =>
            manhi <= conv_std_logic_vector(1648,24);
            manlo <= conv_std_logic_vector(21727943,28);
      WHEN "0001101000" =>
            manhi <= conv_std_logic_vector(1664,24);
            manlo <= conv_std_logic_vector(22151900,28);
      WHEN "0001101001" =>
            manhi <= conv_std_logic_vector(1680,24);
            manlo <= conv_std_logic_vector(22579954,28);
      WHEN "0001101010" =>
            manhi <= conv_std_logic_vector(1696,24);
            manlo <= conv_std_logic_vector(23012103,28);
      WHEN "0001101011" =>
            manhi <= conv_std_logic_vector(1712,24);
            manlo <= conv_std_logic_vector(23448350,28);
      WHEN "0001101100" =>
            manhi <= conv_std_logic_vector(1728,24);
            manlo <= conv_std_logic_vector(23888692,28);
      WHEN "0001101101" =>
            manhi <= conv_std_logic_vector(1744,24);
            manlo <= conv_std_logic_vector(24333131,28);
      WHEN "0001101110" =>
            manhi <= conv_std_logic_vector(1760,24);
            manlo <= conv_std_logic_vector(24781667,28);
      WHEN "0001101111" =>
            manhi <= conv_std_logic_vector(1776,24);
            manlo <= conv_std_logic_vector(25234298,28);
      WHEN "0001110000" =>
            manhi <= conv_std_logic_vector(1792,24);
            manlo <= conv_std_logic_vector(25691027,28);
      WHEN "0001110001" =>
            manhi <= conv_std_logic_vector(1808,24);
            manlo <= conv_std_logic_vector(26151851,28);
      WHEN "0001110010" =>
            manhi <= conv_std_logic_vector(1824,24);
            manlo <= conv_std_logic_vector(26616773,28);
      WHEN "0001110011" =>
            manhi <= conv_std_logic_vector(1840,24);
            manlo <= conv_std_logic_vector(27085790,28);
      WHEN "0001110100" =>
            manhi <= conv_std_logic_vector(1856,24);
            manlo <= conv_std_logic_vector(27558904,28);
      WHEN "0001110101" =>
            manhi <= conv_std_logic_vector(1872,24);
            manlo <= conv_std_logic_vector(28036115,28);
      WHEN "0001110110" =>
            manhi <= conv_std_logic_vector(1888,24);
            manlo <= conv_std_logic_vector(28517422,28);
      WHEN "0001110111" =>
            manhi <= conv_std_logic_vector(1904,24);
            manlo <= conv_std_logic_vector(29002825,28);
      WHEN "0001111000" =>
            manhi <= conv_std_logic_vector(1920,24);
            manlo <= conv_std_logic_vector(29492325,28);
      WHEN "0001111001" =>
            manhi <= conv_std_logic_vector(1936,24);
            manlo <= conv_std_logic_vector(29985921,28);
      WHEN "0001111010" =>
            manhi <= conv_std_logic_vector(1952,24);
            manlo <= conv_std_logic_vector(30483614,28);
      WHEN "0001111011" =>
            manhi <= conv_std_logic_vector(1968,24);
            manlo <= conv_std_logic_vector(30985404,28);
      WHEN "0001111100" =>
            manhi <= conv_std_logic_vector(1984,24);
            manlo <= conv_std_logic_vector(31491289,28);
      WHEN "0001111101" =>
            manhi <= conv_std_logic_vector(2000,24);
            manlo <= conv_std_logic_vector(32001272,28);
      WHEN "0001111110" =>
            manhi <= conv_std_logic_vector(2016,24);
            manlo <= conv_std_logic_vector(32515350,28);
      WHEN "0001111111" =>
            manhi <= conv_std_logic_vector(2032,24);
            manlo <= conv_std_logic_vector(33033526,28);
      WHEN "0010000000" =>
            manhi <= conv_std_logic_vector(2048,24);
            manlo <= conv_std_logic_vector(33555797,28);
      WHEN "0010000001" =>
            manhi <= conv_std_logic_vector(2064,24);
            manlo <= conv_std_logic_vector(34082166,28);
      WHEN "0010000010" =>
            manhi <= conv_std_logic_vector(2080,24);
            manlo <= conv_std_logic_vector(34612630,28);
      WHEN "0010000011" =>
            manhi <= conv_std_logic_vector(2096,24);
            manlo <= conv_std_logic_vector(35147192,28);
      WHEN "0010000100" =>
            manhi <= conv_std_logic_vector(2112,24);
            manlo <= conv_std_logic_vector(35685849,28);
      WHEN "0010000101" =>
            manhi <= conv_std_logic_vector(2128,24);
            manlo <= conv_std_logic_vector(36228604,28);
      WHEN "0010000110" =>
            manhi <= conv_std_logic_vector(2144,24);
            manlo <= conv_std_logic_vector(36775455,28);
      WHEN "0010000111" =>
            manhi <= conv_std_logic_vector(2160,24);
            manlo <= conv_std_logic_vector(37326402,28);
      WHEN "0010001000" =>
            manhi <= conv_std_logic_vector(2176,24);
            manlo <= conv_std_logic_vector(37881446,28);
      WHEN "0010001001" =>
            manhi <= conv_std_logic_vector(2192,24);
            manlo <= conv_std_logic_vector(38440586,28);
      WHEN "0010001010" =>
            manhi <= conv_std_logic_vector(2208,24);
            manlo <= conv_std_logic_vector(39003823,28);
      WHEN "0010001011" =>
            manhi <= conv_std_logic_vector(2224,24);
            manlo <= conv_std_logic_vector(39571157,28);
      WHEN "0010001100" =>
            manhi <= conv_std_logic_vector(2240,24);
            manlo <= conv_std_logic_vector(40142587,28);
      WHEN "0010001101" =>
            manhi <= conv_std_logic_vector(2256,24);
            manlo <= conv_std_logic_vector(40718113,28);
      WHEN "0010001110" =>
            manhi <= conv_std_logic_vector(2272,24);
            manlo <= conv_std_logic_vector(41297736,28);
      WHEN "0010001111" =>
            manhi <= conv_std_logic_vector(2288,24);
            manlo <= conv_std_logic_vector(41881456,28);
      WHEN "0010010000" =>
            manhi <= conv_std_logic_vector(2304,24);
            manlo <= conv_std_logic_vector(42469272,28);
      WHEN "0010010001" =>
            manhi <= conv_std_logic_vector(2320,24);
            manlo <= conv_std_logic_vector(43061185,28);
      WHEN "0010010010" =>
            manhi <= conv_std_logic_vector(2336,24);
            manlo <= conv_std_logic_vector(43657194,28);
      WHEN "0010010011" =>
            manhi <= conv_std_logic_vector(2352,24);
            manlo <= conv_std_logic_vector(44257300,28);
      WHEN "0010010100" =>
            manhi <= conv_std_logic_vector(2368,24);
            manlo <= conv_std_logic_vector(44861503,28);
      WHEN "0010010101" =>
            manhi <= conv_std_logic_vector(2384,24);
            manlo <= conv_std_logic_vector(45469802,28);
      WHEN "0010010110" =>
            manhi <= conv_std_logic_vector(2400,24);
            manlo <= conv_std_logic_vector(46082197,28);
      WHEN "0010010111" =>
            manhi <= conv_std_logic_vector(2416,24);
            manlo <= conv_std_logic_vector(46698690,28);
      WHEN "0010011000" =>
            manhi <= conv_std_logic_vector(2432,24);
            manlo <= conv_std_logic_vector(47319278,28);
      WHEN "0010011001" =>
            manhi <= conv_std_logic_vector(2448,24);
            manlo <= conv_std_logic_vector(47943964,28);
      WHEN "0010011010" =>
            manhi <= conv_std_logic_vector(2464,24);
            manlo <= conv_std_logic_vector(48572746,28);
      WHEN "0010011011" =>
            manhi <= conv_std_logic_vector(2480,24);
            manlo <= conv_std_logic_vector(49205624,28);
      WHEN "0010011100" =>
            manhi <= conv_std_logic_vector(2496,24);
            manlo <= conv_std_logic_vector(49842600,28);
      WHEN "0010011101" =>
            manhi <= conv_std_logic_vector(2512,24);
            manlo <= conv_std_logic_vector(50483672,28);
      WHEN "0010011110" =>
            manhi <= conv_std_logic_vector(2528,24);
            manlo <= conv_std_logic_vector(51128840,28);
      WHEN "0010011111" =>
            manhi <= conv_std_logic_vector(2544,24);
            manlo <= conv_std_logic_vector(51778105,28);
      WHEN "0010100000" =>
            manhi <= conv_std_logic_vector(2560,24);
            manlo <= conv_std_logic_vector(52431467,28);
      WHEN "0010100001" =>
            manhi <= conv_std_logic_vector(2576,24);
            manlo <= conv_std_logic_vector(53088925,28);
      WHEN "0010100010" =>
            manhi <= conv_std_logic_vector(2592,24);
            manlo <= conv_std_logic_vector(53750480,28);
      WHEN "0010100011" =>
            manhi <= conv_std_logic_vector(2608,24);
            manlo <= conv_std_logic_vector(54416132,28);
      WHEN "0010100100" =>
            manhi <= conv_std_logic_vector(2624,24);
            manlo <= conv_std_logic_vector(55085880,28);
      WHEN "0010100101" =>
            manhi <= conv_std_logic_vector(2640,24);
            manlo <= conv_std_logic_vector(55759725,28);
      WHEN "0010100110" =>
            manhi <= conv_std_logic_vector(2656,24);
            manlo <= conv_std_logic_vector(56437666,28);
      WHEN "0010100111" =>
            manhi <= conv_std_logic_vector(2672,24);
            manlo <= conv_std_logic_vector(57119704,28);
      WHEN "0010101000" =>
            manhi <= conv_std_logic_vector(2688,24);
            manlo <= conv_std_logic_vector(57805839,28);
      WHEN "0010101001" =>
            manhi <= conv_std_logic_vector(2704,24);
            manlo <= conv_std_logic_vector(58496071,28);
      WHEN "0010101010" =>
            manhi <= conv_std_logic_vector(2720,24);
            manlo <= conv_std_logic_vector(59190399,28);
      WHEN "0010101011" =>
            manhi <= conv_std_logic_vector(2736,24);
            manlo <= conv_std_logic_vector(59888823,28);
      WHEN "0010101100" =>
            manhi <= conv_std_logic_vector(2752,24);
            manlo <= conv_std_logic_vector(60591345,28);
      WHEN "0010101101" =>
            manhi <= conv_std_logic_vector(2768,24);
            manlo <= conv_std_logic_vector(61297963,28);
      WHEN "0010101110" =>
            manhi <= conv_std_logic_vector(2784,24);
            manlo <= conv_std_logic_vector(62008678,28);
      WHEN "0010101111" =>
            manhi <= conv_std_logic_vector(2800,24);
            manlo <= conv_std_logic_vector(62723489,28);
      WHEN "0010110000" =>
            manhi <= conv_std_logic_vector(2816,24);
            manlo <= conv_std_logic_vector(63442397,28);
      WHEN "0010110001" =>
            manhi <= conv_std_logic_vector(2832,24);
            manlo <= conv_std_logic_vector(64165402,28);
      WHEN "0010110010" =>
            manhi <= conv_std_logic_vector(2848,24);
            manlo <= conv_std_logic_vector(64892504,28);
      WHEN "0010110011" =>
            manhi <= conv_std_logic_vector(2864,24);
            manlo <= conv_std_logic_vector(65623702,28);
      WHEN "0010110100" =>
            manhi <= conv_std_logic_vector(2880,24);
            manlo <= conv_std_logic_vector(66358997,28);
      WHEN "0010110101" =>
            manhi <= conv_std_logic_vector(2896,24);
            manlo <= conv_std_logic_vector(67098389,28);
      WHEN "0010110110" =>
            manhi <= conv_std_logic_vector(2912,24);
            manlo <= conv_std_logic_vector(67841877,28);
      WHEN "0010110111" =>
            manhi <= conv_std_logic_vector(2928,24);
            manlo <= conv_std_logic_vector(68589462,28);
      WHEN "0010111000" =>
            manhi <= conv_std_logic_vector(2944,24);
            manlo <= conv_std_logic_vector(69341144,28);
      WHEN "0010111001" =>
            manhi <= conv_std_logic_vector(2960,24);
            manlo <= conv_std_logic_vector(70096922,28);
      WHEN "0010111010" =>
            manhi <= conv_std_logic_vector(2976,24);
            manlo <= conv_std_logic_vector(70856798,28);
      WHEN "0010111011" =>
            manhi <= conv_std_logic_vector(2992,24);
            manlo <= conv_std_logic_vector(71620769,28);
      WHEN "0010111100" =>
            manhi <= conv_std_logic_vector(3008,24);
            manlo <= conv_std_logic_vector(72388838,28);
      WHEN "0010111101" =>
            manhi <= conv_std_logic_vector(3024,24);
            manlo <= conv_std_logic_vector(73161004,28);
      WHEN "0010111110" =>
            manhi <= conv_std_logic_vector(3040,24);
            manlo <= conv_std_logic_vector(73937266,28);
      WHEN "0010111111" =>
            manhi <= conv_std_logic_vector(3056,24);
            manlo <= conv_std_logic_vector(74717625,28);
      WHEN "0011000000" =>
            manhi <= conv_std_logic_vector(3072,24);
            manlo <= conv_std_logic_vector(75502080,28);
      WHEN "0011000001" =>
            manhi <= conv_std_logic_vector(3088,24);
            manlo <= conv_std_logic_vector(76290633,28);
      WHEN "0011000010" =>
            manhi <= conv_std_logic_vector(3104,24);
            manlo <= conv_std_logic_vector(77083282,28);
      WHEN "0011000011" =>
            manhi <= conv_std_logic_vector(3120,24);
            manlo <= conv_std_logic_vector(77880028,28);
      WHEN "0011000100" =>
            manhi <= conv_std_logic_vector(3136,24);
            manlo <= conv_std_logic_vector(78680870,28);
      WHEN "0011000101" =>
            manhi <= conv_std_logic_vector(3152,24);
            manlo <= conv_std_logic_vector(79485810,28);
      WHEN "0011000110" =>
            manhi <= conv_std_logic_vector(3168,24);
            manlo <= conv_std_logic_vector(80294846,28);
      WHEN "0011000111" =>
            manhi <= conv_std_logic_vector(3184,24);
            manlo <= conv_std_logic_vector(81107979,28);
      WHEN "0011001000" =>
            manhi <= conv_std_logic_vector(3200,24);
            manlo <= conv_std_logic_vector(81925209,28);
      WHEN "0011001001" =>
            manhi <= conv_std_logic_vector(3216,24);
            manlo <= conv_std_logic_vector(82746535,28);
      WHEN "0011001010" =>
            manhi <= conv_std_logic_vector(3232,24);
            manlo <= conv_std_logic_vector(83571958,28);
      WHEN "0011001011" =>
            manhi <= conv_std_logic_vector(3248,24);
            manlo <= conv_std_logic_vector(84401479,28);
      WHEN "0011001100" =>
            manhi <= conv_std_logic_vector(3264,24);
            manlo <= conv_std_logic_vector(85235095,28);
      WHEN "0011001101" =>
            manhi <= conv_std_logic_vector(3280,24);
            manlo <= conv_std_logic_vector(86072809,28);
      WHEN "0011001110" =>
            manhi <= conv_std_logic_vector(3296,24);
            manlo <= conv_std_logic_vector(86914620,28);
      WHEN "0011001111" =>
            manhi <= conv_std_logic_vector(3312,24);
            manlo <= conv_std_logic_vector(87760527,28);
      WHEN "0011010000" =>
            manhi <= conv_std_logic_vector(3328,24);
            manlo <= conv_std_logic_vector(88610531,28);
      WHEN "0011010001" =>
            manhi <= conv_std_logic_vector(3344,24);
            manlo <= conv_std_logic_vector(89464632,28);
      WHEN "0011010010" =>
            manhi <= conv_std_logic_vector(3360,24);
            manlo <= conv_std_logic_vector(90322830,28);
      WHEN "0011010011" =>
            manhi <= conv_std_logic_vector(3376,24);
            manlo <= conv_std_logic_vector(91185124,28);
      WHEN "0011010100" =>
            manhi <= conv_std_logic_vector(3392,24);
            manlo <= conv_std_logic_vector(92051516,28);
      WHEN "0011010101" =>
            manhi <= conv_std_logic_vector(3408,24);
            manlo <= conv_std_logic_vector(92922004,28);
      WHEN "0011010110" =>
            manhi <= conv_std_logic_vector(3424,24);
            manlo <= conv_std_logic_vector(93796589,28);
      WHEN "0011010111" =>
            manhi <= conv_std_logic_vector(3440,24);
            manlo <= conv_std_logic_vector(94675271,28);
      WHEN "0011011000" =>
            manhi <= conv_std_logic_vector(3456,24);
            manlo <= conv_std_logic_vector(95558049,28);
      WHEN "0011011001" =>
            manhi <= conv_std_logic_vector(3472,24);
            manlo <= conv_std_logic_vector(96444925,28);
      WHEN "0011011010" =>
            manhi <= conv_std_logic_vector(3488,24);
            manlo <= conv_std_logic_vector(97335897,28);
      WHEN "0011011011" =>
            manhi <= conv_std_logic_vector(3504,24);
            manlo <= conv_std_logic_vector(98230967,28);
      WHEN "0011011100" =>
            manhi <= conv_std_logic_vector(3520,24);
            manlo <= conv_std_logic_vector(99130133,28);
      WHEN "0011011101" =>
            manhi <= conv_std_logic_vector(3536,24);
            manlo <= conv_std_logic_vector(100033396,28);
      WHEN "0011011110" =>
            manhi <= conv_std_logic_vector(3552,24);
            manlo <= conv_std_logic_vector(100940755,28);
      WHEN "0011011111" =>
            manhi <= conv_std_logic_vector(3568,24);
            manlo <= conv_std_logic_vector(101852212,28);
      WHEN "0011100000" =>
            manhi <= conv_std_logic_vector(3584,24);
            manlo <= conv_std_logic_vector(102767766,28);
      WHEN "0011100001" =>
            manhi <= conv_std_logic_vector(3600,24);
            manlo <= conv_std_logic_vector(103687416,28);
      WHEN "0011100010" =>
            manhi <= conv_std_logic_vector(3616,24);
            manlo <= conv_std_logic_vector(104611163,28);
      WHEN "0011100011" =>
            manhi <= conv_std_logic_vector(3632,24);
            manlo <= conv_std_logic_vector(105539008,28);
      WHEN "0011100100" =>
            manhi <= conv_std_logic_vector(3648,24);
            manlo <= conv_std_logic_vector(106470949,28);
      WHEN "0011100101" =>
            manhi <= conv_std_logic_vector(3664,24);
            manlo <= conv_std_logic_vector(107406987,28);
      WHEN "0011100110" =>
            manhi <= conv_std_logic_vector(3680,24);
            manlo <= conv_std_logic_vector(108347122,28);
      WHEN "0011100111" =>
            manhi <= conv_std_logic_vector(3696,24);
            manlo <= conv_std_logic_vector(109291353,28);
      WHEN "0011101000" =>
            manhi <= conv_std_logic_vector(3712,24);
            manlo <= conv_std_logic_vector(110239682,28);
      WHEN "0011101001" =>
            manhi <= conv_std_logic_vector(3728,24);
            manlo <= conv_std_logic_vector(111192108,28);
      WHEN "0011101010" =>
            manhi <= conv_std_logic_vector(3744,24);
            manlo <= conv_std_logic_vector(112148630,28);
      WHEN "0011101011" =>
            manhi <= conv_std_logic_vector(3760,24);
            manlo <= conv_std_logic_vector(113109250,28);
      WHEN "0011101100" =>
            manhi <= conv_std_logic_vector(3776,24);
            manlo <= conv_std_logic_vector(114073966,28);
      WHEN "0011101101" =>
            manhi <= conv_std_logic_vector(3792,24);
            manlo <= conv_std_logic_vector(115042779,28);
      WHEN "0011101110" =>
            manhi <= conv_std_logic_vector(3808,24);
            manlo <= conv_std_logic_vector(116015689,28);
      WHEN "0011101111" =>
            manhi <= conv_std_logic_vector(3824,24);
            manlo <= conv_std_logic_vector(116992696,28);
      WHEN "0011110000" =>
            manhi <= conv_std_logic_vector(3840,24);
            manlo <= conv_std_logic_vector(117973801,28);
      WHEN "0011110001" =>
            manhi <= conv_std_logic_vector(3856,24);
            manlo <= conv_std_logic_vector(118959001,28);
      WHEN "0011110010" =>
            manhi <= conv_std_logic_vector(3872,24);
            manlo <= conv_std_logic_vector(119948299,28);
      WHEN "0011110011" =>
            manhi <= conv_std_logic_vector(3888,24);
            manlo <= conv_std_logic_vector(120941694,28);
      WHEN "0011110100" =>
            manhi <= conv_std_logic_vector(3904,24);
            manlo <= conv_std_logic_vector(121939186,28);
      WHEN "0011110101" =>
            manhi <= conv_std_logic_vector(3920,24);
            manlo <= conv_std_logic_vector(122940775,28);
      WHEN "0011110110" =>
            manhi <= conv_std_logic_vector(3936,24);
            manlo <= conv_std_logic_vector(123946461,28);
      WHEN "0011110111" =>
            manhi <= conv_std_logic_vector(3952,24);
            manlo <= conv_std_logic_vector(124956243,28);
      WHEN "0011111000" =>
            manhi <= conv_std_logic_vector(3968,24);
            manlo <= conv_std_logic_vector(125970123,28);
      WHEN "0011111001" =>
            manhi <= conv_std_logic_vector(3984,24);
            manlo <= conv_std_logic_vector(126988100,28);
      WHEN "0011111010" =>
            manhi <= conv_std_logic_vector(4000,24);
            manlo <= conv_std_logic_vector(128010173,28);
      WHEN "0011111011" =>
            manhi <= conv_std_logic_vector(4016,24);
            manlo <= conv_std_logic_vector(129036344,28);
      WHEN "0011111100" =>
            manhi <= conv_std_logic_vector(4032,24);
            manlo <= conv_std_logic_vector(130066611,28);
      WHEN "0011111101" =>
            manhi <= conv_std_logic_vector(4048,24);
            manlo <= conv_std_logic_vector(131100976,28);
      WHEN "0011111110" =>
            manhi <= conv_std_logic_vector(4064,24);
            manlo <= conv_std_logic_vector(132139437,28);
      WHEN "0011111111" =>
            manhi <= conv_std_logic_vector(4080,24);
            manlo <= conv_std_logic_vector(133181996,28);
      WHEN "0100000000" =>
            manhi <= conv_std_logic_vector(4096,24);
            manlo <= conv_std_logic_vector(134228651,28);
      WHEN "0100000001" =>
            manhi <= conv_std_logic_vector(4112,24);
            manlo <= conv_std_logic_vector(135279404,28);
      WHEN "0100000010" =>
            manhi <= conv_std_logic_vector(4128,24);
            manlo <= conv_std_logic_vector(136334253,28);
      WHEN "0100000011" =>
            manhi <= conv_std_logic_vector(4144,24);
            manlo <= conv_std_logic_vector(137393200,28);
      WHEN "0100000100" =>
            manhi <= conv_std_logic_vector(4160,24);
            manlo <= conv_std_logic_vector(138456243,28);
      WHEN "0100000101" =>
            manhi <= conv_std_logic_vector(4176,24);
            manlo <= conv_std_logic_vector(139523384,28);
      WHEN "0100000110" =>
            manhi <= conv_std_logic_vector(4192,24);
            manlo <= conv_std_logic_vector(140594622,28);
      WHEN "0100000111" =>
            manhi <= conv_std_logic_vector(4208,24);
            manlo <= conv_std_logic_vector(141669956,28);
      WHEN "0100001000" =>
            manhi <= conv_std_logic_vector(4224,24);
            manlo <= conv_std_logic_vector(142749388,28);
      WHEN "0100001001" =>
            manhi <= conv_std_logic_vector(4240,24);
            manlo <= conv_std_logic_vector(143832916,28);
      WHEN "0100001010" =>
            manhi <= conv_std_logic_vector(4256,24);
            manlo <= conv_std_logic_vector(144920542,28);
      WHEN "0100001011" =>
            manhi <= conv_std_logic_vector(4272,24);
            manlo <= conv_std_logic_vector(146012265,28);
      WHEN "0100001100" =>
            manhi <= conv_std_logic_vector(4288,24);
            manlo <= conv_std_logic_vector(147108085,28);
      WHEN "0100001101" =>
            manhi <= conv_std_logic_vector(4304,24);
            manlo <= conv_std_logic_vector(148208001,28);
      WHEN "0100001110" =>
            manhi <= conv_std_logic_vector(4320,24);
            manlo <= conv_std_logic_vector(149312015,28);
      WHEN "0100001111" =>
            manhi <= conv_std_logic_vector(4336,24);
            manlo <= conv_std_logic_vector(150420126,28);
      WHEN "0100010000" =>
            manhi <= conv_std_logic_vector(4352,24);
            manlo <= conv_std_logic_vector(151532334,28);
      WHEN "0100010001" =>
            manhi <= conv_std_logic_vector(4368,24);
            manlo <= conv_std_logic_vector(152648639,28);
      WHEN "0100010010" =>
            manhi <= conv_std_logic_vector(4384,24);
            manlo <= conv_std_logic_vector(153769041,28);
      WHEN "0100010011" =>
            manhi <= conv_std_logic_vector(4400,24);
            manlo <= conv_std_logic_vector(154893541,28);
      WHEN "0100010100" =>
            manhi <= conv_std_logic_vector(4416,24);
            manlo <= conv_std_logic_vector(156022137,28);
      WHEN "0100010101" =>
            manhi <= conv_std_logic_vector(4432,24);
            manlo <= conv_std_logic_vector(157154830,28);
      WHEN "0100010110" =>
            manhi <= conv_std_logic_vector(4448,24);
            manlo <= conv_std_logic_vector(158291621,28);
      WHEN "0100010111" =>
            manhi <= conv_std_logic_vector(4464,24);
            manlo <= conv_std_logic_vector(159432508,28);
      WHEN "0100011000" =>
            manhi <= conv_std_logic_vector(4480,24);
            manlo <= conv_std_logic_vector(160577493,28);
      WHEN "0100011001" =>
            manhi <= conv_std_logic_vector(4496,24);
            manlo <= conv_std_logic_vector(161726574,28);
      WHEN "0100011010" =>
            manhi <= conv_std_logic_vector(4512,24);
            manlo <= conv_std_logic_vector(162879753,28);
      WHEN "0100011011" =>
            manhi <= conv_std_logic_vector(4528,24);
            manlo <= conv_std_logic_vector(164037029,28);
      WHEN "0100011100" =>
            manhi <= conv_std_logic_vector(4544,24);
            manlo <= conv_std_logic_vector(165198402,28);
      WHEN "0100011101" =>
            manhi <= conv_std_logic_vector(4560,24);
            manlo <= conv_std_logic_vector(166363872,28);
      WHEN "0100011110" =>
            manhi <= conv_std_logic_vector(4576,24);
            manlo <= conv_std_logic_vector(167533439,28);
      WHEN "0100011111" =>
            manhi <= conv_std_logic_vector(4592,24);
            manlo <= conv_std_logic_vector(168707104,28);
      WHEN "0100100000" =>
            manhi <= conv_std_logic_vector(4608,24);
            manlo <= conv_std_logic_vector(169884865,28);
      WHEN "0100100001" =>
            manhi <= conv_std_logic_vector(4624,24);
            manlo <= conv_std_logic_vector(171066724,28);
      WHEN "0100100010" =>
            manhi <= conv_std_logic_vector(4640,24);
            manlo <= conv_std_logic_vector(172252679,28);
      WHEN "0100100011" =>
            manhi <= conv_std_logic_vector(4656,24);
            manlo <= conv_std_logic_vector(173442732,28);
      WHEN "0100100100" =>
            manhi <= conv_std_logic_vector(4672,24);
            manlo <= conv_std_logic_vector(174636882,28);
      WHEN "0100100101" =>
            manhi <= conv_std_logic_vector(4688,24);
            manlo <= conv_std_logic_vector(175835129,28);
      WHEN "0100100110" =>
            manhi <= conv_std_logic_vector(4704,24);
            manlo <= conv_std_logic_vector(177037474,28);
      WHEN "0100100111" =>
            manhi <= conv_std_logic_vector(4720,24);
            manlo <= conv_std_logic_vector(178243915,28);
      WHEN "0100101000" =>
            manhi <= conv_std_logic_vector(4736,24);
            manlo <= conv_std_logic_vector(179454454,28);
      WHEN "0100101001" =>
            manhi <= conv_std_logic_vector(4752,24);
            manlo <= conv_std_logic_vector(180669089,28);
      WHEN "0100101010" =>
            manhi <= conv_std_logic_vector(4768,24);
            manlo <= conv_std_logic_vector(181887822,28);
      WHEN "0100101011" =>
            manhi <= conv_std_logic_vector(4784,24);
            manlo <= conv_std_logic_vector(183110652,28);
      WHEN "0100101100" =>
            manhi <= conv_std_logic_vector(4800,24);
            manlo <= conv_std_logic_vector(184337579,28);
      WHEN "0100101101" =>
            manhi <= conv_std_logic_vector(4816,24);
            manlo <= conv_std_logic_vector(185568604,28);
      WHEN "0100101110" =>
            manhi <= conv_std_logic_vector(4832,24);
            manlo <= conv_std_logic_vector(186803725,28);
      WHEN "0100101111" =>
            manhi <= conv_std_logic_vector(4848,24);
            manlo <= conv_std_logic_vector(188042944,28);
      WHEN "0100110000" =>
            manhi <= conv_std_logic_vector(4864,24);
            manlo <= conv_std_logic_vector(189286260,28);
      WHEN "0100110001" =>
            manhi <= conv_std_logic_vector(4880,24);
            manlo <= conv_std_logic_vector(190533673,28);
      WHEN "0100110010" =>
            manhi <= conv_std_logic_vector(4896,24);
            manlo <= conv_std_logic_vector(191785183,28);
      WHEN "0100110011" =>
            manhi <= conv_std_logic_vector(4912,24);
            manlo <= conv_std_logic_vector(193040791,28);
      WHEN "0100110100" =>
            manhi <= conv_std_logic_vector(4928,24);
            manlo <= conv_std_logic_vector(194300496,28);
      WHEN "0100110101" =>
            manhi <= conv_std_logic_vector(4944,24);
            manlo <= conv_std_logic_vector(195564298,28);
      WHEN "0100110110" =>
            manhi <= conv_std_logic_vector(4960,24);
            manlo <= conv_std_logic_vector(196832197,28);
      WHEN "0100110111" =>
            manhi <= conv_std_logic_vector(4976,24);
            manlo <= conv_std_logic_vector(198104193,28);
      WHEN "0100111000" =>
            manhi <= conv_std_logic_vector(4992,24);
            manlo <= conv_std_logic_vector(199380286,28);
      WHEN "0100111001" =>
            manhi <= conv_std_logic_vector(5008,24);
            manlo <= conv_std_logic_vector(200660477,28);
      WHEN "0100111010" =>
            manhi <= conv_std_logic_vector(5024,24);
            manlo <= conv_std_logic_vector(201944765,28);
      WHEN "0100111011" =>
            manhi <= conv_std_logic_vector(5040,24);
            manlo <= conv_std_logic_vector(203233150,28);
      WHEN "0100111100" =>
            manhi <= conv_std_logic_vector(5056,24);
            manlo <= conv_std_logic_vector(204525633,28);
      WHEN "0100111101" =>
            manhi <= conv_std_logic_vector(5072,24);
            manlo <= conv_std_logic_vector(205822213,28);
      WHEN "0100111110" =>
            manhi <= conv_std_logic_vector(5088,24);
            manlo <= conv_std_logic_vector(207122889,28);
      WHEN "0100111111" =>
            manhi <= conv_std_logic_vector(5104,24);
            manlo <= conv_std_logic_vector(208427664,28);
      WHEN "0101000000" =>
            manhi <= conv_std_logic_vector(5120,24);
            manlo <= conv_std_logic_vector(209736535,28);
      WHEN "0101000001" =>
            manhi <= conv_std_logic_vector(5136,24);
            manlo <= conv_std_logic_vector(211049504,28);
      WHEN "0101000010" =>
            manhi <= conv_std_logic_vector(5152,24);
            manlo <= conv_std_logic_vector(212366570,28);
      WHEN "0101000011" =>
            manhi <= conv_std_logic_vector(5168,24);
            manlo <= conv_std_logic_vector(213687733,28);
      WHEN "0101000100" =>
            manhi <= conv_std_logic_vector(5184,24);
            manlo <= conv_std_logic_vector(215012993,28);
      WHEN "0101000101" =>
            manhi <= conv_std_logic_vector(5200,24);
            manlo <= conv_std_logic_vector(216342351,28);
      WHEN "0101000110" =>
            manhi <= conv_std_logic_vector(5216,24);
            manlo <= conv_std_logic_vector(217675806,28);
      WHEN "0101000111" =>
            manhi <= conv_std_logic_vector(5232,24);
            manlo <= conv_std_logic_vector(219013358,28);
      WHEN "0101001000" =>
            manhi <= conv_std_logic_vector(5248,24);
            manlo <= conv_std_logic_vector(220355007,28);
      WHEN "0101001001" =>
            manhi <= conv_std_logic_vector(5264,24);
            manlo <= conv_std_logic_vector(221700754,28);
      WHEN "0101001010" =>
            manhi <= conv_std_logic_vector(5280,24);
            manlo <= conv_std_logic_vector(223050598,28);
      WHEN "0101001011" =>
            manhi <= conv_std_logic_vector(5296,24);
            manlo <= conv_std_logic_vector(224404540,28);
      WHEN "0101001100" =>
            manhi <= conv_std_logic_vector(5312,24);
            manlo <= conv_std_logic_vector(225762578,28);
      WHEN "0101001101" =>
            manhi <= conv_std_logic_vector(5328,24);
            manlo <= conv_std_logic_vector(227124714,28);
      WHEN "0101001110" =>
            manhi <= conv_std_logic_vector(5344,24);
            manlo <= conv_std_logic_vector(228490948,28);
      WHEN "0101001111" =>
            manhi <= conv_std_logic_vector(5360,24);
            manlo <= conv_std_logic_vector(229861278,28);
      WHEN "0101010000" =>
            manhi <= conv_std_logic_vector(5376,24);
            manlo <= conv_std_logic_vector(231235706,28);
      WHEN "0101010001" =>
            manhi <= conv_std_logic_vector(5392,24);
            manlo <= conv_std_logic_vector(232614231,28);
      WHEN "0101010010" =>
            manhi <= conv_std_logic_vector(5408,24);
            manlo <= conv_std_logic_vector(233996854,28);
      WHEN "0101010011" =>
            manhi <= conv_std_logic_vector(5424,24);
            manlo <= conv_std_logic_vector(235383573,28);
      WHEN "0101010100" =>
            manhi <= conv_std_logic_vector(5440,24);
            manlo <= conv_std_logic_vector(236774391,28);
      WHEN "0101010101" =>
            manhi <= conv_std_logic_vector(5456,24);
            manlo <= conv_std_logic_vector(238169305,28);
      WHEN "0101010110" =>
            manhi <= conv_std_logic_vector(5472,24);
            manlo <= conv_std_logic_vector(239568317,28);
      WHEN "0101010111" =>
            manhi <= conv_std_logic_vector(5488,24);
            manlo <= conv_std_logic_vector(240971426,28);
      WHEN "0101011000" =>
            manhi <= conv_std_logic_vector(5504,24);
            manlo <= conv_std_logic_vector(242378633,28);
      WHEN "0101011001" =>
            manhi <= conv_std_logic_vector(5520,24);
            manlo <= conv_std_logic_vector(243789936,28);
      WHEN "0101011010" =>
            manhi <= conv_std_logic_vector(5536,24);
            manlo <= conv_std_logic_vector(245205338,28);
      WHEN "0101011011" =>
            manhi <= conv_std_logic_vector(5552,24);
            manlo <= conv_std_logic_vector(246624836,28);
      WHEN "0101011100" =>
            manhi <= conv_std_logic_vector(5568,24);
            manlo <= conv_std_logic_vector(248048432,28);
      WHEN "0101011101" =>
            manhi <= conv_std_logic_vector(5584,24);
            manlo <= conv_std_logic_vector(249476125,28);
      WHEN "0101011110" =>
            manhi <= conv_std_logic_vector(5600,24);
            manlo <= conv_std_logic_vector(250907916,28);
      WHEN "0101011111" =>
            manhi <= conv_std_logic_vector(5616,24);
            manlo <= conv_std_logic_vector(252343804,28);
      WHEN "0101100000" =>
            manhi <= conv_std_logic_vector(5632,24);
            manlo <= conv_std_logic_vector(253783789,28);
      WHEN "0101100001" =>
            manhi <= conv_std_logic_vector(5648,24);
            manlo <= conv_std_logic_vector(255227872,28);
      WHEN "0101100010" =>
            manhi <= conv_std_logic_vector(5664,24);
            manlo <= conv_std_logic_vector(256676052,28);
      WHEN "0101100011" =>
            manhi <= conv_std_logic_vector(5680,24);
            manlo <= conv_std_logic_vector(258128329,28);
      WHEN "0101100100" =>
            manhi <= conv_std_logic_vector(5696,24);
            manlo <= conv_std_logic_vector(259584704,28);
      WHEN "0101100101" =>
            manhi <= conv_std_logic_vector(5712,24);
            manlo <= conv_std_logic_vector(261045176,28);
      WHEN "0101100110" =>
            manhi <= conv_std_logic_vector(5728,24);
            manlo <= conv_std_logic_vector(262509746,28);
      WHEN "0101100111" =>
            manhi <= conv_std_logic_vector(5744,24);
            manlo <= conv_std_logic_vector(263978413,28);
      WHEN "0101101000" =>
            manhi <= conv_std_logic_vector(5760,24);
            manlo <= conv_std_logic_vector(265451178,28);
      WHEN "0101101001" =>
            manhi <= conv_std_logic_vector(5776,24);
            manlo <= conv_std_logic_vector(266928039,28);
      WHEN "0101101010" =>
            manhi <= conv_std_logic_vector(5792,24);
            manlo <= conv_std_logic_vector(268408999,28);
      WHEN "0101101011" =>
            manhi <= conv_std_logic_vector(5809,24);
            manlo <= conv_std_logic_vector(1458599,28);
      WHEN "0101101100" =>
            manhi <= conv_std_logic_vector(5825,24);
            manlo <= conv_std_logic_vector(2947754,28);
      WHEN "0101101101" =>
            manhi <= conv_std_logic_vector(5841,24);
            manlo <= conv_std_logic_vector(4441005,28);
      WHEN "0101101110" =>
            manhi <= conv_std_logic_vector(5857,24);
            manlo <= conv_std_logic_vector(5938354,28);
      WHEN "0101101111" =>
            manhi <= conv_std_logic_vector(5873,24);
            manlo <= conv_std_logic_vector(7439800,28);
      WHEN "0101110000" =>
            manhi <= conv_std_logic_vector(5889,24);
            manlo <= conv_std_logic_vector(8945344,28);
      WHEN "0101110001" =>
            manhi <= conv_std_logic_vector(5905,24);
            manlo <= conv_std_logic_vector(10454985,28);
      WHEN "0101110010" =>
            manhi <= conv_std_logic_vector(5921,24);
            manlo <= conv_std_logic_vector(11968724,28);
      WHEN "0101110011" =>
            manhi <= conv_std_logic_vector(5937,24);
            manlo <= conv_std_logic_vector(13486560,28);
      WHEN "0101110100" =>
            manhi <= conv_std_logic_vector(5953,24);
            manlo <= conv_std_logic_vector(15008494,28);
      WHEN "0101110101" =>
            manhi <= conv_std_logic_vector(5969,24);
            manlo <= conv_std_logic_vector(16534525,28);
      WHEN "0101110110" =>
            manhi <= conv_std_logic_vector(5985,24);
            manlo <= conv_std_logic_vector(18064653,28);
      WHEN "0101110111" =>
            manhi <= conv_std_logic_vector(6001,24);
            manlo <= conv_std_logic_vector(19598879,28);
      WHEN "0101111000" =>
            manhi <= conv_std_logic_vector(6017,24);
            manlo <= conv_std_logic_vector(21137203,28);
      WHEN "0101111001" =>
            manhi <= conv_std_logic_vector(6033,24);
            manlo <= conv_std_logic_vector(22679624,28);
      WHEN "0101111010" =>
            manhi <= conv_std_logic_vector(6049,24);
            manlo <= conv_std_logic_vector(24226142,28);
      WHEN "0101111011" =>
            manhi <= conv_std_logic_vector(6065,24);
            manlo <= conv_std_logic_vector(25776758,28);
      WHEN "0101111100" =>
            manhi <= conv_std_logic_vector(6081,24);
            manlo <= conv_std_logic_vector(27331471,28);
      WHEN "0101111101" =>
            manhi <= conv_std_logic_vector(6097,24);
            manlo <= conv_std_logic_vector(28890282,28);
      WHEN "0101111110" =>
            manhi <= conv_std_logic_vector(6113,24);
            manlo <= conv_std_logic_vector(30453190,28);
      WHEN "0101111111" =>
            manhi <= conv_std_logic_vector(6129,24);
            manlo <= conv_std_logic_vector(32020196,28);
      WHEN "0110000000" =>
            manhi <= conv_std_logic_vector(6145,24);
            manlo <= conv_std_logic_vector(33591299,28);
      WHEN "0110000001" =>
            manhi <= conv_std_logic_vector(6161,24);
            manlo <= conv_std_logic_vector(35166500,28);
      WHEN "0110000010" =>
            manhi <= conv_std_logic_vector(6177,24);
            manlo <= conv_std_logic_vector(36745798,28);
      WHEN "0110000011" =>
            manhi <= conv_std_logic_vector(6193,24);
            manlo <= conv_std_logic_vector(38329194,28);
      WHEN "0110000100" =>
            manhi <= conv_std_logic_vector(6209,24);
            manlo <= conv_std_logic_vector(39916688,28);
      WHEN "0110000101" =>
            manhi <= conv_std_logic_vector(6225,24);
            manlo <= conv_std_logic_vector(41508278,28);
      WHEN "0110000110" =>
            manhi <= conv_std_logic_vector(6241,24);
            manlo <= conv_std_logic_vector(43103967,28);
      WHEN "0110000111" =>
            manhi <= conv_std_logic_vector(6257,24);
            manlo <= conv_std_logic_vector(44703753,28);
      WHEN "0110001000" =>
            manhi <= conv_std_logic_vector(6273,24);
            manlo <= conv_std_logic_vector(46307636,28);
      WHEN "0110001001" =>
            manhi <= conv_std_logic_vector(6289,24);
            manlo <= conv_std_logic_vector(47915617,28);
      WHEN "0110001010" =>
            manhi <= conv_std_logic_vector(6305,24);
            manlo <= conv_std_logic_vector(49527695,28);
      WHEN "0110001011" =>
            manhi <= conv_std_logic_vector(6321,24);
            manlo <= conv_std_logic_vector(51143871,28);
      WHEN "0110001100" =>
            manhi <= conv_std_logic_vector(6337,24);
            manlo <= conv_std_logic_vector(52764145,28);
      WHEN "0110001101" =>
            manhi <= conv_std_logic_vector(6353,24);
            manlo <= conv_std_logic_vector(54388516,28);
      WHEN "0110001110" =>
            manhi <= conv_std_logic_vector(6369,24);
            manlo <= conv_std_logic_vector(56016985,28);
      WHEN "0110001111" =>
            manhi <= conv_std_logic_vector(6385,24);
            manlo <= conv_std_logic_vector(57649551,28);
      WHEN "0110010000" =>
            manhi <= conv_std_logic_vector(6401,24);
            manlo <= conv_std_logic_vector(59286215,28);
      WHEN "0110010001" =>
            manhi <= conv_std_logic_vector(6417,24);
            manlo <= conv_std_logic_vector(60926976,28);
      WHEN "0110010010" =>
            manhi <= conv_std_logic_vector(6433,24);
            manlo <= conv_std_logic_vector(62571835,28);
      WHEN "0110010011" =>
            manhi <= conv_std_logic_vector(6449,24);
            manlo <= conv_std_logic_vector(64220791,28);
      WHEN "0110010100" =>
            manhi <= conv_std_logic_vector(6465,24);
            manlo <= conv_std_logic_vector(65873845,28);
      WHEN "0110010101" =>
            manhi <= conv_std_logic_vector(6481,24);
            manlo <= conv_std_logic_vector(67530997,28);
      WHEN "0110010110" =>
            manhi <= conv_std_logic_vector(6497,24);
            manlo <= conv_std_logic_vector(69192246,28);
      WHEN "0110010111" =>
            manhi <= conv_std_logic_vector(6513,24);
            manlo <= conv_std_logic_vector(70857593,28);
      WHEN "0110011000" =>
            manhi <= conv_std_logic_vector(6529,24);
            manlo <= conv_std_logic_vector(72527037,28);
      WHEN "0110011001" =>
            manhi <= conv_std_logic_vector(6545,24);
            manlo <= conv_std_logic_vector(74200579,28);
      WHEN "0110011010" =>
            manhi <= conv_std_logic_vector(6561,24);
            manlo <= conv_std_logic_vector(75878219,28);
      WHEN "0110011011" =>
            manhi <= conv_std_logic_vector(6577,24);
            manlo <= conv_std_logic_vector(77559956,28);
      WHEN "0110011100" =>
            manhi <= conv_std_logic_vector(6593,24);
            manlo <= conv_std_logic_vector(79245791,28);
      WHEN "0110011101" =>
            manhi <= conv_std_logic_vector(6609,24);
            manlo <= conv_std_logic_vector(80935723,28);
      WHEN "0110011110" =>
            manhi <= conv_std_logic_vector(6625,24);
            manlo <= conv_std_logic_vector(82629753,28);
      WHEN "0110011111" =>
            manhi <= conv_std_logic_vector(6641,24);
            manlo <= conv_std_logic_vector(84327881,28);
      WHEN "0110100000" =>
            manhi <= conv_std_logic_vector(6657,24);
            manlo <= conv_std_logic_vector(86030106,28);
      WHEN "0110100001" =>
            manhi <= conv_std_logic_vector(6673,24);
            manlo <= conv_std_logic_vector(87736429,28);
      WHEN "0110100010" =>
            manhi <= conv_std_logic_vector(6689,24);
            manlo <= conv_std_logic_vector(89446849,28);
      WHEN "0110100011" =>
            manhi <= conv_std_logic_vector(6705,24);
            manlo <= conv_std_logic_vector(91161367,28);
      WHEN "0110100100" =>
            manhi <= conv_std_logic_vector(6721,24);
            manlo <= conv_std_logic_vector(92879983,28);
      WHEN "0110100101" =>
            manhi <= conv_std_logic_vector(6737,24);
            manlo <= conv_std_logic_vector(94602697,28);
      WHEN "0110100110" =>
            manhi <= conv_std_logic_vector(6753,24);
            manlo <= conv_std_logic_vector(96329508,28);
      WHEN "0110100111" =>
            manhi <= conv_std_logic_vector(6769,24);
            manlo <= conv_std_logic_vector(98060416,28);
      WHEN "0110101000" =>
            manhi <= conv_std_logic_vector(6785,24);
            manlo <= conv_std_logic_vector(99795423,28);
      WHEN "0110101001" =>
            manhi <= conv_std_logic_vector(6801,24);
            manlo <= conv_std_logic_vector(101534527,28);
      WHEN "0110101010" =>
            manhi <= conv_std_logic_vector(6817,24);
            manlo <= conv_std_logic_vector(103277728,28);
      WHEN "0110101011" =>
            manhi <= conv_std_logic_vector(6833,24);
            manlo <= conv_std_logic_vector(105025028,28);
      WHEN "0110101100" =>
            manhi <= conv_std_logic_vector(6849,24);
            manlo <= conv_std_logic_vector(106776425,28);
      WHEN "0110101101" =>
            manhi <= conv_std_logic_vector(6865,24);
            manlo <= conv_std_logic_vector(108531919,28);
      WHEN "0110101110" =>
            manhi <= conv_std_logic_vector(6881,24);
            manlo <= conv_std_logic_vector(110291512,28);
      WHEN "0110101111" =>
            manhi <= conv_std_logic_vector(6897,24);
            manlo <= conv_std_logic_vector(112055202,28);
      WHEN "0110110000" =>
            manhi <= conv_std_logic_vector(6913,24);
            manlo <= conv_std_logic_vector(113822989,28);
      WHEN "0110110001" =>
            manhi <= conv_std_logic_vector(6929,24);
            manlo <= conv_std_logic_vector(115594875,28);
      WHEN "0110110010" =>
            manhi <= conv_std_logic_vector(6945,24);
            manlo <= conv_std_logic_vector(117370858,28);
      WHEN "0110110011" =>
            manhi <= conv_std_logic_vector(6961,24);
            manlo <= conv_std_logic_vector(119150939,28);
      WHEN "0110110100" =>
            manhi <= conv_std_logic_vector(6977,24);
            manlo <= conv_std_logic_vector(120935117,28);
      WHEN "0110110101" =>
            manhi <= conv_std_logic_vector(6993,24);
            manlo <= conv_std_logic_vector(122723393,28);
      WHEN "0110110110" =>
            manhi <= conv_std_logic_vector(7009,24);
            manlo <= conv_std_logic_vector(124515767,28);
      WHEN "0110110111" =>
            manhi <= conv_std_logic_vector(7025,24);
            manlo <= conv_std_logic_vector(126312239,28);
      WHEN "0110111000" =>
            manhi <= conv_std_logic_vector(7041,24);
            manlo <= conv_std_logic_vector(128112808,28);
      WHEN "0110111001" =>
            manhi <= conv_std_logic_vector(7057,24);
            manlo <= conv_std_logic_vector(129917475,28);
      WHEN "0110111010" =>
            manhi <= conv_std_logic_vector(7073,24);
            manlo <= conv_std_logic_vector(131726240,28);
      WHEN "0110111011" =>
            manhi <= conv_std_logic_vector(7089,24);
            manlo <= conv_std_logic_vector(133539102,28);
      WHEN "0110111100" =>
            manhi <= conv_std_logic_vector(7105,24);
            manlo <= conv_std_logic_vector(135356063,28);
      WHEN "0110111101" =>
            manhi <= conv_std_logic_vector(7121,24);
            manlo <= conv_std_logic_vector(137177121,28);
      WHEN "0110111110" =>
            manhi <= conv_std_logic_vector(7137,24);
            manlo <= conv_std_logic_vector(139002276,28);
      WHEN "0110111111" =>
            manhi <= conv_std_logic_vector(7153,24);
            manlo <= conv_std_logic_vector(140831530,28);
      WHEN "0111000000" =>
            manhi <= conv_std_logic_vector(7169,24);
            manlo <= conv_std_logic_vector(142664881,28);
      WHEN "0111000001" =>
            manhi <= conv_std_logic_vector(7185,24);
            manlo <= conv_std_logic_vector(144502330,28);
      WHEN "0111000010" =>
            manhi <= conv_std_logic_vector(7201,24);
            manlo <= conv_std_logic_vector(146343877,28);
      WHEN "0111000011" =>
            manhi <= conv_std_logic_vector(7217,24);
            manlo <= conv_std_logic_vector(148189521,28);
      WHEN "0111000100" =>
            manhi <= conv_std_logic_vector(7233,24);
            manlo <= conv_std_logic_vector(150039263,28);
      WHEN "0111000101" =>
            manhi <= conv_std_logic_vector(7249,24);
            manlo <= conv_std_logic_vector(151893103,28);
      WHEN "0111000110" =>
            manhi <= conv_std_logic_vector(7265,24);
            manlo <= conv_std_logic_vector(153751041,28);
      WHEN "0111000111" =>
            manhi <= conv_std_logic_vector(7281,24);
            manlo <= conv_std_logic_vector(155613076,28);
      WHEN "0111001000" =>
            manhi <= conv_std_logic_vector(7297,24);
            manlo <= conv_std_logic_vector(157479210,28);
      WHEN "0111001001" =>
            manhi <= conv_std_logic_vector(7313,24);
            manlo <= conv_std_logic_vector(159349441,28);
      WHEN "0111001010" =>
            manhi <= conv_std_logic_vector(7329,24);
            manlo <= conv_std_logic_vector(161223770,28);
      WHEN "0111001011" =>
            manhi <= conv_std_logic_vector(7345,24);
            manlo <= conv_std_logic_vector(163102196,28);
      WHEN "0111001100" =>
            manhi <= conv_std_logic_vector(7361,24);
            manlo <= conv_std_logic_vector(164984721,28);
      WHEN "0111001101" =>
            manhi <= conv_std_logic_vector(7377,24);
            manlo <= conv_std_logic_vector(166871343,28);
      WHEN "0111001110" =>
            manhi <= conv_std_logic_vector(7393,24);
            manlo <= conv_std_logic_vector(168762063,28);
      WHEN "0111001111" =>
            manhi <= conv_std_logic_vector(7409,24);
            manlo <= conv_std_logic_vector(170656881,28);
      WHEN "0111010000" =>
            manhi <= conv_std_logic_vector(7425,24);
            manlo <= conv_std_logic_vector(172555797,28);
      WHEN "0111010001" =>
            manhi <= conv_std_logic_vector(7441,24);
            manlo <= conv_std_logic_vector(174458810,28);
      WHEN "0111010010" =>
            manhi <= conv_std_logic_vector(7457,24);
            manlo <= conv_std_logic_vector(176365921,28);
      WHEN "0111010011" =>
            manhi <= conv_std_logic_vector(7473,24);
            manlo <= conv_std_logic_vector(178277130,28);
      WHEN "0111010100" =>
            manhi <= conv_std_logic_vector(7489,24);
            manlo <= conv_std_logic_vector(180192437,28);
      WHEN "0111010101" =>
            manhi <= conv_std_logic_vector(7505,24);
            manlo <= conv_std_logic_vector(182111842,28);
      WHEN "0111010110" =>
            manhi <= conv_std_logic_vector(7521,24);
            manlo <= conv_std_logic_vector(184035345,28);
      WHEN "0111010111" =>
            manhi <= conv_std_logic_vector(7537,24);
            manlo <= conv_std_logic_vector(185962945,28);
      WHEN "0111011000" =>
            manhi <= conv_std_logic_vector(7553,24);
            manlo <= conv_std_logic_vector(187894643,28);
      WHEN "0111011001" =>
            manhi <= conv_std_logic_vector(7569,24);
            manlo <= conv_std_logic_vector(189830439,28);
      WHEN "0111011010" =>
            manhi <= conv_std_logic_vector(7585,24);
            manlo <= conv_std_logic_vector(191770333,28);
      WHEN "0111011011" =>
            manhi <= conv_std_logic_vector(7601,24);
            manlo <= conv_std_logic_vector(193714325,28);
      WHEN "0111011100" =>
            manhi <= conv_std_logic_vector(7617,24);
            manlo <= conv_std_logic_vector(195662415,28);
      WHEN "0111011101" =>
            manhi <= conv_std_logic_vector(7633,24);
            manlo <= conv_std_logic_vector(197614602,28);
      WHEN "0111011110" =>
            manhi <= conv_std_logic_vector(7649,24);
            manlo <= conv_std_logic_vector(199570888,28);
      WHEN "0111011111" =>
            manhi <= conv_std_logic_vector(7665,24);
            manlo <= conv_std_logic_vector(201531271,28);
      WHEN "0111100000" =>
            manhi <= conv_std_logic_vector(7681,24);
            manlo <= conv_std_logic_vector(203495752,28);
      WHEN "0111100001" =>
            manhi <= conv_std_logic_vector(7697,24);
            manlo <= conv_std_logic_vector(205464331,28);
      WHEN "0111100010" =>
            manhi <= conv_std_logic_vector(7713,24);
            manlo <= conv_std_logic_vector(207437008,28);
      WHEN "0111100011" =>
            manhi <= conv_std_logic_vector(7729,24);
            manlo <= conv_std_logic_vector(209413783,28);
      WHEN "0111100100" =>
            manhi <= conv_std_logic_vector(7745,24);
            manlo <= conv_std_logic_vector(211394656,28);
      WHEN "0111100101" =>
            manhi <= conv_std_logic_vector(7761,24);
            manlo <= conv_std_logic_vector(213379626,28);
      WHEN "0111100110" =>
            manhi <= conv_std_logic_vector(7777,24);
            manlo <= conv_std_logic_vector(215368695,28);
      WHEN "0111100111" =>
            manhi <= conv_std_logic_vector(7793,24);
            manlo <= conv_std_logic_vector(217361861,28);
      WHEN "0111101000" =>
            manhi <= conv_std_logic_vector(7809,24);
            manlo <= conv_std_logic_vector(219359125,28);
      WHEN "0111101001" =>
            manhi <= conv_std_logic_vector(7825,24);
            manlo <= conv_std_logic_vector(221360487,28);
      WHEN "0111101010" =>
            manhi <= conv_std_logic_vector(7841,24);
            manlo <= conv_std_logic_vector(223365947,28);
      WHEN "0111101011" =>
            manhi <= conv_std_logic_vector(7857,24);
            manlo <= conv_std_logic_vector(225375505,28);
      WHEN "0111101100" =>
            manhi <= conv_std_logic_vector(7873,24);
            manlo <= conv_std_logic_vector(227389161,28);
      WHEN "0111101101" =>
            manhi <= conv_std_logic_vector(7889,24);
            manlo <= conv_std_logic_vector(229406915,28);
      WHEN "0111101110" =>
            manhi <= conv_std_logic_vector(7905,24);
            manlo <= conv_std_logic_vector(231428767,28);
      WHEN "0111101111" =>
            manhi <= conv_std_logic_vector(7921,24);
            manlo <= conv_std_logic_vector(233454716,28);
      WHEN "0111110000" =>
            manhi <= conv_std_logic_vector(7937,24);
            manlo <= conv_std_logic_vector(235484764,28);
      WHEN "0111110001" =>
            manhi <= conv_std_logic_vector(7953,24);
            manlo <= conv_std_logic_vector(237518910,28);
      WHEN "0111110010" =>
            manhi <= conv_std_logic_vector(7969,24);
            manlo <= conv_std_logic_vector(239557153,28);
      WHEN "0111110011" =>
            manhi <= conv_std_logic_vector(7985,24);
            manlo <= conv_std_logic_vector(241599495,28);
      WHEN "0111110100" =>
            manhi <= conv_std_logic_vector(8001,24);
            manlo <= conv_std_logic_vector(243645934,28);
      WHEN "0111110101" =>
            manhi <= conv_std_logic_vector(8017,24);
            manlo <= conv_std_logic_vector(245696471,28);
      WHEN "0111110110" =>
            manhi <= conv_std_logic_vector(8033,24);
            manlo <= conv_std_logic_vector(247751107,28);
      WHEN "0111110111" =>
            manhi <= conv_std_logic_vector(8049,24);
            manlo <= conv_std_logic_vector(249809840,28);
      WHEN "0111111000" =>
            manhi <= conv_std_logic_vector(8065,24);
            manlo <= conv_std_logic_vector(251872671,28);
      WHEN "0111111001" =>
            manhi <= conv_std_logic_vector(8081,24);
            manlo <= conv_std_logic_vector(253939600,28);
      WHEN "0111111010" =>
            manhi <= conv_std_logic_vector(8097,24);
            manlo <= conv_std_logic_vector(256010627,28);
      WHEN "0111111011" =>
            manhi <= conv_std_logic_vector(8113,24);
            manlo <= conv_std_logic_vector(258085753,28);
      WHEN "0111111100" =>
            manhi <= conv_std_logic_vector(8129,24);
            manlo <= conv_std_logic_vector(260164976,28);
      WHEN "0111111101" =>
            manhi <= conv_std_logic_vector(8145,24);
            manlo <= conv_std_logic_vector(262248297,28);
      WHEN "0111111110" =>
            manhi <= conv_std_logic_vector(8161,24);
            manlo <= conv_std_logic_vector(264335716,28);
      WHEN "0111111111" =>
            manhi <= conv_std_logic_vector(8177,24);
            manlo <= conv_std_logic_vector(266427233,28);
      WHEN "1000000000" =>
            manhi <= conv_std_logic_vector(8194,24);
            manlo <= conv_std_logic_vector(87392,28);
      WHEN "1000000001" =>
            manhi <= conv_std_logic_vector(8210,24);
            manlo <= conv_std_logic_vector(2187105,28);
      WHEN "1000000010" =>
            manhi <= conv_std_logic_vector(8226,24);
            manlo <= conv_std_logic_vector(4290916,28);
      WHEN "1000000011" =>
            manhi <= conv_std_logic_vector(8242,24);
            manlo <= conv_std_logic_vector(6398825,28);
      WHEN "1000000100" =>
            manhi <= conv_std_logic_vector(8258,24);
            manlo <= conv_std_logic_vector(8510832,28);
      WHEN "1000000101" =>
            manhi <= conv_std_logic_vector(8274,24);
            manlo <= conv_std_logic_vector(10626938,28);
      WHEN "1000000110" =>
            manhi <= conv_std_logic_vector(8290,24);
            manlo <= conv_std_logic_vector(12747141,28);
      WHEN "1000000111" =>
            manhi <= conv_std_logic_vector(8306,24);
            manlo <= conv_std_logic_vector(14871442,28);
      WHEN "1000001000" =>
            manhi <= conv_std_logic_vector(8322,24);
            manlo <= conv_std_logic_vector(16999841,28);
      WHEN "1000001001" =>
            manhi <= conv_std_logic_vector(8338,24);
            manlo <= conv_std_logic_vector(19132338,28);
      WHEN "1000001010" =>
            manhi <= conv_std_logic_vector(8354,24);
            manlo <= conv_std_logic_vector(21268934,28);
      WHEN "1000001011" =>
            manhi <= conv_std_logic_vector(8370,24);
            manlo <= conv_std_logic_vector(23409627,28);
      WHEN "1000001100" =>
            manhi <= conv_std_logic_vector(8386,24);
            manlo <= conv_std_logic_vector(25554418,28);
      WHEN "1000001101" =>
            manhi <= conv_std_logic_vector(8402,24);
            manlo <= conv_std_logic_vector(27703308,28);
      WHEN "1000001110" =>
            manhi <= conv_std_logic_vector(8418,24);
            manlo <= conv_std_logic_vector(29856295,28);
      WHEN "1000001111" =>
            manhi <= conv_std_logic_vector(8434,24);
            manlo <= conv_std_logic_vector(32013381,28);
      WHEN "1000010000" =>
            manhi <= conv_std_logic_vector(8450,24);
            manlo <= conv_std_logic_vector(34174564,28);
      WHEN "1000010001" =>
            manhi <= conv_std_logic_vector(8466,24);
            manlo <= conv_std_logic_vector(36339846,28);
      WHEN "1000010010" =>
            manhi <= conv_std_logic_vector(8482,24);
            manlo <= conv_std_logic_vector(38509225,28);
      WHEN "1000010011" =>
            manhi <= conv_std_logic_vector(8498,24);
            manlo <= conv_std_logic_vector(40682703,28);
      WHEN "1000010100" =>
            manhi <= conv_std_logic_vector(8514,24);
            manlo <= conv_std_logic_vector(42860279,28);
      WHEN "1000010101" =>
            manhi <= conv_std_logic_vector(8530,24);
            manlo <= conv_std_logic_vector(45041953,28);
      WHEN "1000010110" =>
            manhi <= conv_std_logic_vector(8546,24);
            manlo <= conv_std_logic_vector(47227725,28);
      WHEN "1000010111" =>
            manhi <= conv_std_logic_vector(8562,24);
            manlo <= conv_std_logic_vector(49417595,28);
      WHEN "1000011000" =>
            manhi <= conv_std_logic_vector(8578,24);
            manlo <= conv_std_logic_vector(51611563,28);
      WHEN "1000011001" =>
            manhi <= conv_std_logic_vector(8594,24);
            manlo <= conv_std_logic_vector(53809629,28);
      WHEN "1000011010" =>
            manhi <= conv_std_logic_vector(8610,24);
            manlo <= conv_std_logic_vector(56011794,28);
      WHEN "1000011011" =>
            manhi <= conv_std_logic_vector(8626,24);
            manlo <= conv_std_logic_vector(58218056,28);
      WHEN "1000011100" =>
            manhi <= conv_std_logic_vector(8642,24);
            manlo <= conv_std_logic_vector(60428417,28);
      WHEN "1000011101" =>
            manhi <= conv_std_logic_vector(8658,24);
            manlo <= conv_std_logic_vector(62642876,28);
      WHEN "1000011110" =>
            manhi <= conv_std_logic_vector(8674,24);
            manlo <= conv_std_logic_vector(64861432,28);
      WHEN "1000011111" =>
            manhi <= conv_std_logic_vector(8690,24);
            manlo <= conv_std_logic_vector(67084087,28);
      WHEN "1000100000" =>
            manhi <= conv_std_logic_vector(8706,24);
            manlo <= conv_std_logic_vector(69310840,28);
      WHEN "1000100001" =>
            manhi <= conv_std_logic_vector(8722,24);
            manlo <= conv_std_logic_vector(71541691,28);
      WHEN "1000100010" =>
            manhi <= conv_std_logic_vector(8738,24);
            manlo <= conv_std_logic_vector(73776641,28);
      WHEN "1000100011" =>
            manhi <= conv_std_logic_vector(8754,24);
            manlo <= conv_std_logic_vector(76015688,28);
      WHEN "1000100100" =>
            manhi <= conv_std_logic_vector(8770,24);
            manlo <= conv_std_logic_vector(78258834,28);
      WHEN "1000100101" =>
            manhi <= conv_std_logic_vector(8786,24);
            manlo <= conv_std_logic_vector(80506077,28);
      WHEN "1000100110" =>
            manhi <= conv_std_logic_vector(8802,24);
            manlo <= conv_std_logic_vector(82757419,28);
      WHEN "1000100111" =>
            manhi <= conv_std_logic_vector(8818,24);
            manlo <= conv_std_logic_vector(85012859,28);
      WHEN "1000101000" =>
            manhi <= conv_std_logic_vector(8834,24);
            manlo <= conv_std_logic_vector(87272397,28);
      WHEN "1000101001" =>
            manhi <= conv_std_logic_vector(8850,24);
            manlo <= conv_std_logic_vector(89536034,28);
      WHEN "1000101010" =>
            manhi <= conv_std_logic_vector(8866,24);
            manlo <= conv_std_logic_vector(91803768,28);
      WHEN "1000101011" =>
            manhi <= conv_std_logic_vector(8882,24);
            manlo <= conv_std_logic_vector(94075601,28);
      WHEN "1000101100" =>
            manhi <= conv_std_logic_vector(8898,24);
            manlo <= conv_std_logic_vector(96351532,28);
      WHEN "1000101101" =>
            manhi <= conv_std_logic_vector(8914,24);
            manlo <= conv_std_logic_vector(98631561,28);
      WHEN "1000101110" =>
            manhi <= conv_std_logic_vector(8930,24);
            manlo <= conv_std_logic_vector(100915688,28);
      WHEN "1000101111" =>
            manhi <= conv_std_logic_vector(8946,24);
            manlo <= conv_std_logic_vector(103203913,28);
      WHEN "1000110000" =>
            manhi <= conv_std_logic_vector(8962,24);
            manlo <= conv_std_logic_vector(105496237,28);
      WHEN "1000110001" =>
            manhi <= conv_std_logic_vector(8978,24);
            manlo <= conv_std_logic_vector(107792658,28);
      WHEN "1000110010" =>
            manhi <= conv_std_logic_vector(8994,24);
            manlo <= conv_std_logic_vector(110093178,28);
      WHEN "1000110011" =>
            manhi <= conv_std_logic_vector(9010,24);
            manlo <= conv_std_logic_vector(112397796,28);
      WHEN "1000110100" =>
            manhi <= conv_std_logic_vector(9026,24);
            manlo <= conv_std_logic_vector(114706513,28);
      WHEN "1000110101" =>
            manhi <= conv_std_logic_vector(9042,24);
            manlo <= conv_std_logic_vector(117019327,28);
      WHEN "1000110110" =>
            manhi <= conv_std_logic_vector(9058,24);
            manlo <= conv_std_logic_vector(119336240,28);
      WHEN "1000110111" =>
            manhi <= conv_std_logic_vector(9074,24);
            manlo <= conv_std_logic_vector(121657251,28);
      WHEN "1000111000" =>
            manhi <= conv_std_logic_vector(9090,24);
            manlo <= conv_std_logic_vector(123982360,28);
      WHEN "1000111001" =>
            manhi <= conv_std_logic_vector(9106,24);
            manlo <= conv_std_logic_vector(126311567,28);
      WHEN "1000111010" =>
            manhi <= conv_std_logic_vector(9122,24);
            manlo <= conv_std_logic_vector(128644873,28);
      WHEN "1000111011" =>
            manhi <= conv_std_logic_vector(9138,24);
            manlo <= conv_std_logic_vector(130982277,28);
      WHEN "1000111100" =>
            manhi <= conv_std_logic_vector(9154,24);
            manlo <= conv_std_logic_vector(133323779,28);
      WHEN "1000111101" =>
            manhi <= conv_std_logic_vector(9170,24);
            manlo <= conv_std_logic_vector(135669379,28);
      WHEN "1000111110" =>
            manhi <= conv_std_logic_vector(9186,24);
            manlo <= conv_std_logic_vector(138019077,28);
      WHEN "1000111111" =>
            manhi <= conv_std_logic_vector(9202,24);
            manlo <= conv_std_logic_vector(140372874,28);
      WHEN "1001000000" =>
            manhi <= conv_std_logic_vector(9218,24);
            manlo <= conv_std_logic_vector(142730769,28);
      WHEN "1001000001" =>
            manhi <= conv_std_logic_vector(9234,24);
            manlo <= conv_std_logic_vector(145092762,28);
      WHEN "1001000010" =>
            manhi <= conv_std_logic_vector(9250,24);
            manlo <= conv_std_logic_vector(147458854,28);
      WHEN "1001000011" =>
            manhi <= conv_std_logic_vector(9266,24);
            manlo <= conv_std_logic_vector(149829044,28);
      WHEN "1001000100" =>
            manhi <= conv_std_logic_vector(9282,24);
            manlo <= conv_std_logic_vector(152203332,28);
      WHEN "1001000101" =>
            manhi <= conv_std_logic_vector(9298,24);
            manlo <= conv_std_logic_vector(154581718,28);
      WHEN "1001000110" =>
            manhi <= conv_std_logic_vector(9314,24);
            manlo <= conv_std_logic_vector(156964202,28);
      WHEN "1001000111" =>
            manhi <= conv_std_logic_vector(9330,24);
            manlo <= conv_std_logic_vector(159350785,28);
      WHEN "1001001000" =>
            manhi <= conv_std_logic_vector(9346,24);
            manlo <= conv_std_logic_vector(161741466,28);
      WHEN "1001001001" =>
            manhi <= conv_std_logic_vector(9362,24);
            manlo <= conv_std_logic_vector(164136246,28);
      WHEN "1001001010" =>
            manhi <= conv_std_logic_vector(9378,24);
            manlo <= conv_std_logic_vector(166535123,28);
      WHEN "1001001011" =>
            manhi <= conv_std_logic_vector(9394,24);
            manlo <= conv_std_logic_vector(168938099,28);
      WHEN "1001001100" =>
            manhi <= conv_std_logic_vector(9410,24);
            manlo <= conv_std_logic_vector(171345174,28);
      WHEN "1001001101" =>
            manhi <= conv_std_logic_vector(9426,24);
            manlo <= conv_std_logic_vector(173756346,28);
      WHEN "1001001110" =>
            manhi <= conv_std_logic_vector(9442,24);
            manlo <= conv_std_logic_vector(176171617,28);
      WHEN "1001001111" =>
            manhi <= conv_std_logic_vector(9458,24);
            manlo <= conv_std_logic_vector(178590986,28);
      WHEN "1001010000" =>
            manhi <= conv_std_logic_vector(9474,24);
            manlo <= conv_std_logic_vector(181014454,28);
      WHEN "1001010001" =>
            manhi <= conv_std_logic_vector(9490,24);
            manlo <= conv_std_logic_vector(183442020,28);
      WHEN "1001010010" =>
            manhi <= conv_std_logic_vector(9506,24);
            manlo <= conv_std_logic_vector(185873684,28);
      WHEN "1001010011" =>
            manhi <= conv_std_logic_vector(9522,24);
            manlo <= conv_std_logic_vector(188309446,28);
      WHEN "1001010100" =>
            manhi <= conv_std_logic_vector(9538,24);
            manlo <= conv_std_logic_vector(190749307,28);
      WHEN "1001010101" =>
            manhi <= conv_std_logic_vector(9554,24);
            manlo <= conv_std_logic_vector(193193266,28);
      WHEN "1001010110" =>
            manhi <= conv_std_logic_vector(9570,24);
            manlo <= conv_std_logic_vector(195641323,28);
      WHEN "1001010111" =>
            manhi <= conv_std_logic_vector(9586,24);
            manlo <= conv_std_logic_vector(198093479,28);
      WHEN "1001011000" =>
            manhi <= conv_std_logic_vector(9602,24);
            manlo <= conv_std_logic_vector(200549733,28);
      WHEN "1001011001" =>
            manhi <= conv_std_logic_vector(9618,24);
            manlo <= conv_std_logic_vector(203010086,28);
      WHEN "1001011010" =>
            manhi <= conv_std_logic_vector(9634,24);
            manlo <= conv_std_logic_vector(205474536,28);
      WHEN "1001011011" =>
            manhi <= conv_std_logic_vector(9650,24);
            manlo <= conv_std_logic_vector(207943085,28);
      WHEN "1001011100" =>
            manhi <= conv_std_logic_vector(9666,24);
            manlo <= conv_std_logic_vector(210415733,28);
      WHEN "1001011101" =>
            manhi <= conv_std_logic_vector(9682,24);
            manlo <= conv_std_logic_vector(212892479,28);
      WHEN "1001011110" =>
            manhi <= conv_std_logic_vector(9698,24);
            manlo <= conv_std_logic_vector(215373323,28);
      WHEN "1001011111" =>
            manhi <= conv_std_logic_vector(9714,24);
            manlo <= conv_std_logic_vector(217858266,28);
      WHEN "1001100000" =>
            manhi <= conv_std_logic_vector(9730,24);
            manlo <= conv_std_logic_vector(220347307,28);
      WHEN "1001100001" =>
            manhi <= conv_std_logic_vector(9746,24);
            manlo <= conv_std_logic_vector(222840446,28);
      WHEN "1001100010" =>
            manhi <= conv_std_logic_vector(9762,24);
            manlo <= conv_std_logic_vector(225337684,28);
      WHEN "1001100011" =>
            manhi <= conv_std_logic_vector(9778,24);
            manlo <= conv_std_logic_vector(227839020,28);
      WHEN "1001100100" =>
            manhi <= conv_std_logic_vector(9794,24);
            manlo <= conv_std_logic_vector(230344454,28);
      WHEN "1001100101" =>
            manhi <= conv_std_logic_vector(9810,24);
            manlo <= conv_std_logic_vector(232853987,28);
      WHEN "1001100110" =>
            manhi <= conv_std_logic_vector(9826,24);
            manlo <= conv_std_logic_vector(235367618,28);
      WHEN "1001100111" =>
            manhi <= conv_std_logic_vector(9842,24);
            manlo <= conv_std_logic_vector(237885348,28);
      WHEN "1001101000" =>
            manhi <= conv_std_logic_vector(9858,24);
            manlo <= conv_std_logic_vector(240407176,28);
      WHEN "1001101001" =>
            manhi <= conv_std_logic_vector(9874,24);
            manlo <= conv_std_logic_vector(242933102,28);
      WHEN "1001101010" =>
            manhi <= conv_std_logic_vector(9890,24);
            manlo <= conv_std_logic_vector(245463127,28);
      WHEN "1001101011" =>
            manhi <= conv_std_logic_vector(9906,24);
            manlo <= conv_std_logic_vector(247997251,28);
      WHEN "1001101100" =>
            manhi <= conv_std_logic_vector(9922,24);
            manlo <= conv_std_logic_vector(250535472,28);
      WHEN "1001101101" =>
            manhi <= conv_std_logic_vector(9938,24);
            manlo <= conv_std_logic_vector(253077793,28);
      WHEN "1001101110" =>
            manhi <= conv_std_logic_vector(9954,24);
            manlo <= conv_std_logic_vector(255624211,28);
      WHEN "1001101111" =>
            manhi <= conv_std_logic_vector(9970,24);
            manlo <= conv_std_logic_vector(258174728,28);
      WHEN "1001110000" =>
            manhi <= conv_std_logic_vector(9986,24);
            manlo <= conv_std_logic_vector(260729344,28);
      WHEN "1001110001" =>
            manhi <= conv_std_logic_vector(10002,24);
            manlo <= conv_std_logic_vector(263288057,28);
      WHEN "1001110010" =>
            manhi <= conv_std_logic_vector(10018,24);
            manlo <= conv_std_logic_vector(265850870,28);
      WHEN "1001110011" =>
            manhi <= conv_std_logic_vector(10034,24);
            manlo <= conv_std_logic_vector(268417780,28);
      WHEN "1001110100" =>
            manhi <= conv_std_logic_vector(10051,24);
            manlo <= conv_std_logic_vector(2553334,28);
      WHEN "1001110101" =>
            manhi <= conv_std_logic_vector(10067,24);
            manlo <= conv_std_logic_vector(5128441,28);
      WHEN "1001110110" =>
            manhi <= conv_std_logic_vector(10083,24);
            manlo <= conv_std_logic_vector(7707647,28);
      WHEN "1001110111" =>
            manhi <= conv_std_logic_vector(10099,24);
            manlo <= conv_std_logic_vector(10290952,28);
      WHEN "1001111000" =>
            manhi <= conv_std_logic_vector(10115,24);
            manlo <= conv_std_logic_vector(12878355,28);
      WHEN "1001111001" =>
            manhi <= conv_std_logic_vector(10131,24);
            manlo <= conv_std_logic_vector(15469857,28);
      WHEN "1001111010" =>
            manhi <= conv_std_logic_vector(10147,24);
            manlo <= conv_std_logic_vector(18065457,28);
      WHEN "1001111011" =>
            manhi <= conv_std_logic_vector(10163,24);
            manlo <= conv_std_logic_vector(20665155,28);
      WHEN "1001111100" =>
            manhi <= conv_std_logic_vector(10179,24);
            manlo <= conv_std_logic_vector(23268952,28);
      WHEN "1001111101" =>
            manhi <= conv_std_logic_vector(10195,24);
            manlo <= conv_std_logic_vector(25876847,28);
      WHEN "1001111110" =>
            manhi <= conv_std_logic_vector(10211,24);
            manlo <= conv_std_logic_vector(28488841,28);
      WHEN "1001111111" =>
            manhi <= conv_std_logic_vector(10227,24);
            manlo <= conv_std_logic_vector(31104934,28);
      WHEN "1010000000" =>
            manhi <= conv_std_logic_vector(10243,24);
            manlo <= conv_std_logic_vector(33725125,28);
      WHEN "1010000001" =>
            manhi <= conv_std_logic_vector(10259,24);
            manlo <= conv_std_logic_vector(36349414,28);
      WHEN "1010000010" =>
            manhi <= conv_std_logic_vector(10275,24);
            manlo <= conv_std_logic_vector(38977802,28);
      WHEN "1010000011" =>
            manhi <= conv_std_logic_vector(10291,24);
            manlo <= conv_std_logic_vector(41610288,28);
      WHEN "1010000100" =>
            manhi <= conv_std_logic_vector(10307,24);
            manlo <= conv_std_logic_vector(44246873,28);
      WHEN "1010000101" =>
            manhi <= conv_std_logic_vector(10323,24);
            manlo <= conv_std_logic_vector(46887557,28);
      WHEN "1010000110" =>
            manhi <= conv_std_logic_vector(10339,24);
            manlo <= conv_std_logic_vector(49532339,28);
      WHEN "1010000111" =>
            manhi <= conv_std_logic_vector(10355,24);
            manlo <= conv_std_logic_vector(52181219,28);
      WHEN "1010001000" =>
            manhi <= conv_std_logic_vector(10371,24);
            manlo <= conv_std_logic_vector(54834198,28);
      WHEN "1010001001" =>
            manhi <= conv_std_logic_vector(10387,24);
            manlo <= conv_std_logic_vector(57491276,28);
      WHEN "1010001010" =>
            manhi <= conv_std_logic_vector(10403,24);
            manlo <= conv_std_logic_vector(60152452,28);
      WHEN "1010001011" =>
            manhi <= conv_std_logic_vector(10419,24);
            manlo <= conv_std_logic_vector(62817727,28);
      WHEN "1010001100" =>
            manhi <= conv_std_logic_vector(10435,24);
            manlo <= conv_std_logic_vector(65487100,28);
      WHEN "1010001101" =>
            manhi <= conv_std_logic_vector(10451,24);
            manlo <= conv_std_logic_vector(68160572,28);
      WHEN "1010001110" =>
            manhi <= conv_std_logic_vector(10467,24);
            manlo <= conv_std_logic_vector(70838142,28);
      WHEN "1010001111" =>
            manhi <= conv_std_logic_vector(10483,24);
            manlo <= conv_std_logic_vector(73519811,28);
      WHEN "1010010000" =>
            manhi <= conv_std_logic_vector(10499,24);
            manlo <= conv_std_logic_vector(76205578,28);
      WHEN "1010010001" =>
            manhi <= conv_std_logic_vector(10515,24);
            manlo <= conv_std_logic_vector(78895444,28);
      WHEN "1010010010" =>
            manhi <= conv_std_logic_vector(10531,24);
            manlo <= conv_std_logic_vector(81589409,28);
      WHEN "1010010011" =>
            manhi <= conv_std_logic_vector(10547,24);
            manlo <= conv_std_logic_vector(84287472,28);
      WHEN "1010010100" =>
            manhi <= conv_std_logic_vector(10563,24);
            manlo <= conv_std_logic_vector(86989633,28);
      WHEN "1010010101" =>
            manhi <= conv_std_logic_vector(10579,24);
            manlo <= conv_std_logic_vector(89695894,28);
      WHEN "1010010110" =>
            manhi <= conv_std_logic_vector(10595,24);
            manlo <= conv_std_logic_vector(92406252,28);
      WHEN "1010010111" =>
            manhi <= conv_std_logic_vector(10611,24);
            manlo <= conv_std_logic_vector(95120710,28);
      WHEN "1010011000" =>
            manhi <= conv_std_logic_vector(10627,24);
            manlo <= conv_std_logic_vector(97839266,28);
      WHEN "1010011001" =>
            manhi <= conv_std_logic_vector(10643,24);
            manlo <= conv_std_logic_vector(100561920,28);
      WHEN "1010011010" =>
            manhi <= conv_std_logic_vector(10659,24);
            manlo <= conv_std_logic_vector(103288674,28);
      WHEN "1010011011" =>
            manhi <= conv_std_logic_vector(10675,24);
            manlo <= conv_std_logic_vector(106019525,28);
      WHEN "1010011100" =>
            manhi <= conv_std_logic_vector(10691,24);
            manlo <= conv_std_logic_vector(108754476,28);
      WHEN "1010011101" =>
            manhi <= conv_std_logic_vector(10707,24);
            manlo <= conv_std_logic_vector(111493525,28);
      WHEN "1010011110" =>
            manhi <= conv_std_logic_vector(10723,24);
            manlo <= conv_std_logic_vector(114236673,28);
      WHEN "1010011111" =>
            manhi <= conv_std_logic_vector(10739,24);
            manlo <= conv_std_logic_vector(116983919,28);
      WHEN "1010100000" =>
            manhi <= conv_std_logic_vector(10755,24);
            manlo <= conv_std_logic_vector(119735264,28);
      WHEN "1010100001" =>
            manhi <= conv_std_logic_vector(10771,24);
            manlo <= conv_std_logic_vector(122490707,28);
      WHEN "1010100010" =>
            manhi <= conv_std_logic_vector(10787,24);
            manlo <= conv_std_logic_vector(125250249,28);
      WHEN "1010100011" =>
            manhi <= conv_std_logic_vector(10803,24);
            manlo <= conv_std_logic_vector(128013890,28);
      WHEN "1010100100" =>
            manhi <= conv_std_logic_vector(10819,24);
            manlo <= conv_std_logic_vector(130781629,28);
      WHEN "1010100101" =>
            manhi <= conv_std_logic_vector(10835,24);
            manlo <= conv_std_logic_vector(133553468,28);
      WHEN "1010100110" =>
            manhi <= conv_std_logic_vector(10851,24);
            manlo <= conv_std_logic_vector(136329404,28);
      WHEN "1010100111" =>
            manhi <= conv_std_logic_vector(10867,24);
            manlo <= conv_std_logic_vector(139109440,28);
      WHEN "1010101000" =>
            manhi <= conv_std_logic_vector(10883,24);
            manlo <= conv_std_logic_vector(141893574,28);
      WHEN "1010101001" =>
            manhi <= conv_std_logic_vector(10899,24);
            manlo <= conv_std_logic_vector(144681806,28);
      WHEN "1010101010" =>
            manhi <= conv_std_logic_vector(10915,24);
            manlo <= conv_std_logic_vector(147474137,28);
      WHEN "1010101011" =>
            manhi <= conv_std_logic_vector(10931,24);
            manlo <= conv_std_logic_vector(150270567,28);
      WHEN "1010101100" =>
            manhi <= conv_std_logic_vector(10947,24);
            manlo <= conv_std_logic_vector(153071096,28);
      WHEN "1010101101" =>
            manhi <= conv_std_logic_vector(10963,24);
            manlo <= conv_std_logic_vector(155875723,28);
      WHEN "1010101110" =>
            manhi <= conv_std_logic_vector(10979,24);
            manlo <= conv_std_logic_vector(158684449,28);
      WHEN "1010101111" =>
            manhi <= conv_std_logic_vector(10995,24);
            manlo <= conv_std_logic_vector(161497274,28);
      WHEN "1010110000" =>
            manhi <= conv_std_logic_vector(11011,24);
            manlo <= conv_std_logic_vector(164314197,28);
      WHEN "1010110001" =>
            manhi <= conv_std_logic_vector(11027,24);
            manlo <= conv_std_logic_vector(167135219,28);
      WHEN "1010110010" =>
            manhi <= conv_std_logic_vector(11043,24);
            manlo <= conv_std_logic_vector(169960340,28);
      WHEN "1010110011" =>
            manhi <= conv_std_logic_vector(11059,24);
            manlo <= conv_std_logic_vector(172789560,28);
      WHEN "1010110100" =>
            manhi <= conv_std_logic_vector(11075,24);
            manlo <= conv_std_logic_vector(175622878,28);
      WHEN "1010110101" =>
            manhi <= conv_std_logic_vector(11091,24);
            manlo <= conv_std_logic_vector(178460295,28);
      WHEN "1010110110" =>
            manhi <= conv_std_logic_vector(11107,24);
            manlo <= conv_std_logic_vector(181301810,28);
      WHEN "1010110111" =>
            manhi <= conv_std_logic_vector(11123,24);
            manlo <= conv_std_logic_vector(184147424,28);
      WHEN "1010111000" =>
            manhi <= conv_std_logic_vector(11139,24);
            manlo <= conv_std_logic_vector(186997137,28);
      WHEN "1010111001" =>
            manhi <= conv_std_logic_vector(11155,24);
            manlo <= conv_std_logic_vector(189850949,28);
      WHEN "1010111010" =>
            manhi <= conv_std_logic_vector(11171,24);
            manlo <= conv_std_logic_vector(192708860,28);
      WHEN "1010111011" =>
            manhi <= conv_std_logic_vector(11187,24);
            manlo <= conv_std_logic_vector(195570869,28);
      WHEN "1010111100" =>
            manhi <= conv_std_logic_vector(11203,24);
            manlo <= conv_std_logic_vector(198436977,28);
      WHEN "1010111101" =>
            manhi <= conv_std_logic_vector(11219,24);
            manlo <= conv_std_logic_vector(201307183,28);
      WHEN "1010111110" =>
            manhi <= conv_std_logic_vector(11235,24);
            manlo <= conv_std_logic_vector(204181489,28);
      WHEN "1010111111" =>
            manhi <= conv_std_logic_vector(11251,24);
            manlo <= conv_std_logic_vector(207059893,28);
      WHEN "1011000000" =>
            manhi <= conv_std_logic_vector(11267,24);
            manlo <= conv_std_logic_vector(209942395,28);
      WHEN "1011000001" =>
            manhi <= conv_std_logic_vector(11283,24);
            manlo <= conv_std_logic_vector(212828997,28);
      WHEN "1011000010" =>
            manhi <= conv_std_logic_vector(11299,24);
            manlo <= conv_std_logic_vector(215719697,28);
      WHEN "1011000011" =>
            manhi <= conv_std_logic_vector(11315,24);
            manlo <= conv_std_logic_vector(218614497,28);
      WHEN "1011000100" =>
            manhi <= conv_std_logic_vector(11331,24);
            manlo <= conv_std_logic_vector(221513394,28);
      WHEN "1011000101" =>
            manhi <= conv_std_logic_vector(11347,24);
            manlo <= conv_std_logic_vector(224416391,28);
      WHEN "1011000110" =>
            manhi <= conv_std_logic_vector(11363,24);
            manlo <= conv_std_logic_vector(227323486,28);
      WHEN "1011000111" =>
            manhi <= conv_std_logic_vector(11379,24);
            manlo <= conv_std_logic_vector(230234681,28);
      WHEN "1011001000" =>
            manhi <= conv_std_logic_vector(11395,24);
            manlo <= conv_std_logic_vector(233149974,28);
      WHEN "1011001001" =>
            manhi <= conv_std_logic_vector(11411,24);
            manlo <= conv_std_logic_vector(236069365,28);
      WHEN "1011001010" =>
            manhi <= conv_std_logic_vector(11427,24);
            manlo <= conv_std_logic_vector(238992856,28);
      WHEN "1011001011" =>
            manhi <= conv_std_logic_vector(11443,24);
            manlo <= conv_std_logic_vector(241920445,28);
      WHEN "1011001100" =>
            manhi <= conv_std_logic_vector(11459,24);
            manlo <= conv_std_logic_vector(244852133,28);
      WHEN "1011001101" =>
            manhi <= conv_std_logic_vector(11475,24);
            manlo <= conv_std_logic_vector(247787920,28);
      WHEN "1011001110" =>
            manhi <= conv_std_logic_vector(11491,24);
            manlo <= conv_std_logic_vector(250727806,28);
      WHEN "1011001111" =>
            manhi <= conv_std_logic_vector(11507,24);
            manlo <= conv_std_logic_vector(253671790,28);
      WHEN "1011010000" =>
            manhi <= conv_std_logic_vector(11523,24);
            manlo <= conv_std_logic_vector(256619874,28);
      WHEN "1011010001" =>
            manhi <= conv_std_logic_vector(11539,24);
            manlo <= conv_std_logic_vector(259572056,28);
      WHEN "1011010010" =>
            manhi <= conv_std_logic_vector(11555,24);
            manlo <= conv_std_logic_vector(262528337,28);
      WHEN "1011010011" =>
            manhi <= conv_std_logic_vector(11571,24);
            manlo <= conv_std_logic_vector(265488717,28);
      WHEN "1011010100" =>
            manhi <= conv_std_logic_vector(11588,24);
            manlo <= conv_std_logic_vector(17739,28);
      WHEN "1011010101" =>
            manhi <= conv_std_logic_vector(11604,24);
            manlo <= conv_std_logic_vector(2986317,28);
      WHEN "1011010110" =>
            manhi <= conv_std_logic_vector(11620,24);
            manlo <= conv_std_logic_vector(5958993,28);
      WHEN "1011010111" =>
            manhi <= conv_std_logic_vector(11636,24);
            manlo <= conv_std_logic_vector(8935768,28);
      WHEN "1011011000" =>
            manhi <= conv_std_logic_vector(11652,24);
            manlo <= conv_std_logic_vector(11916642,28);
      WHEN "1011011001" =>
            manhi <= conv_std_logic_vector(11668,24);
            manlo <= conv_std_logic_vector(14901615,28);
      WHEN "1011011010" =>
            manhi <= conv_std_logic_vector(11684,24);
            manlo <= conv_std_logic_vector(17890686,28);
      WHEN "1011011011" =>
            manhi <= conv_std_logic_vector(11700,24);
            manlo <= conv_std_logic_vector(20883857,28);
      WHEN "1011011100" =>
            manhi <= conv_std_logic_vector(11716,24);
            manlo <= conv_std_logic_vector(23881126,28);
      WHEN "1011011101" =>
            manhi <= conv_std_logic_vector(11732,24);
            manlo <= conv_std_logic_vector(26882494,28);
      WHEN "1011011110" =>
            manhi <= conv_std_logic_vector(11748,24);
            manlo <= conv_std_logic_vector(29887961,28);
      WHEN "1011011111" =>
            manhi <= conv_std_logic_vector(11764,24);
            manlo <= conv_std_logic_vector(32897527,28);
      WHEN "1011100000" =>
            manhi <= conv_std_logic_vector(11780,24);
            manlo <= conv_std_logic_vector(35911192,28);
      WHEN "1011100001" =>
            manhi <= conv_std_logic_vector(11796,24);
            manlo <= conv_std_logic_vector(38928956,28);
      WHEN "1011100010" =>
            manhi <= conv_std_logic_vector(11812,24);
            manlo <= conv_std_logic_vector(41950818,28);
      WHEN "1011100011" =>
            manhi <= conv_std_logic_vector(11828,24);
            manlo <= conv_std_logic_vector(44976780,28);
      WHEN "1011100100" =>
            manhi <= conv_std_logic_vector(11844,24);
            manlo <= conv_std_logic_vector(48006840,28);
      WHEN "1011100101" =>
            manhi <= conv_std_logic_vector(11860,24);
            manlo <= conv_std_logic_vector(51040999,28);
      WHEN "1011100110" =>
            manhi <= conv_std_logic_vector(11876,24);
            manlo <= conv_std_logic_vector(54079258,28);
      WHEN "1011100111" =>
            manhi <= conv_std_logic_vector(11892,24);
            manlo <= conv_std_logic_vector(57121615,28);
      WHEN "1011101000" =>
            manhi <= conv_std_logic_vector(11908,24);
            manlo <= conv_std_logic_vector(60168071,28);
      WHEN "1011101001" =>
            manhi <= conv_std_logic_vector(11924,24);
            manlo <= conv_std_logic_vector(63218625,28);
      WHEN "1011101010" =>
            manhi <= conv_std_logic_vector(11940,24);
            manlo <= conv_std_logic_vector(66273279,28);
      WHEN "1011101011" =>
            manhi <= conv_std_logic_vector(11956,24);
            manlo <= conv_std_logic_vector(69332032,28);
      WHEN "1011101100" =>
            manhi <= conv_std_logic_vector(11972,24);
            manlo <= conv_std_logic_vector(72394883,28);
      WHEN "1011101101" =>
            manhi <= conv_std_logic_vector(11988,24);
            manlo <= conv_std_logic_vector(75461834,28);
      WHEN "1011101110" =>
            manhi <= conv_std_logic_vector(12004,24);
            manlo <= conv_std_logic_vector(78532883,28);
      WHEN "1011101111" =>
            manhi <= conv_std_logic_vector(12020,24);
            manlo <= conv_std_logic_vector(81608032,28);
      WHEN "1011110000" =>
            manhi <= conv_std_logic_vector(12036,24);
            manlo <= conv_std_logic_vector(84687279,28);
      WHEN "1011110001" =>
            manhi <= conv_std_logic_vector(12052,24);
            manlo <= conv_std_logic_vector(87770625,28);
      WHEN "1011110010" =>
            manhi <= conv_std_logic_vector(12068,24);
            manlo <= conv_std_logic_vector(90858070,28);
      WHEN "1011110011" =>
            manhi <= conv_std_logic_vector(12084,24);
            manlo <= conv_std_logic_vector(93949615,28);
      WHEN "1011110100" =>
            manhi <= conv_std_logic_vector(12100,24);
            manlo <= conv_std_logic_vector(97045258,28);
      WHEN "1011110101" =>
            manhi <= conv_std_logic_vector(12116,24);
            manlo <= conv_std_logic_vector(100145000,28);
      WHEN "1011110110" =>
            manhi <= conv_std_logic_vector(12132,24);
            manlo <= conv_std_logic_vector(103248841,28);
      WHEN "1011110111" =>
            manhi <= conv_std_logic_vector(12148,24);
            manlo <= conv_std_logic_vector(106356781,28);
      WHEN "1011111000" =>
            manhi <= conv_std_logic_vector(12164,24);
            manlo <= conv_std_logic_vector(109468819,28);
      WHEN "1011111001" =>
            manhi <= conv_std_logic_vector(12180,24);
            manlo <= conv_std_logic_vector(112584957,28);
      WHEN "1011111010" =>
            manhi <= conv_std_logic_vector(12196,24);
            manlo <= conv_std_logic_vector(115705194,28);
      WHEN "1011111011" =>
            manhi <= conv_std_logic_vector(12212,24);
            manlo <= conv_std_logic_vector(118829530,28);
      WHEN "1011111100" =>
            manhi <= conv_std_logic_vector(12228,24);
            manlo <= conv_std_logic_vector(121957965,28);
      WHEN "1011111101" =>
            manhi <= conv_std_logic_vector(12244,24);
            manlo <= conv_std_logic_vector(125090499,28);
      WHEN "1011111110" =>
            manhi <= conv_std_logic_vector(12260,24);
            manlo <= conv_std_logic_vector(128227131,28);
      WHEN "1011111111" =>
            manhi <= conv_std_logic_vector(12276,24);
            manlo <= conv_std_logic_vector(131367863,28);
      WHEN "1100000000" =>
            manhi <= conv_std_logic_vector(12292,24);
            manlo <= conv_std_logic_vector(134512694,28);
      WHEN "1100000001" =>
            manhi <= conv_std_logic_vector(12308,24);
            manlo <= conv_std_logic_vector(137661624,28);
      WHEN "1100000010" =>
            manhi <= conv_std_logic_vector(12324,24);
            manlo <= conv_std_logic_vector(140814653,28);
      WHEN "1100000011" =>
            manhi <= conv_std_logic_vector(12340,24);
            manlo <= conv_std_logic_vector(143971780,28);
      WHEN "1100000100" =>
            manhi <= conv_std_logic_vector(12356,24);
            manlo <= conv_std_logic_vector(147133007,28);
      WHEN "1100000101" =>
            manhi <= conv_std_logic_vector(12372,24);
            manlo <= conv_std_logic_vector(150298333,28);
      WHEN "1100000110" =>
            manhi <= conv_std_logic_vector(12388,24);
            manlo <= conv_std_logic_vector(153467758,28);
      WHEN "1100000111" =>
            manhi <= conv_std_logic_vector(12404,24);
            manlo <= conv_std_logic_vector(156641282,28);
      WHEN "1100001000" =>
            manhi <= conv_std_logic_vector(12420,24);
            manlo <= conv_std_logic_vector(159818905,28);
      WHEN "1100001001" =>
            manhi <= conv_std_logic_vector(12436,24);
            manlo <= conv_std_logic_vector(163000627,28);
      WHEN "1100001010" =>
            manhi <= conv_std_logic_vector(12452,24);
            manlo <= conv_std_logic_vector(166186448,28);
      WHEN "1100001011" =>
            manhi <= conv_std_logic_vector(12468,24);
            manlo <= conv_std_logic_vector(169376368,28);
      WHEN "1100001100" =>
            manhi <= conv_std_logic_vector(12484,24);
            manlo <= conv_std_logic_vector(172570387,28);
      WHEN "1100001101" =>
            manhi <= conv_std_logic_vector(12500,24);
            manlo <= conv_std_logic_vector(175768505,28);
      WHEN "1100001110" =>
            manhi <= conv_std_logic_vector(12516,24);
            manlo <= conv_std_logic_vector(178970722,28);
      WHEN "1100001111" =>
            manhi <= conv_std_logic_vector(12532,24);
            manlo <= conv_std_logic_vector(182177038,28);
      WHEN "1100010000" =>
            manhi <= conv_std_logic_vector(12548,24);
            manlo <= conv_std_logic_vector(185387453,28);
      WHEN "1100010001" =>
            manhi <= conv_std_logic_vector(12564,24);
            manlo <= conv_std_logic_vector(188601968,28);
      WHEN "1100010010" =>
            manhi <= conv_std_logic_vector(12580,24);
            manlo <= conv_std_logic_vector(191820581,28);
      WHEN "1100010011" =>
            manhi <= conv_std_logic_vector(12596,24);
            manlo <= conv_std_logic_vector(195043294,28);
      WHEN "1100010100" =>
            manhi <= conv_std_logic_vector(12612,24);
            manlo <= conv_std_logic_vector(198270105,28);
      WHEN "1100010101" =>
            manhi <= conv_std_logic_vector(12628,24);
            manlo <= conv_std_logic_vector(201501016,28);
      WHEN "1100010110" =>
            manhi <= conv_std_logic_vector(12644,24);
            manlo <= conv_std_logic_vector(204736025,28);
      WHEN "1100010111" =>
            manhi <= conv_std_logic_vector(12660,24);
            manlo <= conv_std_logic_vector(207975134,28);
      WHEN "1100011000" =>
            manhi <= conv_std_logic_vector(12676,24);
            manlo <= conv_std_logic_vector(211218342,28);
      WHEN "1100011001" =>
            manhi <= conv_std_logic_vector(12692,24);
            manlo <= conv_std_logic_vector(214465649,28);
      WHEN "1100011010" =>
            manhi <= conv_std_logic_vector(12708,24);
            manlo <= conv_std_logic_vector(217717055,28);
      WHEN "1100011011" =>
            manhi <= conv_std_logic_vector(12724,24);
            manlo <= conv_std_logic_vector(220972560,28);
      WHEN "1100011100" =>
            manhi <= conv_std_logic_vector(12740,24);
            manlo <= conv_std_logic_vector(224232165,28);
      WHEN "1100011101" =>
            manhi <= conv_std_logic_vector(12756,24);
            manlo <= conv_std_logic_vector(227495868,28);
      WHEN "1100011110" =>
            manhi <= conv_std_logic_vector(12772,24);
            manlo <= conv_std_logic_vector(230763671,28);
      WHEN "1100011111" =>
            manhi <= conv_std_logic_vector(12788,24);
            manlo <= conv_std_logic_vector(234035572,28);
      WHEN "1100100000" =>
            manhi <= conv_std_logic_vector(12804,24);
            manlo <= conv_std_logic_vector(237311573,28);
      WHEN "1100100001" =>
            manhi <= conv_std_logic_vector(12820,24);
            manlo <= conv_std_logic_vector(240591673,28);
      WHEN "1100100010" =>
            manhi <= conv_std_logic_vector(12836,24);
            manlo <= conv_std_logic_vector(243875872,28);
      WHEN "1100100011" =>
            manhi <= conv_std_logic_vector(12852,24);
            manlo <= conv_std_logic_vector(247164170,28);
      WHEN "1100100100" =>
            manhi <= conv_std_logic_vector(12868,24);
            manlo <= conv_std_logic_vector(250456567,28);
      WHEN "1100100101" =>
            manhi <= conv_std_logic_vector(12884,24);
            manlo <= conv_std_logic_vector(253753064,28);
      WHEN "1100100110" =>
            manhi <= conv_std_logic_vector(12900,24);
            manlo <= conv_std_logic_vector(257053659,28);
      WHEN "1100100111" =>
            manhi <= conv_std_logic_vector(12916,24);
            manlo <= conv_std_logic_vector(260358354,28);
      WHEN "1100101000" =>
            manhi <= conv_std_logic_vector(12932,24);
            manlo <= conv_std_logic_vector(263667148,28);
      WHEN "1100101001" =>
            manhi <= conv_std_logic_vector(12948,24);
            manlo <= conv_std_logic_vector(266980041,28);
      WHEN "1100101010" =>
            manhi <= conv_std_logic_vector(12965,24);
            manlo <= conv_std_logic_vector(1861577,28);
      WHEN "1100101011" =>
            manhi <= conv_std_logic_vector(12981,24);
            manlo <= conv_std_logic_vector(5182668,28);
      WHEN "1100101100" =>
            manhi <= conv_std_logic_vector(12997,24);
            manlo <= conv_std_logic_vector(8507859,28);
      WHEN "1100101101" =>
            manhi <= conv_std_logic_vector(13013,24);
            manlo <= conv_std_logic_vector(11837149,28);
      WHEN "1100101110" =>
            manhi <= conv_std_logic_vector(13029,24);
            manlo <= conv_std_logic_vector(15170538,28);
      WHEN "1100101111" =>
            manhi <= conv_std_logic_vector(13045,24);
            manlo <= conv_std_logic_vector(18508026,28);
      WHEN "1100110000" =>
            manhi <= conv_std_logic_vector(13061,24);
            manlo <= conv_std_logic_vector(21849613,28);
      WHEN "1100110001" =>
            manhi <= conv_std_logic_vector(13077,24);
            manlo <= conv_std_logic_vector(25195299,28);
      WHEN "1100110010" =>
            manhi <= conv_std_logic_vector(13093,24);
            manlo <= conv_std_logic_vector(28545085,28);
      WHEN "1100110011" =>
            manhi <= conv_std_logic_vector(13109,24);
            manlo <= conv_std_logic_vector(31898970,28);
      WHEN "1100110100" =>
            manhi <= conv_std_logic_vector(13125,24);
            manlo <= conv_std_logic_vector(35256954,28);
      WHEN "1100110101" =>
            manhi <= conv_std_logic_vector(13141,24);
            manlo <= conv_std_logic_vector(38619037,28);
      WHEN "1100110110" =>
            manhi <= conv_std_logic_vector(13157,24);
            manlo <= conv_std_logic_vector(41985219,28);
      WHEN "1100110111" =>
            manhi <= conv_std_logic_vector(13173,24);
            manlo <= conv_std_logic_vector(45355501,28);
      WHEN "1100111000" =>
            manhi <= conv_std_logic_vector(13189,24);
            manlo <= conv_std_logic_vector(48729882,28);
      WHEN "1100111001" =>
            manhi <= conv_std_logic_vector(13205,24);
            manlo <= conv_std_logic_vector(52108362,28);
      WHEN "1100111010" =>
            manhi <= conv_std_logic_vector(13221,24);
            manlo <= conv_std_logic_vector(55490941,28);
      WHEN "1100111011" =>
            manhi <= conv_std_logic_vector(13237,24);
            manlo <= conv_std_logic_vector(58877620,28);
      WHEN "1100111100" =>
            manhi <= conv_std_logic_vector(13253,24);
            manlo <= conv_std_logic_vector(62268398,28);
      WHEN "1100111101" =>
            manhi <= conv_std_logic_vector(13269,24);
            manlo <= conv_std_logic_vector(65663275,28);
      WHEN "1100111110" =>
            manhi <= conv_std_logic_vector(13285,24);
            manlo <= conv_std_logic_vector(69062251,28);
      WHEN "1100111111" =>
            manhi <= conv_std_logic_vector(13301,24);
            manlo <= conv_std_logic_vector(72465326,28);
      WHEN "1101000000" =>
            manhi <= conv_std_logic_vector(13317,24);
            manlo <= conv_std_logic_vector(75872501,28);
      WHEN "1101000001" =>
            manhi <= conv_std_logic_vector(13333,24);
            manlo <= conv_std_logic_vector(79283775,28);
      WHEN "1101000010" =>
            manhi <= conv_std_logic_vector(13349,24);
            manlo <= conv_std_logic_vector(82699148,28);
      WHEN "1101000011" =>
            manhi <= conv_std_logic_vector(13365,24);
            manlo <= conv_std_logic_vector(86118621,28);
      WHEN "1101000100" =>
            manhi <= conv_std_logic_vector(13381,24);
            manlo <= conv_std_logic_vector(89542193,28);
      WHEN "1101000101" =>
            manhi <= conv_std_logic_vector(13397,24);
            manlo <= conv_std_logic_vector(92969864,28);
      WHEN "1101000110" =>
            manhi <= conv_std_logic_vector(13413,24);
            manlo <= conv_std_logic_vector(96401634,28);
      WHEN "1101000111" =>
            manhi <= conv_std_logic_vector(13429,24);
            manlo <= conv_std_logic_vector(99837503,28);
      WHEN "1101001000" =>
            manhi <= conv_std_logic_vector(13445,24);
            manlo <= conv_std_logic_vector(103277472,28);
      WHEN "1101001001" =>
            manhi <= conv_std_logic_vector(13461,24);
            manlo <= conv_std_logic_vector(106721540,28);
      WHEN "1101001010" =>
            manhi <= conv_std_logic_vector(13477,24);
            manlo <= conv_std_logic_vector(110169708,28);
      WHEN "1101001011" =>
            manhi <= conv_std_logic_vector(13493,24);
            manlo <= conv_std_logic_vector(113621975,28);
      WHEN "1101001100" =>
            manhi <= conv_std_logic_vector(13509,24);
            manlo <= conv_std_logic_vector(117078341,28);
      WHEN "1101001101" =>
            manhi <= conv_std_logic_vector(13525,24);
            manlo <= conv_std_logic_vector(120538806,28);
      WHEN "1101001110" =>
            manhi <= conv_std_logic_vector(13541,24);
            manlo <= conv_std_logic_vector(124003370,28);
      WHEN "1101001111" =>
            manhi <= conv_std_logic_vector(13557,24);
            manlo <= conv_std_logic_vector(127472034,28);
      WHEN "1101010000" =>
            manhi <= conv_std_logic_vector(13573,24);
            manlo <= conv_std_logic_vector(130944798,28);
      WHEN "1101010001" =>
            manhi <= conv_std_logic_vector(13589,24);
            manlo <= conv_std_logic_vector(134421660,28);
      WHEN "1101010010" =>
            manhi <= conv_std_logic_vector(13605,24);
            manlo <= conv_std_logic_vector(137902622,28);
      WHEN "1101010011" =>
            manhi <= conv_std_logic_vector(13621,24);
            manlo <= conv_std_logic_vector(141387683,28);
      WHEN "1101010100" =>
            manhi <= conv_std_logic_vector(13637,24);
            manlo <= conv_std_logic_vector(144876844,28);
      WHEN "1101010101" =>
            manhi <= conv_std_logic_vector(13653,24);
            manlo <= conv_std_logic_vector(148370104,28);
      WHEN "1101010110" =>
            manhi <= conv_std_logic_vector(13669,24);
            manlo <= conv_std_logic_vector(151867463,28);
      WHEN "1101010111" =>
            manhi <= conv_std_logic_vector(13685,24);
            manlo <= conv_std_logic_vector(155368921,28);
      WHEN "1101011000" =>
            manhi <= conv_std_logic_vector(13701,24);
            manlo <= conv_std_logic_vector(158874479,28);
      WHEN "1101011001" =>
            manhi <= conv_std_logic_vector(13717,24);
            manlo <= conv_std_logic_vector(162384136,28);
      WHEN "1101011010" =>
            manhi <= conv_std_logic_vector(13733,24);
            manlo <= conv_std_logic_vector(165897893,28);
      WHEN "1101011011" =>
            manhi <= conv_std_logic_vector(13749,24);
            manlo <= conv_std_logic_vector(169415749,28);
      WHEN "1101011100" =>
            manhi <= conv_std_logic_vector(13765,24);
            manlo <= conv_std_logic_vector(172937704,28);
      WHEN "1101011101" =>
            manhi <= conv_std_logic_vector(13781,24);
            manlo <= conv_std_logic_vector(176463758,28);
      WHEN "1101011110" =>
            manhi <= conv_std_logic_vector(13797,24);
            manlo <= conv_std_logic_vector(179993912,28);
      WHEN "1101011111" =>
            manhi <= conv_std_logic_vector(13813,24);
            manlo <= conv_std_logic_vector(183528166,28);
      WHEN "1101100000" =>
            manhi <= conv_std_logic_vector(13829,24);
            manlo <= conv_std_logic_vector(187066519,28);
      WHEN "1101100001" =>
            manhi <= conv_std_logic_vector(13845,24);
            manlo <= conv_std_logic_vector(190608971,28);
      WHEN "1101100010" =>
            manhi <= conv_std_logic_vector(13861,24);
            manlo <= conv_std_logic_vector(194155522,28);
      WHEN "1101100011" =>
            manhi <= conv_std_logic_vector(13877,24);
            manlo <= conv_std_logic_vector(197706173,28);
      WHEN "1101100100" =>
            manhi <= conv_std_logic_vector(13893,24);
            manlo <= conv_std_logic_vector(201260923,28);
      WHEN "1101100101" =>
            manhi <= conv_std_logic_vector(13909,24);
            manlo <= conv_std_logic_vector(204819773,28);
      WHEN "1101100110" =>
            manhi <= conv_std_logic_vector(13925,24);
            manlo <= conv_std_logic_vector(208382722,28);
      WHEN "1101100111" =>
            manhi <= conv_std_logic_vector(13941,24);
            manlo <= conv_std_logic_vector(211949770,28);
      WHEN "1101101000" =>
            manhi <= conv_std_logic_vector(13957,24);
            manlo <= conv_std_logic_vector(215520918,28);
      WHEN "1101101001" =>
            manhi <= conv_std_logic_vector(13973,24);
            manlo <= conv_std_logic_vector(219096165,28);
      WHEN "1101101010" =>
            manhi <= conv_std_logic_vector(13989,24);
            manlo <= conv_std_logic_vector(222675512,28);
      WHEN "1101101011" =>
            manhi <= conv_std_logic_vector(14005,24);
            manlo <= conv_std_logic_vector(226258958,28);
      WHEN "1101101100" =>
            manhi <= conv_std_logic_vector(14021,24);
            manlo <= conv_std_logic_vector(229846504,28);
      WHEN "1101101101" =>
            manhi <= conv_std_logic_vector(14037,24);
            manlo <= conv_std_logic_vector(233438148,28);
      WHEN "1101101110" =>
            manhi <= conv_std_logic_vector(14053,24);
            manlo <= conv_std_logic_vector(237033893,28);
      WHEN "1101101111" =>
            manhi <= conv_std_logic_vector(14069,24);
            manlo <= conv_std_logic_vector(240633737,28);
      WHEN "1101110000" =>
            manhi <= conv_std_logic_vector(14085,24);
            manlo <= conv_std_logic_vector(244237680,28);
      WHEN "1101110001" =>
            manhi <= conv_std_logic_vector(14101,24);
            manlo <= conv_std_logic_vector(247845722,28);
      WHEN "1101110010" =>
            manhi <= conv_std_logic_vector(14117,24);
            manlo <= conv_std_logic_vector(251457864,28);
      WHEN "1101110011" =>
            manhi <= conv_std_logic_vector(14133,24);
            manlo <= conv_std_logic_vector(255074106,28);
      WHEN "1101110100" =>
            manhi <= conv_std_logic_vector(14149,24);
            manlo <= conv_std_logic_vector(258694447,28);
      WHEN "1101110101" =>
            manhi <= conv_std_logic_vector(14165,24);
            manlo <= conv_std_logic_vector(262318887,28);
      WHEN "1101110110" =>
            manhi <= conv_std_logic_vector(14181,24);
            manlo <= conv_std_logic_vector(265947427,28);
      WHEN "1101110111" =>
            manhi <= conv_std_logic_vector(14198,24);
            manlo <= conv_std_logic_vector(1144611,28);
      WHEN "1101111000" =>
            manhi <= conv_std_logic_vector(14214,24);
            manlo <= conv_std_logic_vector(4781350,28);
      WHEN "1101111001" =>
            manhi <= conv_std_logic_vector(14230,24);
            manlo <= conv_std_logic_vector(8422188,28);
      WHEN "1101111010" =>
            manhi <= conv_std_logic_vector(14246,24);
            manlo <= conv_std_logic_vector(12067126,28);
      WHEN "1101111011" =>
            manhi <= conv_std_logic_vector(14262,24);
            manlo <= conv_std_logic_vector(15716163,28);
      WHEN "1101111100" =>
            manhi <= conv_std_logic_vector(14278,24);
            manlo <= conv_std_logic_vector(19369300,28);
      WHEN "1101111101" =>
            manhi <= conv_std_logic_vector(14294,24);
            manlo <= conv_std_logic_vector(23026536,28);
      WHEN "1101111110" =>
            manhi <= conv_std_logic_vector(14310,24);
            manlo <= conv_std_logic_vector(26687871,28);
      WHEN "1101111111" =>
            manhi <= conv_std_logic_vector(14326,24);
            manlo <= conv_std_logic_vector(30353307,28);
      WHEN "1110000000" =>
            manhi <= conv_std_logic_vector(14342,24);
            manlo <= conv_std_logic_vector(34022841,28);
      WHEN "1110000001" =>
            manhi <= conv_std_logic_vector(14358,24);
            manlo <= conv_std_logic_vector(37696476,28);
      WHEN "1110000010" =>
            manhi <= conv_std_logic_vector(14374,24);
            manlo <= conv_std_logic_vector(41374209,28);
      WHEN "1110000011" =>
            manhi <= conv_std_logic_vector(14390,24);
            manlo <= conv_std_logic_vector(45056043,28);
      WHEN "1110000100" =>
            manhi <= conv_std_logic_vector(14406,24);
            manlo <= conv_std_logic_vector(48741975,28);
      WHEN "1110000101" =>
            manhi <= conv_std_logic_vector(14422,24);
            manlo <= conv_std_logic_vector(52432007,28);
      WHEN "1110000110" =>
            manhi <= conv_std_logic_vector(14438,24);
            manlo <= conv_std_logic_vector(56126139,28);
      WHEN "1110000111" =>
            manhi <= conv_std_logic_vector(14454,24);
            manlo <= conv_std_logic_vector(59824371,28);
      WHEN "1110001000" =>
            manhi <= conv_std_logic_vector(14470,24);
            manlo <= conv_std_logic_vector(63526701,28);
      WHEN "1110001001" =>
            manhi <= conv_std_logic_vector(14486,24);
            manlo <= conv_std_logic_vector(67233132,28);
      WHEN "1110001010" =>
            manhi <= conv_std_logic_vector(14502,24);
            manlo <= conv_std_logic_vector(70943662,28);
      WHEN "1110001011" =>
            manhi <= conv_std_logic_vector(14518,24);
            manlo <= conv_std_logic_vector(74658291,28);
      WHEN "1110001100" =>
            manhi <= conv_std_logic_vector(14534,24);
            manlo <= conv_std_logic_vector(78377020,28);
      WHEN "1110001101" =>
            manhi <= conv_std_logic_vector(14550,24);
            manlo <= conv_std_logic_vector(82099849,28);
      WHEN "1110001110" =>
            manhi <= conv_std_logic_vector(14566,24);
            manlo <= conv_std_logic_vector(85826777,28);
      WHEN "1110001111" =>
            manhi <= conv_std_logic_vector(14582,24);
            manlo <= conv_std_logic_vector(89557804,28);
      WHEN "1110010000" =>
            manhi <= conv_std_logic_vector(14598,24);
            manlo <= conv_std_logic_vector(93292931,28);
      WHEN "1110010001" =>
            manhi <= conv_std_logic_vector(14614,24);
            manlo <= conv_std_logic_vector(97032158,28);
      WHEN "1110010010" =>
            manhi <= conv_std_logic_vector(14630,24);
            manlo <= conv_std_logic_vector(100775484,28);
      WHEN "1110010011" =>
            manhi <= conv_std_logic_vector(14646,24);
            manlo <= conv_std_logic_vector(104522910,28);
      WHEN "1110010100" =>
            manhi <= conv_std_logic_vector(14662,24);
            manlo <= conv_std_logic_vector(108274436,28);
      WHEN "1110010101" =>
            manhi <= conv_std_logic_vector(14678,24);
            manlo <= conv_std_logic_vector(112030061,28);
      WHEN "1110010110" =>
            manhi <= conv_std_logic_vector(14694,24);
            manlo <= conv_std_logic_vector(115789786,28);
      WHEN "1110010111" =>
            manhi <= conv_std_logic_vector(14710,24);
            manlo <= conv_std_logic_vector(119553610,28);
      WHEN "1110011000" =>
            manhi <= conv_std_logic_vector(14726,24);
            manlo <= conv_std_logic_vector(123321534,28);
      WHEN "1110011001" =>
            manhi <= conv_std_logic_vector(14742,24);
            manlo <= conv_std_logic_vector(127093557,28);
      WHEN "1110011010" =>
            manhi <= conv_std_logic_vector(14758,24);
            manlo <= conv_std_logic_vector(130869680,28);
      WHEN "1110011011" =>
            manhi <= conv_std_logic_vector(14774,24);
            manlo <= conv_std_logic_vector(134649903,28);
      WHEN "1110011100" =>
            manhi <= conv_std_logic_vector(14790,24);
            manlo <= conv_std_logic_vector(138434225,28);
      WHEN "1110011101" =>
            manhi <= conv_std_logic_vector(14806,24);
            manlo <= conv_std_logic_vector(142222647,28);
      WHEN "1110011110" =>
            manhi <= conv_std_logic_vector(14822,24);
            manlo <= conv_std_logic_vector(146015168,28);
      WHEN "1110011111" =>
            manhi <= conv_std_logic_vector(14838,24);
            manlo <= conv_std_logic_vector(149811789,28);
      WHEN "1110100000" =>
            manhi <= conv_std_logic_vector(14854,24);
            manlo <= conv_std_logic_vector(153612510,28);
      WHEN "1110100001" =>
            manhi <= conv_std_logic_vector(14870,24);
            manlo <= conv_std_logic_vector(157417330,28);
      WHEN "1110100010" =>
            manhi <= conv_std_logic_vector(14886,24);
            manlo <= conv_std_logic_vector(161226250,28);
      WHEN "1110100011" =>
            manhi <= conv_std_logic_vector(14902,24);
            manlo <= conv_std_logic_vector(165039270,28);
      WHEN "1110100100" =>
            manhi <= conv_std_logic_vector(14918,24);
            manlo <= conv_std_logic_vector(168856389,28);
      WHEN "1110100101" =>
            manhi <= conv_std_logic_vector(14934,24);
            manlo <= conv_std_logic_vector(172677608,28);
      WHEN "1110100110" =>
            manhi <= conv_std_logic_vector(14950,24);
            manlo <= conv_std_logic_vector(176502926,28);
      WHEN "1110100111" =>
            manhi <= conv_std_logic_vector(14966,24);
            manlo <= conv_std_logic_vector(180332344,28);
      WHEN "1110101000" =>
            manhi <= conv_std_logic_vector(14982,24);
            manlo <= conv_std_logic_vector(184165862,28);
      WHEN "1110101001" =>
            manhi <= conv_std_logic_vector(14998,24);
            manlo <= conv_std_logic_vector(188003480,28);
      WHEN "1110101010" =>
            manhi <= conv_std_logic_vector(15014,24);
            manlo <= conv_std_logic_vector(191845197,28);
      WHEN "1110101011" =>
            manhi <= conv_std_logic_vector(15030,24);
            manlo <= conv_std_logic_vector(195691014,28);
      WHEN "1110101100" =>
            manhi <= conv_std_logic_vector(15046,24);
            manlo <= conv_std_logic_vector(199540930,28);
      WHEN "1110101101" =>
            manhi <= conv_std_logic_vector(15062,24);
            manlo <= conv_std_logic_vector(203394946,28);
      WHEN "1110101110" =>
            manhi <= conv_std_logic_vector(15078,24);
            manlo <= conv_std_logic_vector(207253062,28);
      WHEN "1110101111" =>
            manhi <= conv_std_logic_vector(15094,24);
            manlo <= conv_std_logic_vector(211115277,28);
      WHEN "1110110000" =>
            manhi <= conv_std_logic_vector(15110,24);
            manlo <= conv_std_logic_vector(214981593,28);
      WHEN "1110110001" =>
            manhi <= conv_std_logic_vector(15126,24);
            manlo <= conv_std_logic_vector(218852007,28);
      WHEN "1110110010" =>
            manhi <= conv_std_logic_vector(15142,24);
            manlo <= conv_std_logic_vector(222726522,28);
      WHEN "1110110011" =>
            manhi <= conv_std_logic_vector(15158,24);
            manlo <= conv_std_logic_vector(226605136,28);
      WHEN "1110110100" =>
            manhi <= conv_std_logic_vector(15174,24);
            manlo <= conv_std_logic_vector(230487850,28);
      WHEN "1110110101" =>
            manhi <= conv_std_logic_vector(15190,24);
            manlo <= conv_std_logic_vector(234374664,28);
      WHEN "1110110110" =>
            manhi <= conv_std_logic_vector(15206,24);
            manlo <= conv_std_logic_vector(238265577,28);
      WHEN "1110110111" =>
            manhi <= conv_std_logic_vector(15222,24);
            manlo <= conv_std_logic_vector(242160590,28);
      WHEN "1110111000" =>
            manhi <= conv_std_logic_vector(15238,24);
            manlo <= conv_std_logic_vector(246059703,28);
      WHEN "1110111001" =>
            manhi <= conv_std_logic_vector(15254,24);
            manlo <= conv_std_logic_vector(249962916,28);
      WHEN "1110111010" =>
            manhi <= conv_std_logic_vector(15270,24);
            manlo <= conv_std_logic_vector(253870228,28);
      WHEN "1110111011" =>
            manhi <= conv_std_logic_vector(15286,24);
            manlo <= conv_std_logic_vector(257781640,28);
      WHEN "1110111100" =>
            manhi <= conv_std_logic_vector(15302,24);
            manlo <= conv_std_logic_vector(261697152,28);
      WHEN "1110111101" =>
            manhi <= conv_std_logic_vector(15318,24);
            manlo <= conv_std_logic_vector(265616763,28);
      WHEN "1110111110" =>
            manhi <= conv_std_logic_vector(15335,24);
            manlo <= conv_std_logic_vector(1105018,28);
      WHEN "1110111111" =>
            manhi <= conv_std_logic_vector(15351,24);
            manlo <= conv_std_logic_vector(5032829,28);
      WHEN "1111000000" =>
            manhi <= conv_std_logic_vector(15367,24);
            manlo <= conv_std_logic_vector(8964740,28);
      WHEN "1111000001" =>
            manhi <= conv_std_logic_vector(15383,24);
            manlo <= conv_std_logic_vector(12900750,28);
      WHEN "1111000010" =>
            manhi <= conv_std_logic_vector(15399,24);
            manlo <= conv_std_logic_vector(16840860,28);
      WHEN "1111000011" =>
            manhi <= conv_std_logic_vector(15415,24);
            manlo <= conv_std_logic_vector(20785070,28);
      WHEN "1111000100" =>
            manhi <= conv_std_logic_vector(15431,24);
            manlo <= conv_std_logic_vector(24733380,28);
      WHEN "1111000101" =>
            manhi <= conv_std_logic_vector(15447,24);
            manlo <= conv_std_logic_vector(28685790,28);
      WHEN "1111000110" =>
            manhi <= conv_std_logic_vector(15463,24);
            manlo <= conv_std_logic_vector(32642299,28);
      WHEN "1111000111" =>
            manhi <= conv_std_logic_vector(15479,24);
            manlo <= conv_std_logic_vector(36602908,28);
      WHEN "1111001000" =>
            manhi <= conv_std_logic_vector(15495,24);
            manlo <= conv_std_logic_vector(40567617,28);
      WHEN "1111001001" =>
            manhi <= conv_std_logic_vector(15511,24);
            manlo <= conv_std_logic_vector(44536425,28);
      WHEN "1111001010" =>
            manhi <= conv_std_logic_vector(15527,24);
            manlo <= conv_std_logic_vector(48509334,28);
      WHEN "1111001011" =>
            manhi <= conv_std_logic_vector(15543,24);
            manlo <= conv_std_logic_vector(52486342,28);
      WHEN "1111001100" =>
            manhi <= conv_std_logic_vector(15559,24);
            manlo <= conv_std_logic_vector(56467450,28);
      WHEN "1111001101" =>
            manhi <= conv_std_logic_vector(15575,24);
            manlo <= conv_std_logic_vector(60452657,28);
      WHEN "1111001110" =>
            manhi <= conv_std_logic_vector(15591,24);
            manlo <= conv_std_logic_vector(64441965,28);
      WHEN "1111001111" =>
            manhi <= conv_std_logic_vector(15607,24);
            manlo <= conv_std_logic_vector(68435372,28);
      WHEN "1111010000" =>
            manhi <= conv_std_logic_vector(15623,24);
            manlo <= conv_std_logic_vector(72432880,28);
      WHEN "1111010001" =>
            manhi <= conv_std_logic_vector(15639,24);
            manlo <= conv_std_logic_vector(76434487,28);
      WHEN "1111010010" =>
            manhi <= conv_std_logic_vector(15655,24);
            manlo <= conv_std_logic_vector(80440193,28);
      WHEN "1111010011" =>
            manhi <= conv_std_logic_vector(15671,24);
            manlo <= conv_std_logic_vector(84450000,28);
      WHEN "1111010100" =>
            manhi <= conv_std_logic_vector(15687,24);
            manlo <= conv_std_logic_vector(88463906,28);
      WHEN "1111010101" =>
            manhi <= conv_std_logic_vector(15703,24);
            manlo <= conv_std_logic_vector(92481913,28);
      WHEN "1111010110" =>
            manhi <= conv_std_logic_vector(15719,24);
            manlo <= conv_std_logic_vector(96504019,28);
      WHEN "1111010111" =>
            manhi <= conv_std_logic_vector(15735,24);
            manlo <= conv_std_logic_vector(100530225,28);
      WHEN "1111011000" =>
            manhi <= conv_std_logic_vector(15751,24);
            manlo <= conv_std_logic_vector(104560531,28);
      WHEN "1111011001" =>
            manhi <= conv_std_logic_vector(15767,24);
            manlo <= conv_std_logic_vector(108594936,28);
      WHEN "1111011010" =>
            manhi <= conv_std_logic_vector(15783,24);
            manlo <= conv_std_logic_vector(112633442,28);
      WHEN "1111011011" =>
            manhi <= conv_std_logic_vector(15799,24);
            manlo <= conv_std_logic_vector(116676047,28);
      WHEN "1111011100" =>
            manhi <= conv_std_logic_vector(15815,24);
            manlo <= conv_std_logic_vector(120722752,28);
      WHEN "1111011101" =>
            manhi <= conv_std_logic_vector(15831,24);
            manlo <= conv_std_logic_vector(124773557,28);
      WHEN "1111011110" =>
            manhi <= conv_std_logic_vector(15847,24);
            manlo <= conv_std_logic_vector(128828462,28);
      WHEN "1111011111" =>
            manhi <= conv_std_logic_vector(15863,24);
            manlo <= conv_std_logic_vector(132887467,28);
      WHEN "1111100000" =>
            manhi <= conv_std_logic_vector(15879,24);
            manlo <= conv_std_logic_vector(136950572,28);
      WHEN "1111100001" =>
            manhi <= conv_std_logic_vector(15895,24);
            manlo <= conv_std_logic_vector(141017776,28);
      WHEN "1111100010" =>
            manhi <= conv_std_logic_vector(15911,24);
            manlo <= conv_std_logic_vector(145089081,28);
      WHEN "1111100011" =>
            manhi <= conv_std_logic_vector(15927,24);
            manlo <= conv_std_logic_vector(149164485,28);
      WHEN "1111100100" =>
            manhi <= conv_std_logic_vector(15943,24);
            manlo <= conv_std_logic_vector(153243989,28);
      WHEN "1111100101" =>
            manhi <= conv_std_logic_vector(15959,24);
            manlo <= conv_std_logic_vector(157327593,28);
      WHEN "1111100110" =>
            manhi <= conv_std_logic_vector(15975,24);
            manlo <= conv_std_logic_vector(161415297,28);
      WHEN "1111100111" =>
            manhi <= conv_std_logic_vector(15991,24);
            manlo <= conv_std_logic_vector(165507101,28);
      WHEN "1111101000" =>
            manhi <= conv_std_logic_vector(16007,24);
            manlo <= conv_std_logic_vector(169603005,28);
      WHEN "1111101001" =>
            manhi <= conv_std_logic_vector(16023,24);
            manlo <= conv_std_logic_vector(173703009,28);
      WHEN "1111101010" =>
            manhi <= conv_std_logic_vector(16039,24);
            manlo <= conv_std_logic_vector(177807112,28);
      WHEN "1111101011" =>
            manhi <= conv_std_logic_vector(16055,24);
            manlo <= conv_std_logic_vector(181915316,28);
      WHEN "1111101100" =>
            manhi <= conv_std_logic_vector(16071,24);
            manlo <= conv_std_logic_vector(186027619,28);
      WHEN "1111101101" =>
            manhi <= conv_std_logic_vector(16087,24);
            manlo <= conv_std_logic_vector(190144023,28);
      WHEN "1111101110" =>
            manhi <= conv_std_logic_vector(16103,24);
            manlo <= conv_std_logic_vector(194264526,28);
      WHEN "1111101111" =>
            manhi <= conv_std_logic_vector(16119,24);
            manlo <= conv_std_logic_vector(198389129,28);
      WHEN "1111110000" =>
            manhi <= conv_std_logic_vector(16135,24);
            manlo <= conv_std_logic_vector(202517832,28);
      WHEN "1111110001" =>
            manhi <= conv_std_logic_vector(16151,24);
            manlo <= conv_std_logic_vector(206650635,28);
      WHEN "1111110010" =>
            manhi <= conv_std_logic_vector(16167,24);
            manlo <= conv_std_logic_vector(210787538,28);
      WHEN "1111110011" =>
            manhi <= conv_std_logic_vector(16183,24);
            manlo <= conv_std_logic_vector(214928541,28);
      WHEN "1111110100" =>
            manhi <= conv_std_logic_vector(16199,24);
            manlo <= conv_std_logic_vector(219073644,28);
      WHEN "1111110101" =>
            manhi <= conv_std_logic_vector(16215,24);
            manlo <= conv_std_logic_vector(223222847,28);
      WHEN "1111110110" =>
            manhi <= conv_std_logic_vector(16231,24);
            manlo <= conv_std_logic_vector(227376150,28);
      WHEN "1111110111" =>
            manhi <= conv_std_logic_vector(16247,24);
            manlo <= conv_std_logic_vector(231533553,28);
      WHEN "1111111000" =>
            manhi <= conv_std_logic_vector(16263,24);
            manlo <= conv_std_logic_vector(235695056,28);
      WHEN "1111111001" =>
            manhi <= conv_std_logic_vector(16279,24);
            manlo <= conv_std_logic_vector(239860659,28);
      WHEN "1111111010" =>
            manhi <= conv_std_logic_vector(16295,24);
            manlo <= conv_std_logic_vector(244030361,28);
      WHEN "1111111011" =>
            manhi <= conv_std_logic_vector(16311,24);
            manlo <= conv_std_logic_vector(248204164,28);
      WHEN "1111111100" =>
            manhi <= conv_std_logic_vector(16327,24);
            manlo <= conv_std_logic_vector(252382067,28);
      WHEN "1111111101" =>
            manhi <= conv_std_logic_vector(16343,24);
            manlo <= conv_std_logic_vector(256564069,28);
      WHEN "1111111110" =>
            manhi <= conv_std_logic_vector(16359,24);
            manlo <= conv_std_logic_vector(260750172,28);
      WHEN "1111111111" =>
            manhi <= conv_std_logic_vector(16375,24);
            manlo <= conv_std_logic_vector(264940375,28);
      WHEN others =>
           manhi <= conv_std_logic_vector(0,24);
           manlo <= conv_std_logic_vector(0,28);
    END CASE;
  END PROCESS;

END rtl;
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   DP_EXPLUTNEG.VHD                          ***
--***                                             ***
--***   Function: Look Up Table - EXP()           ***
--***                                             ***
--***   Generated by MATLAB Utility               ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_explutneg IS
PORT (
      add : IN STD_LOGIC_VECTOR (10 DOWNTO 1);
      manhi : OUT STD_LOGIC_VECTOR (24 DOWNTO 1);
      manlo : OUT STD_LOGIC_VECTOR (28 DOWNTO 1);
      exponent : OUT STD_LOGIC_VECTOR (11 DOWNTO 1)
     );
END dp_explutneg;

ARCHITECTURE rtl OF dp_explutneg IS

BEGIN

  pca: PROCESS (add)
  BEGIN
    CASE add IS
      WHEN "0000000000" =>
            manhi <= conv_std_logic_vector(0,24);
            manlo <= conv_std_logic_vector(0,28);
            exponent <= conv_std_logic_vector(1023,11);
      WHEN "0000000001" =>
            manhi <= conv_std_logic_vector(7910755,24);
            manlo <= conv_std_logic_vector(103608120,28);
            exponent <= conv_std_logic_vector(1021,11);
      WHEN "0000000010" =>
            manhi <= conv_std_logic_vector(1387178,24);
            manlo <= conv_std_logic_vector(62882252,28);
            exponent <= conv_std_logic_vector(1020,11);
      WHEN "0000000011" =>
            manhi <= conv_std_logic_vector(9952012,24);
            manlo <= conv_std_logic_vector(214872239,28);
            exponent <= conv_std_logic_vector(1018,11);
      WHEN "0000000100" =>
            manhi <= conv_std_logic_vector(2889051,24);
            manlo <= conv_std_logic_vector(136396020,28);
            exponent <= conv_std_logic_vector(1017,11);
      WHEN "0000000101" =>
            manhi <= conv_std_logic_vector(12162046,24);
            manlo <= conv_std_logic_vector(873334,28);
            exponent <= conv_std_logic_vector(1015,11);
      WHEN "0000000110" =>
            manhi <= conv_std_logic_vector(4515103,24);
            manlo <= conv_std_logic_vector(18076886,28);
            exponent <= conv_std_logic_vector(1014,11);
      WHEN "0000000111" =>
            manhi <= conv_std_logic_vector(14554809,24);
            manlo <= conv_std_logic_vector(203729295,28);
            exponent <= conv_std_logic_vector(1012,11);
      WHEN "0000001000" =>
            manhi <= conv_std_logic_vector(6275600,24);
            manlo <= conv_std_logic_vector(68167597,28);
            exponent <= conv_std_logic_vector(1011,11);
      WHEN "0000001001" =>
            manhi <= conv_std_logic_vector(184098,24);
            manlo <= conv_std_logic_vector(86398042,28);
            exponent <= conv_std_logic_vector(1010,11);
      WHEN "0000001010" =>
            manhi <= conv_std_logic_vector(8181659,24);
            manlo <= conv_std_logic_vector(90471578,28);
            exponent <= conv_std_logic_vector(1008,11);
      WHEN "0000001011" =>
            manhi <= conv_std_logic_vector(1586498,24);
            manlo <= conv_std_logic_vector(59729764,28);
            exponent <= conv_std_logic_vector(1007,11);
      WHEN "0000001100" =>
            manhi <= conv_std_logic_vector(10245315,24);
            manlo <= conv_std_logic_vector(188988555,28);
            exponent <= conv_std_logic_vector(1005,11);
      WHEN "0000001101" =>
            manhi <= conv_std_logic_vector(3104851,24);
            manlo <= conv_std_logic_vector(194518424,28);
            exponent <= conv_std_logic_vector(1004,11);
      WHEN "0000001110" =>
            manhi <= conv_std_logic_vector(12479599,24);
            manlo <= conv_std_logic_vector(229643794,28);
            exponent <= conv_std_logic_vector(1002,11);
      WHEN "0000001111" =>
            manhi <= conv_std_logic_vector(4748746,24);
            manlo <= conv_std_logic_vector(36170808,28);
            exponent <= conv_std_logic_vector(1001,11);
      WHEN "0000010000" =>
            manhi <= conv_std_logic_vector(14898619,24);
            manlo <= conv_std_logic_vector(183403979,28);
            exponent <= conv_std_logic_vector(999,11);
      WHEN "0000010001" =>
            manhi <= conv_std_logic_vector(6528561,24);
            manlo <= conv_std_logic_vector(123365533,28);
            exponent <= conv_std_logic_vector(998,11);
      WHEN "0000010010" =>
            manhi <= conv_std_logic_vector(370216,24);
            manlo <= conv_std_logic_vector(208248737,28);
            exponent <= conv_std_logic_vector(997,11);
      WHEN "0000010011" =>
            manhi <= conv_std_logic_vector(8455535,24);
            manlo <= conv_std_logic_vector(254564210,28);
            exponent <= conv_std_logic_vector(995,11);
      WHEN "0000010100" =>
            manhi <= conv_std_logic_vector(1788005,24);
            manlo <= conv_std_logic_vector(99840615,28);
            exponent <= conv_std_logic_vector(994,11);
      WHEN "0000010101" =>
            manhi <= conv_std_logic_vector(10541837,24);
            manlo <= conv_std_logic_vector(14529516,28);
            exponent <= conv_std_logic_vector(992,11);
      WHEN "0000010110" =>
            manhi <= conv_std_logic_vector(3323019,24);
            manlo <= conv_std_logic_vector(252804514,28);
            exponent <= conv_std_logic_vector(991,11);
      WHEN "0000010111" =>
            manhi <= conv_std_logic_vector(12800638,24);
            manlo <= conv_std_logic_vector(70515377,28);
            exponent <= conv_std_logic_vector(989,11);
      WHEN "0000011000" =>
            manhi <= conv_std_logic_vector(4984952,24);
            manlo <= conv_std_logic_vector(266936970,28);
            exponent <= conv_std_logic_vector(988,11);
      WHEN "0000011001" =>
            manhi <= conv_std_logic_vector(15246202,24);
            manlo <= conv_std_logic_vector(73384750,28);
            exponent <= conv_std_logic_vector(986,11);
      WHEN "0000011010" =>
            manhi <= conv_std_logic_vector(6784298,24);
            manlo <= conv_std_logic_vector(117472834,28);
            exponent <= conv_std_logic_vector(985,11);
      WHEN "0000011011" =>
            manhi <= conv_std_logic_vector(558377,24);
            manlo <= conv_std_logic_vector(141983386,28);
            exponent <= conv_std_logic_vector(984,11);
      WHEN "0000011100" =>
            manhi <= conv_std_logic_vector(8732417,24);
            manlo <= conv_std_logic_vector(225268666,28);
            exponent <= conv_std_logic_vector(982,11);
      WHEN "0000011101" =>
            manhi <= conv_std_logic_vector(1991723,24);
            manlo <= conv_std_logic_vector(183207072,28);
            exponent <= conv_std_logic_vector(981,11);
      WHEN "0000011110" =>
            manhi <= conv_std_logic_vector(10841612,24);
            manlo <= conv_std_logic_vector(44859253,28);
            exponent <= conv_std_logic_vector(979,11);
      WHEN "0000011111" =>
            manhi <= conv_std_logic_vector(3543582,24);
            manlo <= conv_std_logic_vector(38615994,28);
            exponent <= conv_std_logic_vector(978,11);
      WHEN "0000100000" =>
            manhi <= conv_std_logic_vector(13125199,24);
            manlo <= conv_std_logic_vector(123823208,28);
            exponent <= conv_std_logic_vector(976,11);
      WHEN "0000100001" =>
            manhi <= conv_std_logic_vector(5223751,24);
            manlo <= conv_std_logic_vector(209149352,28);
            exponent <= conv_std_logic_vector(975,11);
      WHEN "0000100010" =>
            manhi <= conv_std_logic_vector(15597598,24);
            manlo <= conv_std_logic_vector(248916640,28);
            exponent <= conv_std_logic_vector(973,11);
      WHEN "0000100011" =>
            manhi <= conv_std_logic_vector(7042841,24);
            manlo <= conv_std_logic_vector(173666528,28);
            exponent <= conv_std_logic_vector(972,11);
      WHEN "0000100100" =>
            manhi <= conv_std_logic_vector(748602,24);
            manlo <= conv_std_logic_vector(266199140,28);
            exponent <= conv_std_logic_vector(971,11);
      WHEN "0000100101" =>
            manhi <= conv_std_logic_vector(9012337,24);
            manlo <= conv_std_logic_vector(264921173,28);
            exponent <= conv_std_logic_vector(969,11);
      WHEN "0000100110" =>
            manhi <= conv_std_logic_vector(2197677,24);
            manlo <= conv_std_logic_vector(112079619,28);
            exponent <= conv_std_logic_vector(968,11);
      WHEN "0000100111" =>
            manhi <= conv_std_logic_vector(11144676,24);
            manlo <= conv_std_logic_vector(200497976,28);
            exponent <= conv_std_logic_vector(966,11);
      WHEN "0000101000" =>
            manhi <= conv_std_logic_vector(3766564,24);
            manlo <= conv_std_logic_vector(161159716,28);
            exponent <= conv_std_logic_vector(965,11);
      WHEN "0000101001" =>
            manhi <= conv_std_logic_vector(13453322,24);
            manlo <= conv_std_logic_vector(28788768,28);
            exponent <= conv_std_logic_vector(963,11);
      WHEN "0000101010" =>
            manhi <= conv_std_logic_vector(5465170,24);
            manlo <= conv_std_logic_vector(249755484,28);
            exponent <= conv_std_logic_vector(962,11);
      WHEN "0000101011" =>
            manhi <= conv_std_logic_vector(15952851,24);
            manlo <= conv_std_logic_vector(133443390,28);
            exponent <= conv_std_logic_vector(960,11);
      WHEN "0000101100" =>
            manhi <= conv_std_logic_vector(7304221,24);
            manlo <= conv_std_logic_vector(236407020,28);
            exponent <= conv_std_logic_vector(959,11);
      WHEN "0000101101" =>
            manhi <= conv_std_logic_vector(940915,24);
            manlo <= conv_std_logic_vector(220198205,28);
            exponent <= conv_std_logic_vector(958,11);
      WHEN "0000101110" =>
            manhi <= conv_std_logic_vector(9295329,24);
            manlo <= conv_std_logic_vector(196124030,28);
            exponent <= conv_std_logic_vector(956,11);
      WHEN "0000101111" =>
            manhi <= conv_std_logic_vector(2405891,24);
            manlo <= conv_std_logic_vector(28613594,28);
            exponent <= conv_std_logic_vector(955,11);
      WHEN "0000110000" =>
            manhi <= conv_std_logic_vector(11451066,24);
            manlo <= conv_std_logic_vector(238698933,28);
            exponent <= conv_std_logic_vector(953,11);
      WHEN "0000110001" =>
            manhi <= conv_std_logic_vector(3991993,24);
            manlo <= conv_std_logic_vector(233279365,28);
            exponent <= conv_std_logic_vector(952,11);
      WHEN "0000110010" =>
            manhi <= conv_std_logic_vector(13785045,24);
            manlo <= conv_std_logic_vector(75368511,28);
            exponent <= conv_std_logic_vector(950,11);
      WHEN "0000110011" =>
            manhi <= conv_std_logic_vector(5709239,24);
            manlo <= conv_std_logic_vector(54173026,28);
            exponent <= conv_std_logic_vector(949,11);
      WHEN "0000110100" =>
            manhi <= conv_std_logic_vector(16312002,24);
            manlo <= conv_std_logic_vector(78993710,28);
            exponent <= conv_std_logic_vector(947,11);
      WHEN "0000110101" =>
            manhi <= conv_std_logic_vector(7568470,24);
            manlo <= conv_std_logic_vector(72422582,28);
            exponent <= conv_std_logic_vector(946,11);
      WHEN "0000110110" =>
            manhi <= conv_std_logic_vector(1135338,24);
            manlo <= conv_std_logic_vector(246889480,28);
            exponent <= conv_std_logic_vector(945,11);
      WHEN "0000110111" =>
            manhi <= conv_std_logic_vector(9581426,24);
            manlo <= conv_std_logic_vector(208117876,28);
            exponent <= conv_std_logic_vector(943,11);
      WHEN "0000111000" =>
            manhi <= conv_std_logic_vector(2616389,24);
            manlo <= conv_std_logic_vector(147217980,28);
            exponent <= conv_std_logic_vector(942,11);
      WHEN "0000111001" =>
            manhi <= conv_std_logic_vector(11760819,24);
            manlo <= conv_std_logic_vector(23037889,28);
            exponent <= conv_std_logic_vector(940,11);
      WHEN "0000111010" =>
            manhi <= conv_std_logic_vector(4219896,24);
            manlo <= conv_std_logic_vector(214481816,28);
            exponent <= conv_std_logic_vector(939,11);
      WHEN "0000111011" =>
            manhi <= conv_std_logic_vector(14120408,24);
            manlo <= conv_std_logic_vector(131761485,28);
            exponent <= conv_std_logic_vector(937,11);
      WHEN "0000111100" =>
            manhi <= conv_std_logic_vector(5955985,24);
            manlo <= conv_std_logic_vector(177821786,28);
            exponent <= conv_std_logic_vector(936,11);
      WHEN "0000111101" =>
            manhi <= conv_std_logic_vector(16675094,24);
            manlo <= conv_std_logic_vector(25356748,28);
            exponent <= conv_std_logic_vector(934,11);
      WHEN "0000111110" =>
            manhi <= conv_std_logic_vector(7835618,24);
            manlo <= conv_std_logic_vector(77011020,28);
            exponent <= conv_std_logic_vector(933,11);
      WHEN "0000111111" =>
            manhi <= conv_std_logic_vector(1331895,24);
            manlo <= conv_std_logic_vector(119779026,28);
            exponent <= conv_std_logic_vector(932,11);
      WHEN "0001000000" =>
            manhi <= conv_std_logic_vector(9870663,24);
            manlo <= conv_std_logic_vector(52552908,28);
            exponent <= conv_std_logic_vector(930,11);
      WHEN "0001000001" =>
            manhi <= conv_std_logic_vector(2829197,24);
            manlo <= conv_std_logic_vector(218477336,28);
            exponent <= conv_std_logic_vector(929,11);
      WHEN "0001000010" =>
            manhi <= conv_std_logic_vector(12073970,24);
            manlo <= conv_std_logic_vector(61450731,28);
            exponent <= conv_std_logic_vector(927,11);
      WHEN "0001000011" =>
            manhi <= conv_std_logic_vector(4450300,24);
            manlo <= conv_std_logic_vector(143360086,28);
            exponent <= conv_std_logic_vector(926,11);
      WHEN "0001000100" =>
            manhi <= conv_std_logic_vector(14459451,24);
            manlo <= conv_std_logic_vector(182543396,28);
            exponent <= conv_std_logic_vector(924,11);
      WHEN "0001000101" =>
            manhi <= conv_std_logic_vector(6205439,24);
            manlo <= conv_std_logic_vector(188004913,28);
            exponent <= conv_std_logic_vector(923,11);
      WHEN "0001000110" =>
            manhi <= conv_std_logic_vector(132477,24);
            manlo <= conv_std_logic_vector(19160299,28);
            exponent <= conv_std_logic_vector(922,11);
      WHEN "0001000111" =>
            manhi <= conv_std_logic_vector(8105697,24);
            manlo <= conv_std_logic_vector(201304075,28);
            exponent <= conv_std_logic_vector(920,11);
      WHEN "0001001000" =>
            manhi <= conv_std_logic_vector(1530608,24);
            manlo <= conv_std_logic_vector(217452229,28);
            exponent <= conv_std_logic_vector(919,11);
      WHEN "0001001001" =>
            manhi <= conv_std_logic_vector(10163073,24);
            manlo <= conv_std_logic_vector(118320126,28);
            exponent <= conv_std_logic_vector(917,11);
      WHEN "0001001010" =>
            manhi <= conv_std_logic_vector(3044341,24);
            manlo <= conv_std_logic_vector(66824260,28);
            exponent <= conv_std_logic_vector(916,11);
      WHEN "0001001011" =>
            manhi <= conv_std_logic_vector(12390557,24);
            manlo <= conv_std_logic_vector(165235674,28);
            exponent <= conv_std_logic_vector(914,11);
      WHEN "0001001100" =>
            manhi <= conv_std_logic_vector(4683232,24);
            manlo <= conv_std_logic_vector(138461149,28);
            exponent <= conv_std_logic_vector(913,11);
      WHEN "0001001101" =>
            manhi <= conv_std_logic_vector(14802215,24);
            manlo <= conv_std_logic_vector(61508170,28);
            exponent <= conv_std_logic_vector(911,11);
      WHEN "0001001110" =>
            manhi <= conv_std_logic_vector(6457631,24);
            manlo <= conv_std_logic_vector(7025744,28);
            exponent <= conv_std_logic_vector(910,11);
      WHEN "0001001111" =>
            manhi <= conv_std_logic_vector(318029,24);
            manlo <= conv_std_logic_vector(21309721,28);
            exponent <= conv_std_logic_vector(909,11);
      WHEN "0001010000" =>
            manhi <= conv_std_logic_vector(8378740,24);
            manlo <= conv_std_logic_vector(221720132,28);
            exponent <= conv_std_logic_vector(907,11);
      WHEN "0001010001" =>
            manhi <= conv_std_logic_vector(1731502,24);
            manlo <= conv_std_logic_vector(182144977,28);
            exponent <= conv_std_logic_vector(906,11);
      WHEN "0001010010" =>
            manhi <= conv_std_logic_vector(10458692,24);
            manlo <= conv_std_logic_vector(90475423,28);
            exponent <= conv_std_logic_vector(904,11);
      WHEN "0001010011" =>
            manhi <= conv_std_logic_vector(3261845,24);
            manlo <= conv_std_logic_vector(128220642,28);
            exponent <= conv_std_logic_vector(903,11);
      WHEN "0001010100" =>
            manhi <= conv_std_logic_vector(12710618,24);
            manlo <= conv_std_logic_vector(255552070,28);
            exponent <= conv_std_logic_vector(901,11);
      WHEN "0001010101" =>
            manhi <= conv_std_logic_vector(4918720,24);
            manlo <= conv_std_logic_vector(130727832,28);
            exponent <= conv_std_logic_vector(900,11);
      WHEN "0001010110" =>
            manhi <= conv_std_logic_vector(15148739,24);
            manlo <= conv_std_logic_vector(258265342,28);
            exponent <= conv_std_logic_vector(898,11);
      WHEN "0001010111" =>
            manhi <= conv_std_logic_vector(6712589,24);
            manlo <= conv_std_logic_vector(181573149,28);
            exponent <= conv_std_logic_vector(897,11);
      WHEN "0001011000" =>
            manhi <= conv_std_logic_vector(505617,24);
            manlo <= conv_std_logic_vector(45883390,28);
            exponent <= conv_std_logic_vector(896,11);
      WHEN "0001011001" =>
            manhi <= conv_std_logic_vector(8654780,24);
            manlo <= conv_std_logic_vector(9428106,28);
            exponent <= conv_std_logic_vector(894,11);
      WHEN "0001011010" =>
            manhi <= conv_std_logic_vector(1934600,24);
            manlo <= conv_std_logic_vector(262677610,28);
            exponent <= conv_std_logic_vector(893,11);
      WHEN "0001011011" =>
            manhi <= conv_std_logic_vector(10757555,24);
            manlo <= conv_std_logic_vector(25094861,28);
            exponent <= conv_std_logic_vector(891,11);
      WHEN "0001011100" =>
            manhi <= conv_std_logic_vector(3481736,24);
            manlo <= conv_std_logic_vector(108799619,28);
            exponent <= conv_std_logic_vector(890,11);
      WHEN "0001011101" =>
            manhi <= conv_std_logic_vector(13034192,24);
            manlo <= conv_std_logic_vector(96190464,28);
            exponent <= conv_std_logic_vector(888,11);
      WHEN "0001011110" =>
            manhi <= conv_std_logic_vector(5156792,24);
            manlo <= conv_std_logic_vector(132821234,28);
            exponent <= conv_std_logic_vector(887,11);
      WHEN "0001011111" =>
            manhi <= conv_std_logic_vector(15499067,24);
            manlo <= conv_std_logic_vector(40497064,28);
            exponent <= conv_std_logic_vector(885,11);
      WHEN "0001100000" =>
            manhi <= conv_std_logic_vector(6970346,24);
            manlo <= conv_std_logic_vector(4633646,28);
            exponent <= conv_std_logic_vector(884,11);
      WHEN "0001100001" =>
            manhi <= conv_std_logic_vector(695263,24);
            manlo <= conv_std_logic_vector(184734272,28);
            exponent <= conv_std_logic_vector(883,11);
      WHEN "0001100010" =>
            manhi <= conv_std_logic_vector(8933848,24);
            manlo <= conv_std_logic_vector(68258056,28);
            exponent <= conv_std_logic_vector(881,11);
      WHEN "0001100011" =>
            manhi <= conv_std_logic_vector(2139927,24);
            manlo <= conv_std_logic_vector(241478077,28);
            exponent <= conv_std_logic_vector(880,11);
      WHEN "0001100100" =>
            manhi <= conv_std_logic_vector(11059697,24);
            manlo <= conv_std_logic_vector(81964893,28);
            exponent <= conv_std_logic_vector(878,11);
      WHEN "0001100101" =>
            manhi <= conv_std_logic_vector(3704040,24);
            manlo <= conv_std_logic_vector(59435624,28);
            exponent <= conv_std_logic_vector(877,11);
      WHEN "0001100110" =>
            manhi <= conv_std_logic_vector(13361316,24);
            manlo <= conv_std_logic_vector(100097713,28);
            exponent <= conv_std_logic_vector(875,11);
      WHEN "0001100111" =>
            manhi <= conv_std_logic_vector(5397476,24);
            manlo <= conv_std_logic_vector(240017437,28);
            exponent <= conv_std_logic_vector(874,11);
      WHEN "0001101000" =>
            manhi <= conv_std_logic_vector(15853238,24);
            manlo <= conv_std_logic_vector(139632179,28);
            exponent <= conv_std_logic_vector(872,11);
      WHEN "0001101001" =>
            manhi <= conv_std_logic_vector(7230930,24);
            manlo <= conv_std_logic_vector(200816807,28);
            exponent <= conv_std_logic_vector(871,11);
      WHEN "0001101010" =>
            manhi <= conv_std_logic_vector(886991,24);
            manlo <= conv_std_logic_vector(58654941,28);
            exponent <= conv_std_logic_vector(870,11);
      WHEN "0001101011" =>
            manhi <= conv_std_logic_vector(9215978,24);
            manlo <= conv_std_logic_vector(193575030,28);
            exponent <= conv_std_logic_vector(868,11);
      WHEN "0001101100" =>
            manhi <= conv_std_logic_vector(2347507,24);
            manlo <= conv_std_logic_vector(240661664,28);
            exponent <= conv_std_logic_vector(867,11);
      WHEN "0001101101" =>
            manhi <= conv_std_logic_vector(11365154,24);
            manlo <= conv_std_logic_vector(257284930,28);
            exponent <= conv_std_logic_vector(865,11);
      WHEN "0001101110" =>
            manhi <= conv_std_logic_vector(3928783,24);
            manlo <= conv_std_logic_vector(108146246,28);
            exponent <= conv_std_logic_vector(864,11);
      WHEN "0001101111" =>
            manhi <= conv_std_logic_vector(13692029,24);
            manlo <= conv_std_logic_vector(256867284,28);
            exponent <= conv_std_logic_vector(862,11);
      WHEN "0001110000" =>
            manhi <= conv_std_logic_vector(5640802,24);
            manlo <= conv_std_logic_vector(94243132,28);
            exponent <= conv_std_logic_vector(861,11);
      WHEN "0001110001" =>
            manhi <= conv_std_logic_vector(16211296,24);
            manlo <= conv_std_logic_vector(67825654,28);
            exponent <= conv_std_logic_vector(859,11);
      WHEN "0001110010" =>
            manhi <= conv_std_logic_vector(7494374,24);
            manlo <= conv_std_logic_vector(242982196,28);
            exponent <= conv_std_logic_vector(858,11);
      WHEN "0001110011" =>
            manhi <= conv_std_logic_vector(1080822,24);
            manlo <= conv_std_logic_vector(160277009,28);
            exponent <= conv_std_logic_vector(857,11);
      WHEN "0001110100" =>
            manhi <= conv_std_logic_vector(9501205,24);
            manlo <= conv_std_logic_vector(10212621,28);
            exponent <= conv_std_logic_vector(855,11);
      WHEN "0001110101" =>
            manhi <= conv_std_logic_vector(2557365,24);
            manlo <= conv_std_logic_vector(185941944,28);
            exponent <= conv_std_logic_vector(854,11);
      WHEN "0001110110" =>
            manhi <= conv_std_logic_vector(11673964,24);
            manlo <= conv_std_logic_vector(116382402,28);
            exponent <= conv_std_logic_vector(852,11);
      WHEN "0001110111" =>
            manhi <= conv_std_logic_vector(4155992,24);
            manlo <= conv_std_logic_vector(192503267,28);
            exponent <= conv_std_logic_vector(851,11);
      WHEN "0001111000" =>
            manhi <= conv_std_logic_vector(14026372,24);
            manlo <= conv_std_logic_vector(133984890,28);
            exponent <= conv_std_logic_vector(849,11);
      WHEN "0001111001" =>
            manhi <= conv_std_logic_vector(5886797,24);
            manlo <= conv_std_logic_vector(227169396,28);
            exponent <= conv_std_logic_vector(848,11);
      WHEN "0001111010" =>
            manhi <= conv_std_logic_vector(16573282,24);
            manlo <= conv_std_logic_vector(266790864,28);
            exponent <= conv_std_logic_vector(846,11);
      WHEN "0001111011" =>
            manhi <= conv_std_logic_vector(7760709,24);
            manlo <= conv_std_logic_vector(232279832,28);
            exponent <= conv_std_logic_vector(845,11);
      WHEN "0001111100" =>
            manhi <= conv_std_logic_vector(1276780,24);
            manlo <= conv_std_logic_vector(244188460,28);
            exponent <= conv_std_logic_vector(844,11);
      WHEN "0001111101" =>
            manhi <= conv_std_logic_vector(9789561,24);
            manlo <= conv_std_logic_vector(47289108,28);
            exponent <= conv_std_logic_vector(842,11);
      WHEN "0001111110" =>
            manhi <= conv_std_logic_vector(2769526,24);
            manlo <= conv_std_logic_vector(75856665,28);
            exponent <= conv_std_logic_vector(841,11);
      WHEN "0001111111" =>
            manhi <= conv_std_logic_vector(11986162,24);
            manlo <= conv_std_logic_vector(137053172,28);
            exponent <= conv_std_logic_vector(839,11);
      WHEN "0010000000" =>
            manhi <= conv_std_logic_vector(4385695,24);
            manlo <= conv_std_logic_vector(60488459,28);
            exponent <= conv_std_logic_vector(838,11);
      WHEN "0010000001" =>
            manhi <= conv_std_logic_vector(14364383,24);
            manlo <= conv_std_logic_vector(220265084,28);
            exponent <= conv_std_logic_vector(836,11);
      WHEN "0010000010" =>
            manhi <= conv_std_logic_vector(6135492,24);
            manlo <= conv_std_logic_vector(182090040,28);
            exponent <= conv_std_logic_vector(835,11);
      WHEN "0010000011" =>
            manhi <= conv_std_logic_vector(81012,24);
            manlo <= conv_std_logic_vector(249275143,28);
            exponent <= conv_std_logic_vector(834,11);
      WHEN "0010000100" =>
            manhi <= conv_std_logic_vector(8029967,24);
            manlo <= conv_std_logic_vector(93846972,28);
            exponent <= conv_std_logic_vector(832,11);
      WHEN "0010000101" =>
            manhi <= conv_std_logic_vector(1474889,24);
            manlo <= conv_std_logic_vector(132978099,28);
            exponent <= conv_std_logic_vector(831,11);
      WHEN "0010000110" =>
            manhi <= conv_std_logic_vector(10081081,24);
            manlo <= conv_std_logic_vector(128680817,28);
            exponent <= conv_std_logic_vector(829,11);
      WHEN "0010000111" =>
            manhi <= conv_std_logic_vector(2984014,24);
            manlo <= conv_std_logic_vector(251002315,28);
            exponent <= conv_std_logic_vector(828,11);
      WHEN "0010001000" =>
            manhi <= conv_std_logic_vector(12301786,24);
            manlo <= conv_std_logic_vector(100124707,28);
            exponent <= conv_std_logic_vector(826,11);
      WHEN "0010001001" =>
            manhi <= conv_std_logic_vector(4617918,24);
            manlo <= conv_std_logic_vector(76665129,28);
            exponent <= conv_std_logic_vector(825,11);
      WHEN "0010001010" =>
            manhi <= conv_std_logic_vector(14706104,24);
            manlo <= conv_std_logic_vector(48076192,28);
            exponent <= conv_std_logic_vector(823,11);
      WHEN "0010001011" =>
            manhi <= conv_std_logic_vector(6386916,24);
            manlo <= conv_std_logic_vector(125471070,28);
            exponent <= conv_std_logic_vector(822,11);
      WHEN "0010001100" =>
            manhi <= conv_std_logic_vector(266000,24);
            manlo <= conv_std_logic_vector(57624675,28);
            exponent <= conv_std_logic_vector(821,11);
      WHEN "0010001101" =>
            manhi <= conv_std_logic_vector(8302179,24);
            manlo <= conv_std_logic_vector(114693198,28);
            exponent <= conv_std_logic_vector(819,11);
      WHEN "0010001110" =>
            manhi <= conv_std_logic_vector(1675171,24);
            manlo <= conv_std_logic_vector(254852645,28);
            exponent <= conv_std_logic_vector(818,11);
      WHEN "0010001111" =>
            manhi <= conv_std_logic_vector(10375800,24);
            manlo <= conv_std_logic_vector(179426511,28);
            exponent <= conv_std_logic_vector(816,11);
      WHEN "0010010000" =>
            manhi <= conv_std_logic_vector(3200857,24);
            manlo <= conv_std_logic_vector(52664716,28);
            exponent <= conv_std_logic_vector(815,11);
      WHEN "0010010001" =>
            manhi <= conv_std_logic_vector(12620873,24);
            manlo <= conv_std_logic_vector(164386702,28);
            exponent <= conv_std_logic_vector(813,11);
      WHEN "0010010010" =>
            manhi <= conv_std_logic_vector(4852689,24);
            manlo <= conv_std_logic_vector(149310968,28);
            exponent <= conv_std_logic_vector(812,11);
      WHEN "0010010011" =>
            manhi <= conv_std_logic_vector(15051574,24);
            manlo <= conv_std_logic_vector(73675604,28);
            exponent <= conv_std_logic_vector(810,11);
      WHEN "0010010100" =>
            manhi <= conv_std_logic_vector(6641099,24);
            manlo <= conv_std_logic_vector(42591307,28);
            exponent <= conv_std_logic_vector(809,11);
      WHEN "0010010101" =>
            manhi <= conv_std_logic_vector(453017,24);
            manlo <= conv_std_logic_vector(104016801,28);
            exponent <= conv_std_logic_vector(808,11);
      WHEN "0010010110" =>
            manhi <= conv_std_logic_vector(8577378,24);
            manlo <= conv_std_logic_vector(139419332,28);
            exponent <= conv_std_logic_vector(806,11);
      WHEN "0010010111" =>
            manhi <= conv_std_logic_vector(1877652,24);
            manlo <= conv_std_logic_vector(33778363,28);
            exponent <= conv_std_logic_vector(805,11);
      WHEN "0010011000" =>
            manhi <= conv_std_logic_vector(10673753,24);
            manlo <= conv_std_logic_vector(226837452,28);
            exponent <= conv_std_logic_vector(803,11);
      WHEN "0010011001" =>
            manhi <= conv_std_logic_vector(3420078,24);
            manlo <= conv_std_logic_vector(239554874,28);
            exponent <= conv_std_logic_vector(802,11);
      WHEN "0010011010" =>
            manhi <= conv_std_logic_vector(12943462,24);
            manlo <= conv_std_logic_vector(62486566,28);
            exponent <= conv_std_logic_vector(800,11);
      WHEN "0010011011" =>
            manhi <= conv_std_logic_vector(5090036,24);
            manlo <= conv_std_logic_vector(268173235,28);
            exponent <= conv_std_logic_vector(799,11);
      WHEN "0010011100" =>
            manhi <= conv_std_logic_vector(15400835,24);
            manlo <= conv_std_logic_vector(67898261,28);
            exponent <= conv_std_logic_vector(797,11);
      WHEN "0010011101" =>
            manhi <= conv_std_logic_vector(6898071,24);
            manlo <= conv_std_logic_vector(6935226,28);
            exponent <= conv_std_logic_vector(796,11);
      WHEN "0010011110" =>
            manhi <= conv_std_logic_vector(642086,24);
            manlo <= conv_std_logic_vector(193616024,28);
            exponent <= conv_std_logic_vector(795,11);
      WHEN "0010011111" =>
            manhi <= conv_std_logic_vector(8855597,24);
            manlo <= conv_std_logic_vector(108124901,28);
            exponent <= conv_std_logic_vector(793,11);
      WHEN "0010100000" =>
            manhi <= conv_std_logic_vector(2082354,24);
            manlo <= conv_std_logic_vector(37727361,28);
            exponent <= conv_std_logic_vector(792,11);
      WHEN "0010100001" =>
            manhi <= conv_std_logic_vector(10974976,24);
            manlo <= conv_std_logic_vector(133184200,28);
            exponent <= conv_std_logic_vector(790,11);
      WHEN "0010100010" =>
            manhi <= conv_std_logic_vector(3641706,24);
            manlo <= conv_std_logic_vector(35844662,28);
            exponent <= conv_std_logic_vector(789,11);
      WHEN "0010100011" =>
            manhi <= conv_std_logic_vector(13269590,24);
            manlo <= conv_std_logic_vector(175886280,28);
            exponent <= conv_std_logic_vector(787,11);
      WHEN "0010100100" =>
            manhi <= conv_std_logic_vector(5329988,24);
            manlo <= conv_std_logic_vector(236927280,28);
            exponent <= conv_std_logic_vector(786,11);
      WHEN "0010100101" =>
            manhi <= conv_std_logic_vector(15753928,24);
            manlo <= conv_std_logic_vector(191213976,28);
            exponent <= conv_std_logic_vector(784,11);
      WHEN "0010100110" =>
            manhi <= conv_std_logic_vector(7157862,24);
            manlo <= conv_std_logic_vector(181160855,28);
            exponent <= conv_std_logic_vector(783,11);
      WHEN "0010100111" =>
            manhi <= conv_std_logic_vector(833230,24);
            manlo <= conv_std_logic_vector(197197075,28);
            exponent <= conv_std_logic_vector(782,11);
      WHEN "0010101000" =>
            manhi <= conv_std_logic_vector(9136869,24);
            manlo <= conv_std_logic_vector(57456047,28);
            exponent <= conv_std_logic_vector(780,11);
      WHEN "0010101001" =>
            manhi <= conv_std_logic_vector(2289302,24);
            manlo <= conv_std_logic_vector(100400411,28);
            exponent <= conv_std_logic_vector(779,11);
      WHEN "0010101010" =>
            manhi <= conv_std_logic_vector(11279504,24);
            manlo <= conv_std_logic_vector(133702078,28);
            exponent <= conv_std_logic_vector(777,11);
      WHEN "0010101011" =>
            manhi <= conv_std_logic_vector(3865765,24);
            manlo <= conv_std_logic_vector(84791606,28);
            exponent <= conv_std_logic_vector(776,11);
      WHEN "0010101100" =>
            manhi <= conv_std_logic_vector(13599297,24);
            manlo <= conv_std_logic_vector(193913492,28);
            exponent <= conv_std_logic_vector(774,11);
      WHEN "0010101101" =>
            manhi <= conv_std_logic_vector(5572573,24);
            manlo <= conv_std_logic_vector(210951234,28);
            exponent <= conv_std_logic_vector(773,11);
      WHEN "0010101110" =>
            manhi <= conv_std_logic_vector(16110896,24);
            manlo <= conv_std_logic_vector(189751005,28);
            exponent <= conv_std_logic_vector(771,11);
      WHEN "0010101111" =>
            manhi <= conv_std_logic_vector(7420505,24);
            manlo <= conv_std_logic_vector(12771910,28);
            exponent <= conv_std_logic_vector(770,11);
      WHEN "0010110000" =>
            manhi <= conv_std_logic_vector(1026472,24);
            manlo <= conv_std_logic_vector(51864863,28);
            exponent <= conv_std_logic_vector(769,11);
      WHEN "0010110001" =>
            manhi <= conv_std_logic_vector(9421227,24);
            manlo <= conv_std_logic_vector(121664951,28);
            exponent <= conv_std_logic_vector(767,11);
      WHEN "0010110010" =>
            manhi <= conv_std_logic_vector(2498521,24);
            manlo <= conv_std_logic_vector(127312793,28);
            exponent <= conv_std_logic_vector(766,11);
      WHEN "0010110011" =>
            manhi <= conv_std_logic_vector(11587374,24);
            manlo <= conv_std_logic_vector(32431827,28);
            exponent <= conv_std_logic_vector(764,11);
      WHEN "0010110100" =>
            manhi <= conv_std_logic_vector(4092283,24);
            manlo <= conv_std_logic_vector(33663701,28);
            exponent <= conv_std_logic_vector(763,11);
      WHEN "0010110101" =>
            manhi <= conv_std_logic_vector(13932622,24);
            manlo <= conv_std_logic_vector(188745186,28);
            exponent <= conv_std_logic_vector(761,11);
      WHEN "0010110110" =>
            manhi <= conv_std_logic_vector(5817820,24);
            manlo <= conv_std_logic_vector(161368804,28);
            exponent <= conv_std_logic_vector(760,11);
      WHEN "0010110111" =>
            manhi <= conv_std_logic_vector(16471781,24);
            manlo <= conv_std_logic_vector(201946939,28);
            exponent <= conv_std_logic_vector(758,11);
      WHEN "0010111000" =>
            manhi <= conv_std_logic_vector(7686029,24);
            manlo <= conv_std_logic_vector(114155240,28);
            exponent <= conv_std_logic_vector(757,11);
      WHEN "0010111001" =>
            manhi <= conv_std_logic_vector(1221834,24);
            manlo <= conv_std_logic_vector(30217784,28);
            exponent <= conv_std_logic_vector(756,11);
      WHEN "0010111010" =>
            manhi <= conv_std_logic_vector(9708705,24);
            manlo <= conv_std_logic_vector(265245416,28);
            exponent <= conv_std_logic_vector(754,11);
      WHEN "0010111011" =>
            manhi <= conv_std_logic_vector(2710036,24);
            manlo <= conv_std_logic_vector(96582323,28);
            exponent <= conv_std_logic_vector(753,11);
      WHEN "0010111100" =>
            manhi <= conv_std_logic_vector(11898622,24);
            manlo <= conv_std_logic_vector(8685564,28);
            exponent <= conv_std_logic_vector(751,11);
      WHEN "0010111101" =>
            manhi <= conv_std_logic_vector(4321286,24);
            manlo <= conv_std_logic_vector(145205332,28);
            exponent <= conv_std_logic_vector(750,11);
      WHEN "0010111110" =>
            manhi <= conv_std_logic_vector(14269605,24);
            manlo <= conv_std_logic_vector(79792252,28);
            exponent <= conv_std_logic_vector(748,11);
      WHEN "0010111111" =>
            manhi <= conv_std_logic_vector(6065758,24);
            manlo <= conv_std_logic_vector(144408455,28);
            exponent <= conv_std_logic_vector(747,11);
      WHEN "0011000000" =>
            manhi <= conv_std_logic_vector(29705,24);
            manlo <= conv_std_logic_vector(111518540,28);
            exponent <= conv_std_logic_vector(746,11);
      WHEN "0011000001" =>
            manhi <= conv_std_logic_vector(7954467,24);
            manlo <= conv_std_logic_vector(116097284,28);
            exponent <= conv_std_logic_vector(744,11);
      WHEN "0011000010" =>
            manhi <= conv_std_logic_vector(1419339,24);
            manlo <= conv_std_logic_vector(204212637,28);
            exponent <= conv_std_logic_vector(743,11);
      WHEN "0011000011" =>
            manhi <= conv_std_logic_vector(9999339,24);
            manlo <= conv_std_logic_vector(15580207,28);
            exponent <= conv_std_logic_vector(741,11);
      WHEN "0011000100" =>
            manhi <= conv_std_logic_vector(2923872,24);
            manlo <= conv_std_logic_vector(59726033,28);
            exponent <= conv_std_logic_vector(740,11);
      WHEN "0011000101" =>
            manhi <= conv_std_logic_vector(12213285,24);
            manlo <= conv_std_logic_vector(81348195,28);
            exponent <= conv_std_logic_vector(738,11);
      WHEN "0011000110" =>
            manhi <= conv_std_logic_vector(4552802,24);
            manlo <= conv_std_logic_vector(224758002,28);
            exponent <= conv_std_logic_vector(737,11);
      WHEN "0011000111" =>
            manhi <= conv_std_logic_vector(14610285,24);
            manlo <= conv_std_logic_vector(171839647,28);
            exponent <= conv_std_logic_vector(735,11);
      WHEN "0011001000" =>
            manhi <= conv_std_logic_vector(6316417,24);
            manlo <= conv_std_logic_vector(33901818,28);
            exponent <= conv_std_logic_vector(734,11);
      WHEN "0011001001" =>
            manhi <= conv_std_logic_vector(214129,24);
            manlo <= conv_std_logic_vector(187432044,28);
            exponent <= conv_std_logic_vector(733,11);
      WHEN "0011001010" =>
            manhi <= conv_std_logic_vector(8225851,24);
            manlo <= conv_std_logic_vector(10972428,28);
            exponent <= conv_std_logic_vector(731,11);
      WHEN "0011001011" =>
            manhi <= conv_std_logic_vector(1619012,24);
            manlo <= conv_std_logic_vector(177473085,28);
            exponent <= conv_std_logic_vector(730,11);
      WHEN "0011001100" =>
            manhi <= conv_std_logic_vector(10293161,24);
            manlo <= conv_std_logic_vector(74648462,28);
            exponent <= conv_std_logic_vector(728,11);
      WHEN "0011001101" =>
            manhi <= conv_std_logic_vector(3140054,24);
            manlo <= conv_std_logic_vector(142465582,28);
            exponent <= conv_std_logic_vector(727,11);
      WHEN "0011001110" =>
            manhi <= conv_std_logic_vector(12531401,24);
            manlo <= conv_std_logic_vector(110062606,28);
            exponent <= conv_std_logic_vector(725,11);
      WHEN "0011001111" =>
            manhi <= conv_std_logic_vector(4786859,24);
            manlo <= conv_std_logic_vector(158003247,28);
            exponent <= conv_std_logic_vector(724,11);
      WHEN "0011010000" =>
            manhi <= conv_std_logic_vector(14954704,24);
            manlo <= conv_std_logic_vector(82587752,28);
            exponent <= conv_std_logic_vector(722,11);
      WHEN "0011010001" =>
            manhi <= conv_std_logic_vector(6569826,24);
            manlo <= conv_std_logic_vector(59098716,28);
            exponent <= conv_std_logic_vector(721,11);
      WHEN "0011010010" =>
            manhi <= conv_std_logic_vector(400577,24);
            manlo <= conv_std_logic_vector(185198176,28);
            exponent <= conv_std_logic_vector(720,11);
      WHEN "0011010011" =>
            manhi <= conv_std_logic_vector(8500212,24);
            manlo <= conv_std_logic_vector(153765179,28);
            exponent <= conv_std_logic_vector(718,11);
      WHEN "0011010100" =>
            manhi <= conv_std_logic_vector(1820876,24);
            manlo <= conv_std_logic_vector(159783545,28);
            exponent <= conv_std_logic_vector(717,11);
      WHEN "0011010101" =>
            manhi <= conv_std_logic_vector(10590207,24);
            manlo <= conv_std_logic_vector(172648734,28);
            exponent <= conv_std_logic_vector(715,11);
      WHEN "0011010110" =>
            manhi <= conv_std_logic_vector(3358609,24);
            manlo <= conv_std_logic_vector(8670608,28);
            exponent <= conv_std_logic_vector(714,11);
      WHEN "0011010111" =>
            manhi <= conv_std_logic_vector(12853008,24);
            manlo <= conv_std_logic_vector(64863304,28);
            exponent <= conv_std_logic_vector(712,11);
      WHEN "0011011000" =>
            manhi <= conv_std_logic_vector(5023484,24);
            manlo <= conv_std_logic_vector(180279682,28);
            exponent <= conv_std_logic_vector(711,11);
      WHEN "0011011001" =>
            manhi <= conv_std_logic_vector(15302902,24);
            manlo <= conv_std_logic_vector(86126918,28);
            exponent <= conv_std_logic_vector(709,11);
      WHEN "0011011010" =>
            manhi <= conv_std_logic_vector(6826016,24);
            manlo <= conv_std_logic_vector(315265,28);
            exponent <= conv_std_logic_vector(708,11);
      WHEN "0011011011" =>
            manhi <= conv_std_logic_vector(589071,24);
            manlo <= conv_std_logic_vector(160219440,28);
            exponent <= conv_std_logic_vector(707,11);
      WHEN "0011011100" =>
            manhi <= conv_std_logic_vector(8777584,24);
            manlo <= conv_std_logic_vector(189361726,28);
            exponent <= conv_std_logic_vector(705,11);
      WHEN "0011011101" =>
            manhi <= conv_std_logic_vector(2024955,24);
            manlo <= conv_std_logic_vector(162543151,28);
            exponent <= conv_std_logic_vector(704,11);
      WHEN "0011011110" =>
            manhi <= conv_std_logic_vector(10890513,24);
            manlo <= conv_std_logic_vector(142859647,28);
            exponent <= conv_std_logic_vector(702,11);
      WHEN "0011011111" =>
            manhi <= conv_std_logic_vector(3579561,24);
            manlo <= conv_std_logic_vector(203359193,28);
            exponent <= conv_std_logic_vector(701,11);
      WHEN "0011100000" =>
            manhi <= conv_std_logic_vector(13178144,24);
            manlo <= conv_std_logic_vector(27387766,28);
            exponent <= conv_std_logic_vector(699,11);
      WHEN "0011100001" =>
            manhi <= conv_std_logic_vector(5262706,24);
            manlo <= conv_std_logic_vector(72167880,28);
            exponent <= conv_std_logic_vector(698,11);
      WHEN "0011100010" =>
            manhi <= conv_std_logic_vector(15654921,24);
            manlo <= conv_std_logic_vector(40507130,28);
            exponent <= conv_std_logic_vector(696,11);
      WHEN "0011100011" =>
            manhi <= conv_std_logic_vector(7085016,24);
            manlo <= conv_std_logic_vector(263640644,28);
            exponent <= conv_std_logic_vector(695,11);
      WHEN "0011100100" =>
            manhi <= conv_std_logic_vector(779633,24);
            manlo <= conv_std_logic_vector(233308885,28);
            exponent <= conv_std_logic_vector(694,11);
      WHEN "0011100101" =>
            manhi <= conv_std_logic_vector(9058000,24);
            manlo <= conv_std_logic_vector(127336500,28);
            exponent <= conv_std_logic_vector(692,11);
      WHEN "0011100110" =>
            manhi <= conv_std_logic_vector(2231273,24);
            manlo <= conv_std_logic_vector(267969878,28);
            exponent <= conv_std_logic_vector(691,11);
      WHEN "0011100111" =>
            manhi <= conv_std_logic_vector(11194114,24);
            manlo <= conv_std_logic_vector(191206462,28);
            exponent <= conv_std_logic_vector(689,11);
      WHEN "0011101000" =>
            manhi <= conv_std_logic_vector(3802939,24);
            manlo <= conv_std_logic_vector(6046440,28);
            exponent <= conv_std_logic_vector(688,11);
      WHEN "0011101001" =>
            manhi <= conv_std_logic_vector(13506847,24);
            manlo <= conv_std_logic_vector(192101060,28);
            exponent <= conv_std_logic_vector(686,11);
      WHEN "0011101010" =>
            manhi <= conv_std_logic_vector(5504552,24);
            manlo <= conv_std_logic_vector(234133234,28);
            exponent <= conv_std_logic_vector(685,11);
      WHEN "0011101011" =>
            manhi <= conv_std_logic_vector(16010802,24);
            manlo <= conv_std_logic_vector(194370273,28);
            exponent <= conv_std_logic_vector(683,11);
      WHEN "0011101100" =>
            manhi <= conv_std_logic_vector(7346860,24);
            manlo <= conv_std_logic_vector(2864438,28);
            exponent <= conv_std_logic_vector(682,11);
      WHEN "0011101101" =>
            manhi <= conv_std_logic_vector(972287,24);
            manlo <= conv_std_logic_vector(54536955,28);
            exponent <= conv_std_logic_vector(681,11);
      WHEN "0011101110" =>
            manhi <= conv_std_logic_vector(9341493,24);
            manlo <= conv_std_logic_vector(74572905,28);
            exponent <= conv_std_logic_vector(679,11);
      WHEN "0011101111" =>
            manhi <= conv_std_logic_vector(2439856,24);
            manlo <= conv_std_logic_vector(93006730,28);
            exponent <= conv_std_logic_vector(678,11);
      WHEN "0011110000" =>
            manhi <= conv_std_logic_vector(11501047,24);
            manlo <= conv_std_logic_vector(92098230,28);
            exponent <= conv_std_logic_vector(676,11);
      WHEN "0011110001" =>
            manhi <= conv_std_logic_vector(4028767,24);
            manlo <= conv_std_logic_vector(115940390,28);
            exponent <= conv_std_logic_vector(675,11);
      WHEN "0011110010" =>
            manhi <= conv_std_logic_vector(13839158,24);
            manlo <= conv_std_logic_vector(62227559,28);
            exponent <= conv_std_logic_vector(673,11);
      WHEN "0011110011" =>
            manhi <= conv_std_logic_vector(5749053,24);
            manlo <= conv_std_logic_vector(76824142,28);
            exponent <= conv_std_logic_vector(672,11);
      WHEN "0011110100" =>
            manhi <= conv_std_logic_vector(16370589,24);
            manlo <= conv_std_logic_vector(114548734,28);
            exponent <= conv_std_logic_vector(670,11);
      WHEN "0011110101" =>
            manhi <= conv_std_logic_vector(7611576,24);
            manlo <= conv_std_logic_vector(73252889,28);
            exponent <= conv_std_logic_vector(669,11);
      WHEN "0011110110" =>
            manhi <= conv_std_logic_vector(1167054,24);
            manlo <= conv_std_logic_vector(146134399,28);
            exponent <= conv_std_logic_vector(668,11);
      WHEN "0011110111" =>
            manhi <= conv_std_logic_vector(9628096,24);
            manlo <= conv_std_logic_vector(236331104,28);
            exponent <= conv_std_logic_vector(666,11);
      WHEN "0011111000" =>
            manhi <= conv_std_logic_vector(2650727,24);
            manlo <= conv_std_logic_vector(132284651,28);
            exponent <= conv_std_logic_vector(665,11);
      WHEN "0011111001" =>
            manhi <= conv_std_logic_vector(11811347,24);
            manlo <= conv_std_logic_vector(263325685,28);
            exponent <= conv_std_logic_vector(663,11);
      WHEN "0011111010" =>
            manhi <= conv_std_logic_vector(4257073,24);
            manlo <= conv_std_logic_vector(236873507,28);
            exponent <= conv_std_logic_vector(662,11);
      WHEN "0011111011" =>
            manhi <= conv_std_logic_vector(14175115,24);
            manlo <= conv_std_logic_vector(61615323,28);
            exponent <= conv_std_logic_vector(660,11);
      WHEN "0011111100" =>
            manhi <= conv_std_logic_vector(5996236,24);
            manlo <= conv_std_logic_vector(169476567,28);
            exponent <= conv_std_logic_vector(659,11);
      WHEN "0011111101" =>
            manhi <= conv_std_logic_vector(16734324,24);
            manlo <= conv_std_logic_vector(29597837,28);
            exponent <= conv_std_logic_vector(657,11);
      WHEN "0011111110" =>
            manhi <= conv_std_logic_vector(7879197,24);
            manlo <= conv_std_logic_vector(79755942,28);
            exponent <= conv_std_logic_vector(656,11);
      WHEN "0011111111" =>
            manhi <= conv_std_logic_vector(1363959,24);
            manlo <= conv_std_logic_vector(24177677,28);
            exponent <= conv_std_logic_vector(655,11);
      WHEN "0100000000" =>
            manhi <= conv_std_logic_vector(9917845,24);
            manlo <= conv_std_logic_vector(112021148,28);
            exponent <= conv_std_logic_vector(653,11);
      WHEN "0100000001" =>
            manhi <= conv_std_logic_vector(2863912,24);
            manlo <= conv_std_logic_vector(148304045,28);
            exponent <= conv_std_logic_vector(652,11);
      WHEN "0100000010" =>
            manhi <= conv_std_logic_vector(12125053,24);
            manlo <= conv_std_logic_vector(156617262,28);
            exponent <= conv_std_logic_vector(650,11);
      WHEN "0100000011" =>
            manhi <= conv_std_logic_vector(4487885,24);
            manlo <= conv_std_logic_vector(151904422,28);
            exponent <= conv_std_logic_vector(649,11);
      WHEN "0100000100" =>
            manhi <= conv_std_logic_vector(14514758,24);
            manlo <= conv_std_logic_vector(193824214,28);
            exponent <= conv_std_logic_vector(647,11);
      WHEN "0100000101" =>
            manhi <= conv_std_logic_vector(6246132,24);
            manlo <= conv_std_logic_vector(93361418,28);
            exponent <= conv_std_logic_vector(646,11);
      WHEN "0100000110" =>
            manhi <= conv_std_logic_vector(162417,24);
            manlo <= conv_std_logic_vector(12929741,28);
            exponent <= conv_std_logic_vector(645,11);
      WHEN "0100000111" =>
            manhi <= conv_std_logic_vector(8149754,24);
            manlo <= conv_std_logic_vector(257063442,28);
            exponent <= conv_std_logic_vector(643,11);
      WHEN "0100001000" =>
            manhi <= conv_std_logic_vector(1563024,24);
            manlo <= conv_std_logic_vector(78378796,28);
            exponent <= conv_std_logic_vector(642,11);
      WHEN "0100001001" =>
            manhi <= conv_std_logic_vector(10210773,24);
            manlo <= conv_std_logic_vector(106907060,28);
            exponent <= conv_std_logic_vector(640,11);
      WHEN "0100001010" =>
            manhi <= conv_std_logic_vector(3079436,24);
            manlo <= conv_std_logic_vector(245979562,28);
            exponent <= conv_std_logic_vector(639,11);
      WHEN "0100001011" =>
            manhi <= conv_std_logic_vector(12442201,24);
            manlo <= conv_std_logic_vector(137868870,28);
            exponent <= conv_std_logic_vector(637,11);
      WHEN "0100001100" =>
            manhi <= conv_std_logic_vector(4721229,24);
            manlo <= conv_std_logic_vector(261058204,28);
            exponent <= conv_std_logic_vector(636,11);
      WHEN "0100001101" =>
            manhi <= conv_std_logic_vector(14858129,24);
            manlo <= conv_std_logic_vector(43405174,28);
            exponent <= conv_std_logic_vector(634,11);
      WHEN "0100001110" =>
            manhi <= conv_std_logic_vector(6498770,24);
            manlo <= conv_std_logic_vector(53338521,28);
            exponent <= conv_std_logic_vector(633,11);
      WHEN "0100001111" =>
            manhi <= conv_std_logic_vector(348297,24);
            manlo <= conv_std_logic_vector(158641329,28);
            exponent <= conv_std_logic_vector(632,11);
      WHEN "0100010000" =>
            manhi <= conv_std_logic_vector(8423281,24);
            manlo <= conv_std_logic_vector(128446906,28);
            exponent <= conv_std_logic_vector(630,11);
      WHEN "0100010001" =>
            manhi <= conv_std_logic_vector(1764273,24);
            manlo <= conv_std_logic_vector(230657816,28);
            exponent <= conv_std_logic_vector(629,11);
      WHEN "0100010010" =>
            manhi <= conv_std_logic_vector(10506915,24);
            manlo <= conv_std_logic_vector(191032874,28);
            exponent <= conv_std_logic_vector(627,11);
      WHEN "0100010011" =>
            manhi <= conv_std_logic_vector(3297326,24);
            manlo <= conv_std_logic_vector(68145509,28);
            exponent <= conv_std_logic_vector(626,11);
      WHEN "0100010100" =>
            manhi <= conv_std_logic_vector(12762829,24);
            manlo <= conv_std_logic_vector(146161159,28);
            exponent <= conv_std_logic_vector(624,11);
      WHEN "0100010101" =>
            manhi <= conv_std_logic_vector(4957134,24);
            manlo <= conv_std_logic_vector(240027976,28);
            exponent <= conv_std_logic_vector(623,11);
      WHEN "0100010110" =>
            manhi <= conv_std_logic_vector(15205267,24);
            manlo <= conv_std_logic_vector(119370809,28);
            exponent <= conv_std_logic_vector(621,11);
      WHEN "0100010111" =>
            manhi <= conv_std_logic_vector(6754180,24);
            manlo <= conv_std_logic_vector(73501816,28);
            exponent <= conv_std_logic_vector(620,11);
      WHEN "0100011000" =>
            manhi <= conv_std_logic_vector(536217,24);
            manlo <= conv_std_logic_vector(220758658,28);
            exponent <= conv_std_logic_vector(619,11);
      WHEN "0100011001" =>
            manhi <= conv_std_logic_vector(8699809,24);
            manlo <= conv_std_logic_vector(117402516,28);
            exponent <= conv_std_logic_vector(617,11);
      WHEN "0100011010" =>
            manhi <= conv_std_logic_vector(1967731,24);
            manlo <= conv_std_logic_vector(204336317,28);
            exponent <= conv_std_logic_vector(616,11);
      WHEN "0100011011" =>
            manhi <= conv_std_logic_vector(10806307,24);
            manlo <= conv_std_logic_vector(168773516,28);
            exponent <= conv_std_logic_vector(614,11);
      WHEN "0100011100" =>
            manhi <= conv_std_logic_vector(3517606,24);
            manlo <= conv_std_logic_vector(138553816,28);
            exponent <= conv_std_logic_vector(613,11);
      WHEN "0100011101" =>
            manhi <= conv_std_logic_vector(13086975,24);
            manlo <= conv_std_logic_vector(231838082,28);
            exponent <= conv_std_logic_vector(611,11);
      WHEN "0100011110" =>
            manhi <= conv_std_logic_vector(5195628,24);
            manlo <= conv_std_logic_vector(114805284,28);
            exponent <= conv_std_logic_vector(610,11);
      WHEN "0100011111" =>
            manhi <= conv_std_logic_vector(15556214,24);
            manlo <= conv_std_logic_vector(245890169,28);
            exponent <= conv_std_logic_vector(608,11);
      WHEN "0100100000" =>
            manhi <= conv_std_logic_vector(7012392,24);
            manlo <= conv_std_logic_vector(266576824,28);
            exponent <= conv_std_logic_vector(607,11);
      WHEN "0100100001" =>
            manhi <= conv_std_logic_vector(726200,24);
            manlo <= conv_std_logic_vector(33318175,28);
            exponent <= conv_std_logic_vector(606,11);
      WHEN "0100100010" =>
            manhi <= conv_std_logic_vector(8979371,24);
            manlo <= conv_std_logic_vector(206515377,28);
            exponent <= conv_std_logic_vector(604,11);
      WHEN "0100100011" =>
            manhi <= conv_std_logic_vector(2173422,24);
            manlo <= conv_std_logic_vector(61774637,28);
            exponent <= conv_std_logic_vector(603,11);
      WHEN "0100100100" =>
            manhi <= conv_std_logic_vector(11108984,24);
            manlo <= conv_std_logic_vector(216833386,28);
            exponent <= conv_std_logic_vector(601,11);
      WHEN "0100100101" =>
            manhi <= conv_std_logic_vector(3740303,24);
            manlo <= conv_std_logic_vector(252090990,28);
            exponent <= conv_std_logic_vector(600,11);
      WHEN "0100100110" =>
            manhi <= conv_std_logic_vector(13414679,24);
            manlo <= conv_std_logic_vector(20856890,28);
            exponent <= conv_std_logic_vector(598,11);
      WHEN "0100100111" =>
            manhi <= conv_std_logic_vector(5436738,24);
            manlo <= conv_std_logic_vector(262578382,28);
            exponent <= conv_std_logic_vector(597,11);
      WHEN "0100101000" =>
            manhi <= conv_std_logic_vector(15911013,24);
            manlo <= conv_std_logic_vector(100481506,28);
            exponent <= conv_std_logic_vector(595,11);
      WHEN "0100101001" =>
            manhi <= conv_std_logic_vector(7273439,24);
            manlo <= conv_std_logic_vector(29586843,28);
            exponent <= conv_std_logic_vector(594,11);
      WHEN "0100101010" =>
            manhi <= conv_std_logic_vector(918267,24);
            manlo <= conv_std_logic_vector(33154287,28);
            exponent <= conv_std_logic_vector(593,11);
      WHEN "0100101011" =>
            manhi <= conv_std_logic_vector(9262001,24);
            manlo <= conv_std_logic_vector(206947959,28);
            exponent <= conv_std_logic_vector(591,11);
      WHEN "0100101100" =>
            manhi <= conv_std_logic_vector(2381369,24);
            manlo <= conv_std_logic_vector(205146615,28);
            exponent <= conv_std_logic_vector(590,11);
      WHEN "0100101101" =>
            manhi <= conv_std_logic_vector(11414983,24);
            manlo <= conv_std_logic_vector(80080029,28);
            exponent <= conv_std_logic_vector(588,11);
      WHEN "0100101110" =>
            manhi <= conv_std_logic_vector(3965445,24);
            manlo <= conv_std_logic_vector(12487826,28);
            exponent <= conv_std_logic_vector(587,11);
      WHEN "0100101111" =>
            manhi <= conv_std_logic_vector(13745978,24);
            manlo <= conv_std_logic_vector(58199715,28);
            exponent <= conv_std_logic_vector(585,11);
      WHEN "0100110000" =>
            manhi <= conv_std_logic_vector(5680495,24);
            manlo <= conv_std_logic_vector(70463110,28);
            exponent <= conv_std_logic_vector(584,11);
      WHEN "0100110001" =>
            manhi <= conv_std_logic_vector(16269705,24);
            manlo <= conv_std_logic_vector(20654997,28);
            exponent <= conv_std_logic_vector(582,11);
      WHEN "0100110010" =>
            manhi <= conv_std_logic_vector(7537349,24);
            manlo <= conv_std_logic_vector(192319832,28);
            exponent <= conv_std_logic_vector(581,11);
      WHEN "0100110011" =>
            manhi <= conv_std_logic_vector(1112441,24);
            manlo <= conv_std_logic_vector(186880957,28);
            exponent <= conv_std_logic_vector(580,11);
      WHEN "0100110100" =>
            manhi <= conv_std_logic_vector(9547733,24);
            manlo <= conv_std_logic_vector(27940083,28);
            exponent <= conv_std_logic_vector(578,11);
      WHEN "0100110101" =>
            manhi <= conv_std_logic_vector(2591599,24);
            manlo <= conv_std_logic_vector(35045549,28);
            exponent <= conv_std_logic_vector(577,11);
      WHEN "0100110110" =>
            manhi <= conv_std_logic_vector(11724339,24);
            manlo <= conv_std_logic_vector(146438512,28);
            exponent <= conv_std_logic_vector(575,11);
      WHEN "0100110111" =>
            manhi <= conv_std_logic_vector(4193056,24);
            manlo <= conv_std_logic_vector(175344679,28);
            exponent <= conv_std_logic_vector(574,11);
      WHEN "0100111000" =>
            manhi <= conv_std_logic_vector(14080912,24);
            manlo <= conv_std_logic_vector(198508677,28);
            exponent <= conv_std_logic_vector(572,11);
      WHEN "0100111001" =>
            manhi <= conv_std_logic_vector(5926926,24);
            manlo <= conv_std_logic_vector(83904648,28);
            exponent <= conv_std_logic_vector(571,11);
      WHEN "0100111010" =>
            manhi <= conv_std_logic_vector(16632332,24);
            manlo <= conv_std_logic_vector(199957404,28);
            exponent <= conv_std_logic_vector(569,11);
      WHEN "0100111011" =>
            manhi <= conv_std_logic_vector(7804156,24);
            manlo <= conv_std_logic_vector(65532420,28);
            exponent <= conv_std_logic_vector(568,11);
      WHEN "0100111100" =>
            manhi <= conv_std_logic_vector(1308746,24);
            manlo <= conv_std_logic_vector(260058525,28);
            exponent <= conv_std_logic_vector(567,11);
      WHEN "0100111101" =>
            manhi <= conv_std_logic_vector(9836599,24);
            manlo <= conv_std_logic_vector(214756046,28);
            exponent <= conv_std_logic_vector(565,11);
      WHEN "0100111110" =>
            manhi <= conv_std_logic_vector(2804135,24);
            manlo <= conv_std_logic_vector(98759674,28);
            exponent <= conv_std_logic_vector(564,11);
      WHEN "0100111111" =>
            manhi <= conv_std_logic_vector(12037090,24);
            manlo <= conv_std_logic_vector(105879341,28);
            exponent <= conv_std_logic_vector(562,11);
      WHEN "0101000000" =>
            manhi <= conv_std_logic_vector(4423165,24);
            manlo <= conv_std_logic_vector(233069674,28);
            exponent <= conv_std_logic_vector(561,11);
      WHEN "0101000001" =>
            manhi <= conv_std_logic_vector(14419522,24);
            manlo <= conv_std_logic_vector(144218340,28);
            exponent <= conv_std_logic_vector(559,11);
      WHEN "0101000010" =>
            manhi <= conv_std_logic_vector(6176061,24);
            manlo <= conv_std_logic_vector(128557517,28);
            exponent <= conv_std_logic_vector(558,11);
      WHEN "0101000011" =>
            manhi <= conv_std_logic_vector(110861,24);
            manlo <= conv_std_logic_vector(210451229,28);
            exponent <= conv_std_logic_vector(557,11);
      WHEN "0101000100" =>
            manhi <= conv_std_logic_vector(8073890,24);
            manlo <= conv_std_logic_vector(126309403,28);
            exponent <= conv_std_logic_vector(555,11);
      WHEN "0101000101" =>
            manhi <= conv_std_logic_vector(1507206,24);
            manlo <= conv_std_logic_vector(86368556,28);
            exponent <= conv_std_logic_vector(554,11);
      WHEN "0101000110" =>
            manhi <= conv_std_logic_vector(10128636,24);
            manlo <= conv_std_logic_vector(70724454,28);
            exponent <= conv_std_logic_vector(552,11);
      WHEN "0101000111" =>
            manhi <= conv_std_logic_vector(3019003,24);
            manlo <= conv_std_logic_vector(212024500,28);
            exponent <= conv_std_logic_vector(551,11);
      WHEN "0101001000" =>
            manhi <= conv_std_logic_vector(12353273,24);
            manlo <= conv_std_logic_vector(25338267,28);
            exponent <= conv_std_logic_vector(549,11);
      WHEN "0101001001" =>
            manhi <= conv_std_logic_vector(4655800,24);
            manlo <= conv_std_logic_vector(26358145,28);
            exponent <= conv_std_logic_vector(548,11);
      WHEN "0101001010" =>
            manhi <= conv_std_logic_vector(14761847,24);
            manlo <= conv_std_logic_vector(252137457,28);
            exponent <= conv_std_logic_vector(546,11);
      WHEN "0101001011" =>
            manhi <= conv_std_logic_vector(6427930,24);
            manlo <= conv_std_logic_vector(116530320,28);
            exponent <= conv_std_logic_vector(545,11);
      WHEN "0101001100" =>
            manhi <= conv_std_logic_vector(296176,24);
            manlo <= conv_std_logic_vector(162393576,28);
            exponent <= conv_std_logic_vector(544,11);
      WHEN "0101001101" =>
            manhi <= conv_std_logic_vector(8346584,24);
            manlo <= conv_std_logic_vector(140031506,28);
            exponent <= conv_std_logic_vector(542,11);
      WHEN "0101001110" =>
            manhi <= conv_std_logic_vector(1707843,24);
            manlo <= conv_std_logic_vector(105232250,28);
            exponent <= conv_std_logic_vector(541,11);
      WHEN "0101001111" =>
            manhi <= conv_std_logic_vector(10423877,24);
            manlo <= conv_std_logic_vector(74257288,28);
            exponent <= conv_std_logic_vector(539,11);
      WHEN "0101010000" =>
            manhi <= conv_std_logic_vector(3236229,24);
            manlo <= conv_std_logic_vector(265138481,28);
            exponent <= conv_std_logic_vector(538,11);
      WHEN "0101010001" =>
            manhi <= conv_std_logic_vector(12672925,24);
            manlo <= conv_std_logic_vector(81471742,28);
            exponent <= conv_std_logic_vector(536,11);
      WHEN "0101010010" =>
            manhi <= conv_std_logic_vector(4890987,24);
            manlo <= conv_std_logic_vector(13504322,28);
            exponent <= conv_std_logic_vector(535,11);
      WHEN "0101010011" =>
            manhi <= conv_std_logic_vector(15107929,24);
            manlo <= conv_std_logic_vector(192561070,28);
            exponent <= conv_std_logic_vector(533,11);
      WHEN "0101010100" =>
            manhi <= conv_std_logic_vector(6682563,24);
            manlo <= conv_std_logic_vector(47334412,28);
            exponent <= conv_std_logic_vector(532,11);
      WHEN "0101010101" =>
            manhi <= conv_std_logic_vector(483524,24);
            manlo <= conv_std_logic_vector(243414774,28);
            exponent <= conv_std_logic_vector(531,11);
      WHEN "0101010110" =>
            manhi <= conv_std_logic_vector(8622270,24);
            manlo <= conv_std_logic_vector(235144322,28);
            exponent <= conv_std_logic_vector(529,11);
      WHEN "0101010111" =>
            manhi <= conv_std_logic_vector(1910682,24);
            manlo <= conv_std_logic_vector(20388866,28);
            exponent <= conv_std_logic_vector(528,11);
      WHEN "0101011000" =>
            manhi <= conv_std_logic_vector(10722358,24);
            manlo <= conv_std_logic_vector(913747,28);
            exponent <= conv_std_logic_vector(526,11);
      WHEN "0101011001" =>
            manhi <= conv_std_logic_vector(3455839,24);
            manlo <= conv_std_logic_vector(223781205,28);
            exponent <= conv_std_logic_vector(525,11);
      WHEN "0101011010" =>
            manhi <= conv_std_logic_vector(12996085,24);
            manlo <= conv_std_logic_vector(24989984,28);
            exponent <= conv_std_logic_vector(523,11);
      WHEN "0101011011" =>
            manhi <= conv_std_logic_vector(5128754,24);
            manlo <= conv_std_logic_vector(197545335,28);
            exponent <= conv_std_logic_vector(522,11);
      WHEN "0101011100" =>
            manhi <= conv_std_logic_vector(15457809,24);
            manlo <= conv_std_logic_vector(24315860,28);
            exponent <= conv_std_logic_vector(520,11);
      WHEN "0101011101" =>
            manhi <= conv_std_logic_vector(6939990,24);
            manlo <= conv_std_logic_vector(8842978,28);
            exponent <= conv_std_logic_vector(519,11);
      WHEN "0101011110" =>
            manhi <= conv_std_logic_vector(672929,24);
            manlo <= conv_std_logic_vector(830489,28);
            exponent <= conv_std_logic_vector(518,11);
      WHEN "0101011111" =>
            manhi <= conv_std_logic_vector(8900982,24);
            manlo <= conv_std_logic_vector(98890321,28);
            exponent <= conv_std_logic_vector(516,11);
      WHEN "0101100000" =>
            manhi <= conv_std_logic_vector(2115746,24);
            manlo <= conv_std_logic_vector(142837003,28);
            exponent <= conv_std_logic_vector(515,11);
      WHEN "0101100001" =>
            manhi <= conv_std_logic_vector(11024113,24);
            manlo <= conv_std_logic_vector(266701758,28);
            exponent <= conv_std_logic_vector(513,11);
      WHEN "0101100010" =>
            manhi <= conv_std_logic_vector(3677859,24);
            manlo <= conv_std_logic_vector(129840563,28);
            exponent <= conv_std_logic_vector(512,11);
      WHEN "0101100011" =>
            manhi <= conv_std_logic_vector(13322790,24);
            manlo <= conv_std_logic_vector(255615990,28);
            exponent <= conv_std_logic_vector(510,11);
      WHEN "0101100100" =>
            manhi <= conv_std_logic_vector(5369131,24);
            manlo <= conv_std_logic_vector(127156783,28);
            exponent <= conv_std_logic_vector(509,11);
      WHEN "0101100101" =>
            manhi <= conv_std_logic_vector(15811527,24);
            manlo <= conv_std_logic_vector(196077973,28);
            exponent <= conv_std_logic_vector(507,11);
      WHEN "0101100110" =>
            manhi <= conv_std_logic_vector(7200241,24);
            manlo <= conv_std_logic_vector(178260644,28);
            exponent <= conv_std_logic_vector(506,11);
      WHEN "0101100111" =>
            manhi <= conv_std_logic_vector(864411,24);
            manlo <= conv_std_logic_vector(121424610,28);
            exponent <= conv_std_logic_vector(505,11);
      WHEN "0101101000" =>
            manhi <= conv_std_logic_vector(9182752,24);
            manlo <= conv_std_logic_vector(52100447,28);
            exponent <= conv_std_logic_vector(503,11);
      WHEN "0101101001" =>
            manhi <= conv_std_logic_vector(2323061,24);
            manlo <= conv_std_logic_vector(49429697,28);
            exponent <= conv_std_logic_vector(502,11);
      WHEN "0101101010" =>
            manhi <= conv_std_logic_vector(11329181,24);
            manlo <= conv_std_logic_vector(50166358,28);
            exponent <= conv_std_logic_vector(500,11);
      WHEN "0101101011" =>
            manhi <= conv_std_logic_vector(3902315,24);
            manlo <= conv_std_logic_vector(102248985,28);
            exponent <= conv_std_logic_vector(499,11);
      WHEN "0101101100" =>
            manhi <= conv_std_logic_vector(13653081,24);
            manlo <= conv_std_logic_vector(212703346,28);
            exponent <= conv_std_logic_vector(497,11);
      WHEN "0101101101" =>
            manhi <= conv_std_logic_vector(5612145,24);
            manlo <= conv_std_logic_vector(239735388,28);
            exponent <= conv_std_logic_vector(496,11);
      WHEN "0101101110" =>
            manhi <= conv_std_logic_vector(16169127,24);
            manlo <= conv_std_logic_vector(205528034,28);
            exponent <= conv_std_logic_vector(494,11);
      WHEN "0101101111" =>
            manhi <= conv_std_logic_vector(7463349,24);
            manlo <= conv_std_logic_vector(17797346,28);
            exponent <= conv_std_logic_vector(493,11);
      WHEN "0101110000" =>
            manhi <= conv_std_logic_vector(1057995,24);
            manlo <= conv_std_logic_vector(16251369,28);
            exponent <= conv_std_logic_vector(492,11);
      WHEN "0101110001" =>
            manhi <= conv_std_logic_vector(9467613,24);
            manlo <= conv_std_logic_vector(244949044,28);
            exponent <= conv_std_logic_vector(490,11);
      WHEN "0101110010" =>
            manhi <= conv_std_logic_vector(2532650,24);
            manlo <= conv_std_logic_vector(194268012,28);
            exponent <= conv_std_logic_vector(489,11);
      WHEN "0101110011" =>
            manhi <= conv_std_logic_vector(11637595,24);
            manlo <= conv_std_logic_vector(246328755,28);
            exponent <= conv_std_logic_vector(487,11);
      WHEN "0101110100" =>
            manhi <= conv_std_logic_vector(4129234,24);
            manlo <= conv_std_logic_vector(69393408,28);
            exponent <= conv_std_logic_vector(486,11);
      WHEN "0101110101" =>
            manhi <= conv_std_logic_vector(13986996,24);
            manlo <= conv_std_logic_vector(255528468,28);
            exponent <= conv_std_logic_vector(484,11);
      WHEN "0101110110" =>
            manhi <= conv_std_logic_vector(5857826,24);
            manlo <= conv_std_logic_vector(251701587,28);
            exponent <= conv_std_logic_vector(483,11);
      WHEN "0101110111" =>
            manhi <= conv_std_logic_vector(16530651,24);
            manlo <= conv_std_logic_vector(211310789,28);
            exponent <= conv_std_logic_vector(481,11);
      WHEN "0101111000" =>
            manhi <= conv_std_logic_vector(7729343,24);
            manlo <= conv_std_logic_vector(154707528,28);
            exponent <= conv_std_logic_vector(480,11);
      WHEN "0101111001" =>
            manhi <= conv_std_logic_vector(1253702,24);
            manlo <= conv_std_logic_vector(237283577,28);
            exponent <= conv_std_logic_vector(479,11);
      WHEN "0101111010" =>
            manhi <= conv_std_logic_vector(9755601,24);
            manlo <= conv_std_logic_vector(121155884,28);
            exponent <= conv_std_logic_vector(477,11);
      WHEN "0101111011" =>
            manhi <= conv_std_logic_vector(2744540,24);
            manlo <= conv_std_logic_vector(30442277,28);
            exponent <= conv_std_logic_vector(476,11);
      WHEN "0101111100" =>
            manhi <= conv_std_logic_vector(11949394,24);
            manlo <= conv_std_logic_vector(246622503,28);
            exponent <= conv_std_logic_vector(474,11);
      WHEN "0101111101" =>
            manhi <= conv_std_logic_vector(4358643,24);
            manlo <= conv_std_logic_vector(38405425,28);
            exponent <= conv_std_logic_vector(473,11);
      WHEN "0101111110" =>
            manhi <= conv_std_logic_vector(14324576,24);
            manlo <= conv_std_logic_vector(53935566,28);
            exponent <= conv_std_logic_vector(471,11);
      WHEN "0101111111" =>
            manhi <= conv_std_logic_vector(6106203,24);
            manlo <= conv_std_logic_vector(233166714,28);
            exponent <= conv_std_logic_vector(470,11);
      WHEN "0110000000" =>
            manhi <= conv_std_logic_vector(59463,24);
            manlo <= conv_std_logic_vector(114545214,28);
            exponent <= conv_std_logic_vector(469,11);
      WHEN "0110000001" =>
            manhi <= conv_std_logic_vector(7998256,24);
            manlo <= conv_std_logic_vector(234808364,28);
            exponent <= conv_std_logic_vector(467,11);
      WHEN "0110000010" =>
            manhi <= conv_std_logic_vector(1451558,24);
            manlo <= conv_std_logic_vector(62230667,28);
            exponent <= conv_std_logic_vector(466,11);
      WHEN "0110000011" =>
            manhi <= conv_std_logic_vector(10046749,24);
            manlo <= conv_std_logic_vector(29683609,28);
            exponent <= conv_std_logic_vector(464,11);
      WHEN "0110000100" =>
            manhi <= conv_std_logic_vector(2958754,24);
            manlo <= conv_std_logic_vector(158313814,28);
            exponent <= conv_std_logic_vector(463,11);
      WHEN "0110000101" =>
            manhi <= conv_std_logic_vector(12264615,24);
            manlo <= conv_std_logic_vector(87551554,28);
            exponent <= conv_std_logic_vector(461,11);
      WHEN "0110000110" =>
            manhi <= conv_std_logic_vector(4590569,24);
            manlo <= conv_std_logic_vector(96025360,28);
            exponent <= conv_std_logic_vector(460,11);
      WHEN "0110000111" =>
            manhi <= conv_std_logic_vector(14665859,24);
            manlo <= conv_std_logic_vector(200220878,28);
            exponent <= conv_std_logic_vector(458,11);
      WHEN "0110001000" =>
            manhi <= conv_std_logic_vector(6357306,24);
            manlo <= conv_std_logic_vector(71997608,28);
            exponent <= conv_std_logic_vector(457,11);
      WHEN "0110001001" =>
            manhi <= conv_std_logic_vector(244214,24);
            manlo <= conv_std_logic_vector(66463607,28);
            exponent <= conv_std_logic_vector(456,11);
      WHEN "0110001010" =>
            manhi <= conv_std_logic_vector(8270120,24);
            manlo <= conv_std_logic_vector(265669912,28);
            exponent <= conv_std_logic_vector(454,11);
      WHEN "0110001011" =>
            manhi <= conv_std_logic_vector(1651584,24);
            manlo <= conv_std_logic_vector(179638473,28);
            exponent <= conv_std_logic_vector(453,11);
      WHEN "0110001100" =>
            manhi <= conv_std_logic_vector(10341091,24);
            manlo <= conv_std_logic_vector(152092530,28);
            exponent <= conv_std_logic_vector(451,11);
      WHEN "0110001101" =>
            manhi <= conv_std_logic_vector(3175319,24);
            manlo <= conv_std_logic_vector(178838140,28);
            exponent <= conv_std_logic_vector(450,11);
      WHEN "0110001110" =>
            manhi <= conv_std_logic_vector(12583294,24);
            manlo <= conv_std_logic_vector(183442082,28);
            exponent <= conv_std_logic_vector(448,11);
      WHEN "0110001111" =>
            manhi <= conv_std_logic_vector(4825040,24);
            manlo <= conv_std_logic_vector(141040370,28);
            exponent <= conv_std_logic_vector(447,11);
      WHEN "0110010000" =>
            manhi <= conv_std_logic_vector(15010888,24);
            manlo <= conv_std_logic_vector(62934477,28);
            exponent <= conv_std_logic_vector(445,11);
      WHEN "0110010001" =>
            manhi <= conv_std_logic_vector(6611164,24);
            manlo <= conv_std_logic_vector(11633311,28);
            exponent <= conv_std_logic_vector(444,11);
      WHEN "0110010010" =>
            manhi <= conv_std_logic_vector(430992,24);
            manlo <= conv_std_logic_vector(96770068,28);
            exponent <= conv_std_logic_vector(443,11);
      WHEN "0110010011" =>
            manhi <= conv_std_logic_vector(8544968,24);
            manlo <= conv_std_logic_vector(80768180,28);
            exponent <= conv_std_logic_vector(441,11);
      WHEN "0110010100" =>
            manhi <= conv_std_logic_vector(1853806,24);
            manlo <= conv_std_logic_vector(5288079,28);
            exponent <= conv_std_logic_vector(440,11);
      WHEN "0110010101" =>
            manhi <= conv_std_logic_vector(10638663,24);
            manlo <= conv_std_logic_vector(235213815,28);
            exponent <= conv_std_logic_vector(438,11);
      WHEN "0110010110" =>
            manhi <= conv_std_logic_vector(3394261,24);
            manlo <= conv_std_logic_vector(36557939,28);
            exponent <= conv_std_logic_vector(437,11);
      WHEN "0110010111" =>
            manhi <= conv_std_logic_vector(12905470,24);
            manlo <= conv_std_logic_vector(253900977,28);
            exponent <= conv_std_logic_vector(435,11);
      WHEN "0110011000" =>
            manhi <= conv_std_logic_vector(5062084,24);
            manlo <= conv_std_logic_vector(153603034,28);
            exponent <= conv_std_logic_vector(434,11);
      WHEN "0110011001" =>
            manhi <= conv_std_logic_vector(15359702,24);
            manlo <= conv_std_logic_vector(204098933,28);
            exponent <= conv_std_logic_vector(432,11);
      WHEN "0110011010" =>
            manhi <= conv_std_logic_vector(6867807,24);
            manlo <= conv_std_logic_vector(115170312,28);
            exponent <= conv_std_logic_vector(431,11);
      WHEN "0110011011" =>
            manhi <= conv_std_logic_vector(619820,24);
            manlo <= conv_std_logic_vector(2986045,28);
            exponent <= conv_std_logic_vector(430,11);
      WHEN "0110011100" =>
            manhi <= conv_std_logic_vector(8822831,24);
            manlo <= conv_std_logic_vector(145826716,28);
            exponent <= conv_std_logic_vector(428,11);
      WHEN "0110011101" =>
            manhi <= conv_std_logic_vector(2058246,24);
            manlo <= conv_std_logic_vector(98876593,28);
            exponent <= conv_std_logic_vector(427,11);
      WHEN "0110011110" =>
            manhi <= conv_std_logic_vector(10939501,24);
            manlo <= conv_std_logic_vector(129141213,28);
            exponent <= conv_std_logic_vector(425,11);
      WHEN "0110011111" =>
            manhi <= conv_std_logic_vector(3615605,24);
            manlo <= conv_std_logic_vector(20427716,28);
            exponent <= conv_std_logic_vector(424,11);
      WHEN "0110100000" =>
            manhi <= conv_std_logic_vector(13231182,24);
            manlo <= conv_std_logic_vector(130335695,28);
            exponent <= conv_std_logic_vector(422,11);
      WHEN "0110100001" =>
            manhi <= conv_std_logic_vector(5301729,24);
            manlo <= conv_std_logic_vector(196124198,28);
            exponent <= conv_std_logic_vector(421,11);
      WHEN "0110100010" =>
            manhi <= conv_std_logic_vector(15712344,24);
            manlo <= conv_std_logic_vector(233039482,28);
            exponent <= conv_std_logic_vector(419,11);
      WHEN "0110100011" =>
            manhi <= conv_std_logic_vector(7127266,24);
            manlo <= conv_std_logic_vector(266329205,28);
            exponent <= conv_std_logic_vector(418,11);
      WHEN "0110100100" =>
            manhi <= conv_std_logic_vector(810719,24);
            manlo <= conv_std_logic_vector(185030259,28);
            exponent <= conv_std_logic_vector(417,11);
      WHEN "0110100101" =>
            manhi <= conv_std_logic_vector(9103743,24);
            manlo <= conv_std_logic_vector(217685905,28);
            exponent <= conv_std_logic_vector(415,11);
      WHEN "0110100110" =>
            manhi <= conv_std_logic_vector(2264930,24);
            manlo <= conv_std_logic_vector(17303531,28);
            exponent <= conv_std_logic_vector(414,11);
      WHEN "0110100111" =>
            manhi <= conv_std_logic_vector(11243640,24);
            manlo <= conv_std_logic_vector(56799625,28);
            exponent <= conv_std_logic_vector(412,11);
      WHEN "0110101000" =>
            manhi <= conv_std_logic_vector(3839377,24);
            manlo <= conv_std_logic_vector(227776580,28);
            exponent <= conv_std_logic_vector(411,11);
      WHEN "0110101001" =>
            manhi <= conv_std_logic_vector(13560468,24);
            manlo <= conv_std_logic_vector(25616516,28);
            exponent <= conv_std_logic_vector(409,11);
      WHEN "0110101010" =>
            manhi <= conv_std_logic_vector(5544004,24);
            manlo <= conv_std_logic_vector(145740137,28);
            exponent <= conv_std_logic_vector(408,11);
      WHEN "0110101011" =>
            manhi <= conv_std_logic_vector(16068856,24);
            manlo <= conv_std_logic_vector(149889545,28);
            exponent <= conv_std_logic_vector(406,11);
      WHEN "0110101100" =>
            manhi <= conv_std_logic_vector(7389573,24);
            manlo <= conv_std_logic_vector(170431948,28);
            exponent <= conv_std_logic_vector(405,11);
      WHEN "0110101101" =>
            manhi <= conv_std_logic_vector(1003714,24);
            manlo <= conv_std_logic_vector(35324999,28);
            exponent <= conv_std_logic_vector(404,11);
      WHEN "0110101110" =>
            manhi <= conv_std_logic_vector(9387738,24);
            manlo <= conv_std_logic_vector(150667400,28);
            exponent <= conv_std_logic_vector(402,11);
      WHEN "0110101111" =>
            manhi <= conv_std_logic_vector(2473881,24);
            manlo <= conv_std_logic_vector(194497484,28);
            exponent <= conv_std_logic_vector(401,11);
      WHEN "0110110000" =>
            manhi <= conv_std_logic_vector(11551116,24);
            manlo <= conv_std_logic_vector(78219737,28);
            exponent <= conv_std_logic_vector(399,11);
      WHEN "0110110001" =>
            manhi <= conv_std_logic_vector(4065606,24);
            manlo <= conv_std_logic_vector(28280174,28);
            exponent <= conv_std_logic_vector(398,11);
      WHEN "0110110010" =>
            manhi <= conv_std_logic_vector(13893366,24);
            manlo <= conv_std_logic_vector(266881350,28);
            exponent <= conv_std_logic_vector(396,11);
      WHEN "0110110011" =>
            manhi <= conv_std_logic_vector(5788937,24);
            manlo <= conv_std_logic_vector(232096008,28);
            exponent <= conv_std_logic_vector(395,11);
      WHEN "0110110100" =>
            manhi <= conv_std_logic_vector(16429280,24);
            manlo <= conv_std_logic_vector(78498076,28);
            exponent <= conv_std_logic_vector(393,11);
      WHEN "0110110101" =>
            manhi <= conv_std_logic_vector(7654758,24);
            manlo <= conv_std_logic_vector(160696217,28);
            exponent <= conv_std_logic_vector(392,11);
      WHEN "0110110110" =>
            manhi <= conv_std_logic_vector(1198826,24);
            manlo <= conv_std_logic_vector(87006684,28);
            exponent <= conv_std_logic_vector(391,11);
      WHEN "0110110111" =>
            manhi <= conv_std_logic_vector(9674849,24);
            manlo <= conv_std_logic_vector(166079254,28);
            exponent <= conv_std_logic_vector(389,11);
      WHEN "0110111000" =>
            manhi <= conv_std_logic_vector(2685126,24);
            manlo <= conv_std_logic_vector(63154951,28);
            exponent <= conv_std_logic_vector(388,11);
      WHEN "0110111001" =>
            manhi <= conv_std_logic_vector(11861966,24);
            manlo <= conv_std_logic_vector(91696135,28);
            exponent <= conv_std_logic_vector(386,11);
      WHEN "0110111010" =>
            manhi <= conv_std_logic_vector(4294316,24);
            manlo <= conv_std_logic_vector(212296424,28);
            exponent <= conv_std_logic_vector(385,11);
      WHEN "0110111011" =>
            manhi <= conv_std_logic_vector(14229918,24);
            manlo <= conv_std_logic_vector(223047784,28);
            exponent <= conv_std_logic_vector(383,11);
      WHEN "0110111100" =>
            manhi <= conv_std_logic_vector(6036558,24);
            manlo <= conv_std_logic_vector(232962025,28);
            exponent <= conv_std_logic_vector(382,11);
      WHEN "0110111101" =>
            manhi <= conv_std_logic_vector(8221,24);
            manlo <= conv_std_logic_vector(133893557,28);
            exponent <= conv_std_logic_vector(381,11);
      WHEN "0110111110" =>
            manhi <= conv_std_logic_vector(7922853,24);
            manlo <= conv_std_logic_vector(125492404,28);
            exponent <= conv_std_logic_vector(379,11);
      WHEN "0110111111" =>
            manhi <= conv_std_logic_vector(1396079,24);
            manlo <= conv_std_logic_vector(135612572,28);
            exponent <= conv_std_logic_vector(378,11);
      WHEN "0111000000" =>
            manhi <= conv_std_logic_vector(9965111,24);
            manlo <= conv_std_logic_vector(47990958,28);
            exponent <= conv_std_logic_vector(376,11);
      WHEN "0111000001" =>
            manhi <= conv_std_logic_vector(2898688,24);
            manlo <= conv_std_logic_vector(203019642,28);
            exponent <= conv_std_logic_vector(375,11);
      WHEN "0111000010" =>
            manhi <= conv_std_logic_vector(12176227,24);
            manlo <= conv_std_logic_vector(103393586,28);
            exponent <= conv_std_logic_vector(373,11);
      WHEN "0111000011" =>
            manhi <= conv_std_logic_vector(4525537,24);
            manlo <= conv_std_logic_vector(38936964,28);
            exponent <= conv_std_logic_vector(372,11);
      WHEN "0111000100" =>
            manhi <= conv_std_logic_vector(14570163,24);
            manlo <= conv_std_logic_vector(185128905,28);
            exponent <= conv_std_logic_vector(370,11);
      WHEN "0111000101" =>
            manhi <= conv_std_logic_vector(6286897,24);
            manlo <= conv_std_logic_vector(12037044,28);
            exponent <= conv_std_logic_vector(369,11);
      WHEN "0111000110" =>
            manhi <= conv_std_logic_vector(192410,24);
            manlo <= conv_std_logic_vector(9691196,28);
            exponent <= conv_std_logic_vector(368,11);
      WHEN "0111000111" =>
            manhi <= conv_std_logic_vector(8193890,24);
            manlo <= conv_std_logic_vector(46224319,28);
            exponent <= conv_std_logic_vector(366,11);
      WHEN "0111001000" =>
            manhi <= conv_std_logic_vector(1595497,24);
            manlo <= conv_std_logic_vector(45130080,28);
            exponent <= conv_std_logic_vector(365,11);
      WHEN "0111001001" =>
            manhi <= conv_std_logic_vector(10258557,24);
            manlo <= conv_std_logic_vector(218068546,28);
            exponent <= conv_std_logic_vector(363,11);
      WHEN "0111001010" =>
            manhi <= conv_std_logic_vector(3114594,24);
            manlo <= conv_std_logic_vector(194203222,28);
            exponent <= conv_std_logic_vector(362,11);
      WHEN "0111001011" =>
            manhi <= conv_std_logic_vector(12493936,24);
            manlo <= conv_std_logic_vector(228530713,28);
            exponent <= conv_std_logic_vector(360,11);
      WHEN "0111001100" =>
            manhi <= conv_std_logic_vector(4759294,24);
            manlo <= conv_std_logic_vector(189728046,28);
            exponent <= conv_std_logic_vector(359,11);
      WHEN "0111001101" =>
            manhi <= conv_std_logic_vector(14914142,24);
            manlo <= conv_std_logic_vector(25337562,28);
            exponent <= conv_std_logic_vector(357,11);
      WHEN "0111001110" =>
            manhi <= conv_std_logic_vector(6539982,24);
            manlo <= conv_std_logic_vector(56762382,28);
            exponent <= conv_std_logic_vector(356,11);
      WHEN "0111001111" =>
            manhi <= conv_std_logic_vector(378619,24);
            manlo <= conv_std_logic_vector(186677702,28);
            exponent <= conv_std_logic_vector(355,11);
      WHEN "0111010000" =>
            manhi <= conv_std_logic_vector(8467900,24);
            manlo <= conv_std_logic_vector(266785510,28);
            exponent <= conv_std_logic_vector(353,11);
      WHEN "0111010001" =>
            manhi <= conv_std_logic_vector(1797103,24);
            manlo <= conv_std_logic_vector(17183357,28);
            exponent <= conv_std_logic_vector(352,11);
      WHEN "0111010010" =>
            manhi <= conv_std_logic_vector(10555224,24);
            manlo <= conv_std_logic_vector(126067134,28);
            exponent <= conv_std_logic_vector(350,11);
      WHEN "0111010011" =>
            manhi <= conv_std_logic_vector(3332869,24);
            manlo <= conv_std_logic_vector(228611260,28);
            exponent <= conv_std_logic_vector(349,11);
      WHEN "0111010100" =>
            manhi <= conv_std_logic_vector(12815132,24);
            manlo <= conv_std_logic_vector(155705738,28);
            exponent <= conv_std_logic_vector(347,11);
      WHEN "0111010101" =>
            manhi <= conv_std_logic_vector(4995617,24);
            manlo <= conv_std_logic_vector(85136440,28);
            exponent <= conv_std_logic_vector(346,11);
      WHEN "0111010110" =>
            manhi <= conv_std_logic_vector(15261895,24);
            manlo <= conv_std_logic_vector(3688335,28);
            exponent <= conv_std_logic_vector(344,11);
      WHEN "0111010111" =>
            manhi <= conv_std_logic_vector(6795844,24);
            manlo <= conv_std_logic_vector(137097782,28);
            exponent <= conv_std_logic_vector(343,11);
      WHEN "0111011000" =>
            manhi <= conv_std_logic_vector(566872,24);
            manlo <= conv_std_logic_vector(175764875,28);
            exponent <= conv_std_logic_vector(342,11);
      WHEN "0111011001" =>
            manhi <= conv_std_logic_vector(8744918,24);
            manlo <= conv_std_logic_vector(152414052,28);
            exponent <= conv_std_logic_vector(340,11);
      WHEN "0111011010" =>
            manhi <= conv_std_logic_vector(2000921,24);
            manlo <= conv_std_logic_vector(54921723,28);
            exponent <= conv_std_logic_vector(339,11);
      WHEN "0111011011" =>
            manhi <= conv_std_logic_vector(10855146,24);
            manlo <= conv_std_logic_vector(129996510,28);
            exponent <= conv_std_logic_vector(337,11);
      WHEN "0111011100" =>
            manhi <= conv_std_logic_vector(3553540,24);
            manlo <= conv_std_logic_vector(37023540,28);
            exponent <= conv_std_logic_vector(336,11);
      WHEN "0111011101" =>
            manhi <= conv_std_logic_vector(13139852,24);
            manlo <= conv_std_logic_vector(221848100,28);
            exponent <= conv_std_logic_vector(334,11);
      WHEN "0111011110" =>
            manhi <= conv_std_logic_vector(5234533,24);
            manlo <= conv_std_logic_vector(32943194,28);
            exponent <= conv_std_logic_vector(333,11);
      WHEN "0111011111" =>
            manhi <= conv_std_logic_vector(15613463,24);
            manlo <= conv_std_logic_vector(232436445,28);
            exponent <= conv_std_logic_vector(331,11);
      WHEN "0111100000" =>
            manhi <= conv_std_logic_vector(7054514,24);
            manlo <= conv_std_logic_vector(111791498,28);
            exponent <= conv_std_logic_vector(330,11);
      WHEN "0111100001" =>
            manhi <= conv_std_logic_vector(757191,24);
            manlo <= conv_std_logic_vector(90062360,28);
            exponent <= conv_std_logic_vector(329,11);
      WHEN "0111100010" =>
            manhi <= conv_std_logic_vector(9024975,24);
            manlo <= conv_std_logic_vector(238219590,28);
            exponent <= conv_std_logic_vector(327,11);
      WHEN "0111100011" =>
            manhi <= conv_std_logic_vector(2206975,24);
            manlo <= conv_std_logic_vector(232222812,28);
            exponent <= conv_std_logic_vector(326,11);
      WHEN "0111100100" =>
            manhi <= conv_std_logic_vector(11158359,24);
            manlo <= conv_std_logic_vector(155073518,28);
            exponent <= conv_std_logic_vector(324,11);
      WHEN "0111100101" =>
            manhi <= conv_std_logic_vector(3776631,24);
            manlo <= conv_std_logic_vector(232102510,28);
            exponent <= conv_std_logic_vector(323,11);
      WHEN "0111100110" =>
            manhi <= conv_std_logic_vector(13468136,24);
            manlo <= conv_std_logic_vector(71264246,28);
            exponent <= conv_std_logic_vector(321,11);
      WHEN "0111100111" =>
            manhi <= conv_std_logic_vector(5476070,24);
            manlo <= conv_std_logic_vector(155401688,28);
            exponent <= conv_std_logic_vector(320,11);
      WHEN "0111101000" =>
            manhi <= conv_std_logic_vector(15968890,24);
            manlo <= conv_std_logic_vector(140531032,28);
            exponent <= conv_std_logic_vector(318,11);
      WHEN "0111101001" =>
            manhi <= conv_std_logic_vector(7316022,24);
            manlo <= conv_std_logic_vector(197790036,28);
            exponent <= conv_std_logic_vector(317,11);
      WHEN "0111101010" =>
            manhi <= conv_std_logic_vector(949598,24);
            manlo <= conv_std_logic_vector(108723575,28);
            exponent <= conv_std_logic_vector(316,11);
      WHEN "0111101011" =>
            manhi <= conv_std_logic_vector(9308106,24);
            manlo <= conv_std_logic_vector(82754530,28);
            exponent <= conv_std_logic_vector(314,11);
      WHEN "0111101100" =>
            manhi <= conv_std_logic_vector(2415291,24);
            manlo <= conv_std_logic_vector(157597766,28);
            exponent <= conv_std_logic_vector(313,11);
      WHEN "0111101101" =>
            manhi <= conv_std_logic_vector(11464899,24);
            manlo <= conv_std_logic_vector(231735034,28);
            exponent <= conv_std_logic_vector(311,11);
      WHEN "0111101110" =>
            manhi <= conv_std_logic_vector(4002171,24);
            manlo <= conv_std_logic_vector(161749904,28);
            exponent <= conv_std_logic_vector(310,11);
      WHEN "0111101111" =>
            manhi <= conv_std_logic_vector(13800021,24);
            manlo <= conv_std_logic_vector(267486845,28);
            exponent <= conv_std_logic_vector(308,11);
      WHEN "0111110000" =>
            manhi <= conv_std_logic_vector(5720258,24);
            manlo <= conv_std_logic_vector(121711942,28);
            exponent <= conv_std_logic_vector(307,11);
      WHEN "0111110001" =>
            manhi <= conv_std_logic_vector(16328217,24);
            manlo <= conv_std_logic_vector(85566619,28);
            exponent <= conv_std_logic_vector(305,11);
      WHEN "0111110010" =>
            manhi <= conv_std_logic_vector(7580400,24);
            manlo <= conv_std_logic_vector(165916765,28);
            exponent <= conv_std_logic_vector(304,11);
      WHEN "0111110011" =>
            manhi <= conv_std_logic_vector(1144116,24);
            manlo <= conv_std_logic_vector(209234965,28);
            exponent <= conv_std_logic_vector(303,11);
      WHEN "0111110100" =>
            manhi <= conv_std_logic_vector(9594343,24);
            manlo <= conv_std_logic_vector(148128653,28);
            exponent <= conv_std_logic_vector(301,11);
      WHEN "0111110101" =>
            manhi <= conv_std_logic_vector(2625893,24);
            manlo <= conv_std_logic_vector(48717694,28);
            exponent <= conv_std_logic_vector(300,11);
      WHEN "0111110110" =>
            manhi <= conv_std_logic_vector(11774803,24);
            manlo <= conv_std_logic_vector(228357100,28);
            exponent <= conv_std_logic_vector(298,11);
      WHEN "0111110111" =>
            manhi <= conv_std_logic_vector(4230186,24);
            manlo <= conv_std_logic_vector(57439900,28);
            exponent <= conv_std_logic_vector(297,11);
      WHEN "0111111000" =>
            manhi <= conv_std_logic_vector(14135549,24);
            manlo <= conv_std_logic_vector(147041206,28);
            exponent <= conv_std_logic_vector(295,11);
      WHEN "0111111001" =>
            manhi <= conv_std_logic_vector(5967125,24);
            manlo <= conv_std_logic_vector(222682176,28);
            exponent <= conv_std_logic_vector(294,11);
      WHEN "0111111010" =>
            manhi <= conv_std_logic_vector(16691487,24);
            manlo <= conv_std_logic_vector(12959237,28);
            exponent <= conv_std_logic_vector(292,11);
      WHEN "0111111011" =>
            manhi <= conv_std_logic_vector(7847679,24);
            manlo <= conv_std_logic_vector(147174066,28);
            exponent <= conv_std_logic_vector(291,11);
      WHEN "0111111100" =>
            manhi <= conv_std_logic_vector(1340769,24);
            manlo <= conv_std_logic_vector(168148656,28);
            exponent <= conv_std_logic_vector(290,11);
      WHEN "0111111101" =>
            manhi <= conv_std_logic_vector(9883721,24);
            manlo <= conv_std_logic_vector(190474495,28);
            exponent <= conv_std_logic_vector(288,11);
      WHEN "0111111110" =>
            manhi <= conv_std_logic_vector(2838805,24);
            manlo <= conv_std_logic_vector(196335986,28);
            exponent <= conv_std_logic_vector(287,11);
      WHEN "0111111111" =>
            manhi <= conv_std_logic_vector(12088108,24);
            manlo <= conv_std_logic_vector(120857634,28);
            exponent <= conv_std_logic_vector(285,11);
      WHEN "1000000000" =>
            manhi <= conv_std_logic_vector(4460702,24);
            manlo <= conv_std_logic_vector(229771569,28);
            exponent <= conv_std_logic_vector(284,11);
      WHEN "1000000001" =>
            manhi <= conv_std_logic_vector(14474758,24);
            manlo <= conv_std_logic_vector(236628147,28);
            exponent <= conv_std_logic_vector(282,11);
      WHEN "1000000010" =>
            manhi <= conv_std_logic_vector(6216702,24);
            manlo <= conv_std_logic_vector(29481361,28);
            exponent <= conv_std_logic_vector(281,11);
      WHEN "1000000011" =>
            manhi <= conv_std_logic_vector(140763,24);
            manlo <= conv_std_logic_vector(131310533,28);
            exponent <= conv_std_logic_vector(280,11);
      WHEN "1000000100" =>
            manhi <= conv_std_logic_vector(8117891,24);
            manlo <= conv_std_logic_vector(96879140,28);
            exponent <= conv_std_logic_vector(278,11);
      WHEN "1000000101" =>
            manhi <= conv_std_logic_vector(1539580,24);
            manlo <= conv_std_logic_vector(98694067,28);
            exponent <= conv_std_logic_vector(277,11);
      WHEN "1000000110" =>
            manhi <= conv_std_logic_vector(10176275,24);
            manlo <= conv_std_logic_vector(66343668,28);
            exponent <= conv_std_logic_vector(275,11);
      WHEN "1000000111" =>
            manhi <= conv_std_logic_vector(3054054,24);
            manlo <= conv_std_logic_vector(159783892,28);
            exponent <= conv_std_logic_vector(274,11);
      WHEN "1000001000" =>
            manhi <= conv_std_logic_vector(12404850,24);
            manlo <= conv_std_logic_vector(262311967,28);
            exponent <= conv_std_logic_vector(272,11);
      WHEN "1000001001" =>
            manhi <= conv_std_logic_vector(4693748,24);
            manlo <= conv_std_logic_vector(264030756,28);
            exponent <= conv_std_logic_vector(271,11);
      WHEN "1000001010" =>
            manhi <= conv_std_logic_vector(14817690,24);
            manlo <= conv_std_logic_vector(106917994,28);
            exponent <= conv_std_logic_vector(269,11);
      WHEN "1000001011" =>
            manhi <= conv_std_logic_vector(6469017,24);
            manlo <= conv_std_logic_vector(5191992,28);
            exponent <= conv_std_logic_vector(268,11);
      WHEN "1000001100" =>
            manhi <= conv_std_logic_vector(326406,24);
            manlo <= conv_std_logic_vector(114083215,28);
            exponent <= conv_std_logic_vector(267,11);
      WHEN "1000001101" =>
            manhi <= conv_std_logic_vector(8391068,24);
            manlo <= conv_std_logic_vector(64117214,28);
            exponent <= conv_std_logic_vector(265,11);
      WHEN "1000001110" =>
            manhi <= conv_std_logic_vector(1740572,24);
            manlo <= conv_std_logic_vector(183091279,28);
            exponent <= conv_std_logic_vector(264,11);
      WHEN "1000001111" =>
            manhi <= conv_std_logic_vector(10472039,24);
            manlo <= conv_std_logic_vector(2244224,28);
            exponent <= conv_std_logic_vector(262,11);
      WHEN "1000010000" =>
            manhi <= conv_std_logic_vector(3271665,24);
            manlo <= conv_std_logic_vector(109958542,28);
            exponent <= conv_std_logic_vector(261,11);
      WHEN "1000010001" =>
            manhi <= conv_std_logic_vector(12725069,24);
            manlo <= conv_std_logic_vector(41968573,28);
            exponent <= conv_std_logic_vector(259,11);
      WHEN "1000010010" =>
            manhi <= conv_std_logic_vector(4929352,24);
            manlo <= conv_std_logic_vector(94809674,28);
            exponent <= conv_std_logic_vector(258,11);
      WHEN "1000010011" =>
            manhi <= conv_std_logic_vector(15164384,24);
            manlo <= conv_std_logic_vector(252890425,28);
            exponent <= conv_std_logic_vector(256,11);
      WHEN "1000010100" =>
            manhi <= conv_std_logic_vector(6724100,24);
            manlo <= conv_std_logic_vector(163583158,28);
            exponent <= conv_std_logic_vector(255,11);
      WHEN "1000010101" =>
            manhi <= conv_std_logic_vector(514086,24);
            manlo <= conv_std_logic_vector(118679222,28);
            exponent <= conv_std_logic_vector(254,11);
      WHEN "1000010110" =>
            manhi <= conv_std_logic_vector(8667242,24);
            manlo <= conv_std_logic_vector(192770478,28);
            exponent <= conv_std_logic_vector(252,11);
      WHEN "1000010111" =>
            manhi <= conv_std_logic_vector(1943770,24);
            manlo <= conv_std_logic_vector(136437165,28);
            exponent <= conv_std_logic_vector(251,11);
      WHEN "1000011000" =>
            manhi <= conv_std_logic_vector(10771048,24);
            manlo <= conv_std_logic_vector(58883744,28);
            exponent <= conv_std_logic_vector(249,11);
      WHEN "1000011001" =>
            manhi <= conv_std_logic_vector(3491664,24);
            manlo <= conv_std_logic_vector(24836209,28);
            exponent <= conv_std_logic_vector(248,11);
      WHEN "1000011010" =>
            manhi <= conv_std_logic_vector(13048801,24);
            manlo <= conv_std_logic_vector(33938829,28);
            exponent <= conv_std_logic_vector(246,11);
      WHEN "1000011011" =>
            manhi <= conv_std_logic_vector(5167541,24);
            manlo <= conv_std_logic_vector(6894318,28);
            exponent <= conv_std_logic_vector(245,11);
      WHEN "1000011100" =>
            manhi <= conv_std_logic_vector(15514883,24);
            manlo <= conv_std_logic_vector(216092120,28);
            exponent <= conv_std_logic_vector(243,11);
      WHEN "1000011101" =>
            manhi <= conv_std_logic_vector(6981983,24);
            manlo <= conv_std_logic_vector(70071320,28);
            exponent <= conv_std_logic_vector(242,11);
      WHEN "1000011110" =>
            manhi <= conv_std_logic_vector(703825,24);
            manlo <= conv_std_logic_vector(239890498,28);
            exponent <= conv_std_logic_vector(241,11);
      WHEN "1000011111" =>
            manhi <= conv_std_logic_vector(8946447,24);
            manlo <= conv_std_logic_vector(185687386,28);
            exponent <= conv_std_logic_vector(239,11);
      WHEN "1000100000" =>
            manhi <= conv_std_logic_vector(2149198,24);
            manlo <= conv_std_logic_vector(12777107,28);
            exponent <= conv_std_logic_vector(238,11);
      WHEN "1000100001" =>
            manhi <= conv_std_logic_vector(11073338,24);
            manlo <= conv_std_logic_vector(132295567,28);
            exponent <= conv_std_logic_vector(236,11);
      WHEN "1000100010" =>
            manhi <= conv_std_logic_vector(3714076,24);
            manlo <= conv_std_logic_vector(227171857,28);
            exponent <= conv_std_logic_vector(235,11);
      WHEN "1000100011" =>
            manhi <= conv_std_logic_vector(13376085,24);
            manlo <= conv_std_logic_vector(119368169,28);
            exponent <= conv_std_logic_vector(233,11);
      WHEN "1000100100" =>
            manhi <= conv_std_logic_vector(5408343,24);
            manlo <= conv_std_logic_vector(99290689,28);
            exponent <= conv_std_logic_vector(232,11);
      WHEN "1000100101" =>
            manhi <= conv_std_logic_vector(15869228,24);
            manlo <= conv_std_logic_vector(196569651,28);
            exponent <= conv_std_logic_vector(230,11);
      WHEN "1000100110" =>
            manhi <= conv_std_logic_vector(7242695,24);
            manlo <= conv_std_logic_vector(184868911,28);
            exponent <= conv_std_logic_vector(229,11);
      WHEN "1000100111" =>
            manhi <= conv_std_logic_vector(895647,24);
            manlo <= conv_std_logic_vector(101480846,28);
            exponent <= conv_std_logic_vector(228,11);
      WHEN "1000101000" =>
            manhi <= conv_std_logic_vector(9228716,24);
            manlo <= conv_std_logic_vector(111040654,28);
            exponent <= conv_std_logic_vector(226,11);
      WHEN "1000101001" =>
            manhi <= conv_std_logic_vector(2356879,24);
            manlo <= conv_std_logic_vector(205878747,28);
            exponent <= conv_std_logic_vector(225,11);
      WHEN "1000101010" =>
            manhi <= conv_std_logic_vector(11378945,24);
            manlo <= conv_std_logic_vector(223412824,28);
            exponent <= conv_std_logic_vector(223,11);
      WHEN "1000101011" =>
            manhi <= conv_std_logic_vector(3938930,24);
            manlo <= conv_std_logic_vector(43159582,28);
            exponent <= conv_std_logic_vector(222,11);
      WHEN "1000101100" =>
            manhi <= conv_std_logic_vector(13706961,24);
            manlo <= conv_std_logic_vector(24539717,28);
            exponent <= conv_std_logic_vector(220,11);
      WHEN "1000101101" =>
            manhi <= conv_std_logic_vector(5651788,24);
            manlo <= conv_std_logic_vector(17696328,28);
            exponent <= conv_std_logic_vector(219,11);
      WHEN "1000101110" =>
            manhi <= conv_std_logic_vector(16227461,24);
            manlo <= conv_std_logic_vector(248897772,28);
            exponent <= conv_std_logic_vector(217,11);
      WHEN "1000101111" =>
            manhi <= conv_std_logic_vector(7506268,24);
            manlo <= conv_std_logic_vector(253353585,28);
            exponent <= conv_std_logic_vector(216,11);
      WHEN "1000110000" =>
            manhi <= conv_std_logic_vector(1089573,24);
            manlo <= conv_std_logic_vector(199085712,28);
            exponent <= conv_std_logic_vector(215,11);
      WHEN "1000110001" =>
            manhi <= conv_std_logic_vector(9514082,24);
            manlo <= conv_std_logic_vector(134954983,28);
            exponent <= conv_std_logic_vector(213,11);
      WHEN "1000110010" =>
            manhi <= conv_std_logic_vector(2566840,24);
            manlo <= conv_std_logic_vector(107836942,28);
            exponent <= conv_std_logic_vector(212,11);
      WHEN "1000110011" =>
            manhi <= conv_std_logic_vector(11687906,24);
            manlo <= conv_std_logic_vector(170784064,28);
            exponent <= conv_std_logic_vector(210,11);
      WHEN "1000110100" =>
            manhi <= conv_std_logic_vector(4166250,24);
            manlo <= conv_std_logic_vector(219198631,28);
            exponent <= conv_std_logic_vector(209,11);
      WHEN "1000110101" =>
            manhi <= conv_std_logic_vector(14041467,24);
            manlo <= conv_std_logic_vector(127426909,28);
            exponent <= conv_std_logic_vector(207,11);
      WHEN "1000110110" =>
            manhi <= conv_std_logic_vector(5897904,24);
            manlo <= conv_std_logic_vector(29159081,28);
            exponent <= conv_std_logic_vector(206,11);
      WHEN "1000110111" =>
            manhi <= conv_std_logic_vector(16589626,24);
            manlo <= conv_std_logic_vector(15093248,28);
            exponent <= conv_std_logic_vector(204,11);
      WHEN "1000111000" =>
            manhi <= conv_std_logic_vector(7772734,24);
            manlo <= conv_std_logic_vector(112367334,28);
            exponent <= conv_std_logic_vector(203,11);
      WHEN "1000111001" =>
            manhi <= conv_std_logic_vector(1285628,24);
            manlo <= conv_std_logic_vector(21894417,28);
            exponent <= conv_std_logic_vector(202,11);
      WHEN "1000111010" =>
            manhi <= conv_std_logic_vector(9802579,24);
            manlo <= conv_std_logic_vector(254146435,28);
            exponent <= conv_std_logic_vector(200,11);
      WHEN "1000111011" =>
            manhi <= conv_std_logic_vector(2779104,24);
            manlo <= conv_std_logic_vector(257348234,28);
            exponent <= conv_std_logic_vector(199,11);
      WHEN "1000111100" =>
            manhi <= conv_std_logic_vector(12000257,24);
            manlo <= conv_std_logic_vector(188607876,28);
            exponent <= conv_std_logic_vector(197,11);
      WHEN "1000111101" =>
            manhi <= conv_std_logic_vector(4396065,24);
            manlo <= conv_std_logic_vector(238395052,28);
            exponent <= conv_std_logic_vector(196,11);
      WHEN "1000111110" =>
            manhi <= conv_std_logic_vector(14379644,24);
            manlo <= conv_std_logic_vector(116776141,28);
            exponent <= conv_std_logic_vector(194,11);
      WHEN "1000111111" =>
            manhi <= conv_std_logic_vector(6146720,24);
            manlo <= conv_std_logic_vector(217697734,28);
            exponent <= conv_std_logic_vector(193,11);
      WHEN "1001000000" =>
            manhi <= conv_std_logic_vector(89274,24);
            manlo <= conv_std_logic_vector(34078121,28);
            exponent <= conv_std_logic_vector(192,11);
      WHEN "1001000001" =>
            manhi <= conv_std_logic_vector(8042123,24);
            manlo <= conv_std_logic_vector(228091050,28);
            exponent <= conv_std_logic_vector(190,11);
      WHEN "1001000010" =>
            manhi <= conv_std_logic_vector(1483833,24);
            manlo <= conv_std_logic_vector(200872250,28);
            exponent <= conv_std_logic_vector(189,11);
      WHEN "1001000011" =>
            manhi <= conv_std_logic_vector(10094243,24);
            manlo <= conv_std_logic_vector(28573613,28);
            exponent <= conv_std_logic_vector(187,11);
      WHEN "1001000100" =>
            manhi <= conv_std_logic_vector(2993698,24);
            manlo <= conv_std_logic_vector(193026703,28);
            exponent <= conv_std_logic_vector(186,11);
      WHEN "1001000101" =>
            manhi <= conv_std_logic_vector(12316036,24);
            manlo <= conv_std_logic_vector(62602992,28);
            exponent <= conv_std_logic_vector(184,11);
      WHEN "1001000110" =>
            manhi <= conv_std_logic_vector(4628402,24);
            manlo <= conv_std_logic_vector(200475490,28);
            exponent <= conv_std_logic_vector(183,11);
      WHEN "1001000111" =>
            manhi <= conv_std_logic_vector(14721532,24);
            manlo <= conv_std_logic_vector(67122338,28);
            exponent <= conv_std_logic_vector(181,11);
      WHEN "1001001000" =>
            manhi <= conv_std_logic_vector(6398267,24);
            manlo <= conv_std_logic_vector(216803728,28);
            exponent <= conv_std_logic_vector(180,11);
      WHEN "1001001001" =>
            manhi <= conv_std_logic_vector(274352,24);
            manlo <= conv_std_logic_vector(17200594,28);
            exponent <= conv_std_logic_vector(179,11);
      WHEN "1001001010" =>
            manhi <= conv_std_logic_vector(8314469,24);
            manlo <= conv_std_logic_vector(86446456,28);
            exponent <= conv_std_logic_vector(177,11);
      WHEN "1001001011" =>
            manhi <= conv_std_logic_vector(1684214,24);
            manlo <= conv_std_logic_vector(93587914,28);
            exponent <= conv_std_logic_vector(176,11);
      WHEN "1001001100" =>
            manhi <= conv_std_logic_vector(10389106,24);
            manlo <= conv_std_logic_vector(193148951,28);
            exponent <= conv_std_logic_vector(174,11);
      WHEN "1001001101" =>
            manhi <= conv_std_logic_vector(3210647,24);
            manlo <= conv_std_logic_vector(64824977,28);
            exponent <= conv_std_logic_vector(173,11);
      WHEN "1001001110" =>
            manhi <= conv_std_logic_vector(12635279,24);
            manlo <= conv_std_logic_vector(224939505,28);
            exponent <= conv_std_logic_vector(171,11);
      WHEN "1001001111" =>
            manhi <= conv_std_logic_vector(4863289,24);
            manlo <= conv_std_logic_vector(17355920,28);
            exponent <= conv_std_logic_vector(170,11);
      WHEN "1001010000" =>
            manhi <= conv_std_logic_vector(15067171,24);
            manlo <= conv_std_logic_vector(171641236,28);
            exponent <= conv_std_logic_vector(168,11);
      WHEN "1001010001" =>
            manhi <= conv_std_logic_vector(6652575,24);
            manlo <= conv_std_logic_vector(15694991,28);
            exponent <= conv_std_logic_vector(167,11);
      WHEN "1001010010" =>
            manhi <= conv_std_logic_vector(461460,24);
            manlo <= conv_std_logic_vector(236949593,28);
            exponent <= conv_std_logic_vector(166,11);
      WHEN "1001010011" =>
            manhi <= conv_std_logic_vector(8589803,24);
            manlo <= conv_std_logic_vector(73170085,28);
            exponent <= conv_std_logic_vector(164,11);
      WHEN "1001010100" =>
            manhi <= conv_std_logic_vector(1886793,24);
            manlo <= conv_std_logic_vector(200887360,28);
            exponent <= conv_std_logic_vector(163,11);
      WHEN "1001010101" =>
            manhi <= conv_std_logic_vector(10687205,24);
            manlo <= conv_std_logic_vector(242930225,28);
            exponent <= conv_std_logic_vector(161,11);
      WHEN "1001010110" =>
            manhi <= conv_std_logic_vector(3429976,24);
            manlo <= conv_std_logic_vector(97980458,28);
            exponent <= conv_std_logic_vector(160,11);
      WHEN "1001010111" =>
            manhi <= conv_std_logic_vector(12958026,24);
            manlo <= conv_std_logic_vector(144828568,28);
            exponent <= conv_std_logic_vector(158,11);
      WHEN "1001011000" =>
            manhi <= conv_std_logic_vector(5100752,24);
            manlo <= conv_std_logic_vector(219332721,28);
            exponent <= conv_std_logic_vector(157,11);
      WHEN "1001011001" =>
            manhi <= conv_std_logic_vector(15416603,24);
            manlo <= conv_std_logic_vector(206580322,28);
            exponent <= conv_std_logic_vector(155,11);
      WHEN "1001011010" =>
            manhi <= conv_std_logic_vector(6909672,24);
            manlo <= conv_std_logic_vector(228709240,28);
            exponent <= conv_std_logic_vector(154,11);
      WHEN "1001011011" =>
            manhi <= conv_std_logic_vector(650622,24);
            manlo <= conv_std_logic_vector(232984198,28);
            exponent <= conv_std_logic_vector(153,11);
      WHEN "1001011100" =>
            manhi <= conv_std_logic_vector(8868158,24);
            manlo <= conv_std_logic_vector(132673062,28);
            exponent <= conv_std_logic_vector(151,11);
      WHEN "1001011101" =>
            manhi <= conv_std_logic_vector(2091596,24);
            manlo <= conv_std_logic_vector(20173170,28);
            exponent <= conv_std_logic_vector(150,11);
      WHEN "1001011110" =>
            manhi <= conv_std_logic_vector(10988576,24);
            manlo <= conv_std_logic_vector(44856082,28);
            exponent <= conv_std_logic_vector(148,11);
      WHEN "1001011111" =>
            manhi <= conv_std_logic_vector(3651712,24);
            manlo <= conv_std_logic_vector(56970522,28);
            exponent <= conv_std_logic_vector(147,11);
      WHEN "1001100000" =>
            manhi <= conv_std_logic_vector(13284314,24);
            manlo <= conv_std_logic_vector(208786223,28);
            exponent <= conv_std_logic_vector(145,11);
      WHEN "1001100001" =>
            manhi <= conv_std_logic_vector(5340822,24);
            manlo <= conv_std_logic_vector(76928898,28);
            exponent <= conv_std_logic_vector(144,11);
      WHEN "1001100010" =>
            manhi <= conv_std_logic_vector(15769870,24);
            manlo <= conv_std_logic_vector(69445892,28);
            exponent <= conv_std_logic_vector(142,11);
      WHEN "1001100011" =>
            manhi <= conv_std_logic_vector(7169591,24);
            manlo <= conv_std_logic_vector(217224162,28);
            exponent <= conv_std_logic_vector(141,11);
      WHEN "1001100100" =>
            manhi <= conv_std_logic_vector(841860,24);
            manlo <= conv_std_logic_vector(147476782,28);
            exponent <= conv_std_logic_vector(140,11);
      WHEN "1001100101" =>
            manhi <= conv_std_logic_vector(9149568,24);
            manlo <= conv_std_logic_vector(37524984,28);
            exponent <= conv_std_logic_vector(138,11);
      WHEN "1001100110" =>
            manhi <= conv_std_logic_vector(2298645,24);
            manlo <= conv_std_logic_vector(193659590,28);
            exponent <= conv_std_logic_vector(137,11);
      WHEN "1001100111" =>
            manhi <= conv_std_logic_vector(11293253,24);
            manlo <= conv_std_logic_vector(107316618,28);
            exponent <= conv_std_logic_vector(135,11);
      WHEN "1001101000" =>
            manhi <= conv_std_logic_vector(3875881,24);
            manlo <= conv_std_logic_vector(51654059,28);
            exponent <= conv_std_logic_vector(134,11);
      WHEN "1001101001" =>
            manhi <= conv_std_logic_vector(13614183,24);
            manlo <= conv_std_logic_vector(111249634,28);
            exponent <= conv_std_logic_vector(132,11);
      WHEN "1001101010" =>
            manhi <= conv_std_logic_vector(5583526,24);
            manlo <= conv_std_logic_vector(17717412,28);
            exponent <= conv_std_logic_vector(131,11);
      WHEN "1001101011" =>
            manhi <= conv_std_logic_vector(16127013,24);
            manlo <= conv_std_logic_vector(48769099,28);
            exponent <= conv_std_logic_vector(129,11);
      WHEN "1001101100" =>
            manhi <= conv_std_logic_vector(7432362,24);
            manlo <= conv_std_logic_vector(238120049,28);
            exponent <= conv_std_logic_vector(128,11);
      WHEN "1001101101" =>
            manhi <= conv_std_logic_vector(1035196,24);
            manlo <= conv_std_logic_vector(188962402,28);
            exponent <= conv_std_logic_vector(127,11);
      WHEN "1001101110" =>
            manhi <= conv_std_logic_vector(9434065,24);
            manlo <= conv_std_logic_vector(194820226,28);
            exponent <= conv_std_logic_vector(125,11);
      WHEN "1001101111" =>
            manhi <= conv_std_logic_vector(2507967,24);
            manlo <= conv_std_logic_vector(93233285,28);
            exponent <= conv_std_logic_vector(124,11);
      WHEN "1001110000" =>
            manhi <= conv_std_logic_vector(11601273,24);
            manlo <= conv_std_logic_vector(239123672,28);
            exponent <= conv_std_logic_vector(122,11);
      WHEN "1001110001" =>
            manhi <= conv_std_logic_vector(4102510,24);
            manlo <= conv_std_logic_vector(1244898,28);
            exponent <= conv_std_logic_vector(121,11);
      WHEN "1001110010" =>
            manhi <= conv_std_logic_vector(13947671,24);
            manlo <= conv_std_logic_vector(197996828,28);
            exponent <= conv_std_logic_vector(119,11);
      WHEN "1001110011" =>
            manhi <= conv_std_logic_vector(5828893,24);
            manlo <= conv_std_logic_vector(16622593,28);
            exponent <= conv_std_logic_vector(118,11);
      WHEN "1001110100" =>
            manhi <= conv_std_logic_vector(16488075,24);
            manlo <= conv_std_logic_vector(20144764,28);
            exponent <= conv_std_logic_vector(116,11);
      WHEN "1001110101" =>
            manhi <= conv_std_logic_vector(7698017,24);
            manlo <= conv_std_logic_vector(102592250,28);
            exponent <= conv_std_logic_vector(115,11);
      WHEN "1001110110" =>
            manhi <= conv_std_logic_vector(1230654,24);
            manlo <= conv_std_logic_vector(96196092,28);
            exponent <= conv_std_logic_vector(114,11);
      WHEN "1001110111" =>
            manhi <= conv_std_logic_vector(9721685,24);
            manlo <= conv_std_logic_vector(36636777,28);
            exponent <= conv_std_logic_vector(112,11);
      WHEN "1001111000" =>
            manhi <= conv_std_logic_vector(2719585,24);
            manlo <= conv_std_logic_vector(237160861,28);
            exponent <= conv_std_logic_vector(111,11);
      WHEN "1001111001" =>
            manhi <= conv_std_logic_vector(11912674,24);
            manlo <= conv_std_logic_vector(87541902,28);
            exponent <= conv_std_logic_vector(109,11);
      WHEN "1001111010" =>
            manhi <= conv_std_logic_vector(4331625,24);
            manlo <= conv_std_logic_vector(172036325,28);
            exponent <= conv_std_logic_vector(108,11);
      WHEN "1001111011" =>
            manhi <= conv_std_logic_vector(14284819,24);
            manlo <= conv_std_logic_vector(125225503,28);
            exponent <= conv_std_logic_vector(106,11);
      WHEN "1001111100" =>
            manhi <= conv_std_logic_vector(6076952,24);
            manlo <= conv_std_logic_vector(133715238,28);
            exponent <= conv_std_logic_vector(105,11);
      WHEN "1001111101" =>
            manhi <= conv_std_logic_vector(37941,24);
            manlo <= conv_std_logic_vector(126448851,28);
            exponent <= conv_std_logic_vector(104,11);
      WHEN "1001111110" =>
            manhi <= conv_std_logic_vector(7966586,24);
            manlo <= conv_std_logic_vector(250893596,28);
            exponent <= conv_std_logic_vector(102,11);
      WHEN "1001111111" =>
            manhi <= conv_std_logic_vector(1428256,24);
            manlo <= conv_std_logic_vector(212630882,28);
            exponent <= conv_std_logic_vector(101,11);
      WHEN "1010000000" =>
            manhi <= conv_std_logic_vector(10012460,24);
            manlo <= conv_std_logic_vector(168603206,28);
            exponent <= conv_std_logic_vector(99,11);
      WHEN "1010000001" =>
            manhi <= conv_std_logic_vector(2933526,24);
            manlo <= conv_std_logic_vector(143402282,28);
            exponent <= conv_std_logic_vector(98,11);
      WHEN "1010000010" =>
            manhi <= conv_std_logic_vector(12227491,24);
            manlo <= conv_std_logic_vector(213203509,28);
            exponent <= conv_std_logic_vector(96,11);
      WHEN "1010000011" =>
            manhi <= conv_std_logic_vector(4563255,24);
            manlo <= conv_std_logic_vector(104522224,28);
            exponent <= conv_std_logic_vector(95,11);
      WHEN "1010000100" =>
            manhi <= conv_std_logic_vector(14625666,24);
            manlo <= conv_std_logic_vector(203000190,28);
            exponent <= conv_std_logic_vector(93,11);
      WHEN "1010000101" =>
            manhi <= conv_std_logic_vector(6327733,24);
            manlo <= conv_std_logic_vector(246711469,28);
            exponent <= conv_std_logic_vector(92,11);
      WHEN "1010000110" =>
            manhi <= conv_std_logic_vector(222456,24);
            manlo <= conv_std_logic_vector(34640152,28);
            exponent <= conv_std_logic_vector(91,11);
      WHEN "1010000111" =>
            manhi <= conv_std_logic_vector(8238103,24);
            manlo <= conv_std_logic_vector(142733230,28);
            exponent <= conv_std_logic_vector(89,11);
      WHEN "1010001000" =>
            manhi <= conv_std_logic_vector(1628027,24);
            manlo <= conv_std_logic_vector(144984792,28);
            exponent <= conv_std_logic_vector(88,11);
      WHEN "1010001001" =>
            manhi <= conv_std_logic_vector(10306426,24);
            manlo <= conv_std_logic_vector(223510234,28);
            exponent <= conv_std_logic_vector(86,11);
      WHEN "1010001010" =>
            manhi <= conv_std_logic_vector(3149814,24);
            manlo <= conv_std_logic_vector(209464872,28);
            exponent <= conv_std_logic_vector(85,11);
      WHEN "1010001011" =>
            manhi <= conv_std_logic_vector(12545763,24);
            manlo <= conv_std_logic_vector(212245812,28);
            exponent <= conv_std_logic_vector(83,11);
      WHEN "1010001100" =>
            manhi <= conv_std_logic_vector(4797426,24);
            manlo <= conv_std_logic_vector(224882259,28);
            exponent <= conv_std_logic_vector(82,11);
      WHEN "1010001101" =>
            manhi <= conv_std_logic_vector(14970254,24);
            manlo <= conv_std_logic_vector(54358776,28);
            exponent <= conv_std_logic_vector(80,11);
      WHEN "1010001110" =>
            manhi <= conv_std_logic_vector(6581267,24);
            manlo <= conv_std_logic_vector(51917314,28);
            exponent <= conv_std_logic_vector(79,11);
      WHEN "1010001111" =>
            manhi <= conv_std_logic_vector(408995,24);
            manlo <= conv_std_logic_vector(130890803,28);
            exponent <= conv_std_logic_vector(78,11);
      WHEN "1010010000" =>
            manhi <= conv_std_logic_vector(8512599,24);
            manlo <= conv_std_logic_vector(137347476,28);
            exponent <= conv_std_logic_vector(76,11);
      WHEN "1010010001" =>
            manhi <= conv_std_logic_vector(1829990,24);
            manlo <= conv_std_logic_vector(106170554,28);
            exponent <= conv_std_logic_vector(75,11);
      WHEN "1010010010" =>
            manhi <= conv_std_logic_vector(10603618,24);
            manlo <= conv_std_logic_vector(204595238,28);
            exponent <= conv_std_logic_vector(73,11);
      WHEN "1010010011" =>
            manhi <= conv_std_logic_vector(3368476,24);
            manlo <= conv_std_logic_vector(102605239,28);
            exponent <= conv_std_logic_vector(72,11);
      WHEN "1010010100" =>
            manhi <= conv_std_logic_vector(12867528,24);
            manlo <= conv_std_logic_vector(59687307,28);
            exponent <= conv_std_logic_vector(70,11);
      WHEN "1010010101" =>
            manhi <= conv_std_logic_vector(5034167,24);
            manlo <= conv_std_logic_vector(235251142,28);
            exponent <= conv_std_logic_vector(69,11);
      WHEN "1010010110" =>
            manhi <= conv_std_logic_vector(15318622,24);
            manlo <= conv_std_logic_vector(227223140,28);
            exponent <= conv_std_logic_vector(67,11);
      WHEN "1010010111" =>
            manhi <= conv_std_logic_vector(6837582,24);
            manlo <= conv_std_logic_vector(138925467,28);
            exponent <= conv_std_logic_vector(66,11);
      WHEN "1010011000" =>
            manhi <= conv_std_logic_vector(597581,24);
            manlo <= conv_std_logic_vector(205088968,28);
            exponent <= conv_std_logic_vector(65,11);
      WHEN "1010011001" =>
            manhi <= conv_std_logic_vector(8790107,24);
            manlo <= conv_std_logic_vector(152356460,28);
            exponent <= conv_std_logic_vector(63,11);
      WHEN "1010011010" =>
            manhi <= conv_std_logic_vector(2034169,24);
            manlo <= conv_std_logic_vector(110749946,28);
            exponent <= conv_std_logic_vector(62,11);
      WHEN "1010011011" =>
            manhi <= conv_std_logic_vector(10904071,24);
            manlo <= conv_std_logic_vector(218226183,28);
            exponent <= conv_std_logic_vector(60,11);
      WHEN "1010011100" =>
            manhi <= conv_std_logic_vector(3589537,24);
            manlo <= conv_std_logic_vector(102830143,28);
            exponent <= conv_std_logic_vector(59,11);
      WHEN "1010011101" =>
            manhi <= conv_std_logic_vector(13192823,24);
            manlo <= conv_std_logic_vector(110639602,28);
            exponent <= conv_std_logic_vector(57,11);
      WHEN "1010011110" =>
            manhi <= conv_std_logic_vector(5273506,24);
            manlo <= conv_std_logic_vector(188352155,28);
            exponent <= conv_std_logic_vector(56,11);
      WHEN "1010011111" =>
            manhi <= conv_std_logic_vector(15670814,24);
            manlo <= conv_std_logic_vector(48227643,28);
            exponent <= conv_std_logic_vector(54,11);
      WHEN "1010100000" =>
            manhi <= conv_std_logic_vector(7096710,24);
            manlo <= conv_std_logic_vector(112532514,28);
            exponent <= conv_std_logic_vector(53,11);
      WHEN "1010100001" =>
            manhi <= conv_std_logic_vector(788237,24);
            manlo <= conv_std_logic_vector(112565412,28);
            exponent <= conv_std_logic_vector(52,11);
      WHEN "1010100010" =>
            manhi <= conv_std_logic_vector(9070660,24);
            manlo <= conv_std_logic_vector(201680253,28);
            exponent <= conv_std_logic_vector(50,11);
      WHEN "1010100011" =>
            manhi <= conv_std_logic_vector(2240588,24);
            manlo <= conv_std_logic_vector(244138286,28);
            exponent <= conv_std_logic_vector(49,11);
      WHEN "1010100100" =>
            manhi <= conv_std_logic_vector(11207821,24);
            manlo <= conv_std_logic_vector(206597824,28);
            exponent <= conv_std_logic_vector(47,11);
      WHEN "1010100101" =>
            manhi <= conv_std_logic_vector(3813024,24);
            manlo <= conv_std_logic_vector(29987310,28);
            exponent <= conv_std_logic_vector(46,11);
      WHEN "1010100110" =>
            manhi <= conv_std_logic_vector(13521688,24);
            manlo <= conv_std_logic_vector(27790821,28);
            exponent <= conv_std_logic_vector(44,11);
      WHEN "1010100111" =>
            manhi <= conv_std_logic_vector(5515471,24);
            manlo <= conv_std_logic_vector(219963166,28);
            exponent <= conv_std_logic_vector(43,11);
      WHEN "1010101000" =>
            manhi <= conv_std_logic_vector(16026870,24);
            manlo <= conv_std_logic_vector(39964772,28);
            exponent <= conv_std_logic_vector(41,11);
      WHEN "1010101001" =>
            manhi <= conv_std_logic_vector(7358681,24);
            manlo <= conv_std_logic_vector(204327682,28);
            exponent <= conv_std_logic_vector(40,11);
      WHEN "1010101010" =>
            manhi <= conv_std_logic_vector(980985,24);
            manlo <= conv_std_logic_vector(43247066,28);
            exponent <= conv_std_logic_vector(39,11);
      WHEN "1010101011" =>
            manhi <= conv_std_logic_vector(9354292,24);
            manlo <= conv_std_logic_vector(128160132,28);
            exponent <= conv_std_logic_vector(37,11);
      WHEN "1010101100" =>
            manhi <= conv_std_logic_vector(2449273,24);
            manlo <= conv_std_logic_vector(126511008,28);
            exponent <= conv_std_logic_vector(36,11);
      WHEN "1010101101" =>
            manhi <= conv_std_logic_vector(11514904,24);
            manlo <= conv_std_logic_vector(217311246,28);
            exponent <= conv_std_logic_vector(34,11);
      WHEN "1010101110" =>
            manhi <= conv_std_logic_vector(4038963,24);
            manlo <= conv_std_logic_vector(49913566,28);
            exponent <= conv_std_logic_vector(33,11);
      WHEN "1010101111" =>
            manhi <= conv_std_logic_vector(13854161,24);
            manlo <= conv_std_logic_vector(124821568,28);
            exponent <= conv_std_logic_vector(31,11);
      WHEN "1010110000" =>
            manhi <= conv_std_logic_vector(5760092,24);
            manlo <= conv_std_logic_vector(12957085,28);
            exponent <= conv_std_logic_vector(30,11);
      WHEN "1010110001" =>
            manhi <= conv_std_logic_vector(16386833,24);
            manlo <= conv_std_logic_vector(43278038,28);
            exponent <= conv_std_logic_vector(28,11);
      WHEN "1010110010" =>
            manhi <= conv_std_logic_vector(7623527,24);
            manlo <= conv_std_logic_vector(199937734,28);
            exponent <= conv_std_logic_vector(27,11);
      WHEN "1010110011" =>
            manhi <= conv_std_logic_vector(1175847,24);
            manlo <= conv_std_logic_vector(253947561,28);
            exponent <= conv_std_logic_vector(26,11);
      WHEN "1010110100" =>
            manhi <= conv_std_logic_vector(9641036,24);
            manlo <= conv_std_logic_vector(141497796,28);
            exponent <= conv_std_logic_vector(24,11);
      WHEN "1010110101" =>
            manhi <= conv_std_logic_vector(2660247,24);
            manlo <= conv_std_logic_vector(255766959,28);
            exponent <= conv_std_logic_vector(23,11);
      WHEN "1010110110" =>
            manhi <= conv_std_logic_vector(11825357,24);
            manlo <= conv_std_logic_vector(136095046,28);
            exponent <= conv_std_logic_vector(21,11);
      WHEN "1010110111" =>
            manhi <= conv_std_logic_vector(4267381,24);
            manlo <= conv_std_logic_vector(138414926,28);
            exponent <= conv_std_logic_vector(20,11);
      WHEN "1010111000" =>
            manhi <= conv_std_logic_vector(14190283,24);
            manlo <= conv_std_logic_vector(25479908,28);
            exponent <= conv_std_logic_vector(18,11);
      WHEN "1010111001" =>
            manhi <= conv_std_logic_vector(6007396,24);
            manlo <= conv_std_logic_vector(140400514,28);
            exponent <= conv_std_logic_vector(17,11);
      WHEN "1010111010" =>
            manhi <= conv_std_logic_vector(16750746,24);
            manlo <= conv_std_logic_vector(23924155,28);
            exponent <= conv_std_logic_vector(15,11);
      WHEN "1010111011" =>
            manhi <= conv_std_logic_vector(7891279,24);
            manlo <= conv_std_logic_vector(245330892,28);
            exponent <= conv_std_logic_vector(14,11);
      WHEN "1010111100" =>
            manhi <= conv_std_logic_vector(1372848,24);
            manlo <= conv_std_logic_vector(263794815,28);
            exponent <= conv_std_logic_vector(13,11);
      WHEN "1010111101" =>
            manhi <= conv_std_logic_vector(9930927,24);
            manlo <= conv_std_logic_vector(14029030,28);
            exponent <= conv_std_logic_vector(11,11);
      WHEN "1010111110" =>
            manhi <= conv_std_logic_vector(2873537,24);
            manlo <= conv_std_logic_vector(129274844,28);
            exponent <= conv_std_logic_vector(10,11);
      WHEN "1010111111" =>
            manhi <= conv_std_logic_vector(12139216,24);
            manlo <= conv_std_logic_vector(224845565,28);
            exponent <= conv_std_logic_vector(8,11);
      WHEN "1011000000" =>
            manhi <= conv_std_logic_vector(4498306,24);
            manlo <= conv_std_logic_vector(82126943,28);
            exponent <= conv_std_logic_vector(7,11);
      WHEN "1011000001" =>
            manhi <= conv_std_logic_vector(14530093,24);
            manlo <= conv_std_logic_vector(7024665,28);
            exponent <= conv_std_logic_vector(5,11);
      WHEN "1011000010" =>
            manhi <= conv_std_logic_vector(6257414,24);
            manlo <= conv_std_logic_vector(187437029,28);
            exponent <= conv_std_logic_vector(4,11);
      WHEN "1011000011" =>
            manhi <= conv_std_logic_vector(170718,24);
            manlo <= conv_std_logic_vector(36971864,28);
            exponent <= conv_std_logic_vector(3,11);
      WHEN "1011000100" =>
            manhi <= conv_std_logic_vector(8161970,24);
            manlo <= conv_std_logic_vector(42518955,28);
            exponent <= conv_std_logic_vector(1,11);
      WHEN "1011000101" =>
            manhi <= conv_std_logic_vector(1572011,24);
            manlo <= conv_std_logic_vector(197150320,28);
            exponent <= conv_std_logic_vector(0,11);
      WHEN others =>
           manhi <= conv_std_logic_vector(0,24);
           manlo <= conv_std_logic_vector(0,28);
           exponent <= conv_std_logic_vector(0,11);
    END CASE;
  END PROCESS;

END rtl;
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   DP_EXPLUTPOS.VHD                          ***
--***                                             ***
--***   Function: Look Up Table - EXP()           ***
--***                                             ***
--***   Generated by MATLAB Utility               ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_explutpos IS
PORT (
      add : IN STD_LOGIC_VECTOR (10 DOWNTO 1);
      manhi : OUT STD_LOGIC_VECTOR (24 DOWNTO 1);
      manlo : OUT STD_LOGIC_VECTOR (28 DOWNTO 1);
      exponent : OUT STD_LOGIC_VECTOR (11 DOWNTO 1)
     );
END dp_explutpos;

ARCHITECTURE rtl OF dp_explutpos IS

BEGIN

  pca: PROCESS (add)
  BEGIN
    CASE add IS
      WHEN "0000000000" =>
            manhi <= conv_std_logic_vector(0,24);
            manlo <= conv_std_logic_vector(0,28);
            exponent <= conv_std_logic_vector(1023,11);
      WHEN "0000000001" =>
            manhi <= conv_std_logic_vector(6025384,24);
            manlo <= conv_std_logic_vector(185882474,28);
            exponent <= conv_std_logic_vector(1024,11);
      WHEN "0000000010" =>
            manhi <= conv_std_logic_vector(14214731,24);
            manlo <= conv_std_logic_vector(148168110,28);
            exponent <= conv_std_logic_vector(1025,11);
      WHEN "0000000011" =>
            manhi <= conv_std_logic_vector(4283995,24);
            manlo <= conv_std_logic_vector(258978054,28);
            exponent <= conv_std_logic_vector(1027,11);
      WHEN "0000000100" =>
            manhi <= conv_std_logic_vector(11847938,24);
            manlo <= conv_std_logic_vector(237451864,28);
            exponent <= conv_std_logic_vector(1028,11);
      WHEN "0000000101" =>
            manhi <= conv_std_logic_vector(2675593,24);
            manlo <= conv_std_logic_vector(158348175,28);
            exponent <= conv_std_logic_vector(1030,11);
      WHEN "0000000110" =>
            manhi <= conv_std_logic_vector(9661893,24);
            manlo <= conv_std_logic_vector(110149775,28);
            exponent <= conv_std_logic_vector(1031,11);
      WHEN "0000000111" =>
            manhi <= conv_std_logic_vector(1190021,24);
            manlo <= conv_std_logic_vector(179232170,28);
            exponent <= conv_std_logic_vector(1033,11);
      WHEN "0000001000" =>
            manhi <= conv_std_logic_vector(7642791,24);
            manlo <= conv_std_logic_vector(222760046,28);
            exponent <= conv_std_logic_vector(1034,11);
      WHEN "0000001001" =>
            manhi <= conv_std_logic_vector(16413015,24);
            manlo <= conv_std_logic_vector(205983618,28);
            exponent <= conv_std_logic_vector(1035,11);
      WHEN "0000001010" =>
            manhi <= conv_std_logic_vector(5777884,24);
            manlo <= conv_std_logic_vector(261424480,28);
            exponent <= conv_std_logic_vector(1037,11);
      WHEN "0000001011" =>
            manhi <= conv_std_logic_vector(13878344,24);
            manlo <= conv_std_logic_vector(149835647,28);
            exponent <= conv_std_logic_vector(1038,11);
      WHEN "0000001100" =>
            manhi <= conv_std_logic_vector(4055397,24);
            manlo <= conv_std_logic_vector(80968858,28);
            exponent <= conv_std_logic_vector(1040,11);
      WHEN "0000001101" =>
            manhi <= conv_std_logic_vector(11537241,24);
            manlo <= conv_std_logic_vector(23775573,28);
            exponent <= conv_std_logic_vector(1041,11);
      WHEN "0000001110" =>
            manhi <= conv_std_logic_vector(2464452,24);
            manlo <= conv_std_logic_vector(146736599,28);
            exponent <= conv_std_logic_vector(1043,11);
      WHEN "0000001111" =>
            manhi <= conv_std_logic_vector(9374922,24);
            manlo <= conv_std_logic_vector(263006855,28);
            exponent <= conv_std_logic_vector(1044,11);
      WHEN "0000010000" =>
            manhi <= conv_std_logic_vector(995005,24);
            manlo <= conv_std_logic_vector(11010080,28);
            exponent <= conv_std_logic_vector(1046,11);
      WHEN "0000010001" =>
            manhi <= conv_std_logic_vector(7377736,24);
            manlo <= conv_std_logic_vector(202286329,28);
            exponent <= conv_std_logic_vector(1047,11);
      WHEN "0000010010" =>
            manhi <= conv_std_logic_vector(16052768,24);
            manlo <= conv_std_logic_vector(152649917,28);
            exponent <= conv_std_logic_vector(1048,11);
      WHEN "0000010011" =>
            manhi <= conv_std_logic_vector(5533071,24);
            manlo <= conv_std_logic_vector(166536930,28);
            exponent <= conv_std_logic_vector(1050,11);
      WHEN "0000010100" =>
            manhi <= conv_std_logic_vector(13545608,24);
            manlo <= conv_std_logic_vector(191424516,28);
            exponent <= conv_std_logic_vector(1051,11);
      WHEN "0000010101" =>
            manhi <= conv_std_logic_vector(3829279,24);
            manlo <= conv_std_logic_vector(228519165,28);
            exponent <= conv_std_logic_vector(1053,11);
      WHEN "0000010110" =>
            manhi <= conv_std_logic_vector(11229915,24);
            manlo <= conv_std_logic_vector(163853824,28);
            exponent <= conv_std_logic_vector(1054,11);
      WHEN "0000010111" =>
            manhi <= conv_std_logic_vector(2255603,24);
            manlo <= conv_std_logic_vector(61996481,28);
            exponent <= conv_std_logic_vector(1056,11);
      WHEN "0000011000" =>
            manhi <= conv_std_logic_vector(9091067,24);
            manlo <= conv_std_logic_vector(88563639,28);
            exponent <= conv_std_logic_vector(1057,11);
      WHEN "0000011001" =>
            manhi <= conv_std_logic_vector(802105,24);
            manlo <= conv_std_logic_vector(34169545,28);
            exponent <= conv_std_logic_vector(1059,11);
      WHEN "0000011010" =>
            manhi <= conv_std_logic_vector(7115558,24);
            manlo <= conv_std_logic_vector(157969244,28);
            exponent <= conv_std_logic_vector(1060,11);
      WHEN "0000011011" =>
            manhi <= conv_std_logic_vector(15696431,24);
            manlo <= conv_std_logic_vector(133591837,28);
            exponent <= conv_std_logic_vector(1061,11);
      WHEN "0000011100" =>
            manhi <= conv_std_logic_vector(5290915,24);
            manlo <= conv_std_logic_vector(127285146,28);
            exponent <= conv_std_logic_vector(1063,11);
      WHEN "0000011101" =>
            manhi <= conv_std_logic_vector(13216484,24);
            manlo <= conv_std_logic_vector(103923798,28);
            exponent <= conv_std_logic_vector(1064,11);
      WHEN "0000011110" =>
            manhi <= conv_std_logic_vector(3605616,24);
            manlo <= conv_std_logic_vector(183249133,28);
            exponent <= conv_std_logic_vector(1066,11);
      WHEN "0000011111" =>
            manhi <= conv_std_logic_vector(10925925,24);
            manlo <= conv_std_logic_vector(227336045,28);
            exponent <= conv_std_logic_vector(1067,11);
      WHEN "0000100000" =>
            manhi <= conv_std_logic_vector(2049020,24);
            manlo <= conv_std_logic_vector(206267948,28);
            exponent <= conv_std_logic_vector(1069,11);
      WHEN "0000100001" =>
            manhi <= conv_std_logic_vector(8810292,24);
            manlo <= conv_std_logic_vector(175265666,28);
            exponent <= conv_std_logic_vector(1070,11);
      WHEN "0000100010" =>
            manhi <= conv_std_logic_vector(611298,24);
            manlo <= conv_std_logic_vector(255467255,28);
            exponent <= conv_std_logic_vector(1072,11);
      WHEN "0000100011" =>
            manhi <= conv_std_logic_vector(6856226,24);
            manlo <= conv_std_logic_vector(29134171,28);
            exponent <= conv_std_logic_vector(1073,11);
      WHEN "0000100100" =>
            manhi <= conv_std_logic_vector(15343962,24);
            manlo <= conv_std_logic_vector(30543222,28);
            exponent <= conv_std_logic_vector(1074,11);
      WHEN "0000100101" =>
            manhi <= conv_std_logic_vector(5051387,24);
            manlo <= conv_std_logic_vector(186253338,28);
            exponent <= conv_std_logic_vector(1076,11);
      WHEN "0000100110" =>
            manhi <= conv_std_logic_vector(12890932,24);
            manlo <= conv_std_logic_vector(102222951,28);
            exponent <= conv_std_logic_vector(1077,11);
      WHEN "0000100111" =>
            manhi <= conv_std_logic_vector(3384381,24);
            manlo <= conv_std_logic_vector(42116377,28);
            exponent <= conv_std_logic_vector(1079,11);
      WHEN "0000101000" =>
            manhi <= conv_std_logic_vector(10625235,24);
            manlo <= conv_std_logic_vector(158954218,28);
            exponent <= conv_std_logic_vector(1080,11);
      WHEN "0000101001" =>
            manhi <= conv_std_logic_vector(1844680,24);
            manlo <= conv_std_logic_vector(148858978,28);
            exponent <= conv_std_logic_vector(1082,11);
      WHEN "0000101010" =>
            manhi <= conv_std_logic_vector(8532565,24);
            manlo <= conv_std_logic_vector(136319321,28);
            exponent <= conv_std_logic_vector(1083,11);
      WHEN "0000101011" =>
            manhi <= conv_std_logic_vector(422563,24);
            manlo <= conv_std_logic_vector(211728497,28);
            exponent <= conv_std_logic_vector(1085,11);
      WHEN "0000101100" =>
            manhi <= conv_std_logic_vector(6599708,24);
            manlo <= conv_std_logic_vector(114522162,28);
            exponent <= conv_std_logic_vector(1086,11);
      WHEN "0000101101" =>
            manhi <= conv_std_logic_vector(14995318,24);
            manlo <= conv_std_logic_vector(117328318,28);
            exponent <= conv_std_logic_vector(1087,11);
      WHEN "0000101110" =>
            manhi <= conv_std_logic_vector(4814459,24);
            manlo <= conv_std_logic_vector(201622499,28);
            exponent <= conv_std_logic_vector(1089,11);
      WHEN "0000101111" =>
            manhi <= conv_std_logic_vector(12568913,24);
            manlo <= conv_std_logic_vector(246987638,28);
            exponent <= conv_std_logic_vector(1090,11);
      WHEN "0000110000" =>
            manhi <= conv_std_logic_vector(3165546,24);
            manlo <= conv_std_logic_vector(248128843,28);
            exponent <= conv_std_logic_vector(1092,11);
      WHEN "0000110001" =>
            manhi <= conv_std_logic_vector(10327809,24);
            manlo <= conv_std_logic_vector(8929872,28);
            exponent <= conv_std_logic_vector(1093,11);
      WHEN "0000110010" =>
            manhi <= conv_std_logic_vector(1642558,24);
            manlo <= conv_std_logic_vector(67636037,28);
            exponent <= conv_std_logic_vector(1095,11);
      WHEN "0000110011" =>
            manhi <= conv_std_logic_vector(8257852,24);
            manlo <= conv_std_logic_vector(219235425,28);
            exponent <= conv_std_logic_vector(1096,11);
      WHEN "0000110100" =>
            manhi <= conv_std_logic_vector(235877,24);
            manlo <= conv_std_logic_vector(42862412,28);
            exponent <= conv_std_logic_vector(1098,11);
      WHEN "0000110101" =>
            manhi <= conv_std_logic_vector(6345974,24);
            manlo <= conv_std_logic_vector(265996080,28);
            exponent <= conv_std_logic_vector(1099,11);
      WHEN "0000110110" =>
            manhi <= conv_std_logic_vector(14650458,24);
            manlo <= conv_std_logic_vector(253213243,28);
            exponent <= conv_std_logic_vector(1100,11);
      WHEN "0000110111" =>
            manhi <= conv_std_logic_vector(4580103,24);
            manlo <= conv_std_logic_vector(114693785,28);
            exponent <= conv_std_logic_vector(1102,11);
      WHEN "0000111000" =>
            manhi <= conv_std_logic_vector(12250390,24);
            manlo <= conv_std_logic_vector(174984615,28);
            exponent <= conv_std_logic_vector(1103,11);
      WHEN "0000111001" =>
            manhi <= conv_std_logic_vector(2949087,24);
            manlo <= conv_std_logic_vector(247325089,28);
            exponent <= conv_std_logic_vector(1105,11);
      WHEN "0000111010" =>
            manhi <= conv_std_logic_vector(10033610,24);
            manlo <= conv_std_logic_vector(200264553,28);
            exponent <= conv_std_logic_vector(1106,11);
      WHEN "0000111011" =>
            manhi <= conv_std_logic_vector(1442629,24);
            manlo <= conv_std_logic_vector(211375075,28);
            exponent <= conv_std_logic_vector(1108,11);
      WHEN "0000111100" =>
            manhi <= conv_std_logic_vector(7986121,24);
            manlo <= conv_std_logic_vector(231029862,28);
            exponent <= conv_std_logic_vector(1109,11);
      WHEN "0000111101" =>
            manhi <= conv_std_logic_vector(51216,24);
            manlo <= conv_std_logic_vector(222707863,28);
            exponent <= conv_std_logic_vector(1111,11);
      WHEN "0000111110" =>
            manhi <= conv_std_logic_vector(6094995,24);
            manlo <= conv_std_logic_vector(155999272,28);
            exponent <= conv_std_logic_vector(1112,11);
      WHEN "0000111111" =>
            manhi <= conv_std_logic_vector(14309342,24);
            manlo <= conv_std_logic_vector(150013864,28);
            exponent <= conv_std_logic_vector(1113,11);
      WHEN "0001000000" =>
            manhi <= conv_std_logic_vector(4348290,24);
            manlo <= conv_std_logic_vector(217421773,28);
            exponent <= conv_std_logic_vector(1115,11);
      WHEN "0001000001" =>
            manhi <= conv_std_logic_vector(11935324,24);
            manlo <= conv_std_logic_vector(171597361,28);
            exponent <= conv_std_logic_vector(1116,11);
      WHEN "0001000010" =>
            manhi <= conv_std_logic_vector(2734978,24);
            manlo <= conv_std_logic_vector(98553735,28);
            exponent <= conv_std_logic_vector(1118,11);
      WHEN "0001000011" =>
            manhi <= conv_std_logic_vector(9742605,24);
            manlo <= conv_std_logic_vector(185429986,28);
            exponent <= conv_std_logic_vector(1119,11);
      WHEN "0001000100" =>
            manhi <= conv_std_logic_vector(1244871,24);
            manlo <= conv_std_logic_vector(93685501,28);
            exponent <= conv_std_logic_vector(1121,11);
      WHEN "0001000101" =>
            manhi <= conv_std_logic_vector(7717340,24);
            manlo <= conv_std_logic_vector(74048432,28);
            exponent <= conv_std_logic_vector(1122,11);
      WHEN "0001000110" =>
            manhi <= conv_std_logic_vector(16514337,24);
            manlo <= conv_std_logic_vector(163855108,28);
            exponent <= conv_std_logic_vector(1123,11);
      WHEN "0001000111" =>
            manhi <= conv_std_logic_vector(5846740,24);
            manlo <= conv_std_logic_vector(81895750,28);
            exponent <= conv_std_logic_vector(1125,11);
      WHEN "0001001000" =>
            manhi <= conv_std_logic_vector(13971928,24);
            manlo <= conv_std_logic_vector(176088988,28);
            exponent <= conv_std_logic_vector(1126,11);
      WHEN "0001001001" =>
            manhi <= conv_std_logic_vector(4118994,24);
            manlo <= conv_std_logic_vector(77780251,28);
            exponent <= conv_std_logic_vector(1128,11);
      WHEN "0001001010" =>
            manhi <= conv_std_logic_vector(11623678,24);
            manlo <= conv_std_logic_vector(95871356,28);
            exponent <= conv_std_logic_vector(1129,11);
      WHEN "0001001011" =>
            manhi <= conv_std_logic_vector(2523192,24);
            manlo <= conv_std_logic_vector(204213760,28);
            exponent <= conv_std_logic_vector(1131,11);
      WHEN "0001001100" =>
            manhi <= conv_std_logic_vector(9454759,24);
            manlo <= conv_std_logic_vector(55860552,28);
            exponent <= conv_std_logic_vector(1132,11);
      WHEN "0001001101" =>
            manhi <= conv_std_logic_vector(1049259,24);
            manlo <= conv_std_logic_vector(102861624,28);
            exponent <= conv_std_logic_vector(1134,11);
      WHEN "0001001110" =>
            manhi <= conv_std_logic_vector(7451476,24);
            manlo <= conv_std_logic_vector(13367584,28);
            exponent <= conv_std_logic_vector(1135,11);
      WHEN "0001001111" =>
            manhi <= conv_std_logic_vector(16152990,24);
            manlo <= conv_std_logic_vector(178012490,28);
            exponent <= conv_std_logic_vector(1136,11);
      WHEN "0001010000" =>
            manhi <= conv_std_logic_vector(5601179,24);
            manlo <= conv_std_logic_vector(159708139,28);
            exponent <= conv_std_logic_vector(1138,11);
      WHEN "0001010001" =>
            manhi <= conv_std_logic_vector(13638177,24);
            manlo <= conv_std_logic_vector(12864164,28);
            exponent <= conv_std_logic_vector(1139,11);
      WHEN "0001010010" =>
            manhi <= conv_std_logic_vector(3892186,24);
            manlo <= conv_std_logic_vector(149492240,28);
            exponent <= conv_std_logic_vector(1141,11);
      WHEN "0001010011" =>
            manhi <= conv_std_logic_vector(11315414,24);
            manlo <= conv_std_logic_vector(184620728,28);
            exponent <= conv_std_logic_vector(1142,11);
      WHEN "0001010100" =>
            manhi <= conv_std_logic_vector(2313705,24);
            manlo <= conv_std_logic_vector(235697385,28);
            exponent <= conv_std_logic_vector(1144,11);
      WHEN "0001010101" =>
            manhi <= conv_std_logic_vector(9170037,24);
            manlo <= conv_std_logic_vector(3974263,28);
            exponent <= conv_std_logic_vector(1145,11);
      WHEN "0001010110" =>
            manhi <= conv_std_logic_vector(855770,24);
            manlo <= conv_std_logic_vector(158952336,28);
            exponent <= conv_std_logic_vector(1147,11);
      WHEN "0001010111" =>
            manhi <= conv_std_logic_vector(7188497,24);
            manlo <= conv_std_logic_vector(138900038,28);
            exponent <= conv_std_logic_vector(1148,11);
      WHEN "0001011000" =>
            manhi <= conv_std_logic_vector(15795565,24);
            manlo <= conv_std_logic_vector(209449517,28);
            exponent <= conv_std_logic_vector(1149,11);
      WHEN "0001011001" =>
            manhi <= conv_std_logic_vector(5358284,24);
            manlo <= conv_std_logic_vector(54736896,28);
            exponent <= conv_std_logic_vector(1151,11);
      WHEN "0001011010" =>
            manhi <= conv_std_logic_vector(13308047,24);
            manlo <= conv_std_logic_vector(264159588,28);
            exponent <= conv_std_logic_vector(1152,11);
      WHEN "0001011011" =>
            manhi <= conv_std_logic_vector(3667840,24);
            manlo <= conv_std_logic_vector(160544132,28);
            exponent <= conv_std_logic_vector(1154,11);
      WHEN "0001011100" =>
            manhi <= conv_std_logic_vector(11010496,24);
            manlo <= conv_std_logic_vector(245935181,28);
            exponent <= conv_std_logic_vector(1155,11);
      WHEN "0001011101" =>
            manhi <= conv_std_logic_vector(2106492,24);
            manlo <= conv_std_logic_vector(206325441,28);
            exponent <= conv_std_logic_vector(1157,11);
      WHEN "0001011110" =>
            manhi <= conv_std_logic_vector(8888405,24);
            manlo <= conv_std_logic_vector(53641237,28);
            exponent <= conv_std_logic_vector(1158,11);
      WHEN "0001011111" =>
            manhi <= conv_std_logic_vector(664381,24);
            manlo <= conv_std_logic_vector(249887163,28);
            exponent <= conv_std_logic_vector(1160,11);
      WHEN "0001100000" =>
            manhi <= conv_std_logic_vector(6928373,24);
            manlo <= conv_std_logic_vector(95946938,28);
            exponent <= conv_std_logic_vector(1161,11);
      WHEN "0001100001" =>
            manhi <= conv_std_logic_vector(15442020,24);
            manlo <= conv_std_logic_vector(105121290,28);
            exponent <= conv_std_logic_vector(1162,11);
      WHEN "0001100010" =>
            manhi <= conv_std_logic_vector(5118025,24);
            manlo <= conv_std_logic_vector(54367076,28);
            exponent <= conv_std_logic_vector(1164,11);
      WHEN "0001100011" =>
            manhi <= conv_std_logic_vector(12981502,24);
            manlo <= conv_std_logic_vector(39000129,28);
            exponent <= conv_std_logic_vector(1165,11);
      WHEN "0001100100" =>
            manhi <= conv_std_logic_vector(3445929,24);
            manlo <= conv_std_logic_vector(186063861,28);
            exponent <= conv_std_logic_vector(1167,11);
      WHEN "0001100101" =>
            manhi <= conv_std_logic_vector(10708888,24);
            manlo <= conv_std_logic_vector(194877084,28);
            exponent <= conv_std_logic_vector(1168,11);
      WHEN "0001100110" =>
            manhi <= conv_std_logic_vector(1901528,24);
            manlo <= conv_std_logic_vector(202114223,28);
            exponent <= conv_std_logic_vector(1170,11);
      WHEN "0001100111" =>
            manhi <= conv_std_logic_vector(8609830,24);
            manlo <= conv_std_logic_vector(59099508,28);
            exponent <= conv_std_logic_vector(1171,11);
      WHEN "0001101000" =>
            manhi <= conv_std_logic_vector(475070,24);
            manlo <= conv_std_logic_vector(162304029,28);
            exponent <= conv_std_logic_vector(1173,11);
      WHEN "0001101001" =>
            manhi <= conv_std_logic_vector(6671072,24);
            manlo <= conv_std_logic_vector(157938310,28);
            exponent <= conv_std_logic_vector(1174,11);
      WHEN "0001101010" =>
            manhi <= conv_std_logic_vector(15092312,24);
            manlo <= conv_std_logic_vector(104450792,28);
            exponent <= conv_std_logic_vector(1175,11);
      WHEN "0001101011" =>
            manhi <= conv_std_logic_vector(4880373,24);
            manlo <= conv_std_logic_vector(261837049,28);
            exponent <= conv_std_logic_vector(1177,11);
      WHEN "0001101100" =>
            manhi <= conv_std_logic_vector(12658500,24);
            manlo <= conv_std_logic_vector(171583716,28);
            exponent <= conv_std_logic_vector(1178,11);
      WHEN "0001101101" =>
            manhi <= conv_std_logic_vector(3226427,24);
            manlo <= conv_std_logic_vector(110595717,28);
            exponent <= conv_std_logic_vector(1180,11);
      WHEN "0001101110" =>
            manhi <= conv_std_logic_vector(10410554,24);
            manlo <= conv_std_logic_vector(52320382,28);
            exponent <= conv_std_logic_vector(1181,11);
      WHEN "0001101111" =>
            manhi <= conv_std_logic_vector(1698789,24);
            manlo <= conv_std_logic_vector(112550995,28);
            exponent <= conv_std_logic_vector(1183,11);
      WHEN "0001110000" =>
            manhi <= conv_std_logic_vector(8334278,24);
            manlo <= conv_std_logic_vector(240753534,28);
            exponent <= conv_std_logic_vector(1184,11);
      WHEN "0001110001" =>
            manhi <= conv_std_logic_vector(287814,24);
            manlo <= conv_std_logic_vector(17691391,28);
            exponent <= conv_std_logic_vector(1186,11);
      WHEN "0001110010" =>
            manhi <= conv_std_logic_vector(6416564,24);
            manlo <= conv_std_logic_vector(151700710,28);
            exponent <= conv_std_logic_vector(1187,11);
      WHEN "0001110011" =>
            manhi <= conv_std_logic_vector(14746400,24);
            manlo <= conv_std_logic_vector(32676275,28);
            exponent <= conv_std_logic_vector(1188,11);
      WHEN "0001110100" =>
            manhi <= conv_std_logic_vector(4645302,24);
            manlo <= conv_std_logic_vector(58452725,28);
            exponent <= conv_std_logic_vector(1190,11);
      WHEN "0001110101" =>
            manhi <= conv_std_logic_vector(12339004,24);
            manlo <= conv_std_logic_vector(267247876,28);
            exponent <= conv_std_logic_vector(1191,11);
      WHEN "0001110110" =>
            manhi <= conv_std_logic_vector(3009307,24);
            manlo <= conv_std_logic_vector(164126253,28);
            exponent <= conv_std_logic_vector(1193,11);
      WHEN "0001110111" =>
            manhi <= conv_std_logic_vector(10115457,24);
            manlo <= conv_std_logic_vector(212237584,28);
            exponent <= conv_std_logic_vector(1194,11);
      WHEN "0001111000" =>
            manhi <= conv_std_logic_vector(1498250,24);
            manlo <= conv_std_logic_vector(166684427,28);
            exponent <= conv_std_logic_vector(1196,11);
      WHEN "0001111001" =>
            manhi <= conv_std_logic_vector(8061718,24);
            manlo <= conv_std_logic_vector(110371593,28);
            exponent <= conv_std_logic_vector(1197,11);
      WHEN "0001111010" =>
            manhi <= conv_std_logic_vector(102590,24);
            manlo <= conv_std_logic_vector(3231911,28);
            exponent <= conv_std_logic_vector(1199,11);
      WHEN "0001111011" =>
            manhi <= conv_std_logic_vector(6164818,24);
            manlo <= conv_std_logic_vector(261783833,28);
            exponent <= conv_std_logic_vector(1200,11);
      WHEN "0001111100" =>
            manhi <= conv_std_logic_vector(14404242,24);
            manlo <= conv_std_logic_vector(104825991,28);
            exponent <= conv_std_logic_vector(1201,11);
      WHEN "0001111101" =>
            manhi <= conv_std_logic_vector(4412781,24);
            manlo <= conv_std_logic_vector(250166254,28);
            exponent <= conv_std_logic_vector(1203,11);
      WHEN "0001111110" =>
            manhi <= conv_std_logic_vector(12022977,24);
            manlo <= conv_std_logic_vector(43417082,28);
            exponent <= conv_std_logic_vector(1204,11);
      WHEN "0001111111" =>
            manhi <= conv_std_logic_vector(2794544,24);
            manlo <= conv_std_logic_vector(115942082,28);
            exponent <= conv_std_logic_vector(1206,11);
      WHEN "0010000000" =>
            manhi <= conv_std_logic_vector(9823564,24);
            manlo <= conv_std_logic_vector(98386456,28);
            exponent <= conv_std_logic_vector(1207,11);
      WHEN "0010000001" =>
            manhi <= conv_std_logic_vector(1299888,24);
            manlo <= conv_std_logic_vector(127046227,28);
            exponent <= conv_std_logic_vector(1209,11);
      WHEN "0010000010" =>
            manhi <= conv_std_logic_vector(7792116,24);
            manlo <= conv_std_logic_vector(80649262,28);
            exponent <= conv_std_logic_vector(1210,11);
      WHEN "0010000011" =>
            manhi <= conv_std_logic_vector(16615968,24);
            manlo <= conv_std_logic_vector(205307910,28);
            exponent <= conv_std_logic_vector(1211,11);
      WHEN "0010000100" =>
            manhi <= conv_std_logic_vector(5915805,24);
            manlo <= conv_std_logic_vector(224185017,28);
            exponent <= conv_std_logic_vector(1213,11);
      WHEN "0010000101" =>
            manhi <= conv_std_logic_vector(14065798,24);
            manlo <= conv_std_logic_vector(119094636,28);
            exponent <= conv_std_logic_vector(1214,11);
      WHEN "0010000110" =>
            manhi <= conv_std_logic_vector(4182785,24);
            manlo <= conv_std_logic_vector(113890892,28);
            exponent <= conv_std_logic_vector(1216,11);
      WHEN "0010000111" =>
            manhi <= conv_std_logic_vector(11710379,24);
            manlo <= conv_std_logic_vector(133692518,28);
            exponent <= conv_std_logic_vector(1217,11);
      WHEN "0010001000" =>
            manhi <= conv_std_logic_vector(2582112,24);
            manlo <= conv_std_logic_vector(79109485,28);
            exponent <= conv_std_logic_vector(1219,11);
      WHEN "0010001001" =>
            manhi <= conv_std_logic_vector(9534839,24);
            manlo <= conv_std_logic_vector(42234535,28);
            exponent <= conv_std_logic_vector(1220,11);
      WHEN "0010001010" =>
            manhi <= conv_std_logic_vector(1103679,24);
            manlo <= conv_std_logic_vector(94193887,28);
            exponent <= conv_std_logic_vector(1222,11);
      WHEN "0010001011" =>
            manhi <= conv_std_logic_vector(7525440,24);
            manlo <= conv_std_logic_vector(121994268,28);
            exponent <= conv_std_logic_vector(1223,11);
      WHEN "0010001100" =>
            manhi <= conv_std_logic_vector(16253518,24);
            manlo <= conv_std_logic_vector(191052573,28);
            exponent <= conv_std_logic_vector(1224,11);
      WHEN "0010001101" =>
            manhi <= conv_std_logic_vector(5669495,24);
            manlo <= conv_std_logic_vector(130696997,28);
            exponent <= conv_std_logic_vector(1226,11);
      WHEN "0010001110" =>
            manhi <= conv_std_logic_vector(13731027,24);
            manlo <= conv_std_logic_vector(260846837,28);
            exponent <= conv_std_logic_vector(1227,11);
      WHEN "0010001111" =>
            manhi <= conv_std_logic_vector(3955285,24);
            manlo <= conv_std_logic_vector(80970159,28);
            exponent <= conv_std_logic_vector(1229,11);
      WHEN "0010010000" =>
            manhi <= conv_std_logic_vector(11401174,24);
            manlo <= conv_std_logic_vector(207600506,28);
            exponent <= conv_std_logic_vector(1230,11);
      WHEN "0010010001" =>
            manhi <= conv_std_logic_vector(2371985,24);
            manlo <= conv_std_logic_vector(241221170,28);
            exponent <= conv_std_logic_vector(1232,11);
      WHEN "0010010010" =>
            manhi <= conv_std_logic_vector(9249247,24);
            manlo <= conv_std_logic_vector(208105818,28);
            exponent <= conv_std_logic_vector(1233,11);
      WHEN "0010010011" =>
            manhi <= conv_std_logic_vector(909599,24);
            manlo <= conv_std_logic_vector(237519888,28);
            exponent <= conv_std_logic_vector(1235,11);
      WHEN "0010010100" =>
            manhi <= conv_std_logic_vector(7261659,24);
            manlo <= conv_std_logic_vector(29935335,28);
            exponent <= conv_std_logic_vector(1236,11);
      WHEN "0010010101" =>
            manhi <= conv_std_logic_vector(15895002,24);
            manlo <= conv_std_logic_vector(186862656,28);
            exponent <= conv_std_logic_vector(1237,11);
      WHEN "0010010110" =>
            manhi <= conv_std_logic_vector(5425858,24);
            manlo <= conv_std_logic_vector(159524243,28);
            exponent <= conv_std_logic_vector(1239,11);
      WHEN "0010010111" =>
            manhi <= conv_std_logic_vector(13399891,24);
            manlo <= conv_std_logic_vector(27586577,28);
            exponent <= conv_std_logic_vector(1240,11);
      WHEN "0010011000" =>
            manhi <= conv_std_logic_vector(3730254,24);
            manlo <= conv_std_logic_vector(125689310,28);
            exponent <= conv_std_logic_vector(1242,11);
      WHEN "0010011001" =>
            manhi <= conv_std_logic_vector(11095326,24);
            manlo <= conv_std_logic_vector(43144000,28);
            exponent <= conv_std_logic_vector(1243,11);
      WHEN "0010011010" =>
            manhi <= conv_std_logic_vector(2164140,24);
            manlo <= conv_std_logic_vector(58280992,28);
            exponent <= conv_std_logic_vector(1245,11);
      WHEN "0010011011" =>
            manhi <= conv_std_logic_vector(8966756,24);
            manlo <= conv_std_logic_vector(55210422,28);
            exponent <= conv_std_logic_vector(1246,11);
      WHEN "0010011100" =>
            manhi <= conv_std_logic_vector(717626,24);
            manlo <= conv_std_logic_vector(257633658,28);
            exponent <= conv_std_logic_vector(1248,11);
      WHEN "0010011101" =>
            manhi <= conv_std_logic_vector(7000740,24);
            manlo <= conv_std_logic_vector(229413090,28);
            exponent <= conv_std_logic_vector(1249,11);
      WHEN "0010011110" =>
            manhi <= conv_std_logic_vector(15540378,24);
            manlo <= conv_std_logic_vector(4808337,28);
            exponent <= conv_std_logic_vector(1250,11);
      WHEN "0010011111" =>
            manhi <= conv_std_logic_vector(5184866,24);
            manlo <= conv_std_logic_vector(37474138,28);
            exponent <= conv_std_logic_vector(1252,11);
      WHEN "0010100000" =>
            manhi <= conv_std_logic_vector(13072348,24);
            manlo <= conv_std_logic_vector(106730632,28);
            exponent <= conv_std_logic_vector(1253,11);
      WHEN "0010100001" =>
            manhi <= conv_std_logic_vector(3507666,24);
            manlo <= conv_std_logic_vector(32844500,28);
            exponent <= conv_std_logic_vector(1255,11);
      WHEN "0010100010" =>
            manhi <= conv_std_logic_vector(10792797,24);
            manlo <= conv_std_logic_vector(62496090,28);
            exponent <= conv_std_logic_vector(1256,11);
      WHEN "0010100011" =>
            manhi <= conv_std_logic_vector(1958550,24);
            manlo <= conv_std_logic_vector(132952012,28);
            exponent <= conv_std_logic_vector(1258,11);
      WHEN "0010100100" =>
            manhi <= conv_std_logic_vector(8687330,24);
            manlo <= conv_std_logic_vector(215605290,28);
            exponent <= conv_std_logic_vector(1259,11);
      WHEN "0010100101" =>
            manhi <= conv_std_logic_vector(527737,24);
            manlo <= conv_std_logic_vector(190928911,28);
            exponent <= conv_std_logic_vector(1261,11);
      WHEN "0010100110" =>
            manhi <= conv_std_logic_vector(6742654,24);
            manlo <= conv_std_logic_vector(163162889,28);
            exponent <= conv_std_logic_vector(1262,11);
      WHEN "0010100111" =>
            manhi <= conv_std_logic_vector(15189602,24);
            manlo <= conv_std_logic_vector(118241780,28);
            exponent <= conv_std_logic_vector(1263,11);
      WHEN "0010101000" =>
            manhi <= conv_std_logic_vector(4946489,24);
            manlo <= conv_std_logic_vector(112771062,28);
            exponent <= conv_std_logic_vector(1265,11);
      WHEN "0010101001" =>
            manhi <= conv_std_logic_vector(12748360,24);
            manlo <= conv_std_logic_vector(226864003,28);
            exponent <= conv_std_logic_vector(1266,11);
      WHEN "0010101010" =>
            manhi <= conv_std_logic_vector(3287493,24);
            manlo <= conv_std_logic_vector(202192272,28);
            exponent <= conv_std_logic_vector(1268,11);
      WHEN "0010101011" =>
            manhi <= conv_std_logic_vector(10493551,24);
            manlo <= conv_std_logic_vector(257093553,28);
            exponent <= conv_std_logic_vector(1269,11);
      WHEN "0010101100" =>
            manhi <= conv_std_logic_vector(1755192,24);
            manlo <= conv_std_logic_vector(66281405,28);
            exponent <= conv_std_logic_vector(1271,11);
      WHEN "0010101101" =>
            manhi <= conv_std_logic_vector(8410938,24);
            manlo <= conv_std_logic_vector(77199396,28);
            exponent <= conv_std_logic_vector(1272,11);
      WHEN "0010101110" =>
            manhi <= conv_std_logic_vector(339909,24);
            manlo <= conv_std_logic_vector(140417186,28);
            exponent <= conv_std_logic_vector(1274,11);
      WHEN "0010101111" =>
            manhi <= conv_std_logic_vector(6487369,24);
            manlo <= conv_std_logic_vector(169769464,28);
            exponent <= conv_std_logic_vector(1275,11);
      WHEN "0010110000" =>
            manhi <= conv_std_logic_vector(14842634,24);
            manlo <= conv_std_logic_vector(49834035,28);
            exponent <= conv_std_logic_vector(1276,11);
      WHEN "0010110001" =>
            manhi <= conv_std_logic_vector(4710700,24);
            manlo <= conv_std_logic_vector(11961455,28);
            exponent <= conv_std_logic_vector(1278,11);
      WHEN "0010110010" =>
            manhi <= conv_std_logic_vector(12427889,24);
            manlo <= conv_std_logic_vector(230234502,28);
            exponent <= conv_std_logic_vector(1279,11);
      WHEN "0010110011" =>
            manhi <= conv_std_logic_vector(3069711,24);
            manlo <= conv_std_logic_vector(36989233,28);
            exponent <= conv_std_logic_vector(1281,11);
      WHEN "0010110100" =>
            manhi <= conv_std_logic_vector(10197554,24);
            manlo <= conv_std_logic_vector(186484869,28);
            exponent <= conv_std_logic_vector(1282,11);
      WHEN "0010110101" =>
            manhi <= conv_std_logic_vector(1554041,24);
            manlo <= conv_std_logic_vector(67530342,28);
            exponent <= conv_std_logic_vector(1284,11);
      WHEN "0010110110" =>
            manhi <= conv_std_logic_vector(8137545,24);
            manlo <= conv_std_logic_vector(198608842,28);
            exponent <= conv_std_logic_vector(1285,11);
      WHEN "0010110111" =>
            manhi <= conv_std_logic_vector(154120,24);
            manlo <= conv_std_logic_vector(6569319,28);
            exponent <= conv_std_logic_vector(1287,11);
      WHEN "0010111000" =>
            manhi <= conv_std_logic_vector(6234855,24);
            manlo <= conv_std_logic_vector(140506894,28);
            exponent <= conv_std_logic_vector(1288,11);
      WHEN "0010111001" =>
            manhi <= conv_std_logic_vector(14499431,24);
            manlo <= conv_std_logic_vector(249287529,28);
            exponent <= conv_std_logic_vector(1289,11);
      WHEN "0010111010" =>
            manhi <= conv_std_logic_vector(4477469,24);
            manlo <= conv_std_logic_vector(249618841,28);
            exponent <= conv_std_logic_vector(1291,11);
      WHEN "0010111011" =>
            manhi <= conv_std_logic_vector(12110897,24);
            manlo <= conv_std_logic_vector(71519058,28);
            exponent <= conv_std_logic_vector(1292,11);
      WHEN "0010111100" =>
            manhi <= conv_std_logic_vector(2854292,24);
            manlo <= conv_std_logic_vector(90637320,28);
            exponent <= conv_std_logic_vector(1294,11);
      WHEN "0010111101" =>
            manhi <= conv_std_logic_vector(9904770,24);
            manlo <= conv_std_logic_vector(50932558,28);
            exponent <= conv_std_logic_vector(1295,11);
      WHEN "0010111110" =>
            manhi <= conv_std_logic_vector(1355073,24);
            manlo <= conv_std_logic_vector(148093260,28);
            exponent <= conv_std_logic_vector(1297,11);
      WHEN "0010111111" =>
            manhi <= conv_std_logic_vector(7867120,24);
            manlo <= conv_std_logic_vector(160620741,28);
            exponent <= conv_std_logic_vector(1298,11);
      WHEN "0011000000" =>
            manhi <= conv_std_logic_vector(16717910,24);
            manlo <= conv_std_logic_vector(46942270,28);
            exponent <= conv_std_logic_vector(1299,11);
      WHEN "0011000001" =>
            manhi <= conv_std_logic_vector(5985082,24);
            manlo <= conv_std_logic_vector(55237426,28);
            exponent <= conv_std_logic_vector(1301,11);
      WHEN "0011000010" =>
            manhi <= conv_std_logic_vector(14159954,24);
            manlo <= conv_std_logic_vector(212966668,28);
            exponent <= conv_std_logic_vector(1302,11);
      WHEN "0011000011" =>
            manhi <= conv_std_logic_vector(4246771,24);
            manlo <= conv_std_logic_vector(79962334,28);
            exponent <= conv_std_logic_vector(1304,11);
      WHEN "0011000100" =>
            manhi <= conv_std_logic_vector(11797345,24);
            manlo <= conv_std_logic_vector(85038862,28);
            exponent <= conv_std_logic_vector(1305,11);
      WHEN "0011000101" =>
            manhi <= conv_std_logic_vector(2641211,24);
            manlo <= conv_std_logic_vector(186806322,28);
            exponent <= conv_std_logic_vector(1307,11);
      WHEN "0011000110" =>
            manhi <= conv_std_logic_vector(9615163,24);
            manlo <= conv_std_logic_vector(153415152,28);
            exponent <= conv_std_logic_vector(1308,11);
      WHEN "0011000111" =>
            manhi <= conv_std_logic_vector(1158265,24);
            manlo <= conv_std_logic_vector(120731907,28);
            exponent <= conv_std_logic_vector(1310,11);
      WHEN "0011001000" =>
            manhi <= conv_std_logic_vector(7599630,24);
            manlo <= conv_std_logic_vector(175764921,28);
            exponent <= conv_std_logic_vector(1311,11);
      WHEN "0011001001" =>
            manhi <= conv_std_logic_vector(16354353,24);
            manlo <= conv_std_logic_vector(174054693,28);
            exponent <= conv_std_logic_vector(1312,11);
      WHEN "0011001010" =>
            manhi <= conv_std_logic_vector(5738019,24);
            manlo <= conv_std_logic_vector(249885394,28);
            exponent <= conv_std_logic_vector(1314,11);
      WHEN "0011001011" =>
            manhi <= conv_std_logic_vector(13824162,24);
            manlo <= conv_std_logic_vector(93203713,28);
            exponent <= conv_std_logic_vector(1315,11);
      WHEN "0011001100" =>
            manhi <= conv_std_logic_vector(4018576,24);
            manlo <= conv_std_logic_vector(180323091,28);
            exponent <= conv_std_logic_vector(1317,11);
      WHEN "0011001101" =>
            manhi <= conv_std_logic_vector(11487196,24);
            manlo <= conv_std_logic_vector(178245939,28);
            exponent <= conv_std_logic_vector(1318,11);
      WHEN "0011001110" =>
            manhi <= conv_std_logic_vector(2430443,24);
            manlo <= conv_std_logic_vector(223919964,28);
            exponent <= conv_std_logic_vector(1320,11);
      WHEN "0011001111" =>
            manhi <= conv_std_logic_vector(9328700,24);
            manlo <= conv_std_logic_vector(93205956,28);
            exponent <= conv_std_logic_vector(1321,11);
      WHEN "0011010000" =>
            manhi <= conv_std_logic_vector(963593,24);
            manlo <= conv_std_logic_vector(135688620,28);
            exponent <= conv_std_logic_vector(1323,11);
      WHEN "0011010001" =>
            manhi <= conv_std_logic_vector(7335044,24);
            manlo <= conv_std_logic_vector(13542358,28);
            exponent <= conv_std_logic_vector(1324,11);
      WHEN "0011010010" =>
            manhi <= conv_std_logic_vector(15994743,24);
            manlo <= conv_std_logic_vector(45394459,28);
            exponent <= conv_std_logic_vector(1325,11);
      WHEN "0011010011" =>
            manhi <= conv_std_logic_vector(5493639,24);
            manlo <= conv_std_logic_vector(73308838,28);
            exponent <= conv_std_logic_vector(1327,11);
      WHEN "0011010100" =>
            manhi <= conv_std_logic_vector(13492014,24);
            manlo <= conv_std_logic_vector(160135181,28);
            exponent <= conv_std_logic_vector(1328,11);
      WHEN "0011010101" =>
            manhi <= conv_std_logic_vector(3792858,24);
            manlo <= conv_std_logic_vector(234346738,28);
            exponent <= conv_std_logic_vector(1330,11);
      WHEN "0011010110" =>
            manhi <= conv_std_logic_vector(11180414,24);
            manlo <= conv_std_logic_vector(98964646,28);
            exponent <= conv_std_logic_vector(1331,11);
      WHEN "0011010111" =>
            manhi <= conv_std_logic_vector(2221963,24);
            manlo <= conv_std_logic_vector(174344531,28);
            exponent <= conv_std_logic_vector(1333,11);
      WHEN "0011011000" =>
            manhi <= conv_std_logic_vector(9045346,24);
            manlo <= conv_std_logic_vector(106947534,28);
            exponent <= conv_std_logic_vector(1334,11);
      WHEN "0011011001" =>
            manhi <= conv_std_logic_vector(771034,24);
            manlo <= conv_std_logic_vector(143065990,28);
            exponent <= conv_std_logic_vector(1336,11);
      WHEN "0011011010" =>
            manhi <= conv_std_logic_vector(7073329,24);
            manlo <= conv_std_logic_vector(73148434,28);
            exponent <= conv_std_logic_vector(1337,11);
      WHEN "0011011011" =>
            manhi <= conv_std_logic_vector(15639035,24);
            manlo <= conv_std_logic_vector(243346703,28);
            exponent <= conv_std_logic_vector(1338,11);
      WHEN "0011011100" =>
            manhi <= conv_std_logic_vector(5251911,24);
            manlo <= conv_std_logic_vector(33842377,28);
            exponent <= conv_std_logic_vector(1340,11);
      WHEN "0011011101" =>
            manhi <= conv_std_logic_vector(13163471,24);
            manlo <= conv_std_logic_vector(263552292,28);
            exponent <= conv_std_logic_vector(1341,11);
      WHEN "0011011110" =>
            manhi <= conv_std_logic_vector(3569591,24);
            manlo <= conv_std_logic_vector(4866264,28);
            exponent <= conv_std_logic_vector(1343,11);
      WHEN "0011011111" =>
            manhi <= conv_std_logic_vector(10876961,24);
            manlo <= conv_std_logic_vector(239517036,28);
            exponent <= conv_std_logic_vector(1344,11);
      WHEN "0011100000" =>
            manhi <= conv_std_logic_vector(2015746,24);
            manlo <= conv_std_logic_vector(83586287,28);
            exponent <= conv_std_logic_vector(1346,11);
      WHEN "0011100001" =>
            manhi <= conv_std_logic_vector(8765067,24);
            manlo <= conv_std_logic_vector(262254542,28);
            exponent <= conv_std_logic_vector(1347,11);
      WHEN "0011100010" =>
            manhi <= conv_std_logic_vector(580565,24);
            manlo <= conv_std_logic_vector(160521039,28);
            exponent <= conv_std_logic_vector(1349,11);
      WHEN "0011100011" =>
            manhi <= conv_std_logic_vector(6814455,24);
            manlo <= conv_std_logic_vector(40288155,28);
            exponent <= conv_std_logic_vector(1350,11);
      WHEN "0011100100" =>
            manhi <= conv_std_logic_vector(15287189,24);
            manlo <= conv_std_logic_vector(132910147,28);
            exponent <= conv_std_logic_vector(1351,11);
      WHEN "0011100101" =>
            manhi <= conv_std_logic_vector(5012806,24);
            manlo <= conv_std_logic_vector(187753904,28);
            exponent <= conv_std_logic_vector(1353,11);
      WHEN "0011100110" =>
            manhi <= conv_std_logic_vector(12838495,24);
            manlo <= conv_std_logic_vector(100071648,28);
            exponent <= conv_std_logic_vector(1354,11);
      WHEN "0011100111" =>
            manhi <= conv_std_logic_vector(3348746,24);
            manlo <= conv_std_logic_vector(138348888,28);
            exponent <= conv_std_logic_vector(1356,11);
      WHEN "0011101000" =>
            manhi <= conv_std_logic_vector(10576803,24);
            manlo <= conv_std_logic_vector(24941937,28);
            exponent <= conv_std_logic_vector(1357,11);
      WHEN "0011101001" =>
            manhi <= conv_std_logic_vector(1811767,24);
            manlo <= conv_std_logic_vector(69497619,28);
            exponent <= conv_std_logic_vector(1359,11);
      WHEN "0011101010" =>
            manhi <= conv_std_logic_vector(8487831,24);
            manlo <= conv_std_logic_vector(188199296,28);
            exponent <= conv_std_logic_vector(1360,11);
      WHEN "0011101011" =>
            manhi <= conv_std_logic_vector(392164,24);
            manlo <= conv_std_logic_vector(4096525,28);
            exponent <= conv_std_logic_vector(1362,11);
      WHEN "0011101100" =>
            manhi <= conv_std_logic_vector(6558390,24);
            manlo <= conv_std_logic_vector(228356857,28);
            exponent <= conv_std_logic_vector(1363,11);
      WHEN "0011101101" =>
            manhi <= conv_std_logic_vector(14939162,24);
            manlo <= conv_std_logic_vector(7826265,28);
            exponent <= conv_std_logic_vector(1364,11);
      WHEN "0011101110" =>
            manhi <= conv_std_logic_vector(4776297,24);
            manlo <= conv_std_logic_vector(138324122,28);
            exponent <= conv_std_logic_vector(1366,11);
      WHEN "0011101111" =>
            manhi <= conv_std_logic_vector(12517046,24);
            manlo <= conv_std_logic_vector(17190560,28);
            exponent <= conv_std_logic_vector(1367,11);
      WHEN "0011110000" =>
            manhi <= conv_std_logic_vector(3130299,24);
            manlo <= conv_std_logic_vector(16562242,28);
            exponent <= conv_std_logic_vector(1369,11);
      WHEN "0011110001" =>
            manhi <= conv_std_logic_vector(10279902,24);
            manlo <= conv_std_logic_vector(59323104,28);
            exponent <= conv_std_logic_vector(1370,11);
      WHEN "0011110010" =>
            manhi <= conv_std_logic_vector(1610002,24);
            manlo <= conv_std_logic_vector(53056333,28);
            exponent <= conv_std_logic_vector(1372,11);
      WHEN "0011110011" =>
            manhi <= conv_std_logic_vector(8213604,24);
            manlo <= conv_std_logic_vector(147986337,28);
            exponent <= conv_std_logic_vector(1373,11);
      WHEN "0011110100" =>
            manhi <= conv_std_logic_vector(205807,24);
            manlo <= conv_std_logic_vector(92802035,28);
            exponent <= conv_std_logic_vector(1375,11);
      WHEN "0011110101" =>
            manhi <= conv_std_logic_vector(6305105,24);
            manlo <= conv_std_logic_vector(235277170,28);
            exponent <= conv_std_logic_vector(1376,11);
      WHEN "0011110110" =>
            manhi <= conv_std_logic_vector(14594912,24);
            manlo <= conv_std_logic_vector(15497684,28);
            exponent <= conv_std_logic_vector(1377,11);
      WHEN "0011110111" =>
            manhi <= conv_std_logic_vector(4542355,24);
            manlo <= conv_std_logic_vector(108677892,28);
            exponent <= conv_std_logic_vector(1379,11);
      WHEN "0011111000" =>
            manhi <= conv_std_logic_vector(12199085,24);
            manlo <= conv_std_logic_vector(206743222,28);
            exponent <= conv_std_logic_vector(1380,11);
      WHEN "0011111001" =>
            manhi <= conv_std_logic_vector(2914222,24);
            manlo <= conv_std_logic_vector(171652524,28);
            exponent <= conv_std_logic_vector(1382,11);
      WHEN "0011111010" =>
            manhi <= conv_std_logic_vector(9986223,24);
            manlo <= conv_std_logic_vector(245598061,28);
            exponent <= conv_std_logic_vector(1383,11);
      WHEN "0011111011" =>
            manhi <= conv_std_logic_vector(1410427,24);
            manlo <= conv_std_logic_vector(26024388,28);
            exponent <= conv_std_logic_vector(1385,11);
      WHEN "0011111100" =>
            manhi <= conv_std_logic_vector(7942353,24);
            manlo <= conv_std_logic_vector(232590388,28);
            exponent <= conv_std_logic_vector(1386,11);
      WHEN "0011111101" =>
            manhi <= conv_std_logic_vector(21473,24);
            manlo <= conv_std_logic_vector(105719295,28);
            exponent <= conv_std_logic_vector(1388,11);
      WHEN "0011111110" =>
            manhi <= conv_std_logic_vector(6054570,24);
            manlo <= conv_std_logic_vector(16265786,28);
            exponent <= conv_std_logic_vector(1389,11);
      WHEN "0011111111" =>
            manhi <= conv_std_logic_vector(14254398,24);
            manlo <= conv_std_logic_vector(155662944,28);
            exponent <= conv_std_logic_vector(1390,11);
      WHEN "0100000000" =>
            manhi <= conv_std_logic_vector(4310952,24);
            manlo <= conv_std_logic_vector(135577274,28);
            exponent <= conv_std_logic_vector(1392,11);
      WHEN "0100000001" =>
            manhi <= conv_std_logic_vector(11884576,24);
            manlo <= conv_std_logic_vector(166805756,28);
            exponent <= conv_std_logic_vector(1393,11);
      WHEN "0100000010" =>
            manhi <= conv_std_logic_vector(2700491,24);
            manlo <= conv_std_logic_vector(137829044,28);
            exponent <= conv_std_logic_vector(1395,11);
      WHEN "0100000011" =>
            manhi <= conv_std_logic_vector(9695733,24);
            manlo <= conv_std_logic_vector(52863001,28);
            exponent <= conv_std_logic_vector(1396,11);
      WHEN "0100000100" =>
            manhi <= conv_std_logic_vector(1213018,24);
            manlo <= conv_std_logic_vector(50179603,28);
            exponent <= conv_std_logic_vector(1398,11);
      WHEN "0100000101" =>
            manhi <= conv_std_logic_vector(7674047,24);
            manlo <= conv_std_logic_vector(91276680,28);
            exponent <= conv_std_logic_vector(1399,11);
      WHEN "0100000110" =>
            manhi <= conv_std_logic_vector(16455496,24);
            manlo <= conv_std_logic_vector(110068760,28);
            exponent <= conv_std_logic_vector(1400,11);
      WHEN "0100000111" =>
            manhi <= conv_std_logic_vector(5806753,24);
            manlo <= conv_std_logic_vector(151304445,28);
            exponent <= conv_std_logic_vector(1402,11);
      WHEN "0100001000" =>
            manhi <= conv_std_logic_vector(13917581,24);
            manlo <= conv_std_logic_vector(10650184,28);
            exponent <= conv_std_logic_vector(1403,11);
      WHEN "0100001001" =>
            manhi <= conv_std_logic_vector(4082061,24);
            manlo <= conv_std_logic_vector(68530707,28);
            exponent <= conv_std_logic_vector(1405,11);
      WHEN "0100001010" =>
            manhi <= conv_std_logic_vector(11573481,24);
            manlo <= conv_std_logic_vector(42662756,28);
            exponent <= conv_std_logic_vector(1406,11);
      WHEN "0100001011" =>
            manhi <= conv_std_logic_vector(2489080,24);
            manlo <= conv_std_logic_vector(61154162,28);
            exponent <= conv_std_logic_vector(1408,11);
      WHEN "0100001100" =>
            manhi <= conv_std_logic_vector(9408395,24);
            manlo <= conv_std_logic_vector(125867240,28);
            exponent <= conv_std_logic_vector(1409,11);
      WHEN "0100001101" =>
            manhi <= conv_std_logic_vector(1017751,24);
            manlo <= conv_std_logic_vector(256555705,28);
            exponent <= conv_std_logic_vector(1411,11);
      WHEN "0100001110" =>
            manhi <= conv_std_logic_vector(7408653,24);
            manlo <= conv_std_logic_vector(4309896,28);
            exponent <= conv_std_logic_vector(1412,11);
      WHEN "0100001111" =>
            manhi <= conv_std_logic_vector(16094788,24);
            manlo <= conv_std_logic_vector(33800670,28);
            exponent <= conv_std_logic_vector(1413,11);
      WHEN "0100010000" =>
            manhi <= conv_std_logic_vector(5561626,24);
            manlo <= conv_std_logic_vector(233573192,28);
            exponent <= conv_std_logic_vector(1415,11);
      WHEN "0100010001" =>
            manhi <= conv_std_logic_vector(13584419,24);
            manlo <= conv_std_logic_vector(86257801,28);
            exponent <= conv_std_logic_vector(1416,11);
      WHEN "0100010010" =>
            manhi <= conv_std_logic_vector(3855654,24);
            manlo <= conv_std_logic_vector(105782775,28);
            exponent <= conv_std_logic_vector(1418,11);
      WHEN "0100010011" =>
            manhi <= conv_std_logic_vector(11265762,24);
            manlo <= conv_std_logic_vector(88738762,28);
            exponent <= conv_std_logic_vector(1419,11);
      WHEN "0100010100" =>
            manhi <= conv_std_logic_vector(2279963,24);
            manlo <= conv_std_logic_vector(161858527,28);
            exponent <= conv_std_logic_vector(1421,11);
      WHEN "0100010101" =>
            manhi <= conv_std_logic_vector(9124176,24);
            manlo <= conv_std_logic_vector(136423424,28);
            exponent <= conv_std_logic_vector(1422,11);
      WHEN "0100010110" =>
            manhi <= conv_std_logic_vector(824605,24);
            manlo <= conv_std_logic_vector(39384255,28);
            exponent <= conv_std_logic_vector(1424,11);
      WHEN "0100010111" =>
            manhi <= conv_std_logic_vector(7146139,24);
            manlo <= conv_std_logic_vector(76626123,28);
            exponent <= conv_std_logic_vector(1425,11);
      WHEN "0100011000" =>
            manhi <= conv_std_logic_vector(15737994,24);
            manlo <= conv_std_logic_vector(261485765,28);
            exponent <= conv_std_logic_vector(1426,11);
      WHEN "0100011001" =>
            manhi <= conv_std_logic_vector(5319160,24);
            manlo <= conv_std_logic_vector(210684009,28);
            exponent <= conv_std_logic_vector(1428,11);
      WHEN "0100011010" =>
            manhi <= conv_std_logic_vector(13254873,24);
            manlo <= conv_std_logic_vector(199859160,28);
            exponent <= conv_std_logic_vector(1429,11);
      WHEN "0100011011" =>
            manhi <= conv_std_logic_vector(3631704,24);
            manlo <= conv_std_logic_vector(256571707,28);
            exponent <= conv_std_logic_vector(1431,11);
      WHEN "0100011100" =>
            manhi <= conv_std_logic_vector(10961383,24);
            manlo <= conv_std_logic_vector(130542749,28);
            exponent <= conv_std_logic_vector(1432,11);
      WHEN "0100011101" =>
            manhi <= conv_std_logic_vector(2073116,24);
            manlo <= conv_std_logic_vector(196665136,28);
            exponent <= conv_std_logic_vector(1434,11);
      WHEN "0100011110" =>
            manhi <= conv_std_logic_vector(8843042,24);
            manlo <= conv_std_logic_vector(124490661,28);
            exponent <= conv_std_logic_vector(1435,11);
      WHEN "0100011111" =>
            manhi <= conv_std_logic_vector(633554,24);
            manlo <= conv_std_logic_vector(202834752,28);
            exponent <= conv_std_logic_vector(1437,11);
      WHEN "0100100000" =>
            manhi <= conv_std_logic_vector(6886474,24);
            manlo <= conv_std_logic_vector(236822279,28);
            exponent <= conv_std_logic_vector(1438,11);
      WHEN "0100100001" =>
            manhi <= conv_std_logic_vector(15385074,24);
            manlo <= conv_std_logic_vector(123405487,28);
            exponent <= conv_std_logic_vector(1439,11);
      WHEN "0100100010" =>
            manhi <= conv_std_logic_vector(5079326,24);
            manlo <= conv_std_logic_vector(115311954,28);
            exponent <= conv_std_logic_vector(1441,11);
      WHEN "0100100011" =>
            manhi <= conv_std_logic_vector(12928905,24);
            manlo <= conv_std_logic_vector(16004876,28);
            exponent <= conv_std_logic_vector(1442,11);
      WHEN "0100100100" =>
            manhi <= conv_std_logic_vector(3410186,24);
            manlo <= conv_std_logic_vector(71831800,28);
            exponent <= conv_std_logic_vector(1444,11);
      WHEN "0100100101" =>
            manhi <= conv_std_logic_vector(10660308,24);
            manlo <= conv_std_logic_vector(100367284,28);
            exponent <= conv_std_logic_vector(1445,11);
      WHEN "0100100110" =>
            manhi <= conv_std_logic_vector(1868514,24);
            manlo <= conv_std_logic_vector(263299419,28);
            exponent <= conv_std_logic_vector(1447,11);
      WHEN "0100100111" =>
            manhi <= conv_std_logic_vector(8564959,24);
            manlo <= conv_std_logic_vector(228656810,28);
            exponent <= conv_std_logic_vector(1448,11);
      WHEN "0100101000" =>
            manhi <= conv_std_logic_vector(444578,24);
            manlo <= conv_std_logic_vector(7489141,28);
            exponent <= conv_std_logic_vector(1450,11);
      WHEN "0100101001" =>
            manhi <= conv_std_logic_vector(6629628,24);
            manlo <= conv_std_logic_vector(236156491,28);
            exponent <= conv_std_logic_vector(1451,11);
      WHEN "0100101010" =>
            manhi <= conv_std_logic_vector(15035984,24);
            manlo <= conv_std_logic_vector(147396312,28);
            exponent <= conv_std_logic_vector(1452,11);
      WHEN "0100101011" =>
            manhi <= conv_std_logic_vector(4842095,24);
            manlo <= conv_std_logic_vector(64271882,28);
            exponent <= conv_std_logic_vector(1454,11);
      WHEN "0100101100" =>
            manhi <= conv_std_logic_vector(12606474,24);
            manlo <= conv_std_logic_vector(118909770,28);
            exponent <= conv_std_logic_vector(1455,11);
      WHEN "0100101101" =>
            manhi <= conv_std_logic_vector(3191071,24);
            manlo <= conv_std_logic_vector(253953386,28);
            exponent <= conv_std_logic_vector(1457,11);
      WHEN "0100101110" =>
            manhi <= conv_std_logic_vector(10362501,24);
            manlo <= conv_std_logic_vector(36129498,28);
            exponent <= conv_std_logic_vector(1458,11);
      WHEN "0100101111" =>
            manhi <= conv_std_logic_vector(1666133,24);
            manlo <= conv_std_logic_vector(262830684,28);
            exponent <= conv_std_logic_vector(1460,11);
      WHEN "0100110000" =>
            manhi <= conv_std_logic_vector(8289895,24);
            manlo <= conv_std_logic_vector(148197046,28);
            exponent <= conv_std_logic_vector(1461,11);
      WHEN "0100110001" =>
            manhi <= conv_std_logic_vector(257652,24);
            manlo <= conv_std_logic_vector(122404338,28);
            exponent <= conv_std_logic_vector(1463,11);
      WHEN "0100110010" =>
            manhi <= conv_std_logic_vector(6375570,24);
            manlo <= conv_std_logic_vector(184430245,28);
            exponent <= conv_std_logic_vector(1464,11);
      WHEN "0100110011" =>
            manhi <= conv_std_logic_vector(14690683,24);
            manlo <= conv_std_logic_vector(178457687,28);
            exponent <= conv_std_logic_vector(1465,11);
      WHEN "0100110100" =>
            manhi <= conv_std_logic_vector(4607438,24);
            manlo <= conv_std_logic_vector(257605193,28);
            exponent <= conv_std_logic_vector(1467,11);
      WHEN "0100110101" =>
            manhi <= conv_std_logic_vector(12287543,24);
            manlo <= conv_std_logic_vector(132163446,28);
            exponent <= conv_std_logic_vector(1468,11);
      WHEN "0100110110" =>
            manhi <= conv_std_logic_vector(2974335,24);
            manlo <= conv_std_logic_vector(240020217,28);
            exponent <= conv_std_logic_vector(1470,11);
      WHEN "0100110111" =>
            manhi <= conv_std_logic_vector(10067926,24);
            manlo <= conv_std_logic_vector(80224641,28);
            exponent <= conv_std_logic_vector(1471,11);
      WHEN "0100111000" =>
            manhi <= conv_std_logic_vector(1465949,24);
            manlo <= conv_std_logic_vector(167328478,28);
            exponent <= conv_std_logic_vector(1473,11);
      WHEN "0100111001" =>
            manhi <= conv_std_logic_vector(8017816,24);
            manlo <= conv_std_logic_vector(215756784,28);
            exponent <= conv_std_logic_vector(1474,11);
      WHEN "0100111010" =>
            manhi <= conv_std_logic_vector(72755,24);
            manlo <= conv_std_logic_vector(208473528,28);
            exponent <= conv_std_logic_vector(1476,11);
      WHEN "0100111011" =>
            manhi <= conv_std_logic_vector(6124270,24);
            manlo <= conv_std_logic_vector(12139444,28);
            exponent <= conv_std_logic_vector(1477,11);
      WHEN "0100111100" =>
            manhi <= conv_std_logic_vector(14349130,24);
            manlo <= conv_std_logic_vector(182729110,28);
            exponent <= conv_std_logic_vector(1478,11);
      WHEN "0100111101" =>
            manhi <= conv_std_logic_vector(4375329,24);
            manlo <= conv_std_logic_vector(172370119,28);
            exponent <= conv_std_logic_vector(1480,11);
      WHEN "0100111110" =>
            manhi <= conv_std_logic_vector(11972074,24);
            manlo <= conv_std_logic_vector(59679792,28);
            exponent <= conv_std_logic_vector(1481,11);
      WHEN "0100111111" =>
            manhi <= conv_std_logic_vector(2759952,24);
            manlo <= conv_std_logic_vector(80023302,28);
            exponent <= conv_std_logic_vector(1483,11);
      WHEN "0101000000" =>
            manhi <= conv_std_logic_vector(9776548,24);
            manlo <= conv_std_logic_vector(209956608,28);
            exponent <= conv_std_logic_vector(1484,11);
      WHEN "0101000001" =>
            manhi <= conv_std_logic_vector(1267938,24);
            manlo <= conv_std_logic_vector(19091951,28);
            exponent <= conv_std_logic_vector(1486,11);
      WHEN "0101000010" =>
            manhi <= conv_std_logic_vector(7748691,24);
            manlo <= conv_std_logic_vector(54127000,28);
            exponent <= conv_std_logic_vector(1487,11);
      WHEN "0101000011" =>
            manhi <= conv_std_logic_vector(16556947,24);
            manlo <= conv_std_logic_vector(251347868,28);
            exponent <= conv_std_logic_vector(1488,11);
      WHEN "0101000100" =>
            manhi <= conv_std_logic_vector(5875697,24);
            manlo <= conv_std_logic_vector(6377900,28);
            exponent <= conv_std_logic_vector(1490,11);
      WHEN "0101000101" =>
            manhi <= conv_std_logic_vector(14011284,24);
            manlo <= conv_std_logic_vector(246175281,28);
            exponent <= conv_std_logic_vector(1491,11);
      WHEN "0101000110" =>
            manhi <= conv_std_logic_vector(4145739,24);
            manlo <= conv_std_logic_vector(172360927,28);
            exponent <= conv_std_logic_vector(1493,11);
      WHEN "0101000111" =>
            manhi <= conv_std_logic_vector(11660029,24);
            manlo <= conv_std_logic_vector(16047086,28);
            exponent <= conv_std_logic_vector(1494,11);
      WHEN "0101001000" =>
            manhi <= conv_std_logic_vector(2547895,24);
            manlo <= conv_std_logic_vector(167600151,28);
            exponent <= conv_std_logic_vector(1496,11);
      WHEN "0101001001" =>
            manhi <= conv_std_logic_vector(9488333,24);
            manlo <= conv_std_logic_vector(236416250,28);
            exponent <= conv_std_logic_vector(1497,11);
      WHEN "0101001010" =>
            manhi <= conv_std_logic_vector(1072075,24);
            manlo <= conv_std_logic_vector(198323037,28);
            exponent <= conv_std_logic_vector(1499,11);
      WHEN "0101001011" =>
            manhi <= conv_std_logic_vector(7482486,24);
            manlo <= conv_std_logic_vector(185820926,28);
            exponent <= conv_std_logic_vector(1500,11);
      WHEN "0101001100" =>
            manhi <= conv_std_logic_vector(16195138,24);
            manlo <= conv_std_logic_vector(133160968,28);
            exponent <= conv_std_logic_vector(1501,11);
      WHEN "0101001101" =>
            manhi <= conv_std_logic_vector(5629822,24);
            manlo <= conv_std_logic_vector(4574050,28);
            exponent <= conv_std_logic_vector(1503,11);
      WHEN "0101001110" =>
            manhi <= conv_std_logic_vector(13677106,24);
            manlo <= conv_std_logic_vector(36414601,28);
            exponent <= conv_std_logic_vector(1504,11);
      WHEN "0101001111" =>
            manhi <= conv_std_logic_vector(3918641,24);
            manlo <= conv_std_logic_vector(165046798,28);
            exponent <= conv_std_logic_vector(1506,11);
      WHEN "0101010000" =>
            manhi <= conv_std_logic_vector(11351370,24);
            manlo <= conv_std_logic_vector(225326735,28);
            exponent <= conv_std_logic_vector(1507,11);
      WHEN "0101010001" =>
            manhi <= conv_std_logic_vector(2338140,24);
            manlo <= conv_std_logic_vector(165476611,28);
            exponent <= conv_std_logic_vector(1509,11);
      WHEN "0101010010" =>
            manhi <= conv_std_logic_vector(9203247,24);
            manlo <= conv_std_logic_vector(71807303,28);
            exponent <= conv_std_logic_vector(1510,11);
      WHEN "0101010011" =>
            manhi <= conv_std_logic_vector(878339,24);
            manlo <= conv_std_logic_vector(80195176,28);
            exponent <= conv_std_logic_vector(1512,11);
      WHEN "0101010100" =>
            manhi <= conv_std_logic_vector(7219171,24);
            manlo <= conv_std_logic_vector(153001068,28);
            exponent <= conv_std_logic_vector(1513,11);
      WHEN "0101010101" =>
            manhi <= conv_std_logic_vector(15837256,24);
            manlo <= conv_std_logic_vector(37596960,28);
            exponent <= conv_std_logic_vector(1514,11);
      WHEN "0101010110" =>
            manhi <= conv_std_logic_vector(5386615,24);
            manlo <= conv_std_logic_vector(198850796,28);
            exponent <= conv_std_logic_vector(1516,11);
      WHEN "0101010111" =>
            manhi <= conv_std_logic_vector(13346554,24);
            manlo <= conv_std_logic_vector(143609986,28);
            exponent <= conv_std_logic_vector(1517,11);
      WHEN "0101011000" =>
            manhi <= conv_std_logic_vector(3694008,24);
            manlo <= conv_std_logic_vector(137568494,28);
            exponent <= conv_std_logic_vector(1519,11);
      WHEN "0101011001" =>
            manhi <= conv_std_logic_vector(11046062,24);
            manlo <= conv_std_logic_vector(214558683,28);
            exponent <= conv_std_logic_vector(1520,11);
      WHEN "0101011010" =>
            manhi <= conv_std_logic_vector(2130662,24);
            manlo <= conv_std_logic_vector(78401205,28);
            exponent <= conv_std_logic_vector(1522,11);
      WHEN "0101011011" =>
            manhi <= conv_std_logic_vector(8921254,24);
            manlo <= conv_std_logic_vector(265219821,28);
            exponent <= conv_std_logic_vector(1523,11);
      WHEN "0101011100" =>
            manhi <= conv_std_logic_vector(686705,24);
            manlo <= conv_std_logic_vector(181591149,28);
            exponent <= conv_std_logic_vector(1525,11);
      WHEN "0101011101" =>
            manhi <= conv_std_logic_vector(6958714,24);
            manlo <= conv_std_logic_vector(127078273,28);
            exponent <= conv_std_logic_vector(1526,11);
      WHEN "0101011110" =>
            manhi <= conv_std_logic_vector(15483258,24);
            manlo <= conv_std_logic_vector(65420394,28);
            exponent <= conv_std_logic_vector(1527,11);
      WHEN "0101011111" =>
            manhi <= conv_std_logic_vector(5146049,24);
            manlo <= conv_std_logic_vector(61347424,28);
            exponent <= conv_std_logic_vector(1529,11);
      WHEN "0101100000" =>
            manhi <= conv_std_logic_vector(13019590,24);
            manlo <= conv_std_logic_vector(200148168,28);
            exponent <= conv_std_logic_vector(1530,11);
      WHEN "0101100001" =>
            manhi <= conv_std_logic_vector(3471813,24);
            manlo <= conv_std_logic_vector(155873600,28);
            exponent <= conv_std_logic_vector(1532,11);
      WHEN "0101100010" =>
            manhi <= conv_std_logic_vector(10744068,24);
            manlo <= conv_std_logic_vector(154763366,28);
            exponent <= conv_std_logic_vector(1533,11);
      WHEN "0101100011" =>
            manhi <= conv_std_logic_vector(1925435,24);
            manlo <= conv_std_logic_vector(252346422,28);
            exponent <= conv_std_logic_vector(1535,11);
      WHEN "0101100100" =>
            manhi <= conv_std_logic_vector(8642323,24);
            manlo <= conv_std_logic_vector(122496413,28);
            exponent <= conv_std_logic_vector(1536,11);
      WHEN "0101100101" =>
            manhi <= conv_std_logic_vector(497152,24);
            manlo <= conv_std_logic_vector(12881703,28);
            exponent <= conv_std_logic_vector(1538,11);
      WHEN "0101100110" =>
            manhi <= conv_std_logic_vector(6701084,24);
            manlo <= conv_std_logic_vector(102402698,28);
            exponent <= conv_std_logic_vector(1539,11);
      WHEN "0101100111" =>
            manhi <= conv_std_logic_vector(15133102,24);
            manlo <= conv_std_logic_vector(173151546,28);
            exponent <= conv_std_logic_vector(1540,11);
      WHEN "0101101000" =>
            manhi <= conv_std_logic_vector(4908093,24);
            manlo <= conv_std_logic_vector(222341698,28);
            exponent <= conv_std_logic_vector(1542,11);
      WHEN "0101101001" =>
            manhi <= conv_std_logic_vector(12696175,24);
            manlo <= conv_std_logic_vector(221558290,28);
            exponent <= conv_std_logic_vector(1543,11);
      WHEN "0101101010" =>
            manhi <= conv_std_logic_vector(3252030,24);
            manlo <= conv_std_logic_vector(95425703,28);
            exponent <= conv_std_logic_vector(1545,11);
      WHEN "0101101011" =>
            manhi <= conv_std_logic_vector(10445352,24);
            manlo <= conv_std_logic_vector(54472775,28);
            exponent <= conv_std_logic_vector(1546,11);
      WHEN "0101101100" =>
            manhi <= conv_std_logic_vector(1722437,24);
            manlo <= conv_std_logic_vector(31541381,28);
            exponent <= conv_std_logic_vector(1548,11);
      WHEN "0101101101" =>
            manhi <= conv_std_logic_vector(8366419,24);
            manlo <= conv_std_logic_vector(121077564,28);
            exponent <= conv_std_logic_vector(1549,11);
      WHEN "0101101110" =>
            manhi <= conv_std_logic_vector(309655,24);
            manlo <= conv_std_logic_vector(224679493,28);
            exponent <= conv_std_logic_vector(1551,11);
      WHEN "0101101111" =>
            manhi <= conv_std_logic_vector(6446250,24);
            manlo <= conv_std_logic_vector(163707479,28);
            exponent <= conv_std_logic_vector(1552,11);
      WHEN "0101110000" =>
            manhi <= conv_std_logic_vector(14786747,24);
            manlo <= conv_std_logic_vector(171718440,28);
            exponent <= conv_std_logic_vector(1553,11);
      WHEN "0101110001" =>
            manhi <= conv_std_logic_vector(4672721,24);
            manlo <= conv_std_logic_vector(53414720,28);
            exponent <= conv_std_logic_vector(1555,11);
      WHEN "0101110010" =>
            manhi <= conv_std_logic_vector(12376271,24);
            manlo <= conv_std_logic_vector(68395953,28);
            exponent <= conv_std_logic_vector(1556,11);
      WHEN "0101110011" =>
            manhi <= conv_std_logic_vector(3034632,24);
            manlo <= conv_std_logic_vector(177229210,28);
            exponent <= conv_std_logic_vector(1558,11);
      WHEN "0101110100" =>
            manhi <= conv_std_logic_vector(10149878,24);
            manlo <= conv_std_logic_vector(27015960,28);
            exponent <= conv_std_logic_vector(1559,11);
      WHEN "0101110101" =>
            manhi <= conv_std_logic_vector(1521641,24);
            manlo <= conv_std_logic_vector(173609470,28);
            exponent <= conv_std_logic_vector(1561,11);
      WHEN "0101110110" =>
            manhi <= conv_std_logic_vector(8093510,24);
            manlo <= conv_std_logic_vector(29891310,28);
            exponent <= conv_std_logic_vector(1562,11);
      WHEN "0101110111" =>
            manhi <= conv_std_logic_vector(124194,24);
            manlo <= conv_std_logic_vector(191198183,28);
            exponent <= conv_std_logic_vector(1564,11);
      WHEN "0101111000" =>
            manhi <= conv_std_logic_vector(6194182,24);
            manlo <= conv_std_logic_vector(216692261,28);
            exponent <= conv_std_logic_vector(1565,11);
      WHEN "0101111001" =>
            manhi <= conv_std_logic_vector(14444151,24);
            manlo <= conv_std_logic_vector(261994424,28);
            exponent <= conv_std_logic_vector(1566,11);
      WHEN "0101111010" =>
            manhi <= conv_std_logic_vector(4439903,24);
            manlo <= conv_std_logic_vector(82463931,28);
            exponent <= conv_std_logic_vector(1568,11);
      WHEN "0101111011" =>
            manhi <= conv_std_logic_vector(12059838,24);
            manlo <= conv_std_logic_vector(250318074,28);
            exponent <= conv_std_logic_vector(1569,11);
      WHEN "0101111100" =>
            manhi <= conv_std_logic_vector(2819594,24);
            manlo <= conv_std_logic_vector(161686084,28);
            exponent <= conv_std_logic_vector(1571,11);
      WHEN "0101111101" =>
            manhi <= conv_std_logic_vector(9857611,24);
            manlo <= conv_std_logic_vector(20946108,28);
            exponent <= conv_std_logic_vector(1572,11);
      WHEN "0101111110" =>
            manhi <= conv_std_logic_vector(1323025,24);
            manlo <= conv_std_logic_vector(164440795,28);
            exponent <= conv_std_logic_vector(1574,11);
      WHEN "0101111111" =>
            manhi <= conv_std_logic_vector(7823562,24);
            manlo <= conv_std_logic_vector(250479918,28);
            exponent <= conv_std_logic_vector(1575,11);
      WHEN "0110000000" =>
            manhi <= conv_std_logic_vector(16658709,24);
            manlo <= conv_std_logic_vector(45608811,28);
            exponent <= conv_std_logic_vector(1576,11);
      WHEN "0110000001" =>
            manhi <= conv_std_logic_vector(5944850,24);
            manlo <= conv_std_logic_vector(255488281,28);
            exponent <= conv_std_logic_vector(1578,11);
      WHEN "0110000010" =>
            manhi <= conv_std_logic_vector(14105274,24);
            manlo <= conv_std_logic_vector(228172930,28);
            exponent <= conv_std_logic_vector(1579,11);
      WHEN "0110000011" =>
            manhi <= conv_std_logic_vector(4209612,24);
            manlo <= conv_std_logic_vector(113758652,28);
            exponent <= conv_std_logic_vector(1581,11);
      WHEN "0110000100" =>
            manhi <= conv_std_logic_vector(11746841,24);
            manlo <= conv_std_logic_vector(45816542,28);
            exponent <= conv_std_logic_vector(1582,11);
      WHEN "0110000101" =>
            manhi <= conv_std_logic_vector(2606890,24);
            manlo <= conv_std_logic_vector(153074390,28);
            exponent <= conv_std_logic_vector(1584,11);
      WHEN "0110000110" =>
            manhi <= conv_std_logic_vector(9568516,24);
            manlo <= conv_std_logic_vector(87350878,28);
            exponent <= conv_std_logic_vector(1585,11);
      WHEN "0110000111" =>
            manhi <= conv_std_logic_vector(1126565,24);
            manlo <= conv_std_logic_vector(96475766,28);
            exponent <= conv_std_logic_vector(1587,11);
      WHEN "0110001000" =>
            manhi <= conv_std_logic_vector(7556545,24);
            manlo <= conv_std_logic_vector(205347948,28);
            exponent <= conv_std_logic_vector(1588,11);
      WHEN "0110001001" =>
            manhi <= conv_std_logic_vector(16295795,24);
            manlo <= conv_std_logic_vector(56881285,28);
            exponent <= conv_std_logic_vector(1589,11);
      WHEN "0110001010" =>
            manhi <= conv_std_logic_vector(5698225,24);
            manlo <= conv_std_logic_vector(93263076,28);
            exponent <= conv_std_logic_vector(1591,11);
      WHEN "0110001011" =>
            manhi <= conv_std_logic_vector(13770075,24);
            manlo <= conv_std_logic_vector(241769289,28);
            exponent <= conv_std_logic_vector(1592,11);
      WHEN "0110001100" =>
            manhi <= conv_std_logic_vector(3981821,24);
            manlo <= conv_std_logic_vector(32359920,28);
            exponent <= conv_std_logic_vector(1594,11);
      WHEN "0110001101" =>
            manhi <= conv_std_logic_vector(11437240,24);
            manlo <= conv_std_logic_vector(185367850,28);
            exponent <= conv_std_logic_vector(1595,11);
      WHEN "0110001110" =>
            manhi <= conv_std_logic_vector(2396495,24);
            manlo <= conv_std_logic_vector(61858550,28);
            exponent <= conv_std_logic_vector(1597,11);
      WHEN "0110001111" =>
            manhi <= conv_std_logic_vector(9282559,24);
            manlo <= conv_std_logic_vector(110304027,28);
            exponent <= conv_std_logic_vector(1598,11);
      WHEN "0110010000" =>
            manhi <= conv_std_logic_vector(932237,24);
            manlo <= conv_std_logic_vector(131077892,28);
            exponent <= conv_std_logic_vector(1600,11);
      WHEN "0110010001" =>
            manhi <= conv_std_logic_vector(7292426,24);
            manlo <= conv_std_logic_vector(215982528,28);
            exponent <= conv_std_logic_vector(1601,11);
      WHEN "0110010010" =>
            manhi <= conv_std_logic_vector(15936820,24);
            manlo <= conv_std_logic_vector(87676082,28);
            exponent <= conv_std_logic_vector(1602,11);
      WHEN "0110010011" =>
            manhi <= conv_std_logic_vector(5454276,24);
            manlo <= conv_std_logic_vector(166577430,28);
            exponent <= conv_std_logic_vector(1604,11);
      WHEN "0110010100" =>
            manhi <= conv_std_logic_vector(13438515,24);
            manlo <= conv_std_logic_vector(55023964,28);
            exponent <= conv_std_logic_vector(1605,11);
      WHEN "0110010101" =>
            manhi <= conv_std_logic_vector(3756502,24);
            manlo <= conv_std_logic_vector(71679026,28);
            exponent <= conv_std_logic_vector(1607,11);
      WHEN "0110010110" =>
            manhi <= conv_std_logic_vector(11131000,24);
            manlo <= conv_std_logic_vector(165886683,28);
            exponent <= conv_std_logic_vector(1608,11);
      WHEN "0110010111" =>
            manhi <= conv_std_logic_vector(2188383,24);
            manlo <= conv_std_logic_vector(140750309,28);
            exponent <= conv_std_logic_vector(1610,11);
      WHEN "0110011000" =>
            manhi <= conv_std_logic_vector(8999706,24);
            manlo <= conv_std_logic_vector(74200045,28);
            exponent <= conv_std_logic_vector(1611,11);
      WHEN "0110011001" =>
            manhi <= conv_std_logic_vector(740018,24);
            manlo <= conv_std_logic_vector(229350227,28);
            exponent <= conv_std_logic_vector(1613,11);
      WHEN "0110011010" =>
            manhi <= conv_std_logic_vector(7031174,24);
            manlo <= conv_std_logic_vector(159659309,28);
            exponent <= conv_std_logic_vector(1614,11);
      WHEN "0110011011" =>
            manhi <= conv_std_logic_vector(15581741,24);
            manlo <= conv_std_logic_vector(203828183,28);
            exponent <= conv_std_logic_vector(1615,11);
      WHEN "0110011100" =>
            manhi <= conv_std_logic_vector(5212975,24);
            manlo <= conv_std_logic_vector(192268981,28);
            exponent <= conv_std_logic_vector(1617,11);
      WHEN "0110011101" =>
            manhi <= conv_std_logic_vector(13110553,24);
            manlo <= conv_std_logic_vector(73367990,28);
            exponent <= conv_std_logic_vector(1618,11);
      WHEN "0110011110" =>
            manhi <= conv_std_logic_vector(3533629,24);
            manlo <= conv_std_logic_vector(7303751,28);
            exponent <= conv_std_logic_vector(1620,11);
      WHEN "0110011111" =>
            manhi <= conv_std_logic_vector(10828084,24);
            manlo <= conv_std_logic_vector(128595197,28);
            exponent <= conv_std_logic_vector(1621,11);
      WHEN "0110100000" =>
            manhi <= conv_std_logic_vector(1982530,24);
            manlo <= conv_std_logic_vector(178601213,28);
            exponent <= conv_std_logic_vector(1623,11);
      WHEN "0110100001" =>
            manhi <= conv_std_logic_vector(8719923,24);
            manlo <= conv_std_logic_vector(62665264,28);
            exponent <= conv_std_logic_vector(1624,11);
      WHEN "0110100010" =>
            manhi <= conv_std_logic_vector(549886,24);
            manlo <= conv_std_logic_vector(151395401,28);
            exponent <= conv_std_logic_vector(1626,11);
      WHEN "0110100011" =>
            manhi <= conv_std_logic_vector(6772758,24);
            manlo <= conv_std_logic_vector(5307652,28);
            exponent <= conv_std_logic_vector(1627,11);
      WHEN "0110100100" =>
            manhi <= conv_std_logic_vector(15230517,24);
            manlo <= conv_std_logic_vector(58871965,28);
            exponent <= conv_std_logic_vector(1628,11);
      WHEN "0110100101" =>
            manhi <= conv_std_logic_vector(4974293,24);
            manlo <= conv_std_logic_vector(240265124,28);
            exponent <= conv_std_logic_vector(1630,11);
      WHEN "0110100110" =>
            manhi <= conv_std_logic_vector(12786151,24);
            manlo <= conv_std_logic_vector(11983156,28);
            exponent <= conv_std_logic_vector(1631,11);
      WHEN "0110100111" =>
            manhi <= conv_std_logic_vector(3313174,24);
            manlo <= conv_std_logic_vector(229882212,28);
            exponent <= conv_std_logic_vector(1633,11);
      WHEN "0110101000" =>
            manhi <= conv_std_logic_vector(10528456,24);
            manlo <= conv_std_logic_vector(52550536,28);
            exponent <= conv_std_logic_vector(1634,11);
      WHEN "0110101001" =>
            manhi <= conv_std_logic_vector(1778912,24);
            manlo <= conv_std_logic_vector(36481057,28);
            exponent <= conv_std_logic_vector(1636,11);
      WHEN "0110101010" =>
            manhi <= conv_std_logic_vector(8443176,24);
            manlo <= conv_std_logic_vector(257480801,28);
            exponent <= conv_std_logic_vector(1637,11);
      WHEN "0110101011" =>
            manhi <= conv_std_logic_vector(361817,24);
            manlo <= conv_std_logic_vector(260890045,28);
            exponent <= conv_std_logic_vector(1639,11);
      WHEN "0110101100" =>
            manhi <= conv_std_logic_vector(6517146,24);
            manlo <= conv_std_logic_vector(80951272,28);
            exponent <= conv_std_logic_vector(1640,11);
      WHEN "0110101101" =>
            manhi <= conv_std_logic_vector(14883104,24);
            manlo <= conv_std_logic_vector(234866389,28);
            exponent <= conv_std_logic_vector(1641,11);
      WHEN "0110101110" =>
            manhi <= conv_std_logic_vector(4738202,24);
            manlo <= conv_std_logic_vector(195793257,28);
            exponent <= conv_std_logic_vector(1643,11);
      WHEN "0110101111" =>
            manhi <= conv_std_logic_vector(12465269,24);
            manlo <= conv_std_logic_vector(236730454,28);
            exponent <= conv_std_logic_vector(1644,11);
      WHEN "0110110000" =>
            manhi <= conv_std_logic_vector(3095113,24);
            manlo <= conv_std_logic_vector(133661452,28);
            exponent <= conv_std_logic_vector(1646,11);
      WHEN "0110110001" =>
            manhi <= conv_std_logic_vector(10232080,24);
            manlo <= conv_std_logic_vector(21926822,28);
            exponent <= conv_std_logic_vector(1647,11);
      WHEN "0110110010" =>
            manhi <= conv_std_logic_vector(1577503,24);
            manlo <= conv_std_logic_vector(183764948,28);
            exponent <= conv_std_logic_vector(1649,11);
      WHEN "0110110011" =>
            manhi <= conv_std_logic_vector(8169434,24);
            manlo <= conv_std_logic_vector(132210812,28);
            exponent <= conv_std_logic_vector(1650,11);
      WHEN "0110110100" =>
            manhi <= conv_std_logic_vector(175790,24);
            manlo <= conv_std_logic_vector(182183516,28);
            exponent <= conv_std_logic_vector(1652,11);
      WHEN "0110110101" =>
            manhi <= conv_std_logic_vector(6264308,24);
            manlo <= conv_std_logic_vector(267417858,28);
            exponent <= conv_std_logic_vector(1653,11);
      WHEN "0110110110" =>
            manhi <= conv_std_logic_vector(14539463,24);
            manlo <= conv_std_logic_vector(93573944,28);
            exponent <= conv_std_logic_vector(1654,11);
      WHEN "0110110111" =>
            manhi <= conv_std_logic_vector(4504674,24);
            manlo <= conv_std_logic_vector(26907375,28);
            exponent <= conv_std_logic_vector(1656,11);
      WHEN "0110111000" =>
            manhi <= conv_std_logic_vector(12147871,24);
            manlo <= conv_std_logic_vector(152302066,28);
            exponent <= conv_std_logic_vector(1657,11);
      WHEN "0110111001" =>
            manhi <= conv_std_logic_vector(2879418,24);
            manlo <= conv_std_logic_vector(263131635,28);
            exponent <= conv_std_logic_vector(1659,11);
      WHEN "0110111010" =>
            manhi <= conv_std_logic_vector(9938920,24);
            manlo <= conv_std_logic_vector(224874222,28);
            exponent <= conv_std_logic_vector(1660,11);
      WHEN "0110111011" =>
            manhi <= conv_std_logic_vector(1378281,24);
            manlo <= conv_std_logic_vector(86745210,28);
            exponent <= conv_std_logic_vector(1662,11);
      WHEN "0110111100" =>
            manhi <= conv_std_logic_vector(7898663,24);
            manlo <= conv_std_logic_vector(61761420,28);
            exponent <= conv_std_logic_vector(1663,11);
      WHEN "0110111101" =>
            manhi <= conv_std_logic_vector(16760781,24);
            manlo <= conv_std_logic_vector(15082626,28);
            exponent <= conv_std_logic_vector(1664,11);
      WHEN "0110111110" =>
            manhi <= conv_std_logic_vector(6014215,24);
            manlo <= conv_std_logic_vector(265801199,28);
            exponent <= conv_std_logic_vector(1666,11);
      WHEN "0110111111" =>
            manhi <= conv_std_logic_vector(14199551,24);
            manlo <= conv_std_logic_vector(191056853,28);
            exponent <= conv_std_logic_vector(1667,11);
      WHEN "0111000000" =>
            manhi <= conv_std_logic_vector(4273680,24);
            manlo <= conv_std_logic_vector(52024524,28);
            exponent <= conv_std_logic_vector(1669,11);
      WHEN "0111000001" =>
            manhi <= conv_std_logic_vector(11833918,24);
            manlo <= conv_std_logic_vector(80047690,28);
            exponent <= conv_std_logic_vector(1670,11);
      WHEN "0111000010" =>
            manhi <= conv_std_logic_vector(2666065,24);
            manlo <= conv_std_logic_vector(164712049,28);
            exponent <= conv_std_logic_vector(1672,11);
      WHEN "0111000011" =>
            manhi <= conv_std_logic_vector(9648943,24);
            manlo <= conv_std_logic_vector(147084012,28);
            exponent <= conv_std_logic_vector(1673,11);
      WHEN "0111000100" =>
            manhi <= conv_std_logic_vector(1181221,24);
            manlo <= conv_std_logic_vector(86912647,28);
            exponent <= conv_std_logic_vector(1675,11);
      WHEN "0111000101" =>
            manhi <= conv_std_logic_vector(7630830,24);
            manlo <= conv_std_logic_vector(247596521,28);
            exponent <= conv_std_logic_vector(1676,11);
      WHEN "0111000110" =>
            manhi <= conv_std_logic_vector(16396759,24);
            manlo <= conv_std_logic_vector(56002502,28);
            exponent <= conv_std_logic_vector(1677,11);
      WHEN "0111000111" =>
            manhi <= conv_std_logic_vector(5766837,24);
            manlo <= conv_std_logic_vector(133369322,28);
            exponent <= conv_std_logic_vector(1679,11);
      WHEN "0111001000" =>
            manhi <= conv_std_logic_vector(13863329,24);
            manlo <= conv_std_logic_vector(128884889,28);
            exponent <= conv_std_logic_vector(1680,11);
      WHEN "0111001001" =>
            manhi <= conv_std_logic_vector(4045193,24);
            manlo <= conv_std_logic_vector(133729186,28);
            exponent <= conv_std_logic_vector(1682,11);
      WHEN "0111001010" =>
            manhi <= conv_std_logic_vector(11523372,24);
            manlo <= conv_std_logic_vector(183024104,28);
            exponent <= conv_std_logic_vector(1683,11);
      WHEN "0111001011" =>
            manhi <= conv_std_logic_vector(2455027,24);
            manlo <= conv_std_logic_vector(264977965,28);
            exponent <= conv_std_logic_vector(1685,11);
      WHEN "0111001100" =>
            manhi <= conv_std_logic_vector(9362113,24);
            manlo <= conv_std_logic_vector(181285013,28);
            exponent <= conv_std_logic_vector(1686,11);
      WHEN "0111001101" =>
            manhi <= conv_std_logic_vector(986300,24);
            manlo <= conv_std_logic_vector(58020653,28);
            exponent <= conv_std_logic_vector(1688,11);
      WHEN "0111001110" =>
            manhi <= conv_std_logic_vector(7365905,24);
            manlo <= conv_std_logic_vector(179835810,28);
            exponent <= conv_std_logic_vector(1689,11);
      WHEN "0111001111" =>
            manhi <= conv_std_logic_vector(16036688,24);
            manlo <= conv_std_logic_vector(123168298,28);
            exponent <= conv_std_logic_vector(1690,11);
      WHEN "0111010000" =>
            manhi <= conv_std_logic_vector(5522144,24);
            manlo <= conv_std_logic_vector(14176725,28);
            exponent <= conv_std_logic_vector(1692,11);
      WHEN "0111010001" =>
            manhi <= conv_std_logic_vector(13530756,24);
            manlo <= conv_std_logic_vector(163453775,28);
            exponent <= conv_std_logic_vector(1693,11);
      WHEN "0111010010" =>
            manhi <= conv_std_logic_vector(3819186,24);
            manlo <= conv_std_logic_vector(214764608,28);
            exponent <= conv_std_logic_vector(1695,11);
      WHEN "0111010011" =>
            manhi <= conv_std_logic_vector(11216197,24);
            manlo <= conv_std_logic_vector(196364225,28);
            exponent <= conv_std_logic_vector(1696,11);
      WHEN "0111010100" =>
            manhi <= conv_std_logic_vector(2246280,24);
            manlo <= conv_std_logic_vector(259235483,28);
            exponent <= conv_std_logic_vector(1698,11);
      WHEN "0111010101" =>
            manhi <= conv_std_logic_vector(9078397,24);
            manlo <= conv_std_logic_vector(15526664,28);
            exponent <= conv_std_logic_vector(1699,11);
      WHEN "0111010110" =>
            manhi <= conv_std_logic_vector(793494,24);
            manlo <= conv_std_logic_vector(210641201,28);
            exponent <= conv_std_logic_vector(1701,11);
      WHEN "0111010111" =>
            manhi <= conv_std_logic_vector(7103855,24);
            manlo <= conv_std_logic_vector(246847656,28);
            exponent <= conv_std_logic_vector(1702,11);
      WHEN "0111011000" =>
            manhi <= conv_std_logic_vector(15680525,24);
            manlo <= conv_std_logic_vector(247378795,28);
            exponent <= conv_std_logic_vector(1703,11);
      WHEN "0111011001" =>
            manhi <= conv_std_logic_vector(5280106,24);
            manlo <= conv_std_logic_vector(138122391,28);
            exponent <= conv_std_logic_vector(1705,11);
      WHEN "0111011010" =>
            manhi <= conv_std_logic_vector(13201793,24);
            manlo <= conv_std_logic_vector(130963079,28);
            exponent <= conv_std_logic_vector(1706,11);
      WHEN "0111011011" =>
            manhi <= conv_std_logic_vector(3595633,24);
            manlo <= conv_std_logic_vector(48727293,28);
            exponent <= conv_std_logic_vector(1708,11);
      WHEN "0111011100" =>
            manhi <= conv_std_logic_vector(10912356,24);
            manlo <= conv_std_logic_vector(231400966,28);
            exponent <= conv_std_logic_vector(1709,11);
      WHEN "0111011101" =>
            manhi <= conv_std_logic_vector(2039799,24);
            manlo <= conv_std_logic_vector(184459756,28);
            exponent <= conv_std_logic_vector(1711,11);
      WHEN "0111011110" =>
            manhi <= conv_std_logic_vector(8797759,24);
            manlo <= conv_std_logic_vector(242699544,28);
            exponent <= conv_std_logic_vector(1712,11);
      WHEN "0111011111" =>
            manhi <= conv_std_logic_vector(602782,24);
            manlo <= conv_std_logic_vector(17680793,28);
            exponent <= conv_std_logic_vector(1714,11);
      WHEN "0111100000" =>
            manhi <= conv_std_logic_vector(6844650,24);
            manlo <= conv_std_logic_vector(123627565,28);
            exponent <= conv_std_logic_vector(1715,11);
      WHEN "0111100001" =>
            manhi <= conv_std_logic_vector(15328229,24);
            manlo <= conv_std_logic_vector(47512453,28);
            exponent <= conv_std_logic_vector(1716,11);
      WHEN "0111100010" =>
            manhi <= conv_std_logic_vector(5040696,24);
            manlo <= conv_std_logic_vector(14711664,28);
            exponent <= conv_std_logic_vector(1718,11);
      WHEN "0111100011" =>
            manhi <= conv_std_logic_vector(12876400,24);
            manlo <= conv_std_logic_vector(251456186,28);
            exponent <= conv_std_logic_vector(1719,11);
      WHEN "0111100100" =>
            manhi <= conv_std_logic_vector(3374506,24);
            manlo <= conv_std_logic_vector(4512772,28);
            exponent <= conv_std_logic_vector(1721,11);
      WHEN "0111100101" =>
            manhi <= conv_std_logic_vector(10611813,24);
            manlo <= conv_std_logic_vector(237626642,28);
            exponent <= conv_std_logic_vector(1722,11);
      WHEN "0111100110" =>
            manhi <= conv_std_logic_vector(1835559,24);
            manlo <= conv_std_logic_vector(150064655,28);
            exponent <= conv_std_logic_vector(1724,11);
      WHEN "0111100111" =>
            manhi <= conv_std_logic_vector(8520168,24);
            manlo <= conv_std_logic_vector(211971382,28);
            exponent <= conv_std_logic_vector(1725,11);
      WHEN "0111101000" =>
            manhi <= conv_std_logic_vector(414139,24);
            manlo <= conv_std_logic_vector(92694471,28);
            exponent <= conv_std_logic_vector(1727,11);
      WHEN "0111101001" =>
            manhi <= conv_std_logic_vector(6588258,24);
            manlo <= conv_std_logic_vector(112977613,28);
            exponent <= conv_std_logic_vector(1728,11);
      WHEN "0111101010" =>
            manhi <= conv_std_logic_vector(14979756,24);
            manlo <= conv_std_logic_vector(71348470,28);
            exponent <= conv_std_logic_vector(1729,11);
      WHEN "0111101011" =>
            manhi <= conv_std_logic_vector(4803884,24);
            manlo <= conv_std_logic_vector(42747344,28);
            exponent <= conv_std_logic_vector(1731,11);
      WHEN "0111101100" =>
            manhi <= conv_std_logic_vector(12554540,24);
            manlo <= conv_std_logic_vector(53825836,28);
            exponent <= conv_std_logic_vector(1732,11);
      WHEN "0111101101" =>
            manhi <= conv_std_logic_vector(3155778,24);
            manlo <= conv_std_logic_vector(260157975,28);
            exponent <= conv_std_logic_vector(1734,11);
      WHEN "0111101110" =>
            manhi <= conv_std_logic_vector(10314533,24);
            manlo <= conv_std_logic_vector(1535990,28);
            exponent <= conv_std_logic_vector(1735,11);
      WHEN "0111101111" =>
            manhi <= conv_std_logic_vector(1633536,24);
            manlo <= conv_std_logic_vector(68681060,28);
            exponent <= conv_std_logic_vector(1737,11);
      WHEN "0111110000" =>
            manhi <= conv_std_logic_vector(8245590,24);
            manlo <= conv_std_logic_vector(175202070,28);
            exponent <= conv_std_logic_vector(1738,11);
      WHEN "0111110001" =>
            manhi <= conv_std_logic_vector(227544,24);
            manlo <= conv_std_logic_vector(41675965,28);
            exponent <= conv_std_logic_vector(1740,11);
      WHEN "0111110010" =>
            manhi <= conv_std_logic_vector(6334649,24);
            manlo <= conv_std_logic_vector(70777607,28);
            exponent <= conv_std_logic_vector(1741,11);
      WHEN "0111110011" =>
            manhi <= conv_std_logic_vector(14635065,24);
            manlo <= conv_std_logic_vector(183612561,28);
            exponent <= conv_std_logic_vector(1742,11);
      WHEN "0111110100" =>
            manhi <= conv_std_logic_vector(4569642,24);
            manlo <= conv_std_logic_vector(167240760,28);
            exponent <= conv_std_logic_vector(1744,11);
      WHEN "0111110101" =>
            manhi <= conv_std_logic_vector(12236172,24);
            manlo <= conv_std_logic_vector(253623266,28);
            exponent <= conv_std_logic_vector(1745,11);
      WHEN "0111110110" =>
            manhi <= conv_std_logic_vector(2939425,24);
            manlo <= conv_std_logic_vector(265128301,28);
            exponent <= conv_std_logic_vector(1747,11);
      WHEN "0111110111" =>
            manhi <= conv_std_logic_vector(10020478,24);
            manlo <= conv_std_logic_vector(219223569,28);
            exponent <= conv_std_logic_vector(1748,11);
      WHEN "0111111000" =>
            manhi <= conv_std_logic_vector(1433705,24);
            manlo <= conv_std_logic_vector(192250058,28);
            exponent <= conv_std_logic_vector(1750,11);
      WHEN "0111111001" =>
            manhi <= conv_std_logic_vector(7973992,24);
            manlo <= conv_std_logic_vector(212144821,28);
            exponent <= conv_std_logic_vector(1751,11);
      WHEN "0111111010" =>
            manhi <= conv_std_logic_vector(42974,24);
            manlo <= conv_std_logic_vector(72952107,28);
            exponent <= conv_std_logic_vector(1753,11);
      WHEN "0111111011" =>
            manhi <= conv_std_logic_vector(6083792,24);
            manlo <= conv_std_logic_vector(210315148,28);
            exponent <= conv_std_logic_vector(1754,11);
      WHEN "0111111100" =>
            manhi <= conv_std_logic_vector(14294116,24);
            manlo <= conv_std_logic_vector(101520926,28);
            exponent <= conv_std_logic_vector(1755,11);
      WHEN "0111111101" =>
            manhi <= conv_std_logic_vector(4337943,24);
            manlo <= conv_std_logic_vector(146945490,28);
            exponent <= conv_std_logic_vector(1757,11);
      WHEN "0111111110" =>
            manhi <= conv_std_logic_vector(11921261,24);
            manlo <= conv_std_logic_vector(67478049,28);
            exponent <= conv_std_logic_vector(1758,11);
      WHEN "0111111111" =>
            manhi <= conv_std_logic_vector(2725421,24);
            manlo <= conv_std_logic_vector(81662013,28);
            exponent <= conv_std_logic_vector(1760,11);
      WHEN "1000000000" =>
            manhi <= conv_std_logic_vector(9729616,24);
            manlo <= conv_std_logic_vector(79332654,28);
            exponent <= conv_std_logic_vector(1761,11);
      WHEN "1000000001" =>
            manhi <= conv_std_logic_vector(1236044,24);
            manlo <= conv_std_logic_vector(37511845,28);
            exponent <= conv_std_logic_vector(1763,11);
      WHEN "1000000010" =>
            manhi <= conv_std_logic_vector(7705342,24);
            manlo <= conv_std_logic_vector(229400607,28);
            exponent <= conv_std_logic_vector(1764,11);
      WHEN "1000000011" =>
            manhi <= conv_std_logic_vector(16498031,24);
            manlo <= conv_std_logic_vector(113896411,28);
            exponent <= conv_std_logic_vector(1765,11);
      WHEN "1000000100" =>
            manhi <= conv_std_logic_vector(5835659,24);
            manlo <= conv_std_logic_vector(27578100,28);
            exponent <= conv_std_logic_vector(1767,11);
      WHEN "1000000101" =>
            manhi <= conv_std_logic_vector(13956867,24);
            manlo <= conv_std_logic_vector(198774093,28);
            exponent <= conv_std_logic_vector(1768,11);
      WHEN "1000000110" =>
            manhi <= conv_std_logic_vector(4108759,24);
            manlo <= conv_std_logic_vector(90336304,28);
            exponent <= conv_std_logic_vector(1770,11);
      WHEN "1000000111" =>
            manhi <= conv_std_logic_vector(11609767,24);
            manlo <= conv_std_logic_vector(164675818,28);
            exponent <= conv_std_logic_vector(1771,11);
      WHEN "1000001000" =>
            manhi <= conv_std_logic_vector(2513739,24);
            manlo <= conv_std_logic_vector(115510945,28);
            exponent <= conv_std_logic_vector(1773,11);
      WHEN "1000001001" =>
            manhi <= conv_std_logic_vector(9441910,24);
            manlo <= conv_std_logic_vector(214725537,28);
            exponent <= conv_std_logic_vector(1774,11);
      WHEN "1000001010" =>
            manhi <= conv_std_logic_vector(1040527,24);
            manlo <= conv_std_logic_vector(264292986,28);
            exponent <= conv_std_logic_vector(1776,11);
      WHEN "1000001011" =>
            manhi <= conv_std_logic_vector(7439608,24);
            manlo <= conv_std_logic_vector(227819416,28);
            exponent <= conv_std_logic_vector(1777,11);
      WHEN "1000001100" =>
            manhi <= conv_std_logic_vector(16136861,24);
            manlo <= conv_std_logic_vector(124712281,28);
            exponent <= conv_std_logic_vector(1778,11);
      WHEN "1000001101" =>
            manhi <= conv_std_logic_vector(5590218,24);
            manlo <= conv_std_logic_vector(179347558,28);
            exponent <= conv_std_logic_vector(1780,11);
      WHEN "1000001110" =>
            manhi <= conv_std_logic_vector(13623279,24);
            manlo <= conv_std_logic_vector(162081347,28);
            exponent <= conv_std_logic_vector(1781,11);
      WHEN "1000001111" =>
            manhi <= conv_std_logic_vector(3882062,24);
            manlo <= conv_std_logic_vector(186291443,28);
            exponent <= conv_std_logic_vector(1783,11);
      WHEN "1000010000" =>
            manhi <= conv_std_logic_vector(11301654,24);
            manlo <= conv_std_logic_vector(250040022,28);
            exponent <= conv_std_logic_vector(1784,11);
      WHEN "1000010001" =>
            manhi <= conv_std_logic_vector(2304355,24);
            manlo <= conv_std_logic_vector(41383777,28);
            exponent <= conv_std_logic_vector(1786,11);
      WHEN "1000010010" =>
            manhi <= conv_std_logic_vector(9157328,24);
            manlo <= conv_std_logic_vector(17021400,28);
            exponent <= conv_std_logic_vector(1787,11);
      WHEN "1000010011" =>
            manhi <= conv_std_logic_vector(847133,24);
            manlo <= conv_std_logic_vector(258834653,28);
            exponent <= conv_std_logic_vector(1789,11);
      WHEN "1000010100" =>
            manhi <= conv_std_logic_vector(7176759,24);
            manlo <= conv_std_logic_vector(33041815,28);
            exponent <= conv_std_logic_vector(1790,11);
      WHEN "1000010101" =>
            manhi <= conv_std_logic_vector(15779611,24);
            manlo <= conv_std_logic_vector(174007449,28);
            exponent <= conv_std_logic_vector(1791,11);
      WHEN "1000010110" =>
            manhi <= conv_std_logic_vector(5347442,24);
            manlo <= conv_std_logic_vector(66333886,28);
            exponent <= conv_std_logic_vector(1793,11);
      WHEN "1000010111" =>
            manhi <= conv_std_logic_vector(13293312,24);
            manlo <= conv_std_logic_vector(63618366,28);
            exponent <= conv_std_logic_vector(1794,11);
      WHEN "1000011000" =>
            manhi <= conv_std_logic_vector(3657826,24);
            manlo <= conv_std_logic_vector(166348998,28);
            exponent <= conv_std_logic_vector(1796,11);
      WHEN "1000011001" =>
            manhi <= conv_std_logic_vector(10996886,24);
            manlo <= conv_std_logic_vector(136487624,28);
            exponent <= conv_std_logic_vector(1797,11);
      WHEN "1000011010" =>
            manhi <= conv_std_logic_vector(2097243,24);
            manlo <= conv_std_logic_vector(144317262,28);
            exponent <= conv_std_logic_vector(1799,11);
      WHEN "1000011011" =>
            manhi <= conv_std_logic_vector(8875834,24);
            manlo <= conv_std_logic_vector(51419886,28);
            exponent <= conv_std_logic_vector(1800,11);
      WHEN "1000011100" =>
            manhi <= conv_std_logic_vector(655839,24);
            manlo <= conv_std_logic_vector(12096311,28);
            exponent <= conv_std_logic_vector(1802,11);
      WHEN "1000011101" =>
            manhi <= conv_std_logic_vector(6916762,24);
            manlo <= conv_std_logic_vector(99793437,28);
            exponent <= conv_std_logic_vector(1803,11);
      WHEN "1000011110" =>
            manhi <= conv_std_logic_vector(15426239,24);
            manlo <= conv_std_logic_vector(114334116,28);
            exponent <= conv_std_logic_vector(1804,11);
      WHEN "1000011111" =>
            manhi <= conv_std_logic_vector(5107300,24);
            manlo <= conv_std_logic_vector(248161218,28);
            exponent <= conv_std_logic_vector(1806,11);
      WHEN "1000100000" =>
            manhi <= conv_std_logic_vector(12966926,24);
            manlo <= conv_std_logic_vector(91321506,28);
            exponent <= conv_std_logic_vector(1807,11);
      WHEN "1000100001" =>
            manhi <= conv_std_logic_vector(3436024,24);
            manlo <= conv_std_logic_vector(109150055,28);
            exponent <= conv_std_logic_vector(1809,11);
      WHEN "1000100010" =>
            manhi <= conv_std_logic_vector(10695426,24);
            manlo <= conv_std_logic_vector(12291314,28);
            exponent <= conv_std_logic_vector(1810,11);
      WHEN "1000100011" =>
            manhi <= conv_std_logic_vector(1892379,24);
            manlo <= conv_std_logic_vector(245137096,28);
            exponent <= conv_std_logic_vector(1812,11);
      WHEN "1000100100" =>
            manhi <= conv_std_logic_vector(8597395,24);
            manlo <= conv_std_logic_vector(176569250,28);
            exponent <= conv_std_logic_vector(1813,11);
      WHEN "1000100101" =>
            manhi <= conv_std_logic_vector(466620,24);
            manlo <= conv_std_logic_vector(119019308,28);
            exponent <= conv_std_logic_vector(1815,11);
      WHEN "1000100110" =>
            manhi <= conv_std_logic_vector(6659587,24);
            manlo <= conv_std_logic_vector(168706814,28);
            exponent <= conv_std_logic_vector(1816,11);
      WHEN "1000100111" =>
            manhi <= conv_std_logic_vector(15076702,24);
            manlo <= conv_std_logic_vector(190651618,28);
            exponent <= conv_std_logic_vector(1817,11);
      WHEN "1000101000" =>
            manhi <= conv_std_logic_vector(4869766,24);
            manlo <= conv_std_logic_vector(26523901,28);
            exponent <= conv_std_logic_vector(1819,11);
      WHEN "1000101001" =>
            manhi <= conv_std_logic_vector(12644083,24);
            manlo <= conv_std_logic_vector(10760420,28);
            exponent <= conv_std_logic_vector(1820,11);
      WHEN "1000101010" =>
            manhi <= conv_std_logic_vector(3216629,24);
            manlo <= conv_std_logic_vector(171149379,28);
            exponent <= conv_std_logic_vector(1822,11);
      WHEN "1000101011" =>
            manhi <= conv_std_logic_vector(10397237,24);
            manlo <= conv_std_logic_vector(171483537,28);
            exponent <= conv_std_logic_vector(1823,11);
      WHEN "1000101100" =>
            manhi <= conv_std_logic_vector(1689739,24);
            manlo <= conv_std_logic_vector(236540182,28);
            exponent <= conv_std_logic_vector(1825,11);
      WHEN "1000101101" =>
            manhi <= conv_std_logic_vector(8321979,24);
            manlo <= conv_std_logic_vector(80365386,28);
            exponent <= conv_std_logic_vector(1826,11);
      WHEN "1000101110" =>
            manhi <= conv_std_logic_vector(279455,24);
            manlo <= conv_std_logic_vector(167185714,28);
            exponent <= conv_std_logic_vector(1828,11);
      WHEN "1000101111" =>
            manhi <= conv_std_logic_vector(6405204,24);
            manlo <= conv_std_logic_vector(70637708,28);
            exponent <= conv_std_logic_vector(1829,11);
      WHEN "1000110000" =>
            manhi <= conv_std_logic_vector(14730959,24);
            manlo <= conv_std_logic_vector(233674466,28);
            exponent <= conv_std_logic_vector(1830,11);
      WHEN "1000110001" =>
            manhi <= conv_std_logic_vector(4634809,24);
            manlo <= conv_std_logic_vector(128626627,28);
            exponent <= conv_std_logic_vector(1832,11);
      WHEN "1000110010" =>
            manhi <= conv_std_logic_vector(12324743,24);
            manlo <= conv_std_logic_vector(237637056,28);
            exponent <= conv_std_logic_vector(1833,11);
      WHEN "1000110011" =>
            manhi <= conv_std_logic_vector(2999616,24);
            manlo <= conv_std_logic_vector(48899908,28);
            exponent <= conv_std_logic_vector(1835,11);
      WHEN "1000110100" =>
            manhi <= conv_std_logic_vector(10102285,24);
            manlo <= conv_std_logic_vector(207402206,28);
            exponent <= conv_std_logic_vector(1836,11);
      WHEN "1000110101" =>
            manhi <= conv_std_logic_vector(1489299,24);
            manlo <= conv_std_logic_vector(82314533,28);
            exponent <= conv_std_logic_vector(1838,11);
      WHEN "1000110110" =>
            manhi <= conv_std_logic_vector(8049552,24);
            manlo <= conv_std_logic_vector(84197942,28);
            exponent <= conv_std_logic_vector(1839,11);
      WHEN "1000110111" =>
            manhi <= conv_std_logic_vector(94322,24);
            manlo <= conv_std_logic_vector(78275083,28);
            exponent <= conv_std_logic_vector(1841,11);
      WHEN "1000111000" =>
            manhi <= conv_std_logic_vector(6153581,24);
            manlo <= conv_std_logic_vector(262556746,28);
            exponent <= conv_std_logic_vector(1842,11);
      WHEN "1000111001" =>
            manhi <= conv_std_logic_vector(14388969,24);
            manlo <= conv_std_logic_vector(195412276,28);
            exponent <= conv_std_logic_vector(1843,11);
      WHEN "1000111010" =>
            manhi <= conv_std_logic_vector(4402403,24);
            manlo <= conv_std_logic_vector(21925377,28);
            exponent <= conv_std_logic_vector(1845,11);
      WHEN "1000111011" =>
            manhi <= conv_std_logic_vector(12008870,24);
            manlo <= conv_std_logic_vector(225943576,28);
            exponent <= conv_std_logic_vector(1846,11);
      WHEN "1000111100" =>
            manhi <= conv_std_logic_vector(2784958,24);
            manlo <= conv_std_logic_vector(51959162,28);
            exponent <= conv_std_logic_vector(1848,11);
      WHEN "1000111101" =>
            manhi <= conv_std_logic_vector(9810535,24);
            manlo <= conv_std_logic_vector(85297068,28);
            exponent <= conv_std_logic_vector(1849,11);
      WHEN "1000111110" =>
            manhi <= conv_std_logic_vector(1291034,24);
            manlo <= conv_std_logic_vector(85003113,28);
            exponent <= conv_std_logic_vector(1851,11);
      WHEN "1000111111" =>
            manhi <= conv_std_logic_vector(7780082,24);
            manlo <= conv_std_logic_vector(68159752,28);
            exponent <= conv_std_logic_vector(1852,11);
      WHEN "1001000000" =>
            manhi <= conv_std_logic_vector(16599612,24);
            manlo <= conv_std_logic_vector(214703512,28);
            exponent <= conv_std_logic_vector(1853,11);
      WHEN "1001000001" =>
            manhi <= conv_std_logic_vector(5904690,24);
            manlo <= conv_std_logic_vector(215968023,28);
            exponent <= conv_std_logic_vector(1855,11);
      WHEN "1001000010" =>
            manhi <= conv_std_logic_vector(14050691,24);
            manlo <= conv_std_logic_vector(147853227,28);
            exponent <= conv_std_logic_vector(1856,11);
      WHEN "1001000011" =>
            manhi <= conv_std_logic_vector(4172519,24);
            manlo <= conv_std_logic_vector(60716388,28);
            exponent <= conv_std_logic_vector(1858,11);
      WHEN "1001000100" =>
            manhi <= conv_std_logic_vector(11696426,24);
            manlo <= conv_std_logic_vector(77359100,28);
            exponent <= conv_std_logic_vector(1859,11);
      WHEN "1001000101" =>
            manhi <= conv_std_logic_vector(2572630,24);
            manlo <= conv_std_logic_vector(28321055,28);
            exponent <= conv_std_logic_vector(1861,11);
      WHEN "1001000110" =>
            manhi <= conv_std_logic_vector(9521951,24);
            manlo <= conv_std_logic_vector(141206574,28);
            exponent <= conv_std_logic_vector(1862,11);
      WHEN "1001000111" =>
            manhi <= conv_std_logic_vector(1094921,24);
            manlo <= conv_std_logic_vector(79834212,28);
            exponent <= conv_std_logic_vector(1864,11);
      WHEN "1001001000" =>
            manhi <= conv_std_logic_vector(7513537,24);
            manlo <= conv_std_logic_vector(6880382,28);
            exponent <= conv_std_logic_vector(1865,11);
      WHEN "1001001001" =>
            manhi <= conv_std_logic_vector(16237340,24);
            manlo <= conv_std_logic_vector(73707069,28);
            exponent <= conv_std_logic_vector(1866,11);
      WHEN "1001001010" =>
            manhi <= conv_std_logic_vector(5658501,24);
            manlo <= conv_std_logic_vector(26563701,28);
            exponent <= conv_std_logic_vector(1868,11);
      WHEN "1001001011" =>
            manhi <= conv_std_logic_vector(13716085,24);
            manlo <= conv_std_logic_vector(13226359,28);
            exponent <= conv_std_logic_vector(1869,11);
      WHEN "1001001100" =>
            manhi <= conv_std_logic_vector(3945130,24);
            manlo <= conv_std_logic_vector(143073903,28);
            exponent <= conv_std_logic_vector(1871,11);
      WHEN "1001001101" =>
            manhi <= conv_std_logic_vector(11387373,24);
            manlo <= conv_std_logic_vector(3175990,28);
            exponent <= conv_std_logic_vector(1872,11);
      WHEN "1001001110" =>
            manhi <= conv_std_logic_vector(2362606,24);
            manlo <= conv_std_logic_vector(168904878,28);
            exponent <= conv_std_logic_vector(1874,11);
      WHEN "1001001111" =>
            manhi <= conv_std_logic_vector(9236500,24);
            manlo <= conv_std_logic_vector(7105104,28);
            exponent <= conv_std_logic_vector(1875,11);
      WHEN "1001010000" =>
            manhi <= conv_std_logic_vector(900936,24);
            manlo <= conv_std_logic_vector(239272854,28);
            exponent <= conv_std_logic_vector(1877,11);
      WHEN "1001010001" =>
            manhi <= conv_std_logic_vector(7249884,24);
            manlo <= conv_std_logic_vector(236935482,28);
            exponent <= conv_std_logic_vector(1878,11);
      WHEN "1001010010" =>
            manhi <= conv_std_logic_vector(15878999,24);
            manlo <= conv_std_logic_vector(230836932,28);
            exponent <= conv_std_logic_vector(1879,11);
      WHEN "1001010011" =>
            manhi <= conv_std_logic_vector(5414983,24);
            manlo <= conv_std_logic_vector(144840810,28);
            exponent <= conv_std_logic_vector(1881,11);
      WHEN "1001010100" =>
            manhi <= conv_std_logic_vector(13385110,24);
            manlo <= conv_std_logic_vector(99584369,28);
            exponent <= conv_std_logic_vector(1882,11);
      WHEN "1001010101" =>
            manhi <= conv_std_logic_vector(3720209,24);
            manlo <= conv_std_logic_vector(246845719,28);
            exponent <= conv_std_logic_vector(1884,11);
      WHEN "1001010110" =>
            manhi <= conv_std_logic_vector(11081674,24);
            manlo <= conv_std_logic_vector(54674652,28);
            exponent <= conv_std_logic_vector(1885,11);
      WHEN "1001010111" =>
            manhi <= conv_std_logic_vector(2154862,24);
            manlo <= conv_std_logic_vector(201440422,28);
            exponent <= conv_std_logic_vector(1887,11);
      WHEN "1001011000" =>
            manhi <= conv_std_logic_vector(8954146,24);
            manlo <= conv_std_logic_vector(220416825,28);
            exponent <= conv_std_logic_vector(1888,11);
      WHEN "1001011001" =>
            manhi <= conv_std_logic_vector(709057,24);
            manlo <= conv_std_logic_vector(266967657,28);
            exponent <= conv_std_logic_vector(1890,11);
      WHEN "1001011010" =>
            manhi <= conv_std_logic_vector(6989094,24);
            manlo <= conv_std_logic_vector(113654547,28);
            exponent <= conv_std_logic_vector(1891,11);
      WHEN "1001011011" =>
            manhi <= conv_std_logic_vector(15524548,24);
            manlo <= conv_std_logic_vector(235342013,28);
            exponent <= conv_std_logic_vector(1892,11);
      WHEN "1001011100" =>
            manhi <= conv_std_logic_vector(5174109,24);
            manlo <= conv_std_logic_vector(32986511,28);
            exponent <= conv_std_logic_vector(1894,11);
      WHEN "1001011101" =>
            manhi <= conv_std_logic_vector(13057728,24);
            manlo <= conv_std_logic_vector(25787653,28);
            exponent <= conv_std_logic_vector(1895,11);
      WHEN "1001011110" =>
            manhi <= conv_std_logic_vector(3497730,24);
            manlo <= conv_std_logic_vector(160351868,28);
            exponent <= conv_std_logic_vector(1897,11);
      WHEN "1001011111" =>
            manhi <= conv_std_logic_vector(10779293,24);
            manlo <= conv_std_logic_vector(121946709,28);
            exponent <= conv_std_logic_vector(1898,11);
      WHEN "1001100000" =>
            manhi <= conv_std_logic_vector(1949373,24);
            manlo <= conv_std_logic_vector(194974600,28);
            exponent <= conv_std_logic_vector(1900,11);
      WHEN "1001100001" =>
            manhi <= conv_std_logic_vector(8674858,24);
            manlo <= conv_std_logic_vector(75445083,28);
            exponent <= conv_std_logic_vector(1901,11);
      WHEN "1001100010" =>
            manhi <= conv_std_logic_vector(519261,24);
            manlo <= conv_std_logic_vector(202318540,28);
            exponent <= conv_std_logic_vector(1903,11);
      WHEN "1001100011" =>
            manhi <= conv_std_logic_vector(6731134,24);
            manlo <= conv_std_logic_vector(157600610,28);
            exponent <= conv_std_logic_vector(1904,11);
      WHEN "1001100100" =>
            manhi <= conv_std_logic_vector(15173945,24);
            manlo <= conv_std_logic_vector(29256816,28);
            exponent <= conv_std_logic_vector(1905,11);
      WHEN "1001100101" =>
            manhi <= conv_std_logic_vector(4935849,24);
            manlo <= conv_std_logic_vector(42999013,28);
            exponent <= conv_std_logic_vector(1907,11);
      WHEN "1001100110" =>
            manhi <= conv_std_logic_vector(12733899,24);
            manlo <= conv_std_logic_vector(62421287,28);
            exponent <= conv_std_logic_vector(1908,11);
      WHEN "1001100111" =>
            manhi <= conv_std_logic_vector(3277666,24);
            manlo <= conv_std_logic_vector(18399062,28);
            exponent <= conv_std_logic_vector(1910,11);
      WHEN "1001101000" =>
            manhi <= conv_std_logic_vector(10480194,24);
            manlo <= conv_std_logic_vector(201166396,28);
            exponent <= conv_std_logic_vector(1911,11);
      WHEN "1001101001" =>
            manhi <= conv_std_logic_vector(1746115,24);
            manlo <= conv_std_logic_vector(22209480,28);
            exponent <= conv_std_logic_vector(1913,11);
      WHEN "1001101010" =>
            manhi <= conv_std_logic_vector(8398601,24);
            manlo <= conv_std_logic_vector(38216343,28);
            exponent <= conv_std_logic_vector(1914,11);
      WHEN "1001101011" =>
            manhi <= conv_std_logic_vector(331525,24);
            manlo <= conv_std_logic_vector(151310615,28);
            exponent <= conv_std_logic_vector(1916,11);
      WHEN "1001101100" =>
            manhi <= conv_std_logic_vector(6475974,24);
            manlo <= conv_std_logic_vector(174528998,28);
            exponent <= conv_std_logic_vector(1917,11);
      WHEN "1001101101" =>
            manhi <= conv_std_logic_vector(14827146,24);
            manlo <= conv_std_logic_vector(214487191,28);
            exponent <= conv_std_logic_vector(1918,11);
      WHEN "1001101110" =>
            manhi <= conv_std_logic_vector(4700175,24);
            manlo <= conv_std_logic_vector(73593076,28);
            exponent <= conv_std_logic_vector(1920,11);
      WHEN "1001101111" =>
            manhi <= conv_std_logic_vector(12413585,24);
            manlo <= conv_std_logic_vector(56806573,28);
            exponent <= conv_std_logic_vector(1921,11);
      WHEN "1001110000" =>
            manhi <= conv_std_logic_vector(3059990,24);
            manlo <= conv_std_logic_vector(32998071,28);
            exponent <= conv_std_logic_vector(1923,11);
      WHEN "1001110001" =>
            manhi <= conv_std_logic_vector(10184342,24);
            manlo <= conv_std_logic_vector(125003687,28);
            exponent <= conv_std_logic_vector(1924,11);
      WHEN "1001110010" =>
            manhi <= conv_std_logic_vector(1545062,24);
            manlo <= conv_std_logic_vector(164026180,28);
            exponent <= conv_std_logic_vector(1926,11);
      WHEN "1001110011" =>
            manhi <= conv_std_logic_vector(8125342,24);
            manlo <= conv_std_logic_vector(134803968,28);
            exponent <= conv_std_logic_vector(1927,11);
      WHEN "1001110100" =>
            manhi <= conv_std_logic_vector(145827,24);
            manlo <= conv_std_logic_vector(17356019,28);
            exponent <= conv_std_logic_vector(1929,11);
      WHEN "1001110101" =>
            manhi <= conv_std_logic_vector(6223584,24);
            manlo <= conv_std_logic_vector(59711433,28);
            exponent <= conv_std_logic_vector(1930,11);
      WHEN "1001110110" =>
            manhi <= conv_std_logic_vector(14484112,24);
            manlo <= conv_std_logic_vector(172427100,28);
            exponent <= conv_std_logic_vector(1931,11);
      WHEN "1001110111" =>
            manhi <= conv_std_logic_vector(4467059,24);
            manlo <= conv_std_logic_vector(106163660,28);
            exponent <= conv_std_logic_vector(1933,11);
      WHEN "1001111000" =>
            manhi <= conv_std_logic_vector(12096747,24);
            manlo <= conv_std_logic_vector(237074316,28);
            exponent <= conv_std_logic_vector(1934,11);
      WHEN "1001111001" =>
            manhi <= conv_std_logic_vector(2844676,24);
            manlo <= conv_std_logic_vector(224090291,28);
            exponent <= conv_std_logic_vector(1936,11);
      WHEN "1001111010" =>
            manhi <= conv_std_logic_vector(9891701,24);
            manlo <= conv_std_logic_vector(98356275,28);
            exponent <= conv_std_logic_vector(1937,11);
      WHEN "1001111011" =>
            manhi <= conv_std_logic_vector(1346192,24);
            manlo <= conv_std_logic_vector(98098154,28);
            exponent <= conv_std_logic_vector(1939,11);
      WHEN "1001111100" =>
            manhi <= conv_std_logic_vector(7855049,24);
            manlo <= conv_std_logic_vector(218711727,28);
            exponent <= conv_std_logic_vector(1940,11);
      WHEN "1001111101" =>
            manhi <= conv_std_logic_vector(16701504,24);
            manlo <= conv_std_logic_vector(74899902,28);
            exponent <= conv_std_logic_vector(1941,11);
      WHEN "1001111110" =>
            manhi <= conv_std_logic_vector(5973933,24);
            manlo <= conv_std_logic_vector(65399866,28);
            exponent <= conv_std_logic_vector(1943,11);
      WHEN "1001111111" =>
            manhi <= conv_std_logic_vector(14144801,24);
            manlo <= conv_std_logic_vector(210121699,28);
            exponent <= conv_std_logic_vector(1944,11);
      WHEN "1010000000" =>
            manhi <= conv_std_logic_vector(4236473,24);
            manlo <= conv_std_logic_vector(203888522,28);
            exponent <= conv_std_logic_vector(1946,11);
      WHEN "1010000001" =>
            manhi <= conv_std_logic_vector(11783349,24);
            manlo <= conv_std_logic_vector(137203293,28);
            exponent <= conv_std_logic_vector(1947,11);
      WHEN "1010000010" =>
            manhi <= conv_std_logic_vector(2631700,24);
            manlo <= conv_std_logic_vector(150283410,28);
            exponent <= conv_std_logic_vector(1949,11);
      WHEN "1010000011" =>
            manhi <= conv_std_logic_vector(9602236,24);
            manlo <= conv_std_logic_vector(160352104,28);
            exponent <= conv_std_logic_vector(1950,11);
      WHEN "1010000100" =>
            manhi <= conv_std_logic_vector(1149480,24);
            manlo <= conv_std_logic_vector(177173803,28);
            exponent <= conv_std_logic_vector(1952,11);
      WHEN "1010000101" =>
            manhi <= conv_std_logic_vector(7587690,24);
            manlo <= conv_std_logic_vector(238268718,28);
            exponent <= conv_std_logic_vector(1953,11);
      WHEN "1010000110" =>
            manhi <= conv_std_logic_vector(16338125,24);
            manlo <= conv_std_logic_vector(220749839,28);
            exponent <= conv_std_logic_vector(1954,11);
      WHEN "1010000111" =>
            manhi <= conv_std_logic_vector(5726991,24);
            manlo <= conv_std_logic_vector(262994505,28);
            exponent <= conv_std_logic_vector(1956,11);
      WHEN "1010001000" =>
            manhi <= conv_std_logic_vector(13809173,24);
            manlo <= conv_std_logic_vector(216783842,28);
            exponent <= conv_std_logic_vector(1957,11);
      WHEN "1010001001" =>
            manhi <= conv_std_logic_vector(4008390,24);
            manlo <= conv_std_logic_vector(242405077,28);
            exponent <= conv_std_logic_vector(1959,11);
      WHEN "1010001010" =>
            manhi <= conv_std_logic_vector(11473352,24);
            manlo <= conv_std_logic_vector(206426515,28);
            exponent <= conv_std_logic_vector(1960,11);
      WHEN "1010001011" =>
            manhi <= conv_std_logic_vector(2421035,24);
            manlo <= conv_std_logic_vector(250208807,28);
            exponent <= conv_std_logic_vector(1962,11);
      WHEN "1010001100" =>
            manhi <= conv_std_logic_vector(9315913,24);
            manlo <= conv_std_logic_vector(183235034,28);
            exponent <= conv_std_logic_vector(1963,11);
      WHEN "1010001101" =>
            manhi <= conv_std_logic_vector(954904,24);
            manlo <= conv_std_logic_vector(17706469,28);
            exponent <= conv_std_logic_vector(1965,11);
      WHEN "1010001110" =>
            manhi <= conv_std_logic_vector(7323233,24);
            manlo <= conv_std_logic_vector(235600136,28);
            exponent <= conv_std_logic_vector(1966,11);
      WHEN "1010001111" =>
            manhi <= conv_std_logic_vector(15978691,24);
            manlo <= conv_std_logic_vector(128873524,28);
            exponent <= conv_std_logic_vector(1967,11);
      WHEN "1010010000" =>
            manhi <= conv_std_logic_vector(5482731,24);
            manlo <= conv_std_logic_vector(5222268,28);
            exponent <= conv_std_logic_vector(1969,11);
      WHEN "1010010001" =>
            manhi <= conv_std_logic_vector(13477188,24);
            manlo <= conv_std_logic_vector(199372940,28);
            exponent <= conv_std_logic_vector(1970,11);
      WHEN "1010010010" =>
            manhi <= conv_std_logic_vector(3782783,24);
            manlo <= conv_std_logic_vector(177367827,28);
            exponent <= conv_std_logic_vector(1972,11);
      WHEN "1010010011" =>
            manhi <= conv_std_logic_vector(11166720,24);
            manlo <= conv_std_logic_vector(197425116,28);
            exponent <= conv_std_logic_vector(1973,11);
      WHEN "1010010100" =>
            manhi <= conv_std_logic_vector(2212657,24);
            manlo <= conv_std_logic_vector(231097832,28);
            exponent <= conv_std_logic_vector(1975,11);
      WHEN "1010010101" =>
            manhi <= conv_std_logic_vector(9032698,24);
            manlo <= conv_std_logic_vector(139698050,28);
            exponent <= conv_std_logic_vector(1976,11);
      WHEN "1010010110" =>
            manhi <= conv_std_logic_vector(762439,24);
            manlo <= conv_std_logic_vector(109718127,28);
            exponent <= conv_std_logic_vector(1978,11);
      WHEN "1010010111" =>
            manhi <= conv_std_logic_vector(7061647,24);
            manlo <= conv_std_logic_vector(77173752,28);
            exponent <= conv_std_logic_vector(1979,11);
      WHEN "1010011000" =>
            manhi <= conv_std_logic_vector(15623158,24);
            manlo <= conv_std_logic_vector(118851961,28);
            exponent <= conv_std_logic_vector(1980,11);
      WHEN "1010011001" =>
            manhi <= conv_std_logic_vector(5241121,24);
            manlo <= conv_std_logic_vector(72680114,28);
            exponent <= conv_std_logic_vector(1982,11);
      WHEN "1010011010" =>
            manhi <= conv_std_logic_vector(13148807,24);
            manlo <= conv_std_logic_vector(12881486,28);
            exponent <= conv_std_logic_vector(1983,11);
      WHEN "1010011011" =>
            manhi <= conv_std_logic_vector(3559625,24);
            manlo <= conv_std_logic_vector(43579850,28);
            exponent <= conv_std_logic_vector(1985,11);
      WHEN "1010011100" =>
            manhi <= conv_std_logic_vector(10863416,24);
            manlo <= conv_std_logic_vector(238889758,28);
            exponent <= conv_std_logic_vector(1986,11);
      WHEN "1010011101" =>
            manhi <= conv_std_logic_vector(2006541,24);
            manlo <= conv_std_logic_vector(141721451,28);
            exponent <= conv_std_logic_vector(1988,11);
      WHEN "1010011110" =>
            manhi <= conv_std_logic_vector(8752557,24);
            manlo <= conv_std_logic_vector(101792997,28);
            exponent <= conv_std_logic_vector(1989,11);
      WHEN "1010011111" =>
            manhi <= conv_std_logic_vector(572063,24);
            manlo <= conv_std_logic_vector(205445723,28);
            exponent <= conv_std_logic_vector(1991,11);
      WHEN "1010100000" =>
            manhi <= conv_std_logic_vector(6802899,24);
            manlo <= conv_std_logic_vector(258099270,28);
            exponent <= conv_std_logic_vector(1992,11);
      WHEN "1010100001" =>
            manhi <= conv_std_logic_vector(15271484,24);
            manlo <= conv_std_logic_vector(98124990,28);
            exponent <= conv_std_logic_vector(1993,11);
      WHEN "1010100010" =>
            manhi <= conv_std_logic_vector(5002133,24);
            manlo <= conv_std_logic_vector(256985826,28);
            exponent <= conv_std_logic_vector(1995,11);
      WHEN "1010100011" =>
            manhi <= conv_std_logic_vector(12823989,24);
            manlo <= conv_std_logic_vector(164377270,28);
            exponent <= conv_std_logic_vector(1996,11);
      WHEN "1010100100" =>
            manhi <= conv_std_logic_vector(3338888,24);
            manlo <= conv_std_logic_vector(222569178,28);
            exponent <= conv_std_logic_vector(1998,11);
      WHEN "1010100101" =>
            manhi <= conv_std_logic_vector(10563405,24);
            manlo <= conv_std_logic_vector(29046646,28);
            exponent <= conv_std_logic_vector(1999,11);
      WHEN "1010100110" =>
            manhi <= conv_std_logic_vector(1802662,24);
            manlo <= conv_std_logic_vector(103161316,28);
            exponent <= conv_std_logic_vector(2001,11);
      WHEN "1010100111" =>
            manhi <= conv_std_logic_vector(8475456,24);
            manlo <= conv_std_logic_vector(239852126,28);
            exponent <= conv_std_logic_vector(2002,11);
      WHEN "1010101000" =>
            manhi <= conv_std_logic_vector(383754,24);
            manlo <= conv_std_logic_vector(123914668,28);
            exponent <= conv_std_logic_vector(2004,11);
      WHEN "1010101001" =>
            manhi <= conv_std_logic_vector(6546961,24);
            manlo <= conv_std_logic_vector(22084044,28);
            exponent <= conv_std_logic_vector(2005,11);
      WHEN "1010101010" =>
            manhi <= conv_std_logic_vector(14923627,24);
            manlo <= conv_std_logic_vector(97508377,28);
            exponent <= conv_std_logic_vector(2006,11);
      WHEN "1010101011" =>
            manhi <= conv_std_logic_vector(4765740,24);
            manlo <= conv_std_logic_vector(165164368,28);
            exponent <= conv_std_logic_vector(2008,11);
      WHEN "1010101100" =>
            manhi <= conv_std_logic_vector(12502697,24);
            manlo <= conv_std_logic_vector(201140216,28);
            exponent <= conv_std_logic_vector(2009,11);
      WHEN "1010101101" =>
            manhi <= conv_std_logic_vector(3120548,24);
            manlo <= conv_std_logic_vector(99561759,28);
            exponent <= conv_std_logic_vector(2011,11);
      WHEN "1010101110" =>
            manhi <= conv_std_logic_vector(10266649,24);
            manlo <= conv_std_logic_vector(176679877,28);
            exponent <= conv_std_logic_vector(2012,11);
      WHEN "1010101111" =>
            manhi <= conv_std_logic_vector(1600996,24);
            manlo <= conv_std_logic_vector(39589446,28);
            exponent <= conv_std_logic_vector(2014,11);
      WHEN "1010110000" =>
            manhi <= conv_std_logic_vector(8201364,24);
            manlo <= conv_std_logic_vector(16114999,28);
            exponent <= conv_std_logic_vector(2015,11);
      WHEN "1010110001" =>
            manhi <= conv_std_logic_vector(197489,24);
            manlo <= conv_std_logic_vector(18649371,28);
            exponent <= conv_std_logic_vector(2017,11);
      WHEN "1010110010" =>
            manhi <= conv_std_logic_vector(6293800,24);
            manlo <= conv_std_logic_vector(44802372,28);
            exponent <= conv_std_logic_vector(2018,11);
      WHEN "1010110011" =>
            manhi <= conv_std_logic_vector(14579546,24);
            manlo <= conv_std_logic_vector(1419236,28);
            exponent <= conv_std_logic_vector(2019,11);
      WHEN "1010110100" =>
            manhi <= conv_std_logic_vector(4531913,24);
            manlo <= conv_std_logic_vector(24044223,28);
            exponent <= conv_std_logic_vector(2021,11);
      WHEN "1010110101" =>
            manhi <= conv_std_logic_vector(12184893,24);
            manlo <= conv_std_logic_vector(51602800,28);
            exponent <= conv_std_logic_vector(2022,11);
      WHEN "1010110110" =>
            manhi <= conv_std_logic_vector(2904577,24);
            manlo <= conv_std_logic_vector(210124577,28);
            exponent <= conv_std_logic_vector(2024,11);
      WHEN "1010110111" =>
            manhi <= conv_std_logic_vector(9973115,24);
            manlo <= conv_std_logic_vector(52505388,28);
            exponent <= conv_std_logic_vector(2025,11);
      WHEN "1010111000" =>
            manhi <= conv_std_logic_vector(1401518,24);
            manlo <= conv_std_logic_vector(214362802,28);
            exponent <= conv_std_logic_vector(2027,11);
      WHEN "1010111001" =>
            manhi <= conv_std_logic_vector(7930246,24);
            manlo <= conv_std_logic_vector(62721516,28);
            exponent <= conv_std_logic_vector(2028,11);
      WHEN "1010111010" =>
            manhi <= conv_std_logic_vector(13245,24);
            manlo <= conv_std_logic_vector(108520727,28);
            exponent <= conv_std_logic_vector(2030,11);
      WHEN "1010111011" =>
            manhi <= conv_std_logic_vector(6043387,24);
            manlo <= conv_std_logic_vector(17001813,28);
            exponent <= conv_std_logic_vector(2031,11);
      WHEN "1010111100" =>
            manhi <= conv_std_logic_vector(14239199,24);
            manlo <= conv_std_logic_vector(83422350,28);
            exponent <= conv_std_logic_vector(2032,11);
      WHEN "1010111101" =>
            manhi <= conv_std_logic_vector(4300623,24);
            manlo <= conv_std_logic_vector(142486326,28);
            exponent <= conv_std_logic_vector(2034,11);
      WHEN "1010111110" =>
            manhi <= conv_std_logic_vector(11870538,24);
            manlo <= conv_std_logic_vector(24126621,28);
            exponent <= conv_std_logic_vector(2035,11);
      WHEN "1010111111" =>
            manhi <= conv_std_logic_vector(2690951,24);
            manlo <= conv_std_logic_vector(91850592,28);
            exponent <= conv_std_logic_vector(2037,11);
      WHEN "1011000000" =>
            manhi <= conv_std_logic_vector(9682766,24);
            manlo <= conv_std_logic_vector(203960059,28);
            exponent <= conv_std_logic_vector(2038,11);
      WHEN "1011000001" =>
            manhi <= conv_std_logic_vector(1204206,24);
            manlo <= conv_std_logic_vector(155513539,28);
            exponent <= conv_std_logic_vector(2040,11);
      WHEN "1011000010" =>
            manhi <= conv_std_logic_vector(7662071,24);
            manlo <= conv_std_logic_vector(33184566,28);
            exponent <= conv_std_logic_vector(2041,11);
      WHEN "1011000011" =>
            manhi <= conv_std_logic_vector(16439219,24);
            manlo <= conv_std_logic_vector(11896414,28);
            exponent <= conv_std_logic_vector(2042,11);
      WHEN "1011000100" =>
            manhi <= conv_std_logic_vector(5795691,24);
            manlo <= conv_std_logic_vector(254151921,28);
            exponent <= conv_std_logic_vector(2044,11);
      WHEN "1011000101" =>
            manhi <= conv_std_logic_vector(13902546,24);
            manlo <= conv_std_logic_vector(199613595,28);
            exponent <= conv_std_logic_vector(2045,11);
      WHEN others =>
           manhi <= conv_std_logic_vector(0,24);
           manlo <= conv_std_logic_vector(0,28);
           exponent <= conv_std_logic_vector(0,11);
    END CASE;
  END PROCESS;

END rtl;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   DP_EXPNORND.VHD                           ***
--***                                             ***
--***   Function: DP Exponent Output Block -      ***
--***   Simple                                    ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_expnornd IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentexp : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaexp : IN STD_LOGIC_VECTOR (53 DOWNTO 1); -- includes roundbit
      nanin : IN STD_LOGIC;
      rangeerror : IN STD_LOGIC;

		signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
      --------------------------------------------------
      nanout : OUT STD_LOGIC;
      overflowout : OUT STD_LOGIC;
      underflowout : OUT STD_LOGIC
		);
END dp_expnornd;

ARCHITECTURE rtl OF dp_expnornd IS

  constant expwidth : positive := 11;
  constant manwidth : positive := 52;
  
  signal nanff : STD_LOGIC;
  signal overflownode, underflownode : STD_LOGIC;
  signal overflowff, underflowff : STD_LOGIC;  
  signal mantissaff : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal exponentff : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  
  signal infinitygen : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal zerogen : STD_LOGIC_VECTOR (expwidth DOWNTO 1);  
  signal setmanzero, setmanmax : STD_LOGIC;
  signal setexpzero, setexpmax : STD_LOGIC;

BEGIN

  pra: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN
        
      nanff <= '0';
      overflowff <= '0';
      underflowff <= '0';
      FOR k IN 1 TO manwidth LOOP
        mantissaff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        exponentff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF(enable = '1') THEN 
      
        nanff <= nanin;
        overflowff <= overflownode;
        underflowff <= underflownode;

        -- nan takes precedence (set max)  
        FOR k IN 1 TO manwidth LOOP
          mantissaff(k) <= (mantissaexp(k+1) AND setmanzero) OR setmanmax;
        END LOOP;
               
        FOR k IN 1 TO expwidth LOOP
          exponentff(k) <= (exponentexp(k) AND setexpzero) OR setexpmax;
        END LOOP;
      
      END IF;
             
    END IF;
      
  END PROCESS;
                                                  
--**********************************
--*** CHECK GENERATED CONDITIONS ***   
--**********************************

  -- infinity if exponent == 255
  infinitygen(1) <= exponentexp(1);
  gia: FOR k IN 2 TO expwidth GENERATE
    infinitygen(k) <= infinitygen(k-1) AND exponentexp(k);
  END GENERATE;
                         
  -- zero if exponent == 0
  zerogen(1) <= exponentexp(1);
  gza: FOR k IN 2 TO expwidth GENERATE
    zerogen(k) <= zerogen(k-1) OR exponentexp(k);
  END GENERATE;
                    
  -- trap any other overflow errors
  -- when sign = 0 and rangeerror = 1, overflow
  -- when sign = 1 and rangeerror = 1, underflow
  overflownode <= NOT(signin) AND rangeerror;
  underflownode <= signin AND rangeerror;
  
  -- set mantissa to 0 when infinity or zero condition
  setmanzero <= NOT(infinitygen(expwidth)) AND zerogen(expwidth) AND NOT(rangeerror);
  -- setmantissa to "11..11" when nan
  setmanmax <= nanin;
  -- set exponent to 0 when zero condition 
  setexpzero <= zerogen(expwidth);
  -- set exponent to "11..11" when nan, infinity, or divide by 0
  setexpmax <= nanin OR infinitygen(expwidth) OR rangeerror;
                             
--***************
--*** OUTPUTS ***
--***************

  signout <= '0';   
  mantissaout <= mantissaff;
  exponentout <= exponentff; 
  -----------------------------------------------
  nanout <= nanff;
  overflowout <= overflowff;
  underflowout <= underflowff;

END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   DP_EXPRND.VHD                             ***
--***                                             ***
--***   Function: DP Exponent Output Block -      ***
--***   Rounded                                   ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_exprnd IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentexp : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaexp : IN STD_LOGIC_VECTOR (53 DOWNTO 1); -- includes roundbit
      nanin : IN STD_LOGIC;
      rangeerror : IN STD_LOGIC;

		signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
      --------------------------------------------------
      nanout : OUT STD_LOGIC;
      overflowout : OUT STD_LOGIC;
      underflowout : OUT STD_LOGIC
		);
END dp_exprnd;

ARCHITECTURE rtl OF dp_exprnd IS

  constant expwidth : positive := 11;
  constant manwidth : positive := 52;
  
  type exponentfftype IS ARRAY (2 DOWNTO 1) OF STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  
  signal zerovec : STD_LOGIC_VECTOR (manwidth-1 DOWNTO 1);
  signal nanff : STD_LOGIC_VECTOR (2 DOWNTO 1);
  signal rangeerrorff : STD_LOGIC;
  signal overflownode, underflownode : STD_LOGIC;
  signal overflowff, underflowff : STD_LOGIC_VECTOR (2 DOWNTO 1);
  signal manoverflowbitff : STD_LOGIC; 
  signal roundmantissaff, mantissaff : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal exponentnode : STD_LOGIC_VECTOR (expwidth+2 DOWNTO 1);
  signal exponentoneff : STD_LOGIC_VECTOR (expwidth+2 DOWNTO 1);
  signal exponenttwoff : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
    
  signal manoverflow : STD_LOGIC_VECTOR (manwidth+1 DOWNTO 1);
  signal infinitygen : STD_LOGIC_VECTOR (expwidth+1 DOWNTO 1);
  signal zerogen : STD_LOGIC_VECTOR (expwidth+1 DOWNTO 1);  
  signal setmanzero, setmanmax : STD_LOGIC;
  signal setexpzero, setexpmax : STD_LOGIC;

BEGIN
    
  gzv: FOR k IN 1 TO manwidth-1 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  pra: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN
        
      nanff <= "00";
      rangeerrorff <= '0';
      overflowff <= "00";
      underflowff <= "00";
      manoverflowbitff <= '0';
      FOR k IN 1 TO manwidth LOOP
        roundmantissaff(k) <= '0';
        mantissaff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth+2 LOOP
        exponentoneff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        exponenttwoff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF(enable = '1') THEN 
      
        nanff(1) <= nanin;
        nanff(2) <= nanff(1);
        rangeerrorff <= rangeerror;
        overflowff(1) <= overflownode;
        overflowff(2) <= overflowff(1);
        underflowff(1) <= underflownode;
        underflowff(2) <= underflowff(1);
        
        manoverflowbitff <= manoverflow(manwidth+1);
        
        roundmantissaff <= mantissaexp(manwidth+1 DOWNTO 2) + (zerovec & mantissaexp(1));
        
        -- nan takes precedence (set max)
        -- nan takes precedence (set max)  
        FOR k IN 1 TO manwidth LOOP
          mantissaff(k) <= (roundmantissaff(k) AND setmanzero) OR setmanmax;
        END LOOP;
        
        exponentoneff(expwidth+2 DOWNTO 1) <= "00" & exponentexp;                 
        FOR k IN 1 TO expwidth LOOP
          exponenttwoff(k) <= (exponentnode(k) AND setexpzero) OR setexpmax;
        END LOOP;
      
      END IF;
             
    END IF;
      
  END PROCESS;
  
  exponentnode <= exponentoneff(expwidth+2 DOWNTO 1) + 
                 (zerovec(expwidth+1 DOWNTO 1) & manoverflowbitff);

--*********************************
--*** PREDICT MANTISSA OVERFLOW ***   
--*********************************
     
  manoverflow(1) <= mantissaexp(1);
  gmoa: FOR k IN 2 TO manwidth+1 GENERATE
    manoverflow(k) <= manoverflow(k-1) AND mantissaexp(k);
  END GENERATE; 
                                                                 
--**********************************
--*** CHECK GENERATED CONDITIONS ***   
--**********************************

  -- infinity if exponent == 255
  infinitygen(1) <= exponentnode(1);
  gia: FOR k IN 2 TO expwidth GENERATE
    infinitygen(k) <= infinitygen(k-1) AND exponentnode(k);
  END GENERATE;
  infinitygen(expwidth+1) <= infinitygen(expwidth) OR 
                            (exponentnode(expwidth+1) AND 
                             NOT(exponentnode(expwidth+2))); -- '1' if infinity
                                                    
  -- zero if exponent == 0
  zerogen(1) <= exponentnode(1);
  gza: FOR k IN 2 TO expwidth GENERATE
    zerogen(k) <= zerogen(k-1) OR exponentnode(k);
  END GENERATE;
  zerogen(expwidth+1) <= zerogen(expwidth) AND 
                         NOT(exponentnode(expwidth+2)); -- '0' if zero
                                           
  -- trap any other overflow errors
  -- when sign = 0 and rangeerror = 1, overflow
  -- when sign = 1 and rangeerror = 1, underflow
  overflownode <= NOT(signin) AND rangeerror;
  underflownode <= signin AND rangeerror;
  
  -- set mantissa to 0 when infinity or zero condition
  setmanzero <= NOT(infinitygen(expwidth+1)) AND zerogen(expwidth+1) AND NOT(rangeerrorff);
  -- setmantissa to "11..11" when nan
  setmanmax <= nanff(1);
  -- set exponent to 0 when zero condition 
  setexpzero <= zerogen(expwidth+1);
  -- set exponent to "11..11" when nan, infinity, or divide by 0
  setexpmax <= nanff(1) OR infinitygen(expwidth+1) OR rangeerrorff;
                             
--***************
--*** OUTPUTS ***
--***************
  
  signout <= '0';   
  mantissaout <= mantissaff;
  exponentout <= exponenttwoff; 
  -----------------------------------------------
  nanout <= nanff(2);
  overflowout <= overflowff(2);
  underflowout <= underflowff(2);

END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   DP_EXPRNDPIPE.VHD                         ***
--***                                             ***
--***   Function: DP Exponent Output Block -      ***
--***   Rounded, Pipelined Add                    ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_exprndpipe IS 
GENERIC (synthesize : integer := 1); 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentexp : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaexp : IN STD_LOGIC_VECTOR (53 DOWNTO 1); -- includes roundbit
      nanin : IN STD_LOGIC;
      rangeerror : IN STD_LOGIC;

		signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
      --------------------------------------------------
      nanout : OUT STD_LOGIC;
      overflowout : OUT STD_LOGIC;
      underflowout : OUT STD_LOGIC
		);
END dp_exprndpipe;

ARCHITECTURE rtl OF dp_exprndpipe IS

  constant expwidth : positive := 11;
  constant manwidth : positive := 52;
  
  type exponentfftype IS ARRAY (3 DOWNTO 1) OF STD_LOGIC_VECTOR (expwidth+2 DOWNTO 1);
  
  signal zerovec : STD_LOGIC_VECTOR (manwidth+1 DOWNTO 1);
  signal nanff : STD_LOGIC_VECTOR (3 DOWNTO 1);
  signal rangeerrorff : STD_LOGIC_VECTOR (2 DOWNTO 1);
  signal overflownode, underflownode : STD_LOGIC; 
  signal overflowff, underflowff : STD_LOGIC_VECTOR (3 DOWNTO 1);  
  signal roundmantissanode : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal mantissaff : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal exponentff : exponentfftype;
       
  signal manoverflow : STD_LOGIC_VECTOR (manwidth+1 DOWNTO 1);
  signal manoverflowff : STD_LOGIC;
  signal infinitygen : STD_LOGIC_VECTOR (expwidth+1 DOWNTO 1);
  signal zerogen : STD_LOGIC_VECTOR (expwidth+1 DOWNTO 1);  
  signal setmanzero, setmanmax : STD_LOGIC;
  signal setexpzero, setexpmax : STD_LOGIC;

  component dp_fxadd 
  GENERIC (
           width : positive := 64;
           pipes : positive := 1;
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
        carryin : IN STD_LOGIC;
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
  end component;
  
BEGIN
    
  gzv: FOR k IN 1 TO manwidth+1 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  pra: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN

      nanff <= "000";
      rangeerrorff <= "00";
      overflowff <= "000";
      underflowff <= "000";
      manoverflowff <= '0';
      FOR k IN 1 TO manwidth LOOP
        mantissaff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        exponentff(1)(k) <= '0';
        exponentff(2)(k) <= '0';
        exponentff(3)(k) <= '0';
      END LOOP;
        
    ELSIF (rising_edge(sysclk)) THEN
    
      IF(enable = '1') THEN 
      
        nanff(1) <= nanin;
        nanff(2) <= nanff(1);
        nanff(3) <= nanff(2);
        rangeerrorff(1) <= rangeerror;
        rangeerrorff(2) <= rangeerrorff(1);
        overflowff(1) <= overflownode;
        overflowff(2) <= overflowff(1);
        overflowff(3) <= overflowff(2);
        underflowff(1) <= underflownode;
        underflowff(2) <= underflowff(1);
        underflowff(3) <= underflowff(2);
        
        manoverflowff <= manoverflow(53);
        
        -- nan takes precedence (set max)
        -- nan takes precedence (set max)  
        FOR k IN 1 TO manwidth LOOP
          mantissaff(k) <= (roundmantissanode(k) AND setmanzero) OR setmanmax;
        END LOOP;
        
        exponentff(1)(expwidth+2 DOWNTO 1) <= "00" & exponentexp(expwidth DOWNTO 1);
        exponentff(2)(expwidth+2 DOWNTO 1) <= (exponentff(1)(expwidth+2 DOWNTO 1)) + 
                                              (zerovec(expwidth+1 DOWNTO 1) & manoverflowff);                 
        FOR k IN 1 TO expwidth LOOP
          exponentff(3)(k) <= (exponentff(2)(k) AND setexpzero) OR setexpmax;
        END LOOP;
      
      END IF;
             
    END IF;
      
  END PROCESS;
       
  rndadd: dp_fxadd 
  GENERIC MAP(width=>manwidth,pipes=>2,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>mantissaexp(manwidth+1 DOWNTO 2),bb=>zerovec(manwidth DOWNTO 1),
            carryin=>mantissaexp(1),
            cc=>roundmantissanode);

--*********************************
--*** PREDICT MANTISSA OVERFLOW ***   
--*********************************
     
  manoverflow(1) <= mantissaexp(1);
  gmoa: FOR k IN 2 TO 53 GENERATE
    manoverflow(k) <= manoverflow(k-1) AND mantissaexp(k);
  END GENERATE;                                           
    
--**********************************
--*** CHECK GENERATED CONDITIONS ***   
--**********************************

  -- infinity if exponent >= 255
  infinitygen(1) <= exponentff(2)(1);
  gia: FOR k IN 2 TO expwidth GENERATE
    infinitygen(k) <= infinitygen(k-1) AND exponentff(2)(k);
  END GENERATE;
  infinitygen(expwidth+1) <= infinitygen(expwidth) OR 
                            (exponentff(2)(expwidth+1) AND 
                             NOT(exponentff(2)(expwidth+2))); -- ;1' if infinity
                         
  -- zero if exponent <= 0
  zerogen(1) <= exponentff(2)(1);
  gza: FOR k IN 2 TO expwidth GENERATE
    zerogen(k) <= zerogen(k-1) OR exponentff(2)(k);
  END GENERATE;
  zerogen(expwidth+1) <= zerogen(expwidth) AND 
                         NOT(exponentff(2)(expwidth+2)); -- '0' if zero
  
    -- trap any other overflow errors
  -- when sign = 0 and rangeerror = 1, overflow
  -- when sign = 1 and rangeerror = 1, underflow
  overflownode <= NOT(signin) AND rangeerror;
  underflownode <= signin AND rangeerror;
                    
  -- set mantissa to 0 when infinity or zero condition
  setmanzero <= NOT(infinitygen(expwidth+1)) AND zerogen(expwidth+1) AND NOT(rangeerrorff(2));
  -- setmantissa to "11..11" when nan
  setmanmax <= nanff(2);
  -- set exponent to 0 when zero condition 
  setexpzero <= zerogen(expwidth+1);
  -- set exponent to "11..11" when nan, infinity, or divide by 0
  setexpmax <= nanff(2) OR infinitygen(expwidth+1) OR rangeerrorff(2);
                             
--***************
--*** OUTPUTS ***
--***************

  signout <= '0';   
  mantissaout <= mantissaff;
  exponentout <= exponentff(3)(expwidth DOWNTO 1); 
  -----------------------------------------------
  nanout <= nanff(3);
  overflowout <= overflowff(3);
  underflowout <= underflowff(3);
  
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   ALTERA FLOATING POINT DATAPATH COMPILER   ***
--***                                             ***
--***   DP_FABS.VHD                               ***
--***                                             ***
--***   Function: Single Precision Absolute Value ***
--***                                             ***
--***   abs(x)                                    ***
--***                                             ***
--***   Created 12/09/09                          ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_fabs IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (52 DOWNTO 1);

		  signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
		  satout, zeroout, nanout : OUT STD_LOGIC
		);
END dp_fabs;

ARCHITECTURE rtl OF dp_fabs IS
 
  signal signff : STD_LOGIC;
  signal exponentff : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal mantissaff : STD_LOGIC_VECTOR (52 DOWNTO 1);
  signal expnode : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal expzerochk, expmaxchk : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal expzero, expmax : STD_LOGIC;
  signal manzerochk : STD_LOGIC_VECTOR (52 DOWNTO 1);
  signal manzero, mannonzero : STD_LOGIC; 

BEGIN
    
  pin: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
    
      signff <= '0';
      FOR k IN 1 TO 11 LOOP
        exponentff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 52 LOOP
        mantissaff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF (enable = '1') THEN
          
        signff <= '0';
        exponentff <= exponentin;
        mantissaff <= mantissain;
        
      END IF;
    
    END IF;  
      
  END PROCESS;

  expzerochk(1) <= exponentff(1);
  expmaxchk(1) <= exponentff(1);
  gxa: FOR k IN 2 TO 11 GENERATE
    expzerochk(k) <= expzerochk(k-1) OR exponentff(k);
    expmaxchk(k) <= expmaxchk(k-1) AND exponentff(k);
  END GENERATE;
  expzero <= NOT(expzerochk(11));
  expmax <= expmaxchk(11);
  
  manzerochk(1) <= mantissaff(1);
  gma: FOR k IN 2 TO 52 GENERATE
    manzerochk(k) <= manzerochk(k-1) OR mantissaff(k);
  END GENERATE;
  manzero <= NOT(manzerochk(52));
  mannonzero <= manzerochk(52);
  
  signout <= signff;
  exponentout <= exponentff;
  mantissaout <= mantissaff;
  satout <= expmax AND manzero;
  zeroout <= expzero;
  nanout <= expmax AND mannonzero;

END rtl;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CONVERSION - TOP LEVEL     ***
--***                                             ***
--***   DP_FIXFLOAT.VHD                           ***
--***                                             ***
--***   Function: Convert Fixed Point to Floating ***
--***   Point Number                              ***
--***                                             ***
--***   01/12/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** LATENCY : unsigned = 3 + 3*speed            ***
--*** LATENCY : signed = 4 + 4*speed              ***
--***************************************************

ENTITY dp_fixfloat IS
GENERIC (
         unsigned : integer := 0; -- unsigned = 0, signed = 1
         decimal : integer := 18;
         fractional : integer := 14;
         precision : integer := 0; -- single = 0, double = 1
         speed : integer := 0 -- low speed = 0, high speed = 1 
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      fixed_number : IN STD_LOGIC_VECTOR (decimal+fractional DOWNTO 1);
      
      sign : OUT STD_LOGIC;
      exponent : OUT STD_LOGIC_VECTOR (8+3*precision DOWNTO 1);
      mantissa : OUT STD_LOGIC_VECTOR (23+29*precision DOWNTO 1)    
     );
END dp_fixfloat;

ARCHITECTURE rtl of dp_fixfloat IS

  constant fixed_width : positive := decimal + fractional;
  -- unsigned has 1 bit less (due to leading 1), signed has 2 less (leading 1 and sign)
  constant fixed_precision : positive := fixed_width - unsigned - 1;
  constant mantissa_width : positive := 23 + 29*precision;
  constant exponent_width : positive := 8 + 3*precision;
  constant exponent_base_number : positive := 126+896*precision+decimal;
   
  -- input stage
  signal zerovec : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal exponentbase : STD_LOGIC_VECTOR (exponent_width DOWNTO 1);
  signal invfixed : STD_LOGIC_VECTOR (fixed_width DOWNTO 1);
  signal absnode, delabsnode : STD_LOGIC_VECTOR (fixed_width DOWNTO 1);
  -- detect range stage
  signal clzinbus : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal count, delcount : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal zerochk, delzerochk : STD_LOGIC;
  signal exponentnode, delexponentnode : STD_LOGIC_VECTOR (exponent_width DOWNTO 1);
  -- normalize stage
  signal shiftinbus : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal shiftnode : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal delshift : STD_LOGIC_VECTOR (fixed_width DOWNTO 1);
  signal shiftvalue : STD_LOGIC_VECTOR (64 DOWNTO 1);
  -- output stage
  signal mantissaroundbit : STD_LOGIC;
  signal exponentoutnode : STD_LOGIC_VECTOR (exponent_width DOWNTO 1);
  signal exponentroundnode : STD_LOGIC_VECTOR (exponent_width DOWNTO 1);
    
  component dp_addpipe IS
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
        carryin : IN STD_LOGIC;
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
  end component;
  
  component dp_clz64 IS
  PORT (
        mantissa : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
        
        leading : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
       );
  end component;
  
  component dp_clzpipe64 IS
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        mantissa : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
        
        leading : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
       );
  end component;
 
  component dp_lsft64 IS
  PORT (
        inbus : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);      
        
        outbus : OUT STD_LOGIC_VECTOR (64 DOWNTO 1)    
       );
  end component;
  
  component dp_lsftpipe64 IS
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        inbus : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);      
        
        outbus : OUT STD_LOGIC_VECTOR (64 DOWNTO 1)    
       );
  end component;
  
  component fp_del IS 
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
 end component;

  component fp_delbit IS 
  GENERIC (
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC; 
      
        cc : OUT STD_LOGIC
       );
 end component;
     
BEGIN
    
  gera : IF NOT((precision = 0) OR 
	             (precision = 1)) GENERATE
	 assert false report "precision must be 0 (single precision) or 1 (double precision)" severity error;
  END GENERATE;
  
  gerb : IF NOT((speed = 0) OR 
	             (speed = 1)) GENERATE
	 assert false report "speed must be 0 or 1" severity error;
  END GENERATE;
  
  gerc : IF NOT((unsigned = 0) OR 
	             (unsigned = 1)) GENERATE
	 assert false report "unsigned must be 0 or 1" severity error;
  END GENERATE;

  gerd : IF (decimal < 1) GENERATE
	 assert false report "decimal must be greater than 1" severity error;
  END GENERATE;
  
  gere : IF (fixed_width > 64) GENERATE
	 assert false report "maximum fixed point precision must be 64 or less" severity error;
  END GENERATE; 
  
  gza: FOR k IN 1 TO 64 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  exponentbase <= conv_std_logic_vector (exponent_base_number,exponent_width);
  
  --*** LEVEL 0 - 2 (ABSNODE) ***
  -- level 0 if unsigned = 0, 
  -- level 1 if signed = 1 & speed = 0, 
  -- level 2 if signed = 1 & speed = 1 
  gabsa: IF (unsigned = 1) GENERATE  
    giva: FOR k IN 1 TO fixed_width GENERATE
      invfixed(k) <= fixed_number(k) XOR fixed_number(fixed_width);
    END GENERATE;
    aabs: dp_addpipe
    GENERIC MAP (width=>fixed_width,pipes=>speed+1)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>invfixed,bb=>zerovec(fixed_width DOWNTO 1),carryin=>fixed_number(fixed_width),
              cc=>absnode);
  END GENERATE;
   
  gabsb: IF (unsigned = 0) GENERATE  
    invfixed <= fixed_number;
    absnode <= invfixed;
  END GENERATE;   
  
  gczc: IF (fixed_width < 64) GENERATE
    clzinbus <= absnode & zerovec(64-fixed_width DOWNTO 1);
  END GENERATE;
  gczd: IF (fixed_width = 64) GENERATE
    clzinbus <= absnode;
  END GENERATE;
  
  --*** LEVEL 1-4 (ABSDELNODE, COUNTFF) ***
  -- level 1 if unsigned = 0 & speed = 0,
  -- level 2 if unsigned = 0 & speed = 1, 
  -- level 2 if signed = 1 & speed = 0, 
  -- level 4 if signed = 1 & speed = 1 
  
  gcca: IF (speed = 0) GENERATE
    cntzip: dp_clz64
    PORT MAP (mantissa=>clzinbus,leading=>count);
  END GENERATE;
  gccb: IF (speed = 1) GENERATE
    cntone: dp_clzpipe64
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              mantissa=>clzinbus,leading=>count);
  END GENERATE;
  
  delabsbus: fp_del
  GENERIC MAP (width=>fixed_width,pipes=>speed+1)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>absnode,cc=>delabsnode);
  
  ddc: fp_del
  GENERIC MAP (width=>6,pipes=>1)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>count,cc=>delcount);
  
  -- check for 0 input - when countff = 0 and absdelnode(64) (unsigned) or 
  -- absdelnode(63) (signed) not '1'
  zerochk <= NOT(delcount(6) OR delcount(5) OR delcount(4) OR delcount(3) OR
                 delcount(2) OR delcount(1) OR delabsnode(fixed_width) OR delabsnode(fixed_width-1));
                 
  delzc: fp_delbit
  GENERIC MAP (pipes=>speed+1)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>zerochk,cc=>delzerochk);
            
  exponentnode <= exponentbase - (zerovec(2+3*precision DOWNTO 1) & delcount);  
  
  delx: fp_del
  GENERIC MAP (width=>exponent_width,pipes=>speed+1)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>exponentnode,cc=>delexponentnode);
            
  --*** LEVEL 2-6 (SHIFTFF) ***
  -- level 2 if unsigned = 0 & speed = 0,
  -- level 3 if unsigned = 0 & speed = 1, 
  -- level 3 if signed = 1 & speed = 0, 
  -- level 6 if signed = 1 & speed = 1 

  gfsc: IF (fixed_width < 64) GENERATE
    shiftinbus <= delabsnode & zerovec(64-fixed_width DOWNTO 1);
  END GENERATE;
  gfsd: IF (fixed_width = 64) GENERATE
    shiftinbus <= delabsnode;
  END GENERATE;

  gssa: IF (speed = 0) GENERATE
    sftzip: dp_lsft64
    PORT MAP (inbus=>shiftinbus,shift=>delcount,
              outbus=>shiftnode);
  END GENERATE;
  gssb: IF (speed = 1) GENERATE
    sftone: dp_lsftpipe64
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              inbus=>shiftinbus,shift=>delcount,
              outbus=>shiftnode);
  END GENERATE;
  
  dels: fp_del
  GENERIC MAP (width=>fixed_width,pipes=>1)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>shiftnode(64 DOWNTO 65-fixed_width),cc=>delshift);

  gsoa: IF (fixed_width = 64) GENERATE
    shiftvalue <= delshift;
  END GENERATE;
  gsob: IF (fixed_width < 64) GENERATE
    shiftvalue <= delshift & zerovec(64-fixed_width DOWNTO 1);
  END GENERATE;
   
  --*** LEVEL 3-8 (OUTPUT) ***
  -- level 3 if unsigned = 0 & speed = 0,
  -- level 5 if unsigned = 0 & speed = 1, 
  -- level 4 if signed = 1 & speed = 0, 
  -- level 8 if signed = 1 & speed = 1 

  -- single precision
  goa: IF (fixed_precision <= 23 AND mantissa_width = 23) GENERATE
    mantissaroundbit <= '0';
    exponentroundnode <= delexponentnode;
    goax: FOR k IN 1 TO 8 GENERATE
      exponentoutnode(k) <= exponentroundnode(k) AND NOT(delzerochk);
    END GENERATE;
  END GENERATE;
  
  gob: IF (fixed_precision > 23 AND mantissa_width = 23) GENERATE
    mantissaroundbit <= ( shiftvalue(41) AND shiftvalue(40) ) OR
                        (NOT(shiftvalue(41)) AND shiftvalue(40) AND
                         (shiftvalue(39) OR shiftvalue(38) OR shiftvalue(37) OR shiftvalue(36) OR 
                          shiftvalue(35) OR shiftvalue(34) OR shiftvalue(33) OR shiftvalue(32) OR 
                          shiftvalue(31) OR shiftvalue(30) OR shiftvalue(29) OR shiftvalue(28)));
    -- check for mantissa overflow here
    exponentroundnode <= delexponentnode;
    gobx: FOR k IN 1 TO 8 GENERATE
      exponentoutnode(k) <= exponentroundnode(k) AND NOT(delzerochk);
    END GENERATE;
  END GENERATE;
  
  -- double precision
  goc: IF (fixed_precision <= 52 AND mantissa_width = 52) GENERATE
    mantissaroundbit <= '0';
    exponentroundnode <= delexponentnode;
    gocx: FOR k IN 1 TO 11 GENERATE
      exponentoutnode(k) <= exponentroundnode(k) AND NOT(delzerochk);
    END GENERATE;
  END GENERATE;
  
  god: IF (fixed_width > 52 AND mantissa_width = 52) GENERATE
    mantissaroundbit <= (shiftvalue(12) AND shiftvalue(11)) OR
                        (NOT(shiftvalue(12)) AND shiftvalue(11) AND
                         (shiftvalue(10) OR shiftvalue(9) OR shiftvalue(8) OR shiftvalue(7) OR 
                          shiftvalue(6) OR shiftvalue(5) OR shiftvalue(4) OR shiftvalue(3) OR 
                          shiftvalue(2) OR shiftvalue(1)));
    -- check for mantissa overflow here
    exponentroundnode <= delexponentnode;
    godx: FOR k IN 1 TO 11 GENERATE
      exponentoutnode(k) <= exponentroundnode(k) AND NOT(delzerochk);
    END GENERATE;
  END GENERATE;
  
  gsgna: IF (unsigned = 0) GENERATE
    sign <= '0';
  END GENERATE;
  gsgnb: IF (unsigned = 1) GENERATE
    delss: fp_delbit
    GENERIC MAP (pipes=>4+4*speed)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>fixed_number(decimal+fractional),cc=>sign);  
  END GENERATE;
  
  mno: dp_addpipe
  GENERIC MAP (width=>mantissa_width,pipes=>speed+1)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>shiftvalue(63 DOWNTO 64-mantissa_width),
            bb=>zerovec(mantissa_width DOWNTO 1),
            carryin=>mantissaroundbit,
            cc=>mantissa);
            
  exo: dp_addpipe
  GENERIC MAP (width=>exponent_width,pipes=>speed+1)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>exponentoutnode,
            bb=>zerovec(exponent_width DOWNTO 1),
            --carryin=>mantissaoverflowbit,
            carryin=>'0',
            cc=>exponent);
                
END rtl;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CONVERSION - TOP LEVEL     ***
--***                                             ***
--***   DP_FLOATFIX.VHD                           ***
--***                                             ***
--***   Function: Convert Floating Point to Fixed ***
--***   Point Number                              ***
--***                                             ***
--***   07/12/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** LATENCY :                                   ***
--***           speed = 0 : 3                     ***
--***           speed = 1 : 5                     ***
--***************************************************

--***************************************************
--*** OUTPUT FORMAT - UNSIGNED                    ***
--*** maximum number is (2^decimal)-1, else       ***
--*** saturate. if input negative, zero output    ***
--*** OUTPUT FORMAT - SIGNED                      ***
--*** maximum number is (2^decimal-1)-1, else     ***
--*** saturate                                    ***
--***************************************************

ENTITY dp_floatfix IS
GENERIC (
         unsigned : integer := 1;  -- unsigned = 0, signed = 1
         decimal : integer := 14;
         fractional : integer := 6;
         precision : integer := 0; -- single = 0, double = 1
         speed : integer := 0 -- low speed = 0, high speed = 1
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      sign : IN STD_LOGIC;
      exponent : IN STD_LOGIC_VECTOR (8+3*precision DOWNTO 1);
      mantissa : IN STD_LOGIC_VECTOR (23+29*precision DOWNTO 1);
      
      fixed_number : OUT STD_LOGIC_VECTOR (decimal+fractional DOWNTO 1)
     );
END dp_floatfix;

ARCHITECTURE rtl of dp_floatfix IS

  constant fixed_width : positive := decimal + fractional;
  constant mantissa_width : positive := 23 + 29*precision;
  constant exponent_width : positive := 8 + 3*precision;
  constant exponent_base_number : positive := 127+896*precision;
  
  -- input stage
  signal zerovec : STD_LOGIC_VECTOR (116 DOWNTO 1);
  signal exponent_base_node : STD_LOGIC_VECTOR (exponent_width+1 DOWNTO 1);
  signal saturate_check : STD_LOGIC_VECTOR (exponent_width+1 DOWNTO 1);
  signal saturate_output, zero_output : STD_LOGIC;
  signal saturate_apply, zero_apply : STD_LOGIC;
  signal sign_apply : STD_LOGIC;
  signal signed_mantissa_node : STD_LOGIC_VECTOR (mantissa_width+2 DOWNTO 1);
  signal signed_mantissa_comp : STD_LOGIC_VECTOR (mantissa_width+2 DOWNTO 1);
  signal signed_mantissa : STD_LOGIC_VECTOR (mantissa_width+2 DOWNTO 1);
  signal input_vector : STD_LOGIC_VECTOR (116 DOWNTO 1);
  signal negexponent : STD_LOGIC_VECTOR (exponent_width DOWNTO 1);
  signal expbase, negexpbase : STD_LOGIC_VECTOR (exponent_width DOWNTO 1);
  signal leftshift, rightshift : STD_LOGIC_VECTOR (exponent_width DOWNTO 1);
  -- shift stage
  signal leftbus, rightbus : STD_LOGIC_VECTOR (116 DOWNTO 1);
  signal shiftbus, shiftbusff : STD_LOGIC_VECTOR (fixed_width DOWNTO 1);
  signal select_bit : STD_LOGIC;
  -- output stage
  signal fixed_numberff : STD_LOGIC_VECTOR (fixed_width DOWNTO 1);
    
  component dp_addpipe IS
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
        carryin : IN STD_LOGIC;
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
  end component;
   
  component dp_lsft64x64 IS
  PORT (
        inbus : IN STD_LOGIC_VECTOR (116 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);      
        
        outbus : OUT STD_LOGIC_VECTOR (116 DOWNTO 1)    
       );
  end component;
  
  component dp_lsftpipe64x64 IS
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        inbus : IN STD_LOGIC_VECTOR (116 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);      
        
        outbus : OUT STD_LOGIC_VECTOR (116 DOWNTO 1)    
       );
  end component;
  
  component dp_rsft64x64 IS
  PORT (
        inbus : IN STD_LOGIC_VECTOR (116 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);      
        
        outbus : OUT STD_LOGIC_VECTOR (116 DOWNTO 1)    
       );
  end component;
  
  component dp_rsftpipe64x64 IS
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        inbus : IN STD_LOGIC_VECTOR (116 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);      
        
        outbus : OUT STD_LOGIC_VECTOR (116 DOWNTO 1)    
       );
  end component;
  
  component fp_delbit IS 
  GENERIC (
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC; 
      
        cc : OUT STD_LOGIC
       );
 end component;
  
BEGIN
  
  gera : IF NOT((unsigned = 0) OR 
	             (unsigned = 1)) GENERATE
	 assert false report "unsigned must be 0 or 1" severity error;
  END GENERATE;
    
  gerb : IF NOT((precision = 0) OR 
	             (precision = 1)) GENERATE
	 assert false report "precision must be 0 (single precision) or 1 (double precision)" severity error;
  END GENERATE;
  
  gerc : IF NOT((speed = 0) OR 
	             (speed = 1)) GENERATE
	 assert false report "speed must be 0 or 1" severity error;
  END GENERATE;
 
  gerd : IF (decimal < 2) GENERATE
	 assert false report "decimal must be greater than 2" severity error;
  END GENERATE;
  
  gere : IF (fixed_width > 64) GENERATE
	 assert false report "maximum fixed point precision must be 64 or less" severity error;
  END GENERATE; 

  gza: FOR k IN 1 TO 116 GENERATE
    zerovec(k) <= '0';
  END GENERATE;

  --*** LEVEL 1-2 ***
  -- level 1 if speed = 0
  -- level 2 if speed = 1
  
  -- check for zero and saturate conditions
  exponent_base_node <= conv_std_logic_vector(exponent_base_number,exponent_width+1);
  
  gzsa: IF (unsigned = 0) GENERATE
    saturate_check <= exponent - exponent_base_node - decimal;
    -- '1' when condition true
    saturate_output <= NOT(saturate_check(exponent_width+1));
    zero_output <= sign;
  END GENERATE;
  
  gzsb: IF (unsigned = 1) GENERATE
    saturate_check <= exponent - exponent_base_node - decimal + 1;
    -- '1' when condition true
    saturate_output <= NOT(saturate_check(exponent_width+1));
    zero_output <= '0';
    
    dss: fp_delbit
    GENERIC MAP (pipes=>2+2*speed)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>sign,
              cc=>sign_apply);
              
  END GENERATE;
  
  ds: fp_delbit
  GENERIC MAP (pipes=>2+2*speed)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>saturate_output,
              cc=>saturate_apply);
              
  dz: fp_delbit
  GENERIC MAP (pipes=>2+2*speed)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>zero_output,
              cc=>zero_apply);
               
  signed_mantissa_node <= "01" & mantissa;
  gsma: FOR k IN 1 TO mantissa_width+2 GENERATE
    signed_mantissa_comp(k) <= signed_mantissa_node(k) XOR sign;
  END GENERATE;
  
  addtop: dp_addpipe
  GENERIC MAP (width=>mantissa_width+2,pipes=>speed+1)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>signed_mantissa_comp,bb=>zerovec(mantissa_width+2 DOWNTO 1),
            carryin=>sign,
            cc=>signed_mantissa);
  
  giva: FOR k IN 116-decimal+3 TO 116 GENERATE
    input_vector(k) <= signed_mantissa(mantissa_width+2);
  END GENERATE;
  input_vector(116-decimal+2 DOWNTO 116-decimal-mantissa_width+1) <= signed_mantissa;
  givb: IF (116-decimal-mantissa_width+1 > 1) GENERATE
    input_vector(116-decimal-mantissa_width DOWNTO 1) <= zerovec(116-decimal-mantissa_width DOWNTO 1);
  END GENERATE;
  
  gcxa: FOR k IN 1 TO exponent_width GENERATE
    negexponent(k) <= NOT(exponent(k));
  END GENERATE;
  gcxb: FOR k IN 1 TO exponent_width-1 GENERATE
    expbase(k) <= '1';
    negexpbase(k) <= '0';
  END GENERATE;
  expbase(exponent_width) <= '0';
  negexpbase(exponent_width) <= '1';
  
  sublx: dp_addpipe
  GENERIC MAP (width=>exponent_width,pipes=>speed+1)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>exponent,bb=>negexpbase,
            carryin=>'1',
            cc=>leftshift);
            
  subrx: dp_addpipe
  GENERIC MAP (width=>exponent_width,pipes=>speed+1)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>negexponent,bb=>expbase,
            carryin=>'1',
            cc=>rightshift);

  --*** LEVEL 2-4 (shiftbusff) ***
  -- level 2 if speed = 0
  -- level 4 if speed = 1
  
  gsfa: IF (speed = 0) GENERATE
    clsc: dp_lsft64x64
    PORT MAP (inbus=>input_vector,shift=>leftshift(6 DOWNTO 1),
              outbus=>leftbus);
            
    crsc: dp_rsft64x64
    PORT MAP (inbus=>input_vector,shift=>rightshift(6 DOWNTO 1),
              outbus=>rightbus);
              
    select_bit <= leftshift(exponent_width);
  END GENERATE;
  
  gsfb: IF (speed = 1) GENERATE
    clsp: dp_lsftpipe64x64
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              inbus=>input_vector,shift=>leftshift(6 DOWNTO 1),
              outbus=>leftbus);
            
    crsp: dp_rsftpipe64x64
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              inbus=>input_vector,shift=>rightshift(6 DOWNTO 1),
              outbus=>rightbus);
              
    db: fp_delbit
    GENERIC MAP (pipes=>1)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>leftshift(exponent_width),
              cc=>select_bit);
  END GENERATE;
    
  gsba: FOR k IN 1 TO fixed_width GENERATE
    shiftbus(k) <= (leftbus(116-fixed_width+k) AND NOT(select_bit)) OR
                   (rightbus(116-fixed_width+k) AND select_bit);
  END GENERATE;
  
  psa: PROCESS (sysclk,reset)
  BEGIN
    IF (reset = '1') THEN
      FOR k IN 1 TO fixed_width LOOP
        shiftbusff(k) <= '0';
      END LOOP; 
    ELSIF (rising_edge(sysclk)) THEN
      IF (enable = '1') THEN
        shiftbusff <= shiftbus;
      END IF;
    END IF;
  END PROCESS;
  
  --*** LEVEL 3-5 ***
  -- level 3 if speed = 0
  -- level 5 if speed = 1

  gou: IF (unsigned = 0) GENERATE
    poa: PROCESS (sysclk,reset)
    BEGIN
      IF (reset = '1') THEN
        FOR k IN 1 TO fixed_width LOOP
          fixed_numberff(k) <= '0';
        END LOOP; 
      ELSIF (rising_edge(sysclk)) THEN
        IF (enable = '1') THEN
          FOR k IN 1 TO fixed_width LOOP    
            fixed_numberff(k) <= (shiftbusff(k) AND NOT(zero_apply)) OR saturate_apply;
          END LOOP;
        END IF;
      END IF;
    END PROCESS;
  END GENERATE;

  gos: IF (unsigned = 1) GENERATE
    pos: PROCESS (sysclk,reset)
    BEGIN
      IF (reset = '1') THEN
        FOR k IN 1 TO fixed_width LOOP
          fixed_numberff(k) <= '0';
        END LOOP; 
      ELSIF (rising_edge(sysclk)) THEN
        IF (enable = '1') THEN
          FOR k IN 1 TO fixed_width-1 LOOP    
            fixed_numberff(k) <= (shiftbusff(k) AND NOT(zero_apply) AND 
                                  NOT(saturate_apply AND sign_apply)) OR
                                 (saturate_apply AND NOT(sign_apply));
          END LOOP;
          fixed_numberff(fixed_width) <= (shiftbusff(fixed_width) AND NOT(zero_apply) AND 
                                          NOT(saturate_apply AND NOT(sign_apply))) OR
                                         (saturate_apply AND sign_apply);
        END IF;
      END IF;
    END PROCESS;
  END GENERATE;
    
  fixed_number <= fixed_numberff;
  
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_FXADD.VHD                              ***
--***                                             ***
--***   Function: Generic Fixed Point Adder       ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_fxadd IS 
GENERIC (
         width : positive := 64;
         pipes : positive := 1;
         synthesize : integer := 0
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      carryin : IN STD_LOGIC;
      
      cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
     );
END dp_fxadd;

ARCHITECTURE rtl OF dp_fxadd IS

  component dp_addb IS
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
        carryin : IN STD_LOGIC;
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
  end component;
  
  component dp_adds IS
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
        carryin : IN STD_LOGIC;
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
  end component;
   
BEGIN
  
  gaa: IF (synthesize = 0) GENERATE
    addone: dp_addb
    GENERIC MAP (width=>width,pipes=>pipes)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>aa,bb=>bb,carryin=>carryin,
              cc=>cc);
  END GENERATE;
  
  gab: IF (synthesize = 1) GENERATE
    addtwo: dp_adds
    GENERIC MAP (width=>width,pipes=>pipes)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>aa,bb=>bb,carryin=>carryin,
              cc=>cc);
  END GENERATE;
       
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_FXSUB.VHD                              ***
--***                                             ***
--***   Function: Generic Fixed Point Subtractor  ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_fxsub IS 
GENERIC (
         width : positive := 64;
         pipes : positive := 1;
         synthesize : integer := 0
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      borrowin : IN STD_LOGIC;
      
      cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
     );
END dp_fxsub;

ARCHITECTURE rtl OF dp_fxsub IS

  component dp_subb IS
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
        borrowin : IN STD_LOGIC;
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
  end component;
  
  component dp_subs IS
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
        borrowin : IN STD_LOGIC;
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
  end component;
   
BEGIN
  
  gaa: IF (synthesize = 0) GENERATE
    addone: dp_subb
    GENERIC MAP (width=>width,pipes=>pipes)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>aa,bb=>bb,borrowin=>borrowin,
              cc=>cc);
  END GENERATE;
  
  gab: IF (synthesize = 1) GENERATE
    addtwo: dp_subs
    GENERIC MAP (width=>width,pipes=>pipes)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>aa,bb=>bb,borrowin=>borrowin,
              cc=>cc);
  END GENERATE;
       
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   DOUBLE PRECISION INVERSE - TOP LEVEL      ***
--***                                             ***
--***   DP_INV.VHD                                ***
--***                                             ***
--***   Function: IEEE754 DP Inverse              ***
--***   (multiplicative iterative algorithm)      ***
--***                                             ***
--***   12/08/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--***                                             ***
--*** Stratix II                                  ***
--*** Latency = 20 + 2*DoubleSpeed +              ***
--***           RoundConvert*(1+DoubleSpeed)      ***
--*** DoubleSpeed = 0, Roundconvert = 0 : 20      ***
--*** DoubleSpeed = 1, Roundconvert = 0 : 22      ***
--*** DoubleSpeed = 0, Roundconvert = 1 : 21      ***
--*** DoubleSpeed = 1, Roundconvert = 1 : 24      ***
--***                                             ***
--*** Stratix III/IV                              ***
--*** Latency = 19 + DoubleSpeed +                ***
--***           Roundconvert*(1+DoubleSpeed)      ***
--*** DoubleSpeed = 0, Roundconvert = 0 : 19      ***
--*** DoubleSpeed = 1, Roundconvert = 0 : 20      ***
--*** DoubleSpeed = 0, Roundconvert = 1 : 20      ***
--*** DoubleSpeed = 1, Roundconvert = 1 : 22      ***
--***                                             ***
--***************************************************

ENTITY dp_inv IS 
GENERIC (
         roundconvert : integer := 0; -- 0 = no round, 1 = round
         doubleaccuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
         doublespeed : integer := 0;   -- 0/1
         device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
         synthesize : integer := 1   -- 0/1    
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (52 DOWNTO 1);

		signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
      --------------------------------------------------
      nanout : OUT STD_LOGIC;
      invalidout : OUT STD_LOGIC;
      dividebyzeroout : OUT STD_LOGIC
		);
END dp_inv;

ARCHITECTURE rtl OF dp_inv IS
  
  constant expwidth : positive := 11;
  constant manwidth : positive := 52;
  
  -- SII Latency = 19 + 2*speed                  
  -- SIII Latency = 18 + speed                   
  constant coredepth : positive := 19+2*doublespeed - device*(1+doublespeed);
  
  type expfftype IS ARRAY (coredepth-1 DOWNTO 1) OF STD_LOGIC_VECTOR (expwidth+2 DOWNTO 1);
  
  signal zerovec : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
    
  signal signinff : STD_LOGIC;
  signal manff : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal expinff : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal expoffset : STD_LOGIC_VECTOR (expwidth+2 DOWNTO 1);
  signal invertnum : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal quotient : STD_LOGIC_VECTOR (55 DOWNTO 1);
  signal signff : STD_LOGIC_VECTOR (coredepth-1 DOWNTO 1);  
  signal expff : expfftype;  

  -- conditions
  signal zeroman : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal zeroexp : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal maxexp : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal zeromaninff : STD_LOGIC;
  signal zeroexpinff : STD_LOGIC;
  signal maxexpinff : STD_LOGIC;
  signal zeroinff : STD_LOGIC;
  signal infinityinff : STD_LOGIC;
  signal naninff : STD_LOGIC;
  signal dividebyzeroff, nanff : STD_LOGIC_VECTOR (coredepth-3 DOWNTO 1);

  component dp_inv_core 
  GENERIC (
           doublespeed : integer := 0;  -- 0/1
           doubleaccuracy : integer := 0;  -- 0/1
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 1      -- 0/1      
          ); 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        divisor : IN STD_LOGIC_VECTOR (54 DOWNTO 1);

		  quotient : OUT STD_LOGIC_VECTOR (55 DOWNTO 1)
		  );
  end component;
  
  component dp_divnornd
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        signin : IN STD_LOGIC;
        exponentdiv : IN STD_LOGIC_VECTOR (13 DOWNTO 1);
        mantissadiv : IN STD_LOGIC_VECTOR (53 DOWNTO 1);
        nanin : IN STD_LOGIC;
        dividebyzeroin : IN STD_LOGIC;

		  signout : OUT STD_LOGIC;
        exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
        mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
        --------------------------------------------------
        nanout : OUT STD_LOGIC;
        invalidout : OUT STD_LOGIC;
        dividebyzeroout : OUT STD_LOGIC
		  );
  end component;
       	
  component dp_divrnd
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        signin : IN STD_LOGIC;
        exponentdiv : IN STD_LOGIC_VECTOR (13 DOWNTO 1);
        mantissadiv : IN STD_LOGIC_VECTOR (53 DOWNTO 1);
        nanin : IN STD_LOGIC;
        dividebyzeroin : IN STD_LOGIC;

		  signout : OUT STD_LOGIC;
        exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
        mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
        --------------------------------------------------
        nanout : OUT STD_LOGIC;
        invalidout : OUT STD_LOGIC;
        dividebyzeroout : OUT STD_LOGIC
		  );
  end component;

  component dp_divrndpipe
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        signin : IN STD_LOGIC;
        exponentdiv : IN STD_LOGIC_VECTOR (13 DOWNTO 1);
        mantissadiv : IN STD_LOGIC_VECTOR (53 DOWNTO 1);
        nanin : IN STD_LOGIC;
        dividebyzeroin : IN STD_LOGIC;

		  signout : OUT STD_LOGIC;
        exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
        mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
        --------------------------------------------------
        nanout : OUT STD_LOGIC;
        invalidout : OUT STD_LOGIC;
        dividebyzeroout : OUT STD_LOGIC
		  );
  end component;
BEGIN
    
  gzva: FOR k IN 1 TO manwidth GENERATE
    zerovec(k) <= '0';
  END GENERATE;

  gxa: FOR k IN 1 TO expwidth-1 GENERATE
    expoffset(k) <= '1';
  END GENERATE;
  expoffset(expwidth+2 DOWNTO expwidth) <= "000";

  pma: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
  
      FOR k IN 1 TO manwidth LOOP
        manff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        expinff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO coredepth-1 LOOP
        signff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO coredepth-1 LOOP
        FOR j IN 1 TO expwidth+2 LOOP
          expff(k)(j) <= '0';
        END LOOP;
      END LOOP;
    
    ELSIF (rising_edge(sysclk)) THEN

      IF (enable = '1') THEN
        
        signinff <= signin;
        manff <= mantissain;
        expinff <= exponentin;

        signff(1) <= signinff;
        FOR k IN 2 TO coredepth-1 LOOP
          signff(k) <= signff(k-1);
        END LOOP;
    
        expff(1)(expwidth+2 DOWNTO 1) <= expoffset - ("00" & expinff);
        expff(2)(expwidth+2 DOWNTO 1) <= expff(1)(expwidth+2 DOWNTO 1) + expoffset;
        FOR k IN 3 TO coredepth-2 LOOP
          expff(k)(expwidth+2 DOWNTO 1) <= expff(k-1)(expwidth+2 DOWNTO 1);
        END LOOP;
        -- quotient always <1, so decrement exponent
        expff(coredepth-1)(expwidth+2 DOWNTO 1) <= expff(coredepth-2)(expwidth+2 DOWNTO 1) - 
                                                  (zerovec(expwidth+1 DOWNTO 1) & '1');   
                                                  
      END IF;
  
    END IF;
  
  END PROCESS;

--********************
--*** CHECK INPUTS ***
--********************

  zeroman(1) <= manff(1);
  gca: FOR k IN 2 TO manwidth GENERATE
    zeroman(k) <= zeroman(k-1) OR manff(k);
  END GENERATE; 
  zeroexp(1) <= expinff(1);
  gcb: FOR k IN 2 TO expwidth GENERATE
    zeroexp(k) <= zeroexp(k-1) OR expinff(k);
  END GENERATE;
  maxexp(1) <= expinff(1);
  gcc: FOR k IN 2 TO expwidth GENERATE
    maxexp(k) <= maxexp(k-1) AND expinff(k);
  END GENERATE;

  pcc: PROCESS (sysclk,reset)
  BEGIN
    
    IF (reset = '1') THEN
      
      zeromaninff <= '0';  
      zeroexpinff <= '0'; 
      maxexpinff <= '0';  
      zeroinff <= '0';
      infinityinff <= '0';
      naninff <= '0';
      FOR k IN 1 TO coredepth-3 LOOP
        dividebyzeroff(k) <= '0';
        nanff(k) <= '0';
      END LOOP;
     
    ELSIF (rising_edge(sysclk)) THEN
            
      IF (enable = '1') THEN
     
        zeromaninff <= zeroman(manwidth);
        zeroexpinff <= zeroexp(expwidth);
        maxexpinff <= maxexp(expwidth);
    
        -- zero when man = 0, exp = 0
        -- infinity when man = 0, exp = max
        -- nan when man != 0, exp = max
    
        -- all ffs '1' when condition true
        zeroinff <= NOT(zeromaninff OR zeroexpinff); 
        infinityinff <= NOT(zeromaninff) AND maxexpinff;
        naninff <= zeromaninff AND maxexpinff;

        -- nan output when nan input
        nanff(1) <= naninff;
        FOR k IN 2 TO coredepth-3 LOOP
          nanff(k) <= nanff(k-1);
        END LOOP;
        
        dividebyzeroff(1) <= zeroinff;
        FOR k IN 2 TO coredepth-3 LOOP
          dividebyzeroff(k) <= dividebyzeroff(k-1);
        END LOOP;
      
      END IF;
   
    END IF;

  END PROCESS;


--*******************
--*** DIVIDE CORE ***
--*******************

  invertnum <= '1' & mantissain & '0';

  invcore: dp_inv_core
  GENERIC MAP (doublespeed=>doublespeed,doubleaccuracy=>doubleaccuracy,
               device=>device,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            divisor=>invertnum,
            quotient=>quotient);
  -- quotient always <1
  
--************************
--*** ROUND AND OUTPUT ***
--************************

  -- in depth coredepth+1 (core + normalff)

  gra: IF (roundconvert = 0) GENERATE

    norndout: dp_divnornd
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              signin=>signff(coredepth-1),
              exponentdiv=>expff(coredepth-1)(expwidth+2 DOWNTO 1),
              mantissadiv=>quotient(53 DOWNTO 1),
              nanin=>nanff(coredepth-3),
              dividebyzeroin=>dividebyzeroff(coredepth-3),

              signout=>signout,exponentout=>exponentout,mantissaout=>mantissaout,
              nanout=>nanout,invalidout=>invalidout,dividebyzeroout=>dividebyzeroout);
            
  END GENERATE;
  
  grb: IF (roundconvert = 1 AND doublespeed = 0) GENERATE

    rndout: dp_divrnd
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              signin=>signff(coredepth-1),
              exponentdiv=>expff(coredepth-1)(expwidth+2 DOWNTO 1),
              mantissadiv=>quotient(53 DOWNTO 1),
              nanin=>nanff(coredepth-3),
              dividebyzeroin=>dividebyzeroff(coredepth-3),

              signout=>signout,exponentout=>exponentout,mantissaout=>mantissaout,
              nanout=>nanout,invalidout=>invalidout,dividebyzeroout=>dividebyzeroout);
            
  END GENERATE;

  grc: IF (roundconvert = 1 AND doublespeed = 1) GENERATE
    
    rndoutpipe: dp_divrndpipe
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              signin=>signff(coredepth-1),
              exponentdiv=>expff(coredepth-1)(expwidth+2 DOWNTO 1),
              mantissadiv=>quotient(53 DOWNTO 1),
              nanin=>nanff(coredepth-3),
              dividebyzeroin=>dividebyzeroff(coredepth-3),

              signout=>signout,exponentout=>exponentout,mantissaout=>mantissaout,
              nanout=>nanout,invalidout=>invalidout,dividebyzeroout=>dividebyzeroout);
            
  END GENERATE;
  
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   DOUBLE PRECISION INVERSE - CORE           ***
--***                                             ***
--***   DP_INV_CORE.VHD                           ***
--***                                             ***
--***   Function: 54 bit Inverse                  ***
--***   (multiplicative iterative algorithm)      ***
--***                                             ***
--***   09/12/07 ML                               ***
--***                                             ***
--***   (c) 2007 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***   24/04/09 - SIII/SIV multiplier support    ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** SII Latency = 19 + 2*doublepeed             ***
--*** SIII Latency = 18 + doublespeed             ***
--***************************************************

ENTITY dp_inv_core IS 
GENERIC (
         doublespeed : integer := 0;  -- 0/1
         doubleaccuracy : integer := 0;  -- 0/1
         device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
         synthesize : integer := 1      -- 0/1      
        ); 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      divisor : IN STD_LOGIC_VECTOR (54 DOWNTO 1);

		quotient : OUT STD_LOGIC_VECTOR (55 DOWNTO 1)
		);
END dp_inv_core;

ARCHITECTURE rtl OF dp_inv_core IS

  --SII mullatency = doublespeed+5, SIII/IV mullatency = 4
  constant mullatency : positive := doublespeed+5 - device*(1+doublespeed);
  
  signal zerovec : STD_LOGIC_VECTOR (54 DOWNTO 1);
  
  signal divisordel : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal invdivisor : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal delinvdivisor : STD_LOGIC_VECTOR (18 DOWNTO 1);
  
  signal scaleden : STD_LOGIC_VECTOR (54 DOWNTO 1);
  
  signal twonode, subscaleden : STD_LOGIC_VECTOR (55 DOWNTO 1);
  signal guessone : STD_LOGIC_VECTOR (55 DOWNTO 1);
  signal guessonevec : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal absoluteval : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal absolutevalff, absoluteff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal abscarryff : STD_LOGIC;
  signal iteratenumnode : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal iteratenum : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal absoluteerror : STD_LOGIC_VECTOR (72 DOWNTO 1);
  signal mulabsguessff : STD_LOGIC_VECTOR (19 DOWNTO 1);
  signal mulabsguess : STD_LOGIC_VECTOR (54 DOWNTO 1);

  signal quotientnode : STD_LOGIC_VECTOR (72 DOWNTO 1);
  
  component fp_div_est IS 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        divisor : IN STD_LOGIC_VECTOR (19 DOWNTO 1);

		  invdivisor : OUT STD_LOGIC_VECTOR (18 DOWNTO 1)
		  );
  end component;
  
  component fp_fxmul IS 
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36;
           pipes : positive := 1;
           accuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1); 
      
        result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
       );
  end component;
  
  component dp_fxadd 
  GENERIC (
           width : positive := 64;
           pipes : positive := 1;
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
        carryin : IN STD_LOGIC;
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
  end component;
  
  component fp_del
  GENERIC (
           width : positive := 64;
           pipes : positive := 2
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
       
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
   end component;  
       
BEGIN
  
  gza: FOR k IN 1 TO 54 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  invcore: fp_div_est
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            divisor=>divisor(54 DOWNTO 36),invdivisor=>invdivisor);
  
  delinone: fp_del
  GENERIC MAP (width=>54,pipes=>5)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>divisor,cc=>divisordel);

  --**********************************
  --*** ITERATION 0 - SCALE INPUTS ***
  --**********************************
  
  -- in level 5, out level 8+speed
  mulscaleone: fp_fxmul
  GENERIC MAP (widthaa=>54,widthbb=>18,widthcc=>54,
               pipes=>3+doublespeed,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>divisordel,databb=>invdivisor,
            result=>scaleden);
              
  --********************
  --*** ITERATION 1  ***
  --********************

  twonode <= '1' & zerovec(54 DOWNTO 1);
  
  gta: FOR k IN 1 TO 54 GENERATE
    subscaleden(k) <= NOT(scaleden(k));
  END GENERATE;
  subscaleden(55) <= '1';
  
  -- in level 8+doublespeed, outlevel 9+2*doublespeed
  addtwoone: dp_fxadd 
  GENERIC MAP (width=>55,pipes=>doublespeed+1,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>twonode,bb=>subscaleden,carryin=>'1',
            cc=>guessone);  
            
  guessonevec <= guessone(54 DOWNTO 1);
  
  -- absolute value of guess lower 36 bits
  -- this is still correct, because (for positive), value will be 1.(17 zeros)error
  -- can also be calculated from guessonevec (code below)
  -- gabs: FOR k IN 1 TO 36 GENERATE
  --   absoluteval(k) <= guessonevec(k) XOR NOT(guessonevec(54));
  -- END GENERATE;
  gabs: FOR k IN 1 TO 36 GENERATE
    absoluteval(k) <= scaleden(k) XOR NOT(scaleden(54));
  END GENERATE;
  
  pta: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN

      FOR k IN 1 TO 36 LOOP
        absolutevalff(k) <= '0';
        absoluteff(k) <= '0';
      END LOOP;
      abscarryff <= '0';
      
    ELSIF (rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN
          
        absolutevalff <= absoluteval; -- out level 9+speed
        abscarryff <= NOT(scaleden(54)); 
        absoluteff <= absolutevalff + (zerovec(35 DOWNTO 1) & abscarryff); -- out level 10+speed
        
      END IF;
    
    END IF;
    
  END PROCESS;

  deloneone: fp_del
  GENERIC MAP (width=>18,pipes=>4+2*doublespeed)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>invdivisor,
            cc=>delinvdivisor);
 
  -- in level 9+2*doublespeed, out level 12+3*doublespeed
  muloneone: fp_fxmul
  GENERIC MAP (widthaa=>54,widthbb=>18,widthcc=>54,
               pipes=>3+doublespeed,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>guessonevec,databb=>delinvdivisor,
            result=>iteratenumnode);
 
  -- in level 10+doublespeed, out level 13+doublespeed
  mulonetwo: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>36,widthcc=>72,
               pipes=>3,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>absoluteff,databb=>absoluteff,
            result=>absoluteerror);
            
  -- if speed = 0, delay absoluteerror 1 clock, else 2
  -- this guess always positive (check??)
  -- change here, error can be [19:1], not [18:1] - this is because (1.[17 zeros].error)^2
  -- gives 1.[34 zeros].error 
  pgaa: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN

      FOR k IN 1 TO 19 LOOP
        mulabsguessff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN
        mulabsguessff <= absoluteerror(72 DOWNTO 54) + 
                        (zerovec(18 DOWNTO 1) & absoluteerror(53));
      END IF;
    
    END IF;
    
  END PROCESS;

  mulabsguess(19 DOWNTO 1) <= mulabsguessff;
  gmga: FOR k IN 20 TO 53 GENERATE
    mulabsguess(k) <= '0';
  END GENERATE;
  mulabsguess(54) <= '1';
  
  -- mulabsguess at 14+doublespeed depth
  -- iteratenum at 12+3*doublespeed depth
  
  -- mulabsguess 5 (5)clocks from absolutevalff
  -- iteratenum 3+2doublespeed (3/5)clocks from abssolutevalff
  -- delay iterate num 
  gdoa: IF (doublespeed = 0) GENERATE
    delonetwo: fp_del
    GENERIC MAP (width=>54,pipes=>2)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>iteratenumnode,
              cc=>iteratenum);
            
  END GENERATE;
  
  gdob: IF (doublespeed = 1) GENERATE
    iteratenum <= iteratenumnode;
  END GENERATE;
  
  --*********************
  --*** OUTPUT SCALE  ***
  --*********************
  
  -- in level 14+doublespeed
  -- SII out level 19+2*doublespeed
  -- SIII/IV out level 18+doublespeed
  mulout: fp_fxmul
  GENERIC MAP (widthaa=>54,widthbb=>54,widthcc=>72,pipes=>mullatency,
               accuracy=>doubleaccuracy,device=>device,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>iteratenum,databb=>mulabsguess,
            result=>quotientnode);
          
  quotient <= quotientnode(71 DOWNTO 17);
                  
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   DOUBLE PRECISION INVERSE SQUARE ROOT      ***
--***              TOP LEVEL                      ***
--***                                             ***
--***   DP_INVSQR.VHD                             ***
--***                                             ***
--***   Function: IEEE754 DP Inverse Square Root  ***
--***   (multiplicative iterative algorithm)      ***
--***                                             ***
--***   11/08/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--***                                             ***
--*** Stratix II                                  ***
--*** Latency = 32 + 2*Speed                      ***
--*** Speed = 0 : 32                              ***
--*** Speed = 1 : 34                              ***
--***                                             ***
--*** Stratix III/IV                              ***
--*** Latency = 31 + Speed                        ***
--*** Speed = 0 : 31                              ***
--*** Speed = 1 : 32                              ***
--***                                             ***
--*************************************************** 
    
ENTITY dp_invsqr IS 
GENERIC (
         doubleaccuracy : integer := 0;  -- 0 = pruned multiplier, 1 = normal multiplier
         doublespeed : integer := 0;  -- 0/1
         device : integer := 0;  -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
         synthesize : integer := 1  -- 0/1    
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin: IN STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (52 DOWNTO 1);

		  signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
      --------------------------------------------------
      nanout : OUT STD_LOGIC;
      invalidout : OUT STD_LOGIC
		);
END dp_invsqr;

ARCHITECTURE rtl OF dp_invsqr IS
  
  constant manwidth : positive := 52;
  constant expwidth : positive := 11;
  
  constant coredepth : positive := 31+2*doublespeed - device*(1+doublespeed);
  
  type expfftype IS ARRAY (coredepth+1 DOWNTO 1) OF STD_LOGIC_VECTOR (expwidth DOWNTO 1);

  signal maninff : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal expinff : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal signff : STD_LOGIC_VECTOR (coredepth+1 DOWNTO 1);
  signal correctff : STD_LOGIC_VECTOR (3 DOWNTO 1);  -- SPR 383712
  signal expff : expfftype;
  signal radicand : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal oddexponent : STD_LOGIC;
  signal invroot : STD_LOGIC_VECTOR (54 DOWNTO 1);
  --signal invroottest : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal manff : STD_LOGIC_VECTOR (manwidth DOWNTO 1); 
  signal zerovec : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal offset : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
    
  -- conditions
  signal nanmanff, nanexpff : STD_LOGIC_VECTOR (coredepth-1 DOWNTO 1);
  signal zeroexpff, zeromanff : STD_LOGIC_VECTOR (coredepth-2 DOWNTO 1); 
  signal expinzero, expinmax : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal maninzero : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal expzero, expmax, manzero : STD_LOGIC;
  signal infinityconditionff, nanconditionff, expzeroff : STD_LOGIC;
  signal correct_powers_of_two : STD_LOGIC;  -- SPR 383712
    
  component dp_invsqr_core IS 
  GENERIC (
           doublespeed : integer := 0;  -- 0/1
           doubleaccuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 1  -- 0/1      
          );         
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        radicand : IN STD_LOGIC_VECTOR (54 DOWNTO 1);
        odd : IN STD_LOGIC;

		  invroot : OUT STD_LOGIC_VECTOR (54 DOWNTO 1)
		  );
  end component;
	
BEGIN
    
  gzva: FOR k IN 1 TO manwidth GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  gxoa: FOR k IN 1 TO expwidth-1 GENERATE
    offset(k) <= '1';
  END GENERATE;
  offset(expwidth) <= '0';

  pma: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN

      FOR k IN 1 TO manwidth LOOP
        maninff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        expinff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO coredepth+1 LOOP
        signff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO coredepth+1 LOOP
        FOR j IN 1 TO expwidth LOOP
          expff(k)(j) <= '0';
        END LOOP;
      END LOOP;
      FOR k IN 1 TO manwidth LOOP
        manff(k) <= '0';
      END LOOP;
	  correctff <= "000";  -- SPR 383712
  
    ELSIF (rising_edge(sysclk)) THEN

      maninff <= mantissain;
      expinff <= exponentin;
    
      signff(1) <= signin;
      FOR k IN 2 TO coredepth+1 LOOP
        signff(k) <= signff(k-1);
      END LOOP;
  
      expff(1)(expwidth DOWNTO 1) <= exponentin;
      expff(2)(expwidth DOWNTO 1) <= expff(1)(expwidth DOWNTO 1) - offset;
      expff(3)(expwidth DOWNTO 1) <= expff(2)(expwidth) & expff(2)(expwidth DOWNTO 2);
      expff(4)(expwidth DOWNTO 1) <= offset - expff(3)(expwidth DOWNTO 1);
      expff(5)(expwidth DOWNTO 1) <= expff(4)(expwidth DOWNTO 1) - 1 + correctff(3);
      FOR k IN 6 TO coredepth LOOP
        expff(k)(expwidth DOWNTO 1) <= expff(k-1)(expwidth DOWNTO 1);
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        expff(coredepth+1)(k) <= (expff(coredepth)(k) AND zeroexpff(coredepth-2)) OR nanexpff(coredepth-2);
      END LOOP;

	  -- SPR 383712
	  correctff(1) <= correct_powers_of_two;
	  correctff(2) <= correctff(1);
	  correctff(3) <= correctff(2);
	  
      FOR k IN 1 TO manwidth LOOP
        manff(k) <= (invroot(k+1) AND zeromanff(coredepth-2)) OR nanmanff(coredepth-2);
      END LOOP;
  
    END IF;
  
  END PROCESS;

--*******************
--*** CONDITIONS ***
--*******************

  pcc: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
      
      FOR k IN 1 TO coredepth-1 LOOP
        nanmanff(k) <= '0';
        nanexpff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO coredepth-2 LOOP
        zeroexpff(k) <= '0';
        zeromanff(k) <= '0';
      END LOOP;
      infinityconditionff <= '0'; 
      nanconditionff <= '0';
      expzeroff <= '0';

    ELSIF (rising_edge(sysclk)) THEN
     
      infinityconditionff <= manzero AND expmax;
      nanconditionff <= signff(1) OR expzero OR (expmax AND manzero);
      expzeroff <= expzero;
 
      nanmanff(1) <= nanconditionff; -- level 3
      nanexpff(1) <= nanconditionff OR infinityconditionff; -- also max exp when infinity
      FOR k IN 2 TO coredepth-1 LOOP
        nanmanff(k) <= nanmanff(k-1);
        nanexpff(k) <= nanexpff(k-1);
      END LOOP;

      zeromanff(1) <= NOT(expzeroff) AND NOT(infinityconditionff); -- level 3
      zeroexpff(1) <= NOT(expzeroff); -- level 3
      FOR k IN 2 TO coredepth-2 LOOP
        zeromanff(k) <= zeromanff(k-1);
        zeroexpff(k) <= zeroexpff(k-1);
      END LOOP;
    
    END IF;
  
  END PROCESS;

--*******************
--*** SQUARE ROOT ***
--*******************
  
  radicand <= '1' & mantissain & '0';
  -- sub 1023, so 1023 (odd) = 2^0 => even
  oddexponent <= NOT(exponentin(1));

  -- does not require rounding, output of core rounded already, LSB always 0
  isqr: dp_invsqr_core
  GENERIC MAP (doublespeed=>doublespeed,doubleaccuracy=>doubleaccuracy,
               device=>device,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            radicand=>radicand,odd=>oddexponent,
            invroot=>invroot);

--*********************
--*** SPECIAL CASES ***
--*********************
-- 1. if negative input, invalid operation, NAN 
-- 2. 0 in, invalid operation, NAN
-- 3. infinity in, invalid operation, infinity out
-- 4. NAN in, invalid operation, NAN

  -- '1' if 0 
  expinzero(1) <= expinff(1);
  gxza: FOR k IN 2 TO expwidth GENERATE
    expinzero(k) <= expinzero(k-1) OR expinff(k);
  END GENERATE;
  expzero <= NOT(expinzero(expwidth)); -- '0' when zero
                 
  -- '1' if nan or infinity
  expinmax(1) <= expinff(1);
  gxia: FOR k IN 2 TO expwidth GENERATE
    expinmax(k) <= expinmax(k-1) AND expinff(k);
  END GENERATE;
  expmax <= expinmax(expwidth); -- '1' when true
          
  -- '1' if zero or infinity
  maninzero(1) <= maninff(1);
  gmza: FOR k IN 2 TO manwidth GENERATE
    maninzero(k) <= maninzero(k-1) OR maninff(k);
  END GENERATE;
  manzero <= NOT(maninzero(manwidth)); 
  -- 09/03/11 ML
  -- if mantissa is 0 and exponent is odd (...123,125,127,129,131...) then dont subtract 1 from offset corrected exponent
  -- '1' is subtracted as any value, no matter how small, in the mantissa will reduce the inverse below the mirrored exponent (around 127)
  -- if the exponent is odd (with mantissa 0) the value is a power of 2 (...0.25,0.5,1,2,4...) and the mirrored exponent is correct
  -- if the exponent is even (with mantissa 0), the inverse square root will have a non zero mantissa and can be handled normally
  correct_powers_of_two <= manzero AND expinff(1);  -- SPR 383712
       
--***************
--*** OUTPUTS ***
--***************

  signout <= signff(coredepth+1);
  exponentout <= expff(coredepth+1)(expwidth DOWNTO 1);   
  mantissaout <= manff;
  -----------------------------------------------
  nanout <= nanmanff(coredepth-1);
  invalidout <= nanmanff(coredepth-1);

END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   DOUBLE PRECISION INVERSE SQUARE ROOT      ***
--***                 CORE                        ***
--***                                             ***
--***   DP_INVSQR_CORE.VHD                        ***
--***                                             ***
--***   Function: 54 bit Inverse Square Root      ***
--***   (multiplicative iterative algorithm)      ***
--***                                             ***
--***   09/12/07 ML                               ***
--***                                             ***
--***   (c) 2007 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***   24/04/09 - SIII/SIV multiplier support    ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** SII Latency = 31 + 2*doublespeed            ***
--*** SIII/IV Latency = 30 + doublespeed          ***
--*** 1. Output is rounded already, LSB always 0  ***
--***************************************************

ENTITY dp_invsqr_core IS 
GENERIC (
         doublespeed : integer := 0;  -- 0/1
         doubleaccuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
         device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
         synthesize : integer := 1  -- 0/1      
        ); 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      radicand : IN STD_LOGIC_VECTOR (54 DOWNTO 1);
      odd : IN STD_LOGIC;

		invroot : OUT STD_LOGIC_VECTOR (54 DOWNTO 1)
		);
END dp_invsqr_core;

ARCHITECTURE rtl OF dp_invsqr_core IS

  --SII mullatency = speed+5, SIII/IV mullatency = 4
  constant mullatency : positive := doublespeed+5 - device*(1+doublespeed);
    
  signal zerovec : STD_LOGIC_VECTOR (54 DOWNTO 1);
  
  signal evennum : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal oddnum : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal guessvec : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal oddff : STD_LOGIC_VECTOR (25+doublespeed DOWNTO 1);
  signal scalenumff : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal guess : STD_LOGIC_VECTOR (18 DOWNTO 1);

  -- 1st iteration
  signal radicanddelone : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal guessdel : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal multoneone : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal multonetwo : STD_LOGIC_VECTOR (37 DOWNTO 1);
  signal multonetwoff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal suboneff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal multonethr : STD_LOGIC_VECTOR (37 DOWNTO 1);
  signal guessonevec : STD_LOGIC_VECTOR (36 DOWNTO 1);
      
  -- 2ns iteration
  signal radicanddeltwo : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal guessonevecdelone : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal guessonevecdeltwo : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal multtwoone : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal multtwotwo : STD_LOGIC_VECTOR (72 DOWNTO 1);
  signal multtwotwoff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal finaladdsub : STD_LOGIC;
  signal finaladdsubff : STD_LOGIC_VECTOR (4 DOWNTO 1);
  signal finaladdff : STD_LOGIC_VECTOR (55 DOWNTO 1);
  signal multtwothr : STD_LOGIC_VECTOR (36 DOWNTO 1);  
  signal finalguessvec : STD_LOGIC_VECTOR (53 DOWNTO 1);
  signal invrootvec : STD_LOGIC_VECTOR (53 DOWNTO 1);

  component fp_invsqr_est IS 
  GENERIC (synthesize : integer := 0); -- 0 = behavioral, 1 = syntheziable
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        radicand : IN STD_LOGIC_VECTOR (19 DOWNTO 1);

		  invroot : OUT STD_LOGIC_VECTOR (18 DOWNTO 1)
		  );
  end component;
  
  component dp_fxadd IS 
  GENERIC (
           width : positive := 64;
           pipes : positive := 1;
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
        carryin : IN STD_LOGIC;
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       ); 
  end component;
  
  component fp_fxmul IS 
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36;
           pipes : positive := 1;
           accuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 0
        );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1); 
      
        result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
       ); 
  end component;
 
  component fp_del 
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
   end component;
   		 
BEGIN
    
  oddnum <= conv_std_logic_vector(185363,18); -- mult by 2^-.5 (odd exp)
  evennum <= conv_std_logic_vector(262143,18); -- mult by 1 (even exp)
  
  gza: FOR k IN 1 TO 54 GENERATE
    zerovec(k) <= '0';
  END GENERATE;

  -- in level 0, out level 5
  look: fp_invsqr_est
  GENERIC MAP (synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            radicand=>radicand(54 DOWNTO 36),invroot=>guessvec);
              
  pta: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN
    
      FOR k IN 1 TO 25+doublespeed LOOP
        oddff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 18 LOOP
        scalenumff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF (enable = '1') THEN
        
        oddff(1) <= odd;
        FOR k IN 2 TO 25+doublespeed LOOP
          oddff(k) <= oddff(k-1);
        END LOOP; 
        
        FOR k IN 1 TO 18 LOOP
          scalenumff(k) <= (oddnum(k) AND oddff(4)) OR (evennum(k) AND NOT(oddff(4)));
        END LOOP;
          
      END IF;
    
    END IF;    
      
  END PROCESS;

  -- in level 5, out level 7
  mulscale: fp_fxmul
  GENERIC MAP (widthaa=>18,widthbb=>18,widthcc=>18,pipes=>2,
               device=>device,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>guessvec,databb=>scalenumff,
            result=>guess);

  --*********************
  --*** ITERATION ONE ***
  --*********************
  --X' = X/2(3-YXX)
  
  deloneone: fp_del
  GENERIC MAP(width=>54,pipes=>9)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>radicand,cc=>radicanddelone);
            
  delonetwo: fp_del
  GENERIC MAP(width=>18,pipes=>7)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>guess,cc=>guessdel);
            
  -- in level 7, out level 9 (18x18=36)
  oneone: fp_fxmul
  GENERIC MAP (widthaa=>18,widthbb=>18,widthcc=>36,pipes=>2,
               device=>device,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>guess,databb=>guess,
            result=>multoneone);
                   
  -- in level 9, out level 12 (36x36=37)
  onetwo: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>36,widthcc=>37,pipes=>3,
               device=>device,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>radicanddelone(54 DOWNTO 19),databb=>multoneone,
            result=>multonetwo);
                   
  -- multonetwo is about 1 - either 1.000000XXX or 0.9999999
  -- mult by 2 if odd exponent (37 DOWNTO 2), otherwise (38 DOWNTO 3)
  -- round bit in position 1 or 2
  pone: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN

      FOR k IN 1 TO 36 LOOP
        multonetwoff(k) <= '0';
        suboneff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF (enable = '1') THEN
        
        --invert here so that borrow can be added in simple expression
        -- level 13
        FOR k IN 1 TO 36 LOOP
          multonetwoff(k) <= NOT((multonetwo(k) AND oddff(12)) OR (multonetwo(k+1) AND NOT(oddff(12))));
        END LOOP;
        -- level 14
        suboneff <= ("11" & zerovec(34 DOWNTO 1)) + 
                    ('1' & multonetwoff(36 DOWNTO 2)) +
                    (zerovec(35 DOWNTO 1) & multonetwoff(1));
          
      END IF;
    
    END IF;    
      
  END PROCESS;    

  -- in level 14, out level 17 (36x18=37)
  onethr: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>18,widthcc=>37,pipes=>3,
               device=>device,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>suboneff,databb=>guessdel,
            result=>multonethr); 
            
  -- mult by 2 - subone is about 1 (1.000 or 0.9999) so will effectively multiply by 0.5
  guessonevec <= multonethr(36 DOWNTO 1);
  
  --************************
  --*** SECOND ITERATION ***
  --************************
  --X' = X/2(3-YXX)
  
  deltwoone: fp_del
  GENERIC MAP(width=>54,pipes=>11)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>radicanddelone,cc=>radicanddeltwo);
            
  -- SII level in 17, level out 26+doublespeed
  -- SIII/IV level in 17, level out 25
  deltwotwo: fp_del
  GENERIC MAP(width=>36,pipes=>(9+doublespeed-device*(1+doublespeed)))
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>guessonevec,cc=>guessonevecdelone);
            
  deltwothr: fp_del
  GENERIC MAP (width=>36,pipes=>4)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>guessonevecdelone,cc=>guessonevecdeltwo);
            
  -- in level 17, out level 20 (36x36=54)
  twoone: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>36,widthcc=>54,pipes=>3,
               accuracy=>doubleaccuracy,device=>device,
               synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>guessonevec,databb=>guessonevec,
            result=>multtwoone); 
            
  -- in level 20, 
  -- SII out level 25/26 - 25+doublespeed
  -- SIII/SIV out level 24   
  twotwo: fp_fxmul
  GENERIC MAP (widthaa=>54,widthbb=>54,widthcc=>72,pipes=>mullatency,
               accuracy=>doubleaccuracy,device=>device,
               synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>multtwoone,databb=>radicanddeltwo,
            result=>multtwotwo); 

  -- multtwotwo is about 1 - either 1.000000XXX or 0.9999999
  -- mult by 2 if odd exponent (55 DOWNTO 2), otherwise (56 DOWNTO 3)
  -- round bit in position 1 or 2
  ptwo: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN

      FOR k IN 1 TO 36 LOOP
        multtwotwoff(k) <= '0';
      END LOOP;
      finaladdsubff <= "0000";
      FOR k IN 1 TO 55 LOOP
        finaladdff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF (enable = '1') THEN
        
        -- SII in level 25+doublespeed, out level 26+doublespeed
        -- SIII in level 24, out level 25
        -- if multwotwo > 1, subtwo negative, subtract multwothr from guessonevec
        -- if multwotwo <= 1, subtwo positive, add multwothr to guessonevec
        FOR k IN 1 TO 36 LOOP
          multtwotwoff(k) <= ((multtwotwo(k+6) AND oddff(25+doublespeed-device*(1+doublespeed))) OR 
                              (multtwotwo(k+7) AND NOT(oddff(25+doublespeed-device*(1+doublespeed))))) XOR finaladdsub;
        END LOOP;
        
        finaladdsubff(1) <= finaladdsub;
        FOR k IN 2 TO 4 LOOP
          finaladdsubff(k) <= finaladdsubff(k-1);
        END LOOP;

        -- makes sure no overflow happens here, for example if less than 30 leading 1s/0s
        -- in multtwotwoff
        -- SII level in 29+doublespeed level out 30+doublespeed
        -- SIII level in 28 level out 29
        FOR k IN 1 TO 26 LOOP
          finaladdff(k) <= multtwothr(k+10) XOR NOT(finaladdsubff(4));
        END LOOP;
        FOR k IN 27 TO 55 LOOP
          finaladdff(k) <= NOT(finaladdsubff(4));
        END LOOP;
          
      END IF;
    
    END IF;    
      
  END PROCESS;  
  
  -- doesnt have to be near msb
  finaladdsub <= multtwotwo(60);  

  -- SII level in (26+doublespeed), level out (29+doublespeed)
  -- SII level in 25, level out 28
  twothr: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>36,widthcc=>36,pipes=>3,
               device=>device,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>multtwotwoff,databb=>guessonevecdelone,
            result=>multtwothr);
                      
  finalguessvec <= guessonevecdeltwo & zerovec(17 DOWNTO 1);
   
  -- SII level in 30+doublespeed, level out 31+2*doublespeed
  -- SIII level in 29, level out 30+doublespeed
  final: dp_fxadd
  GENERIC MAP (width=>53,pipes=>doublespeed+1,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>finalguessvec,bb=>finaladdff(55 DOWNTO 3),carryin=>finaladdff(2),
            cc=>invrootvec);
  
  invroot <= invrootvec & '0';
   
END rtl;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   ALTERA FLOATING POINT DATAPATH COMPILER   ***
--***                                             ***
--***   DP_LDEXP.VHD                              ***
--***                                             ***
--***   Function: Single Precision Load Exponent  ***
--***                                             ***
--***   ldexp(x,n) - x*2^n - IEEE in and out      ***
--***                                             ***
--***   Created 12/09/09                          ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_ldexp IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (52 DOWNTO 1);
      bb : IN STD_LOGIC_VECTOR (32 DOWNTO 1);
      
		  signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
		  satout, zeroout, nanout : OUT STD_LOGIC
		);
END dp_ldexp;

ARCHITECTURE rtl OF dp_ldexp IS
 
  signal signinff : STD_LOGIC;
  signal exponentinff : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal mantissainff : STD_LOGIC_VECTOR (52 DOWNTO 1);
  signal bbff : STD_LOGIC_VECTOR (13 DOWNTO 1);
  signal signoutff : STD_LOGIC;
  signal exponentoutff : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal mantissaoutff : STD_LOGIC_VECTOR (52 DOWNTO 1);
  signal satoutff, zerooutff, nanoutff : STD_LOGIC;
  signal satnode, zeronode, nannode : STD_LOGIC;
  signal expnode : STD_LOGIC_VECTOR (13 DOWNTO 1);
  signal expzeroin, expmaxin : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal expzeronode, expmaxnode : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal expzeroout, expmaxout : STD_LOGIC;
  signal manzeroin : STD_LOGIC_VECTOR (52 DOWNTO 1);
  signal manzero, mannonzero : STD_LOGIC; 

BEGIN
    
  pin: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
    
      signinff <= '0';
      signoutff <= '0';
      FOR k IN 1 TO 11 LOOP
        exponentinff(k) <= '0';
        exponentoutff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 52 LOOP
        mantissainff(k) <= '0';
        mantissaoutff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 13 LOOP
        bbff(k) <= '0';
      END LOOP;
      satoutff <= '0';
      zerooutff <= '0';
      nanoutff <= '0';
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF (enable = '1') THEN

      
        signinff <= signin;
        exponentinff <= exponentin;
        mantissainff <= mantissain;
        
        bbff <= bb(13 DOWNTO 1);
        
        signoutff <= signinff;
        FOR k IN 1 TO 11 LOOP
          exponentoutff(k) <= (expnode(k) AND NOT(zeronode)) OR satnode OR nannode;
        END LOOP;
        FOR k IN 1 TO 52 LOOP
          mantissaoutff(k) <= (mantissainff(k) AND NOT(zeronode) AND NOT(satnode)) OR nannode;
        END LOOP;
        
        satoutff <= satnode;
        zerooutff <= zeronode;
        nanoutff <= nannode;
        
      END IF;
    
    END IF;  
      
  END PROCESS;
  
  expnode <= ("00" & exponentinff) + bbff;
  
  expzeroin(1) <= exponentinff(1);
  expmaxin(1) <= exponentinff(1);
  gxa: FOR k IN 2 TO 11 GENERATE
    expzeroin(k) <= expzeroin(k-1) OR exponentinff(k);
    expmaxin(k) <= expmaxin(k-1) AND exponentinff(k);
  END GENERATE;
  
  expzeronode(1) <= expnode(1);
  expmaxnode(1) <= expnode(1);
  gxb: FOR k IN 2 TO 11 GENERATE
    expzeronode(k) <= expzeronode(k-1) OR expnode(k);
    expmaxnode(k) <= expmaxnode(k-1) AND expnode(k);
  END GENERATE;
  expzeroout <= NOT(expzeroin(11)) OR (NOT(expzeronode(11)) AND NOT(expnode(12))) OR (expnode(13));
  expmaxout <= expmaxin(11) OR (expmaxnode(11) AND NOT(expnode(12))) OR (expnode(12) AND NOT(expnode(13))); 
  
  manzeroin(1) <= mantissainff(1);
  gma: FOR k IN 2 TO 52 GENERATE
    manzeroin(k) <= manzeroin(k-1) OR mantissainff(k);
  END GENERATE;
  manzero <= NOT(manzeroin(52));
  mannonzero <= manzeroin(52);
  
  satnode <= (expmaxin(11) AND NOT(manzeroin(52))) OR expmaxout;
  zeronode <= NOT(expzeroin(11)) OR expzeroout;
  nannode <= expmaxin(11) AND manzeroin(52);
  
	signout <= signoutff;
  exponentout <= exponentoutff;
  mantissaout <= mantissaoutff;
      
  satout <= satoutff;
  zeroout <= zerooutff;
  nanout <= nanoutff;

END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   DOUBLE PRECISION LOG(e) - CORE            ***
--***                                             ***
--***   DP_LN_CORE.VHD                            ***
--***                                             ***
--***   Function: Double Precision LOG (LN) Core  ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***   24/04/09 - SIII/SIV multiplier support    ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** SII/SIII/SIV Latency = 26 + 7*doublespeed   ***
--*** no 54x54 multipliers                        ***
--***************************************************

ENTITY dp_ln_core IS 
GENERIC (
         doublespeed : integer := 0; -- 0/1
         device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
         synthesize : integer := 1 -- 0/1       
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      aaman : IN STD_LOGIC_VECTOR (52 DOWNTO 1); 
      aaexp : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
      
      ccman : OUT STD_LOGIC_VECTOR (53 DOWNTO 1);
      ccexp : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
      ccsgn : OUT STD_LOGIC;
      zeroout : OUT STD_LOGIC
     );
END dp_ln_core;

ARCHITECTURE rtl OF dp_ln_core IS

  signal zerovec : STD_LOGIC_VECTOR (64 DOWNTO 1);
  --*** INPUT BLOCK ***
  signal aamanff : STD_LOGIC_VECTOR (52 DOWNTO 1);
  signal aaexpff : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal aaexpabsff : STD_LOGIC_VECTOR (10 DOWNTO 1);
  signal aaexppos, aaexpneg : STD_LOGIC_VECTOR (12 DOWNTO 1);
  signal aaexpabs : STD_LOGIC_VECTOR (10 DOWNTO 1);
  --*** TABLES ***
  signal lutpowaddff : STD_LOGIC_VECTOR (10 DOWNTO 1);
  signal lutoneaddff, luttwoaddff : STD_LOGIC_VECTOR (9 DOWNTO 1);
  signal lutpowmanff, lutonemanff, luttwomanff : STD_LOGIC_VECTOR (52 DOWNTO 1);
  signal lutpowexpff, lutoneexpff, luttwoexpff : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal lutoneinvff : STD_LOGIC_VECTOR (12 DOWNTO 1); 
  signal luttwoinvff : STD_LOGIC_VECTOR (18 DOWNTO 1);  
  signal lutpowmannode, lutonemannode, luttwomannode : STD_LOGIC_VECTOR (52 DOWNTO 1);
  signal lutpowexpnode, lutoneexpnode, luttwoexpnode : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal lutoneinvnode : STD_LOGIC_VECTOR (12 DOWNTO 1); 
  signal luttwoinvnode : STD_LOGIC_VECTOR (18 DOWNTO 1);   
  signal aanum, aanumdel : STD_LOGIC_VECTOR (54 DOWNTO 1); 
  signal invonenum : STD_LOGIC_VECTOR (18 DOWNTO 1); 
  signal mulonenode : STD_LOGIC_VECTOR (65 DOWNTO 1);
  signal mulonenormff : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal mulonenumdel : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal multwonode : STD_LOGIC_VECTOR (72 DOWNTO 1); 
  signal multwonormff : STD_LOGIC_VECTOR (71 DOWNTO 1);
  --*** SERIES ***
  signal squaredterm : STD_LOGIC_VECTOR (48 DOWNTO 1);
  signal onethird : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal scaledterm, scaledtermdel : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal cubedterm : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal xtermdel : STD_LOGIC_VECTOR (54 DOWNTO 1);   
  signal oneterm, twoterm, thrterm : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal oneplustwoterm : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal seriesterm : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal mantissaseries : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal exponentseries : STD_LOGIC_VECTOR (11 DOWNTO 1);          
  --*** ADD LOGS ***
  signal zeropow, zeroone, zerotwo : STD_LOGIC;
  signal mantissapowernode : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal mantissapower : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal exponentpower : STD_LOGIC_VECTOR (11 DOWNTO 1); 
  signal numberone, numberonedel : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal mantissaone : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal exponentone : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal mantissaaddone : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal exponentaddone : STD_LOGIC_VECTOR (11 DOWNTO 1); 
  signal mantissatwo : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal exponenttwo : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal numbertwo, numbertwodel : STD_LOGIC_VECTOR (75 DOWNTO 1);
  signal mantissaaddtwo : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal exponentaddtwo : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal numberthr, numberthrdel : STD_LOGIC_VECTOR (75 DOWNTO 1);
  signal mantissasum : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal mantissasumabs : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal exponentsum : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal mantissanorm : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal exponentnorm : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal zeronorm : STD_LOGIC;
  signal signff : STD_LOGIC_VECTOR (25+7*doublespeed DOWNTO 1);
  
  component dp_lnlutpow
  PORT (
        add : IN STD_LOGIC_VECTOR (10 DOWNTO 1);
        logman : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
        logexp : OUT STD_LOGIC_VECTOR (11 DOWNTO 1)
       );
  end component;
  
  component dp_lnlut9
  PORT (
        add : IN STD_LOGIC_VECTOR (9 DOWNTO 1);
        inv : OUT STD_LOGIC_VECTOR (12 DOWNTO 1);
        logman : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
        logexp : OUT STD_LOGIC_VECTOR (11 DOWNTO 1)
       );
  end component;

  component dp_lnlut18
  PORT (
        add : IN STD_LOGIC_VECTOR (9 DOWNTO 1);
        inv : OUT STD_LOGIC_VECTOR (18 DOWNTO 1);
        logman : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
        logexp : OUT STD_LOGIC_VECTOR (11 DOWNTO 1)
       );
  end component;
  
  component fp_del
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
  end component;
  
  component dp_fxadd 
  GENERIC (
           width : positive := 64;
           pipes : positive := 1;
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
        carryin : IN STD_LOGIC;
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
  end component;
  
  component dp_fxsub
  GENERIC (
           width : positive := 64;
           pipes : positive := 1;
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
        borrowin : IN STD_LOGIC;
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
  end component;
 
  component fp_fxmul
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36;
           pipes : positive := 1;
           accuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1); 
      
        result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
       );
  end component;
   
  component dp_lnadd
  GENERIC (
           speed : integer := 1; -- '0' for unpiped adder, '1' for piped adder
           synthesize : integer := 1
          ); 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aaman : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
        aaexp : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
        bbman : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
        bbexp : IN STD_LOGIC_VECTOR (11 DOWNTO 1);

	     ccman : OUT STD_LOGIC_VECTOR (64 DOWNTO 1);
	     ccexp : OUT STD_LOGIC_VECTOR (11 DOWNTO 1)
	   );
	end component;
	
  component dp_lnnorm
  GENERIC (
           speed : integer := 1
          ); 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        inman : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
        inexp : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
      
        outman : OUT STD_LOGIC_VECTOR (64 DOWNTO 1);
        outexp : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
        zero : OUT STD_LOGIC
      );	
  end component;
                  
BEGIN
  
  gza: FOR k IN 1 TO 64 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  --*******************
  --*** INPUT BLOCK ***
  --*******************
  
  ppin: PROCESS (sysclk,reset)
  BEGIN
  
    IF (reset = '1') THEN
        
      FOR k IN 1 TO 52 LOOP
        aamanff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 11 LOOP
        aaexpff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 10 LOOP
        aaexpabsff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
     
      IF (enable = '1') THEN       
      
        aamanff <= aaman;  -- level 1
        aaexpff <= aaexp;  -- level 1
      
        aaexpabsff <= aaexpabs;  -- level 2
      
      END IF;
 
    END IF;
    
  END PROCESS;
  
  aaexppos <= ('0' & aaexpff) - "001111111111";
  aaexpneg <= "001111111111" - ('0' & aaexpff);
  gaba: FOR k IN 1 TO 10 GENERATE
    aaexpabs(k) <= (aaexppos(k) AND NOT(aaexppos(12))) OR (aaexpneg(k) AND aaexppos(12));
  END GENERATE;

  --******************************************
  --*** RANGE REDUCTION THROUGH LUT SERIES ***
  --******************************************
    
  plut: PROCESS (sysclk,reset)
  BEGIN
  
    IF (reset = '1') THEN
       
      FOR k IN 1 TO 10 LOOP 
        lutpowaddff(k) <= '0'; 
      END LOOP;
      FOR k IN 1 TO 9 LOOP
        lutoneaddff(k) <= '0';
        luttwoaddff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 52 LOOP
        lutpowmanff(k) <= '0';
        lutonemanff(k) <= '0';
        luttwomanff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 11 LOOP
        lutpowexpff(k) <= '0';
        lutoneexpff(k) <= '0';
        luttwoexpff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 12 LOOP
        lutoneinvff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 18 LOOP
        luttwoinvff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
            
      IF (enable = '1') THEN
          
        lutpowaddff <= aaexpabsff;  -- level 3
        lutoneaddff <= aamanff(52 DOWNTO 44);  -- level 2
        luttwoaddff <= mulonenormff(55 DOWNTO 47);  -- level 8+speed
      
        lutpowmanff <= lutpowmannode;  -- level 4
        lutpowexpff <= lutpowexpnode; -- level 4
      
        lutoneinvff <= lutoneinvnode;  -- level 3
        lutonemanff <= lutonemannode;  -- level 3
        lutoneexpff <= lutoneexpnode; -- level 3
      
        luttwoinvff <= luttwoinvnode;  -- level 9+speed
        luttwomanff <= luttwomannode;  -- level 9+speed
        luttwoexpff <= luttwoexpnode; -- level 9+speed
      
      END IF;
      
    END IF;
    
  END PROCESS;
  
  lutpow: dp_lnlutpow
  PORT MAP (add=>lutpowaddff,
            logman=>lutpowmannode,logexp=>lutpowexpnode);

  lutone: dp_lnlut9
  PORT MAP (add=>lutoneaddff,
            inv=>lutoneinvnode,logman=>lutonemannode,logexp=>lutoneexpnode);
 
  luttwo: dp_lnlut18
  PORT MAP (add=>luttwoaddff,
            inv=>luttwoinvnode,logman=>luttwomannode,logexp=>luttwoexpnode);
           
  aanum <= '1' & aamanff & '0'; 
  
  -- level 1 in, level 3 out
  delone: fp_del
  GENERIC MAP (width=>54,pipes=>2)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>aanum,cc=>aanumdel);
   
  invonenum <= lutoneinvff & "000000";
  
  --mulone <= aanum * invone; -- 53*12 = 65
  
  -- level 3 in, level 6+doublespeed out
  mulone: fp_fxmul
  GENERIC MAP (widthaa=>54,widthbb=>18,widthcc=>65,
               pipes=>3+doublespeed,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>aanumdel,databb=>invonenum,
            result=>mulonenode);

  --multwo <= mulonenorm(64 DOWNTO 11) * invtwo;  -- 54x18=72
  
  -- level 7+speed in, level 9+speed out
  deltwo: fp_del
  GENERIC MAP (width=>54,pipes=>2)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>mulonenormff(64 DOWNTO 11),cc=>mulonenumdel);
  
  -- level 9+doublespeed in, level 12+2*doublespeed out
  multwo: fp_fxmul
  GENERIC MAP (widthaa=>54,widthbb=>18,widthcc=>72,
               pipes=>3+doublespeed,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>mulonenumdel,databb=>luttwoinvff,
            result=>multwonode);

  pmna: PROCESS (sysclk,reset)
  BEGIN
  
    IF (reset = '1') THEN
        
      FOR k IN 1 TO 64 LOOP
        mulonenormff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 71 LOOP
        multwonormff(k) <= '0';
      END LOOP;
   
    ELSIF (rising_edge(sysclk)) THEN
     
      IF (enable = '1') THEN
        
        -- normalize in case input is 1.000000 and inv is 0.5  
        -- level 7+speed
        FOR k IN 1 TO 64 LOOP
          mulonenormff(k) <= (mulonenode(k+1) AND mulonenode(65)) OR 
                             (mulonenode(k) AND NOT(mulonenode(65)));
        END LOOP;
        -- level 13+2*speed
        FOR k IN 1 TO 71 LOOP
          multwonormff(k) <= (multwonode(k+1) AND multwonode(72)) OR 
                             (multwonode(k) AND NOT(multwonode(72)));
        END LOOP;
         
      END IF;       
    END IF;
    
  END PROCESS;  
           
  --************************************
  --*** TAYLOR SERIES OF SMALL RANGE ***
  --************************************
  
  -- taylor series expansion of subrange (36 bits)
  -- x - x*x/2
  -- 16 leading bits, so x*x 16 bits down, +1 bit for 1/2
  -- 36 lower bits in multwo(54:19)
  
  --square <= multwonorm(54 DOWNTO 19) * multwonorm(54 DOWNTO 19);
  
  -- level 13+2*doublespeed in, 16+2*doublespeed out
  multhr: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>36,widthcc=>48,
               pipes=>3,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>multwonormff(54 DOWNTO 19),databb=>multwonormff(54 DOWNTO 19),
            result=>squaredterm);
  
  onethird <= "010101010101010101";
            
  -- level 13+2*doublespeed in, level 15+2*doublespeed out
  mulfor: fp_fxmul
  GENERIC MAP (widthaa=>18,widthbb=>18,widthcc=>18,
               pipes=>2,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>multwonormff(54 DOWNTO 37),databb=>onethird,
            result=>scaledterm);
  
  --level 15+2*doublespeed in, level 16+2*doublespeed out
  delthr: fp_del
  GENERIC MAP (width=>18,pipes=>1)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>scaledterm,cc=>scaledtermdel);
            
  -- level 16+2*doublespeed in, level 18+2*doublespeed out
  mulfiv: fp_fxmul
  GENERIC MAP (widthaa=>18,widthbb=>18,widthcc=>32,
               pipes=>2,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>squaredterm(48 DOWNTO 31),databb=>scaledtermdel,
            result=>cubedterm);
            
  --level 13+2*doublespeed in, level 16+2*doublespeed out
  delfor: fp_del
  GENERIC MAP (width=>54,pipes=>3)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>multwonormff(54 DOWNTO 1),cc=>xtermdel); 
   
  -- level 16+2*doublespeed         
  oneterm <= xtermdel & zerovec(10 DOWNTO 1);
  twoterm <= zerovec(17 DOWNTO 1) & squaredterm(48 DOWNTO 2); -- x*x/2
  -- level 18+2*doublespeed
  thrterm <= zerovec(32 DOWNTO 1) & cubedterm;
  
  --level 16+2*doublespeed in, level 18+2*doublespeed out
  tayone: dp_fxsub
  GENERIC MAP (width=>64,pipes=>2,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>oneterm,bb=>twoterm,borrowin=>'1',
            cc=>oneplustwoterm); 
  
  --level 18+2*doublespeed in, level 19+3*doublespeed out
  taytwo: dp_fxadd
  GENERIC MAP (width=>64,pipes=>1+doublespeed,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>oneplustwoterm,bb=>thrterm,carryin=>'0',
            cc=>seriesterm); 
            
  --mantissaseries <= seriesterm;
  mantissaseries <= '0' & seriesterm(64 DOWNTO 2);
  exponentseries <= conv_std_logic_vector (1006,11); 
            
  --18x18
  --cubed <= square(72 DOWNTO 55) * multwonorm(54 DOWNTO 37);
  --cubedscale <= cubed(36 DOWNTO 19) * onethird;
  
  --**************************
  --*** ADD ALL LOGARITHMS ***
  --**************************
  
  zeropow <= lutpowexpff(11) OR lutpowexpff(10) OR lutpowexpff(9) OR 
             lutpowexpff(8) OR lutpowexpff(7) OR lutpowexpff(6) OR 
             lutpowexpff(5) OR lutpowexpff(4) OR lutpowexpff(3) OR 
             lutpowexpff(2) OR lutpowexpff(1);
             
  -- level 4
  --mantissapower <= zeropow & lutpowmanff & zerovec(11 DOWNTO 1);
  --mantissapower <= '0' & zeropow & lutpowmanff & zerovec(10 DOWNTO 1);
  mantissapowernode <= '0' & zeropow & lutpowmanff & zerovec(10 DOWNTO 1);
  gmpz: FOR k IN 1 TO 64 GENERATE
    mantissapower(k) <= mantissapowernode(k) XOR signff(3);
  END GENERATE;
  exponentpower <= lutpowexpff;
  
  zeroone <= lutoneexpff(11) OR lutoneexpff(10) OR lutoneexpff(9) OR 
             lutoneexpff(8) OR lutoneexpff(7) OR lutoneexpff(6) OR 
             lutoneexpff(5) OR lutoneexpff(4) OR lutoneexpff(3) OR 
             lutoneexpff(2) OR lutoneexpff(1);
             
  -- level 3
  numberone <= zeroone & lutonemanff & lutoneexpff;
  
  -- level 3 in, level 4 out
  delfiv: fp_del
  GENERIC MAP (width=>64,pipes=>1)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>numberone,cc=>numberonedel);
            
  --mantissaone <= numberonedel(64 DOWNTO 12) & zerovec(11 DOWNTO 1);
  mantissaone <= '0' & numberonedel(64 DOWNTO 12) & zerovec(10 DOWNTO 1);
  exponentone <= numberonedel(11 DOWNTO 1); 
  
  -- level 4 in, level 10 out
  addone: dp_lnadd
  GENERIC MAP (speed=>1,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aaman=>mantissapower,aaexp=>exponentpower,
            bbman=>mantissaone,bbexp=>exponentone,
            ccman=>mantissaaddone,ccexp=>exponentaddone);
           
  zerotwo <= luttwoexpff(11) OR luttwoexpff(10) OR luttwoexpff(9) OR 
             luttwoexpff(8) OR luttwoexpff(7) OR luttwoexpff(6) OR 
             luttwoexpff(5) OR luttwoexpff(4) OR luttwoexpff(3) OR 
             luttwoexpff(2) OR luttwoexpff(1);
             
  -- level 9+doublespeed
  --mantissatwo <= zerotwo & luttwomanff & zerovec(11 DOWNTO 1);
  mantissatwo <= '0' & zerotwo & luttwomanff & zerovec(10 DOWNTO 1);
  exponenttwo <= luttwoexpff;

  numbertwo <= mantissatwo & exponenttwo;
    
  gasa: IF (doublespeed = 0) GENERATE
    delsix: fp_del
    GENERIC MAP (width=>75,pipes=>1)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>numbertwo,cc=>numbertwodel);
  END GENERATE;
  gasb: IF (doublespeed = 1) GENERATE
    numbertwodel <= numbertwo;
  END GENERATE;

  -- level 10 in, level 16 out
  addtwo: dp_lnadd
  GENERIC MAP (speed=>1,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aaman=>mantissaaddone,aaexp=>exponentaddone,
            bbman=>numbertwodel(75 DOWNTO 12),bbexp=>numbertwodel(11 DOWNTO 1),
            ccman=>mantissaaddtwo,ccexp=>exponentaddtwo);
            
  numberthr <= mantissaaddtwo & exponentaddtwo;

  -- level 16 in, level 19+3*doublespeed out
  delsev: fp_del
  GENERIC MAP (width=>75,pipes=>3+3*doublespeed)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>numberthr,cc=>numberthrdel);
              
  -- level 19+3*doublespeed in, level 23+5*doublespeed out
  addthr: dp_lnadd
  GENERIC MAP (speed=>doublespeed,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aaman=>mantissaseries,aaexp=>exponentseries,
            bbman=>numberthrdel(75 DOWNTO 12),bbexp=>numberthrdel(11 DOWNTO 1),
            ccman=>mantissasum,ccexp=>exponentsum);            

  gmsa: FOR k IN 1 TO 64 GENERATE
    mantissasumabs(k) <= mantissasum(k) XOR signff(22+5*doublespeed);
  END GENERATE;
  
  -- level 23+5*doublespeed in, level 26+7*doublespeed out
  norm: dp_lnnorm
  GENERIC MAP (speed=>doublespeed)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            inman=>mantissasumabs,inexp=>exponentsum,
            outman=>mantissanorm,outexp=>exponentnorm,
            zero=>zeronorm);
  
  psgna: PROCESS (sysclk, reset)
  BEGIN
      
    IF (reset = '1') THEN
      FOR k IN 1 TO 25+7*doublespeed LOOP
        signff(k) <= '0';
      END LOOP;
    ELSIF (rising_edge(sysclk)) THEN
      signff(1) <= aaexppos(12);
      FOR k IN 2 TO 25+7*doublespeed LOOP
        signff(k) <= signff(k-1);
      END LOOP;    
    END IF;
    
  END PROCESS;

  --***************  
  --*** OUTPUTS ***
  --***************
  
  ccman <= mantissanorm(63 DOWNTO 11);
  ccexp <= exponentnorm;          
  ccsgn <= signff(25+7*doublespeed);
  zeroout <= zeronorm;
  
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   DP_LNADD.VHD                              ***
--***                                             ***
--***   Function: Double Precision Addition of    ***
--***   LN elements                               ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** Latency = 4 + 2*Speed                       ***
--***************************************************

ENTITY dp_lnadd IS 
GENERIC (
         speed : integer := 1; -- '0' for unpiped adder, '1' for piped adder
         synthesize : integer := 1
        ); 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      aaman : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
      aaexp : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
      bbman : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
      bbexp : IN STD_LOGIC_VECTOR (11 DOWNTO 1);

	   ccman : OUT STD_LOGIC_VECTOR (64 DOWNTO 1);
	   ccexp : OUT STD_LOGIC_VECTOR (11 DOWNTO 1)
	 );
END dp_lnadd;

ARCHITECTURE rtl OF dp_lnadd IS
  
  type expbasefftype IS ARRAY (3+2*speed DOWNTO 1) OF STD_LOGIC_VECTOR (13 DOWNTO 1);
  
  signal aamanff, bbmanff : STD_LOGIC_VECTOR (64 DOWNTO 1); 
  signal aaexpff, bbexpff : STD_LOGIC_VECTOR (11 DOWNTO 1);  
  signal manleftff, manrightff : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal aluleftff, alurightff : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal expbaseff : expbasefftype;
  signal shiftff : STD_LOGIC_VECTOR (5 DOWNTO 1);
  signal subexpone, subexptwo : STD_LOGIC_VECTOR (12 DOWNTO 1);
  signal switch : STD_LOGIC;
  signal shiftleftnode, shiftrightnode : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal alunode : STD_LOGIC_VECTOR (64 DOWNTO 1);
  
    component dp_rsft64x5 IS 
  PORT (
        inbus : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (5 DOWNTO 1);
        outbus : OUT STD_LOGIC_VECTOR (64 DOWNTO 1)
      );
  end component;
  
  component dp_rsft64x5pipe IS 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        inbus : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (5 DOWNTO 1);
        outbus : OUT STD_LOGIC_VECTOR (64 DOWNTO 1)
      );
  end component;

  component fp_del
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
  end component;
  
  component dp_fxadd 
  GENERIC (
           width : positive := 64;
           pipes : positive := 1;
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
        carryin : IN STD_LOGIC;
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
  end component;
     
BEGIN
     
  paa: PROCESS (sysclk, reset)
  BEGIN
      
    IF (reset = '1') THEN
       
      FOR k IN 1 TO 64 LOOP 
        aamanff(k) <= '0';
        bbmanff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 11 LOOP 
        aaexpff(k) <= '0';
        bbexpff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 64 LOOP
        manleftff(k) <= '0';
        manrightff(k) <= '0';
        aluleftff(k) <= '0';
        alurightff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 11 LOOP
        FOR j IN 1 TO 3+speed LOOP
          expbaseff(j)(k) <= '0';
        END LOOP;
      END LOOP;
      shiftff <= "00000";
        
    ELSIF (rising_edge(sysclk)) THEN
            
      IF (enable = '1') THEN
          
        --*** LEVEL 1 ***
        aamanff <= aaman;
        bbmanff <= bbman;
        aaexpff <= aaexp;
        bbexpff <= bbexp;
        
        --*** LEVEL 2 ***
        FOR k IN 1 TO 64 LOOP
          manleftff(k) <= (aamanff(k) AND NOT(switch)) OR (bbmanff(k) AND switch);
          manrightff(k) <= (bbmanff(k) AND NOT(switch)) OR (aamanff(k) AND switch);
        END LOOP;
          
        FOR k IN 1 TO 11 LOOP
          expbaseff(1)(k) <= (aaexpff(k) AND NOT(switch)) OR (bbexpff(k) AND switch); 
        END LOOP;
        FOR k IN 2 TO (3+2*speed) LOOP
          expbaseff(k)(11 DOWNTO 1) <= expbaseff(k-1)(11 DOWNTO 1);  -- level 3 to 4/6
        END LOOP;
        
        FOR k IN 1 TO 5 LOOP
          shiftff(k) <= (subexpone(k) AND NOT(switch)) OR (subexptwo(k) AND switch);
        END LOOP;
        
        aluleftff <= shiftleftnode;
        alurightff <= shiftrightnode;
      
      END IF;
        
    END IF;
      
  END PROCESS;
  
  subexpone <= ('0' & aaexpff) - ('0' & bbexpff);
  subexptwo <= ('0' & bbexpff) - ('0' & aaexpff);

  switch <= subexpone(12);

  gsa: IF (speed = 0) GENERATE
  
    shifter: dp_rsft64x5
    PORT MAP (inbus=>manrightff,shift=>shiftff,
              outbus=>shiftrightnode);
              
    shiftleftnode <= manleftff;
              
  END GENERATE;

  gsb: IF (speed = 1) GENERATE
  
    shifter: dp_rsft64x5pipe
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              inbus=>manrightff,shift=>shiftff,
              outbus=>shiftrightnode);
   
    sftdel: fp_del
    GENERIC MAP (width=>64,pipes=>1)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>manleftff,
              cc=>shiftleftnode);

  END GENERATE;

  -- level 3+speed in, level 4+2*speed out
  adder: dp_fxadd
  GENERIC MAP (width=>64,pipes=>speed+1,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>aluleftff,bb=>alurightff,carryin=>'0',
            cc=>alunode);

  --*** OUTPUTS ***
  ccman <= alunode;
  ccexp <= expbaseff(3+2*speed)(11 DOWNTO 1);

END rtl;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   DP_LNCLZ.VHD                              ***
--***                                             ***
--***   Function: Double Precision CLZ (no pipe)  ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_lnclz IS
PORT (
      mantissa : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
      
      leading : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
     );
END dp_lnclz;

ARCHITECTURE rtl of dp_lnclz IS

  type positiontype IS ARRAY (11 DOWNTO 1) OF STD_LOGIC_VECTOR (6 DOWNTO 1);
  
  signal position, positionmux : positiontype;
  signal zerogroup, firstzero : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal lastman : STD_LOGIC_VECTOR (6 DOWNTO 1);
  
  component dp_pos
  GENERIC (start: integer := 0);
  PORT 
       (
        ingroup : IN STD_LOGIC_VECTOR (6 DOWNTO 1); 
        
        position : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
       );
  end component;
  
BEGIN
     
  zerogroup(1) <= mantissa(64) OR mantissa(63) OR mantissa(62) OR mantissa(61) OR mantissa(60) OR mantissa(59);
  zerogroup(2) <= mantissa(58) OR mantissa(57) OR mantissa(56) OR mantissa(55) OR mantissa(54) OR mantissa(53);
  zerogroup(3) <= mantissa(52) OR mantissa(51) OR mantissa(50) OR mantissa(49) OR mantissa(48) OR mantissa(47);
  zerogroup(4) <= mantissa(46) OR mantissa(45) OR mantissa(44) OR mantissa(43) OR mantissa(42) OR mantissa(41);
  zerogroup(5) <= mantissa(40) OR mantissa(39) OR mantissa(38) OR mantissa(37) OR mantissa(36) OR mantissa(35);
  zerogroup(6) <= mantissa(34) OR mantissa(33) OR mantissa(32) OR mantissa(31) OR mantissa(30) OR mantissa(29);
  zerogroup(7) <= mantissa(28) OR mantissa(27) OR mantissa(26) OR mantissa(25) OR mantissa(24) OR mantissa(23);
  zerogroup(8) <= mantissa(22) OR mantissa(21) OR mantissa(20) OR mantissa(19) OR mantissa(18) OR mantissa(17);
  zerogroup(9) <= mantissa(16) OR mantissa(15) OR mantissa(14) OR mantissa(13) OR mantissa(12) OR mantissa(11);
  zerogroup(10) <= mantissa(10) OR mantissa(9) OR mantissa(8) OR mantissa(7) OR mantissa(6) OR mantissa(5);
  zerogroup(11) <= mantissa(4) OR mantissa(3) OR mantissa(2) OR mantissa(1);

  pa: dp_pos 
  GENERIC MAP (start=>0) 
  PORT MAP (ingroup=>mantissa(64 DOWNTO 59),position=>position(1)(6 DOWNTO 1));
  pb: dp_pos 
  GENERIC MAP (start=>6) 
  PORT MAP (ingroup=>mantissa(58 DOWNTO 53),position=>position(2)(6 DOWNTO 1));
  pc: dp_pos 
  GENERIC MAP (start=>12) 
  PORT MAP (ingroup=>mantissa(52 DOWNTO 47),position=>position(3)(6 DOWNTO 1));
  pd: dp_pos 
  GENERIC MAP (start=>18) 
  PORT MAP (ingroup=>mantissa(46 DOWNTO 41),position=>position(4)(6 DOWNTO 1));
  pe: dp_pos 
  GENERIC MAP (start=>24) 
  PORT MAP (ingroup=>mantissa(40 DOWNTO 35),position=>position(5)(6 DOWNTO 1));
  pf: dp_pos 
  GENERIC MAP (start=>30) 
  PORT MAP (ingroup=>mantissa(34 DOWNTO 29),position=>position(6)(6 DOWNTO 1));
  pg: dp_pos 
  GENERIC MAP (start=>36) 
  PORT MAP (ingroup=>mantissa(28 DOWNTO 23),position=>position(7)(6 DOWNTO 1));
  ph: dp_pos 
  GENERIC MAP (start=>42) 
  PORT MAP (ingroup=>mantissa(22 DOWNTO 17),position=>position(8)(6 DOWNTO 1));
  pi: dp_pos 
  GENERIC MAP (start=>48) 
  PORT MAP (ingroup=>mantissa(16 DOWNTO 11),position=>position(9)(6 DOWNTO 1));
  pj: dp_pos 
  GENERIC MAP (start=>54) 
  PORT MAP (ingroup=>mantissa(10 DOWNTO 5),position=>position(10)(6 DOWNTO 1));
  pk: dp_pos 
  GENERIC MAP (start=>60) 
  PORT MAP (ingroup=>lastman,position=>position(11)(6 DOWNTO 1));
      
  lastman <= mantissa(4 DOWNTO 1) & "00";

  firstzero(1) <= zerogroup(1);
  firstzero(2) <= NOT(zerogroup(1)) AND zerogroup(2);
  firstzero(3) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND zerogroup(3);
  firstzero(4) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND zerogroup(4);
  firstzero(5) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND NOT(zerogroup(4)) 
                  AND zerogroup(5);
  firstzero(6) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND NOT(zerogroup(4)) 
                  AND NOT(zerogroup(5)) AND zerogroup(6);                
  firstzero(7) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND NOT(zerogroup(4)) 
                  AND NOT(zerogroup(5)) AND NOT(zerogroup(6)) AND zerogroup(7); 
  firstzero(8) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND NOT(zerogroup(4)) 
                  AND NOT(zerogroup(5)) AND NOT(zerogroup(6)) AND NOT(zerogroup(7)) AND zerogroup(8); 
  firstzero(9) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND NOT(zerogroup(4)) 
                  AND NOT(zerogroup(5)) AND NOT(zerogroup(6)) AND NOT(zerogroup(7)) AND NOT(zerogroup(8)) 
                  AND zerogroup(9); 
  firstzero(10) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND NOT(zerogroup(4)) 
                   AND NOT(zerogroup(5)) AND NOT(zerogroup(6)) AND NOT(zerogroup(7)) AND NOT(zerogroup(8)) 
                   AND NOT(zerogroup(9)) AND zerogroup(10); 
  firstzero(11) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND NOT(zerogroup(4)) 
                   AND NOT(zerogroup(5)) AND NOT(zerogroup(6)) AND NOT(zerogroup(7)) AND NOT(zerogroup(8)) 
                   AND NOT(zerogroup(9)) AND NOT(zerogroup(10)) AND zerogroup(11); 
                
gma: FOR k IN 1 TO 6 GENERATE
  positionmux(1)(k) <= position(1)(k) AND firstzero(1);
  gmb: FOR j IN 2 TO 11 GENERATE
    positionmux(j)(k) <= positionmux(j-1)(k) OR (position(j)(k) AND firstzero(j));
  END GENERATE;
END GENERATE;
  
leading <= positionmux(11)(6 DOWNTO 1);
                                               
END rtl;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   DP_LNCLZPIPE.VHD                          ***
--***                                             ***
--***   Function: Double Precision CLZ pipelined  ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_lnclzpipe IS
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      mantissa : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
      
      leading : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
     );
END dp_lnclzpipe;

ARCHITECTURE rtl of dp_lnclzpipe IS

  type positiontype IS ARRAY (11 DOWNTO 1) OF STD_LOGIC_VECTOR (6 DOWNTO 1);
  
  signal position, positionff, positionmux : positiontype;
  signal zerogroup, zerogroupff, firstzero : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal lastman : STD_LOGIC_VECTOR (6 DOWNTO 1);
  
  component dp_pos
  GENERIC (start: integer := 0);
  PORT 
       (
        ingroup : IN STD_LOGIC_VECTOR (6 DOWNTO 1); 
        
        position : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
       );
  end component;
  
BEGIN
     
  zerogroup(1) <= mantissa(64) OR mantissa(63) OR mantissa(62) OR mantissa(61) OR mantissa(60) OR mantissa(59);
  zerogroup(2) <= mantissa(58) OR mantissa(57) OR mantissa(56) OR mantissa(55) OR mantissa(54) OR mantissa(53);
  zerogroup(3) <= mantissa(52) OR mantissa(51) OR mantissa(50) OR mantissa(49) OR mantissa(48) OR mantissa(47);
  zerogroup(4) <= mantissa(46) OR mantissa(45) OR mantissa(44) OR mantissa(43) OR mantissa(42) OR mantissa(41);
  zerogroup(5) <= mantissa(40) OR mantissa(39) OR mantissa(38) OR mantissa(37) OR mantissa(36) OR mantissa(35);
  zerogroup(6) <= mantissa(34) OR mantissa(33) OR mantissa(32) OR mantissa(31) OR mantissa(30) OR mantissa(29);
  zerogroup(7) <= mantissa(28) OR mantissa(27) OR mantissa(26) OR mantissa(25) OR mantissa(24) OR mantissa(23);
  zerogroup(8) <= mantissa(22) OR mantissa(21) OR mantissa(20) OR mantissa(19) OR mantissa(18) OR mantissa(17);
  zerogroup(9) <= mantissa(16) OR mantissa(15) OR mantissa(14) OR mantissa(13) OR mantissa(12) OR mantissa(11);
  zerogroup(10) <= mantissa(10) OR mantissa(9) OR mantissa(8) OR mantissa(7) OR mantissa(6) OR mantissa(5);
  zerogroup(11) <= mantissa(4) OR mantissa(3) OR mantissa(2) OR mantissa(1);

  pa: dp_pos 
  GENERIC MAP (start=>0) 
  PORT MAP (ingroup=>mantissa(64 DOWNTO 59),position=>position(1)(6 DOWNTO 1));
  pb: dp_pos 
  GENERIC MAP (start=>6) 
  PORT MAP (ingroup=>mantissa(58 DOWNTO 53),position=>position(2)(6 DOWNTO 1));
  pc: dp_pos 
  GENERIC MAP (start=>12) 
  PORT MAP (ingroup=>mantissa(52 DOWNTO 47),position=>position(3)(6 DOWNTO 1));
  pd: dp_pos 
  GENERIC MAP (start=>18) 
  PORT MAP (ingroup=>mantissa(46 DOWNTO 41),position=>position(4)(6 DOWNTO 1));
  pe: dp_pos 
  GENERIC MAP (start=>24) 
  PORT MAP (ingroup=>mantissa(40 DOWNTO 35),position=>position(5)(6 DOWNTO 1));
  pf: dp_pos 
  GENERIC MAP (start=>30) 
  PORT MAP (ingroup=>mantissa(34 DOWNTO 29),position=>position(6)(6 DOWNTO 1));
  pg: dp_pos 
  GENERIC MAP (start=>36) 
  PORT MAP (ingroup=>mantissa(28 DOWNTO 23),position=>position(7)(6 DOWNTO 1));
  ph: dp_pos 
  GENERIC MAP (start=>42) 
  PORT MAP (ingroup=>mantissa(22 DOWNTO 17),position=>position(8)(6 DOWNTO 1));
  pi: dp_pos 
  GENERIC MAP (start=>48) 
  PORT MAP (ingroup=>mantissa(16 DOWNTO 11),position=>position(9)(6 DOWNTO 1));
  pj: dp_pos 
  GENERIC MAP (start=>54) 
  PORT MAP (ingroup=>mantissa(10 DOWNTO 5),position=>position(10)(6 DOWNTO 1));
  pk: dp_pos 
  GENERIC MAP (start=>60) 
  PORT MAP (ingroup=>lastman,position=>position(11)(6 DOWNTO 1));
      
  lastman <= mantissa(4 DOWNTO 1) & "00";

  ppa: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN
        
      FOR k IN 1 TO 11 LOOP
        zerogroupff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 11 LOOP
        FOR j IN 1 TO 6 LOOP
          positionff(k)(j) <= '0';
        END LOOP;
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
    
      zerogroupff <= zerogroup;
      FOR k IN 1 TO 11 LOOP
        positionff(k)(6 DOWNTO 1) <= position(k)(6 DOWNTO 1);
      END LOOP;
              
    END IF;
      
  END PROCESS;
  
  firstzero(1) <= zerogroupff(1);
  firstzero(2) <= NOT(zerogroupff(1)) AND zerogroupff(2);
  firstzero(3) <= NOT(zerogroupff(1)) AND NOT(zerogroupff(2)) AND zerogroupff(3);
  firstzero(4) <= NOT(zerogroupff(1)) AND NOT(zerogroupff(2)) AND NOT(zerogroupff(3)) AND zerogroupff(4);
  firstzero(5) <= NOT(zerogroupff(1)) AND NOT(zerogroupff(2)) AND NOT(zerogroupff(3)) AND 
                  NOT(zerogroupff(4)) AND zerogroupff(5);
  firstzero(6) <= NOT(zerogroupff(1)) AND NOT(zerogroupff(2)) AND NOT(zerogroupff(3)) AND 
                  NOT(zerogroupff(4)) AND NOT(zerogroupff(5)) AND zerogroupff(6);                
  firstzero(7) <= NOT(zerogroupff(1)) AND NOT(zerogroupff(2)) AND NOT(zerogroupff(3)) AND 
                  NOT(zerogroupff(4)) AND NOT(zerogroupff(5)) AND NOT(zerogroupff(6)) AND zerogroupff(7); 
  firstzero(8) <= NOT(zerogroupff(1)) AND NOT(zerogroupff(2)) AND NOT(zerogroupff(3)) AND 
                  NOT(zerogroupff(4)) AND NOT(zerogroupff(5)) AND NOT(zerogroupff(6)) AND 
                  NOT(zerogroupff(7)) AND zerogroupff(8); 
  firstzero(9) <= NOT(zerogroupff(1)) AND NOT(zerogroupff(2)) AND NOT(zerogroupff(3)) AND 
                  NOT(zerogroupff(4)) AND NOT(zerogroupff(5)) AND NOT(zerogroupff(6)) AND 
                  NOT(zerogroupff(7)) AND NOT(zerogroupff(8)) AND zerogroupff(9); 
  firstzero(10) <= NOT(zerogroupff(1)) AND NOT(zerogroupff(2)) AND NOT(zerogroupff(3)) AND 
                   NOT(zerogroupff(4)) AND NOT(zerogroupff(5)) AND NOT(zerogroupff(6)) AND 
                   NOT(zerogroupff(7)) AND NOT(zerogroupff(8)) AND NOT(zerogroupff(9)) AND zerogroupff(10); 
  firstzero(11) <= NOT(zerogroupff(1)) AND NOT(zerogroupff(2)) AND NOT(zerogroupff(3)) AND 
                   NOT(zerogroupff(4)) AND NOT(zerogroupff(5)) AND NOT(zerogroupff(6)) AND 
                   NOT(zerogroupff(7)) AND NOT(zerogroupff(8)) AND NOT(zerogroupff(9)) AND 
                   NOT(zerogroupff(10)) AND zerogroupff(11); 
                
gma: FOR k IN 1 TO 6 GENERATE
  positionmux(1)(k) <= positionff(1)(k) AND firstzero(1);
  gmb: FOR j IN 2 TO 11 GENERATE
    positionmux(j)(k) <= positionmux(j-1)(k) OR (positionff(j)(k) AND firstzero(j));
  END GENERATE;
END GENERATE;
  
leading <= positionmux(11)(6 DOWNTO 1);
                                               
END rtl;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   DP_LNLUT18.VHD                            ***
--***                                             ***
--***   Function: Look Up Table - LN()            ***
--***                                             ***
--***   Generated by MATLAB Utility               ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_lnlut18 IS
PORT (
      add : IN STD_LOGIC_VECTOR (9 DOWNTO 1);
      inv : OUT STD_LOGIC_VECTOR (18 DOWNTO 1);
      logman : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
      logexp : OUT STD_LOGIC_VECTOR (11 DOWNTO 1)
     );
END dp_lnlut18;

ARCHITECTURE rtl OF dp_lnlut18 IS

BEGIN

  pca: PROCESS (add)
  BEGIN
    CASE add IS
      WHEN "000000000" =>
            inv <= conv_std_logic_vector(131072,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(0,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(0,28);
            logexp <= conv_std_logic_vector(0,11);
      WHEN "000000001" =>
            inv <= conv_std_logic_vector(262143,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(31,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(268391765,28);
            logexp <= conv_std_logic_vector(1005,11);
      WHEN "000000010" =>
            inv <= conv_std_logic_vector(262141,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8388752,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(327672,28);
            logexp <= conv_std_logic_vector(1006,11);
      WHEN "000000011" =>
            inv <= conv_std_logic_vector(262139,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4194504,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(666254,28);
            logexp <= conv_std_logic_vector(1007,11);
      WHEN "000000100" =>
            inv <= conv_std_logic_vector(262137,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12583304,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(1889508,28);
            logexp <= conv_std_logic_vector(1007,11);
      WHEN "000000101" =>
            inv <= conv_std_logic_vector(262135,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2097476,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(1982311,28);
            logexp <= conv_std_logic_vector(1008,11);
      WHEN "000000110" =>
            inv <= conv_std_logic_vector(262133,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6291940,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(3642366,28);
            logexp <= conv_std_logic_vector(1008,11);
      WHEN "000000111" =>
            inv <= conv_std_logic_vector(262131,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10486436,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(5990414,28);
            logexp <= conv_std_logic_vector(1008,11);
      WHEN "000001000" =>
            inv <= conv_std_logic_vector(262129,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14680964,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(9223005,28);
            logexp <= conv_std_logic_vector(1008,11);
      WHEN "000001001" =>
            inv <= conv_std_logic_vector(262127,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1049154,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(6702808,28);
            logexp <= conv_std_logic_vector(1009,11);
      WHEN "000001010" =>
            inv <= conv_std_logic_vector(262125,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3146450,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(9367390,28);
            logexp <= conv_std_logic_vector(1009,11);
      WHEN "000001011" =>
            inv <= conv_std_logic_vector(262123,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5243762,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(12637977,28);
            logexp <= conv_std_logic_vector(1009,11);
      WHEN "000001100" =>
            inv <= conv_std_logic_vector(262121,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7341090,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(16612827,28);
            logexp <= conv_std_logic_vector(1009,11);
      WHEN "000001101" =>
            inv <= conv_std_logic_vector(262119,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9438434,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(21341043,28);
            logexp <= conv_std_logic_vector(1009,11);
      WHEN "000001110" =>
            inv <= conv_std_logic_vector(262117,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11535794,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(26871724,28);
            logexp <= conv_std_logic_vector(1009,11);
      WHEN "000001111" =>
            inv <= conv_std_logic_vector(262115,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13633170,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(33303113,28);
            logexp <= conv_std_logic_vector(1009,11);
      WHEN "000010000" =>
            inv <= conv_std_logic_vector(262113,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15730562,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(40684301,28);
            logexp <= conv_std_logic_vector(1009,11);
      WHEN "000010001" =>
            inv <= conv_std_logic_vector(262111,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(525377,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(24532187,28);
            logexp <= conv_std_logic_vector(1010,11);
      WHEN "000010010" =>
            inv <= conv_std_logic_vector(262109,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1574089,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(29270780,28);
            logexp <= conv_std_logic_vector(1010,11);
      WHEN "000010011" =>
            inv <= conv_std_logic_vector(262107,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2622809,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(34582468,28);
            logexp <= conv_std_logic_vector(1010,11);
      WHEN "000010100" =>
            inv <= conv_std_logic_vector(262105,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3671537,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(40499978,28);
            logexp <= conv_std_logic_vector(1010,11);
      WHEN "000010101" =>
            inv <= conv_std_logic_vector(262103,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4720273,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(47056037,28);
            logexp <= conv_std_logic_vector(1010,11);
      WHEN "000010110" =>
            inv <= conv_std_logic_vector(262101,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5769017,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(54283367,28);
            logexp <= conv_std_logic_vector(1010,11);
      WHEN "000010111" =>
            inv <= conv_std_logic_vector(262099,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6817769,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(62214689,28);
            logexp <= conv_std_logic_vector(1010,11);
      WHEN "000011000" =>
            inv <= conv_std_logic_vector(262097,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7866529,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(70882721,28);
            logexp <= conv_std_logic_vector(1010,11);
      WHEN "000011001" =>
            inv <= conv_std_logic_vector(262095,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8915297,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(80328369,28);
            logexp <= conv_std_logic_vector(1010,11);
      WHEN "000011010" =>
            inv <= conv_std_logic_vector(262093,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9964073,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(90567968,28);
            logexp <= conv_std_logic_vector(1010,11);
      WHEN "000011011" =>
            inv <= conv_std_logic_vector(262091,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11012857,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(101650610,28);
            logexp <= conv_std_logic_vector(1010,11);
      WHEN "000011100" =>
            inv <= conv_std_logic_vector(262089,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12061649,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(113592623,28);
            logexp <= conv_std_logic_vector(1010,11);
      WHEN "000011101" =>
            inv <= conv_std_logic_vector(262087,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13110449,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(126443095,28);
            logexp <= conv_std_logic_vector(1010,11);
      WHEN "000011110" =>
            inv <= conv_std_logic_vector(262085,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14159257,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(140226541,28);
            logexp <= conv_std_logic_vector(1010,11);
      WHEN "000011111" =>
            inv <= conv_std_logic_vector(262083,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15208073,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(154975663,28);
            logexp <= conv_std_logic_vector(1010,11);
      WHEN "000100000" =>
            inv <= conv_std_logic_vector(262081,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16256897,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(170731353,28);
            logexp <= conv_std_logic_vector(1010,11);
      WHEN "000100001" =>
            inv <= conv_std_logic_vector(262079,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(264256,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(227972692,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000100010" =>
            inv <= conv_std_logic_vector(262077,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(788676,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(236897961,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000100011" =>
            inv <= conv_std_logic_vector(262075,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1313100,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(246371462,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000100100" =>
            inv <= conv_std_logic_vector(262073,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1837528,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(256409541,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000100101" =>
            inv <= conv_std_logic_vector(262071,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2361960,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(267028543,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000100110" =>
            inv <= conv_std_logic_vector(262069,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2886397,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(9813450,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000100111" =>
            inv <= conv_std_logic_vector(262067,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3410837,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(21647423,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000101000" =>
            inv <= conv_std_logic_vector(262065,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3935281,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(34111345,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000101001" =>
            inv <= conv_std_logic_vector(262063,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4459729,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(47221557,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000101010" =>
            inv <= conv_std_logic_vector(262061,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4984181,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(60998494,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000101011" =>
            inv <= conv_std_logic_vector(262059,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5508637,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(75454397,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000101100" =>
            inv <= conv_std_logic_vector(262057,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6033097,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(90605604,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000101101" =>
            inv <= conv_std_logic_vector(262055,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6557561,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(106472545,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000101110" =>
            inv <= conv_std_logic_vector(262053,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7082029,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(123067460,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000101111" =>
            inv <= conv_std_logic_vector(262051,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7606501,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(140410777,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000110000" =>
            inv <= conv_std_logic_vector(262049,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8130977,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(158510638,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000110001" =>
            inv <= conv_std_logic_vector(262047,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8655457,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(177395659,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000110010" =>
            inv <= conv_std_logic_vector(262045,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9179941,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(197069887,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000110011" =>
            inv <= conv_std_logic_vector(262043,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9704429,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(217561932,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000110100" =>
            inv <= conv_std_logic_vector(262041,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10228921,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(238875840,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000110101" =>
            inv <= conv_std_logic_vector(262039,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10753417,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(261036127,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000110110" =>
            inv <= conv_std_logic_vector(262037,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11277918,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(15623661,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000110111" =>
            inv <= conv_std_logic_vector(262035,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11802422,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(39521584,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000111000" =>
            inv <= conv_std_logic_vector(262033,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12326930,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(64314859,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000111001" =>
            inv <= conv_std_logic_vector(262031,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12851442,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(90015713,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000111010" =>
            inv <= conv_std_logic_vector(262029,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13375958,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(116644561,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000111011" =>
            inv <= conv_std_logic_vector(262027,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13900478,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(144213628,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000111100" =>
            inv <= conv_std_logic_vector(262025,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14425002,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(172743328,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000111101" =>
            inv <= conv_std_logic_vector(262023,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14949530,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(202249979,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000111110" =>
            inv <= conv_std_logic_vector(262021,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15474062,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(232745802,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "000111111" =>
            inv <= conv_std_logic_vector(262019,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15998598,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(264251207,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "001000000" =>
            inv <= conv_std_logic_vector(262017,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16523139,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(28347053,28);
            logexp <= conv_std_logic_vector(1011,11);
      WHEN "001000001" =>
            inv <= conv_std_logic_vector(262015,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(135233,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(165175963,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001000010" =>
            inv <= conv_std_logic_vector(262013,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(397507,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(182491979,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001000011" =>
            inv <= conv_std_logic_vector(262011,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(659783,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(200343364,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001000100" =>
            inv <= conv_std_logic_vector(262009,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(922061,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(218740319,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001000101" =>
            inv <= conv_std_logic_vector(262007,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1184341,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(237688954,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001000110" =>
            inv <= conv_std_logic_vector(262005,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1446623,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(257201513,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001000111" =>
            inv <= conv_std_logic_vector(262003,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1708908,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(8846602,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001001000" =>
            inv <= conv_std_logic_vector(262001,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1971194,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(29507379,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001001001" =>
            inv <= conv_std_logic_vector(261999,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2233482,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(50752445,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001001010" =>
            inv <= conv_std_logic_vector(261997,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2495772,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(72592000,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001001011" =>
            inv <= conv_std_logic_vector(261995,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2758064,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(95036240,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001001100" =>
            inv <= conv_std_logic_vector(261993,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3020358,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(118089223,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001001101" =>
            inv <= conv_std_logic_vector(261991,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3282654,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(141761145,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001001110" =>
            inv <= conv_std_logic_vector(261989,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3544952,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(166062202,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001001111" =>
            inv <= conv_std_logic_vector(261987,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3807252,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(190996450,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001010000" =>
            inv <= conv_std_logic_vector(261985,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4069554,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(216576129,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001010001" =>
            inv <= conv_std_logic_vector(261983,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4331858,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(242805295,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001010010" =>
            inv <= conv_std_logic_vector(261981,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4594165,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(1260730,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001010011" =>
            inv <= conv_std_logic_vector(261979,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4856473,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(28821495,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001010100" =>
            inv <= conv_std_logic_vector(261977,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5118783,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(57056185,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001010101" =>
            inv <= conv_std_logic_vector(261975,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5381095,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(85977038,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001010110" =>
            inv <= conv_std_logic_vector(261973,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5643409,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(115590153,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001010111" =>
            inv <= conv_std_logic_vector(261971,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5905725,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(145903675,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001011000" =>
            inv <= conv_std_logic_vector(261969,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6168043,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(176927792,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001011001" =>
            inv <= conv_std_logic_vector(261967,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6430363,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(208668602,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001011010" =>
            inv <= conv_std_logic_vector(261965,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6692685,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(241134248,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001011011" =>
            inv <= conv_std_logic_vector(261963,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6955010,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(5901507,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001011100" =>
            inv <= conv_std_logic_vector(261961,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7217336,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(39843294,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001011101" =>
            inv <= conv_std_logic_vector(261959,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7479664,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(74536387,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001011110" =>
            inv <= conv_std_logic_vector(261957,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7741994,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(109988926,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001011111" =>
            inv <= conv_std_logic_vector(261955,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8004326,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(146207004,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001100000" =>
            inv <= conv_std_logic_vector(261953,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8266660,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(183200806,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001100001" =>
            inv <= conv_std_logic_vector(261951,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8528996,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(220976425,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001100010" =>
            inv <= conv_std_logic_vector(261949,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8791334,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(259546091,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001100011" =>
            inv <= conv_std_logic_vector(261947,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9053675,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(30478393,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001100100" =>
            inv <= conv_std_logic_vector(261945,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9316017,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(70652380,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001100101" =>
            inv <= conv_std_logic_vector(261943,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9578361,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(111644825,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001100110" =>
            inv <= conv_std_logic_vector(261941,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9840707,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(153461817,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001100111" =>
            inv <= conv_std_logic_vector(261939,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10103055,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(196109445,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001101000" =>
            inv <= conv_std_logic_vector(261937,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10365405,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(239597890,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001101001" =>
            inv <= conv_std_logic_vector(261935,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10627758,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(15499830,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001101010" =>
            inv <= conv_std_logic_vector(261933,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10890112,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(60696356,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001101011" =>
            inv <= conv_std_logic_vector(261931,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11152468,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(106756053,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001101100" =>
            inv <= conv_std_logic_vector(261929,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11414826,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(153689099,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001101101" =>
            inv <= conv_std_logic_vector(261927,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11677186,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(201505673,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001101110" =>
            inv <= conv_std_logic_vector(261925,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11939548,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(250209813,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001101111" =>
            inv <= conv_std_logic_vector(261923,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12201913,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(31378287,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001110000" =>
            inv <= conv_std_logic_vector(261921,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12464279,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(81888089,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001110001" =>
            inv <= conv_std_logic_vector(261919,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12726647,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(133313941,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001110010" =>
            inv <= conv_std_logic_vector(261917,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12989017,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(185659877,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001110011" =>
            inv <= conv_std_logic_vector(261915,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13251389,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(238938120,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001110100" =>
            inv <= conv_std_logic_vector(261913,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13513764,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(24721341,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001110101" =>
            inv <= conv_std_logic_vector(261911,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13776140,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(79886532,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001110110" =>
            inv <= conv_std_logic_vector(261909,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14038518,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(136006365,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001110111" =>
            inv <= conv_std_logic_vector(261907,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14300898,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(193091012,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001111000" =>
            inv <= conv_std_logic_vector(261905,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14563280,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(251146552,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001111001" =>
            inv <= conv_std_logic_vector(261903,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14825665,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(41747701,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001111010" =>
            inv <= conv_std_logic_vector(261901,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15088051,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(101773495,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001111011" =>
            inv <= conv_std_logic_vector(261899,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15350439,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(162796601,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001111100" =>
            inv <= conv_std_logic_vector(261897,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15612829,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(224823097,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001111101" =>
            inv <= conv_std_logic_vector(261895,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15875222,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(19427696,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001111110" =>
            inv <= conv_std_logic_vector(261893,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16137616,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(83489431,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "001111111" =>
            inv <= conv_std_logic_vector(261891,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16400012,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(148578923,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "010000000" =>
            inv <= conv_std_logic_vector(261889,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16662410,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(214708384,28);
            logexp <= conv_std_logic_vector(1012,11);
      WHEN "010000001" =>
            inv <= conv_std_logic_vector(261887,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(73797,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(140941945,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010000010" =>
            inv <= conv_std_logic_vector(261885,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(204998,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(175055756,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010000011" =>
            inv <= conv_std_logic_vector(261883,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(336200,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(209701733,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010000100" =>
            inv <= conv_std_logic_vector(261881,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(467403,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(244882910,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010000101" =>
            inv <= conv_std_logic_vector(261879,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(598608,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(12167891,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010000110" =>
            inv <= conv_std_logic_vector(261877,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(729813,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(48431647,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010000111" =>
            inv <= conv_std_logic_vector(261875,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(861019,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(85243804,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010001000" =>
            inv <= conv_std_logic_vector(261873,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(992226,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(122607396,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010001001" =>
            inv <= conv_std_logic_vector(261871,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1123434,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(160526482,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010001010" =>
            inv <= conv_std_logic_vector(261869,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1254643,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(199006142,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010001011" =>
            inv <= conv_std_logic_vector(261867,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1385853,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(238049411,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010001100" =>
            inv <= conv_std_logic_vector(261865,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1517065,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(9224891,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010001101" =>
            inv <= conv_std_logic_vector(261863,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1648277,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(49409594,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010001110" =>
            inv <= conv_std_logic_vector(261861,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1779490,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(90169054,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010001111" =>
            inv <= conv_std_logic_vector(261859,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1910704,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(131510396,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010010000" =>
            inv <= conv_std_logic_vector(261857,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2041919,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(173435630,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010010001" =>
            inv <= conv_std_logic_vector(261855,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2173135,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(215949833,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010010010" =>
            inv <= conv_std_logic_vector(261853,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2304352,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(259057063,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010010011" =>
            inv <= conv_std_logic_vector(261851,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2435571,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(34325917,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010010100" =>
            inv <= conv_std_logic_vector(261849,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2566790,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(78630340,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010010101" =>
            inv <= conv_std_logic_vector(261847,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2698010,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(123540976,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010010110" =>
            inv <= conv_std_logic_vector(261845,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2829231,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(169060858,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010010111" =>
            inv <= conv_std_logic_vector(261843,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2960453,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(215194037,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010011000" =>
            inv <= conv_std_logic_vector(261841,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3091676,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(261943547,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010011001" =>
            inv <= conv_std_logic_vector(261839,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3222901,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(40881052,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010011010" =>
            inv <= conv_std_logic_vector(261837,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3354126,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(88878449,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010011011" =>
            inv <= conv_std_logic_vector(261835,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3485352,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(137506381,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010011100" =>
            inv <= conv_std_logic_vector(261833,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3616579,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(186767878,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010011101" =>
            inv <= conv_std_logic_vector(261831,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3747807,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(236666992,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010011110" =>
            inv <= conv_std_logic_vector(261829,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3879037,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(18774364,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010011111" =>
            inv <= conv_std_logic_vector(261827,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4010267,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(69961890,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010100000" =>
            inv <= conv_std_logic_vector(261825,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4141498,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(121800212,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010100001" =>
            inv <= conv_std_logic_vector(261823,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4272730,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(174293379,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010100010" =>
            inv <= conv_std_logic_vector(261821,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4403963,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(227445444,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010100011" =>
            inv <= conv_std_logic_vector(261819,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4535198,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(12823978,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010100100" =>
            inv <= conv_std_logic_vector(261817,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4666433,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(67305989,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010100101" =>
            inv <= conv_std_logic_vector(261815,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4797669,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(122458025,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010100110" =>
            inv <= conv_std_logic_vector(261813,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4928906,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(178285160,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010100111" =>
            inv <= conv_std_logic_vector(261811,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5060144,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(234791442,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010101000" =>
            inv <= conv_std_logic_vector(261809,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5191384,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(23545465,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010101001" =>
            inv <= conv_std_logic_vector(261807,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5322624,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(81422190,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010101010" =>
            inv <= conv_std_logic_vector(261805,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5453865,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(139991231,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010101011" =>
            inv <= conv_std_logic_vector(261803,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5585107,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(199255616,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010101100" =>
            inv <= conv_std_logic_vector(261801,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5716350,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(259219392,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010101101" =>
            inv <= conv_std_logic_vector(261799,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5847595,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(51452173,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010101110" =>
            inv <= conv_std_logic_vector(261797,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5978840,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(112827896,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010101111" =>
            inv <= conv_std_logic_vector(261795,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6110086,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(174915153,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010110000" =>
            inv <= conv_std_logic_vector(261793,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6241333,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(237719013,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010110001" =>
            inv <= conv_std_logic_vector(261791,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6372582,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(32808067,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010110010" =>
            inv <= conv_std_logic_vector(261789,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6503831,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(97057274,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010110011" =>
            inv <= conv_std_logic_vector(261787,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6635081,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(162034200,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010110100" =>
            inv <= conv_std_logic_vector(261785,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6766332,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(227743914,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010110101" =>
            inv <= conv_std_logic_vector(261783,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6897585,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(25755007,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010110110" =>
            inv <= conv_std_logic_vector(261781,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7028838,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(92942434,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010110111" =>
            inv <= conv_std_logic_vector(261779,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7160092,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(160875808,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010111000" =>
            inv <= conv_std_logic_vector(261777,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7291347,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(229557128,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010111001" =>
            inv <= conv_std_logic_vector(261775,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7422604,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(30556006,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010111010" =>
            inv <= conv_std_logic_vector(261773,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7553861,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(100748419,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010111011" =>
            inv <= conv_std_logic_vector(261771,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7685119,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(171701934,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010111100" =>
            inv <= conv_std_logic_vector(261769,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7816378,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(243420594,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010111101" =>
            inv <= conv_std_logic_vector(261767,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7947639,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(47474008,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010111110" =>
            inv <= conv_std_logic_vector(261765,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8078900,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(120736110,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "010111111" =>
            inv <= conv_std_logic_vector(261763,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8210162,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(194776508,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011000000" =>
            inv <= conv_std_logic_vector(261761,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8341426,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(1163789,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011000001" =>
            inv <= conv_std_logic_vector(261759,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8472690,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(76771885,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011000010" =>
            inv <= conv_std_logic_vector(261757,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8603955,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(153170403,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011000011" =>
            inv <= conv_std_logic_vector(261755,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8735221,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(230363387,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011000100" =>
            inv <= conv_std_logic_vector(261753,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8866489,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(39919420,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011000101" =>
            inv <= conv_std_logic_vector(261751,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8997757,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(118713456,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011000110" =>
            inv <= conv_std_logic_vector(261749,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9129026,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(198314080,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011000111" =>
            inv <= conv_std_logic_vector(261747,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9260297,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(10289876,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011001000" =>
            inv <= conv_std_logic_vector(261745,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9391568,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(91515797,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011001001" =>
            inv <= conv_std_logic_vector(261743,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9522840,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(173561448,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011001010" =>
            inv <= conv_std_logic_vector(261741,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9654113,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(256429848,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011001011" =>
            inv <= conv_std_logic_vector(261739,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9785388,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(71690601,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011001100" =>
            inv <= conv_std_logic_vector(261737,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9916663,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(156217637,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011001101" =>
            inv <= conv_std_logic_vector(261735,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10047939,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(241580560,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011001110" =>
            inv <= conv_std_logic_vector(261733,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10179217,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(59346931,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011001111" =>
            inv <= conv_std_logic_vector(261731,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10310495,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(146392723,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011010000" =>
            inv <= conv_std_logic_vector(261729,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10441774,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(234286516,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011010001" =>
            inv <= conv_std_logic_vector(261727,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10573055,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(54596894,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011010010" =>
            inv <= conv_std_logic_vector(261725,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10704336,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(144198805,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011010011" =>
            inv <= conv_std_logic_vector(261723,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10835618,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(234660830,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011010100" =>
            inv <= conv_std_logic_vector(261721,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10966902,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(57551551,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011010101" =>
            inv <= conv_std_logic_vector(261719,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11098186,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(149745915,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011010110" =>
            inv <= conv_std_logic_vector(261717,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11229471,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(242812504,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011010111" =>
            inv <= conv_std_logic_vector(261715,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11360758,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(68320919,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011011000" =>
            inv <= conv_std_logic_vector(261713,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11492045,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(163146107,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011011001" =>
            inv <= conv_std_logic_vector(261711,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11623333,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(258854605,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011011010" =>
            inv <= conv_std_logic_vector(261709,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11754623,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(87018057,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011011011" =>
            inv <= conv_std_logic_vector(261707,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11885913,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(184509366,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011011100" =>
            inv <= conv_std_logic_vector(261705,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12017205,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(14462677,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011011101" =>
            inv <= conv_std_logic_vector(261703,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12148497,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(113752937,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011011110" =>
            inv <= conv_std_logic_vector(261701,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12279790,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(213947700,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011011111" =>
            inv <= conv_std_logic_vector(261699,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12411085,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(46617589,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011100000" =>
            inv <= conv_std_logic_vector(261697,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12542380,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(148636528,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011100001" =>
            inv <= conv_std_logic_vector(261695,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12673676,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(251573093,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011100010" =>
            inv <= conv_std_logic_vector(261693,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12804974,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(86995861,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011100011" =>
            inv <= conv_std_logic_vector(261691,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12936272,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(191780799,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011100100" =>
            inv <= conv_std_logic_vector(261689,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13067572,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(29060005,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011100101" =>
            inv <= conv_std_logic_vector(261687,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13198872,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(135708424,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011100110" =>
            inv <= conv_std_logic_vector(261685,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13330173,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(243295652,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011100111" =>
            inv <= conv_std_logic_vector(261683,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13461476,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(83390266,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011101000" =>
            inv <= conv_std_logic_vector(261681,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13592779,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(192867209,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011101001" =>
            inv <= conv_std_logic_vector(261679,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13724084,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(34858577,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011101010" =>
            inv <= conv_std_logic_vector(261677,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13855389,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(146240336,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011101011" =>
            inv <= conv_std_logic_vector(261675,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13986695,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(258581058,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011101100" =>
            inv <= conv_std_logic_vector(261673,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14118003,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(103450342,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011101101" =>
            inv <= conv_std_logic_vector(261671,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14249311,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(217721083,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011101110" =>
            inv <= conv_std_logic_vector(261669,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14380621,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(64528444,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011101111" =>
            inv <= conv_std_logic_vector(261667,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14511931,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(180746345,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011110000" =>
            inv <= conv_std_logic_vector(261665,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14643243,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(29508923,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011110001" =>
            inv <= conv_std_logic_vector(261663,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14774555,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(147690097,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011110010" =>
            inv <= conv_std_logic_vector(261661,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14905868,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(266859463,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011110011" =>
            inv <= conv_std_logic_vector(261659,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15037183,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(118585591,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011110100" =>
            inv <= conv_std_logic_vector(261657,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15168498,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(239742400,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011110101" =>
            inv <= conv_std_logic_vector(261655,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15299815,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(93464027,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011110110" =>
            inv <= conv_std_logic_vector(261653,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15431132,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(216625411,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011110111" =>
            inv <= conv_std_logic_vector(261651,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15562451,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(72360690,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011111000" =>
            inv <= conv_std_logic_vector(261649,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15693770,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(197542758,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011111001" =>
            inv <= conv_std_logic_vector(261647,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15825091,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(55306773,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011111010" =>
            inv <= conv_std_logic_vector(261645,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15956412,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(182526652,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011111011" =>
            inv <= conv_std_logic_vector(261643,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16087735,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(42335507,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011111100" =>
            inv <= conv_std_logic_vector(261641,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16219058,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(171609300,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011111101" =>
            inv <= conv_std_logic_vector(261639,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16350383,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(33481142,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011111110" =>
            inv <= conv_std_logic_vector(261637,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16481708,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(164824949,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "011111111" =>
            inv <= conv_std_logic_vector(261635,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16613035,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(28774856,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "100000000" =>
            inv <= conv_std_logic_vector(261633,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16744362,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(162205798,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "100000001" =>
            inv <= conv_std_logic_vector(261632,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16405,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(97880094,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100000010" =>
            inv <= conv_std_logic_vector(261630,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(82069,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(232492642,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100000011" =>
            inv <= conv_std_logic_vector(261628,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(147734,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(233414771,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100000100" =>
            inv <= conv_std_logic_vector(261626,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(213400,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(100649515,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100000101" =>
            inv <= conv_std_logic_vector(261624,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(279066,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(102634341,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100000110" =>
            inv <= conv_std_logic_vector(261622,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(344732,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(239370238,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100000111" =>
            inv <= conv_std_logic_vector(261620,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(410399,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(242424784,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100001000" =>
            inv <= conv_std_logic_vector(261618,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(476067,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(111799989,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100001001" =>
            inv <= conv_std_logic_vector(261616,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(541735,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(115933322,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100001010" =>
            inv <= conv_std_logic_vector(261614,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(607403,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(254826281,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100001011" =>
            inv <= conv_std_logic_vector(261612,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(673072,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(260045933,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100001100" =>
            inv <= conv_std_logic_vector(261610,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(738742,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(131594288,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100001101" =>
            inv <= conv_std_logic_vector(261608,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(804412,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(137909323,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100001110" =>
            inv <= conv_std_logic_vector(261606,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(870083,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(10556570,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100001111" =>
            inv <= conv_std_logic_vector(261604,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(935754,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(17974519,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100010000" =>
            inv <= conv_std_logic_vector(261602,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1001425,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(160164667,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100010001" =>
            inv <= conv_std_logic_vector(261600,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1067097,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(168694080,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100010010" =>
            inv <= conv_std_logic_vector(261598,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1132770,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(43564256,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100010011" =>
            inv <= conv_std_logic_vector(261596,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1198443,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(53213172,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100010100" =>
            inv <= conv_std_logic_vector(261594,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1264116,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(197642837,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100010101" =>
            inv <= conv_std_logic_vector(261592,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1329790,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(208419294,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100010110" =>
            inv <= conv_std_logic_vector(261590,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1395465,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(85545574,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100010111" =>
            inv <= conv_std_logic_vector(261588,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1461140,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(97458630,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100011000" =>
            inv <= conv_std_logic_vector(261586,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1526815,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(244160472,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100011001" =>
            inv <= conv_std_logic_vector(261584,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1592491,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(257217653,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100011010" =>
            inv <= conv_std_logic_vector(261582,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1658168,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(136632180,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100011011" =>
            inv <= conv_std_logic_vector(261580,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1723845,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(150842541,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100011100" =>
            inv <= conv_std_logic_vector(261578,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1789523,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(31413754,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100011101" =>
            inv <= conv_std_logic_vector(261576,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1855201,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(46784817,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100011110" =>
            inv <= conv_std_logic_vector(261574,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1920879,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(196956715,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100011111" =>
            inv <= conv_std_logic_vector(261572,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1986558,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(213496513,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100100000" =>
            inv <= conv_std_logic_vector(261570,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2052238,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(96406727,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100100001" =>
            inv <= conv_std_logic_vector(261568,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2117918,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(114123801,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100100010" =>
            inv <= conv_std_logic_vector(261566,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2183598,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(266650763,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100100011" =>
            inv <= conv_std_logic_vector(261564,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2249280,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(17118198,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100100100" =>
            inv <= conv_std_logic_vector(261562,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2314961,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(170834480,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100100101" =>
            inv <= conv_std_logic_vector(261560,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2380643,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(190931217,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100100110" =>
            inv <= conv_std_logic_vector(261558,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2446326,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(77410414,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100100111" =>
            inv <= conv_std_logic_vector(261556,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2512009,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(98709023,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100101000" =>
            inv <= conv_std_logic_vector(261554,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2577692,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(254830073,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100101001" =>
            inv <= conv_std_logic_vector(261552,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2643377,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(8903637,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100101010" =>
            inv <= conv_std_logic_vector(261550,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2709061,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(166239111,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100101011" =>
            inv <= conv_std_logic_vector(261548,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2774746,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(189966567,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100101100" =>
            inv <= conv_std_logic_vector(261546,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2840432,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(80089032,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100101101" =>
            inv <= conv_std_logic_vector(261544,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2906118,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(105043970,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100101110" =>
            inv <= conv_std_logic_vector(261542,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2971804,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(264832874,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100101111" =>
            inv <= conv_std_logic_vector(261540,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3037492,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(22586838,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100110000" =>
            inv <= conv_std_logic_vector(261538,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3103179,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(183615258,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100110001" =>
            inv <= conv_std_logic_vector(261536,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3168867,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(211048205,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100110010" =>
            inv <= conv_std_logic_vector(261534,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3234556,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(104888194,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100110011" =>
            inv <= conv_std_logic_vector(261532,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3300245,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(133573199,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100110100" =>
            inv <= conv_std_logic_vector(261530,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3365935,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(28668746,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100110101" =>
            inv <= conv_std_logic_vector(261528,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3431625,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(58613318,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100110110" =>
            inv <= conv_std_logic_vector(261526,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3497315,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(223408408,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100110111" =>
            inv <= conv_std_logic_vector(261524,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3563006,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(254621075,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100111000" =>
            inv <= conv_std_logic_vector(261522,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3628698,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(152253325,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100111001" =>
            inv <= conv_std_logic_vector(261520,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3694390,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(184742106,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100111010" =>
            inv <= conv_std_logic_vector(261518,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3760083,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(83654478,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100111011" =>
            inv <= conv_std_logic_vector(261516,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3825776,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(117428410,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100111100" =>
            inv <= conv_std_logic_vector(261514,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3891470,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(17629430,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100111101" =>
            inv <= conv_std_logic_vector(261512,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3957164,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(52695507,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100111110" =>
            inv <= conv_std_logic_vector(261510,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4022858,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(222629156,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "100111111" =>
            inv <= conv_std_logic_vector(261508,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4088553,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(258996925,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101000000" =>
            inv <= conv_std_logic_vector(261506,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4154249,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(161800305,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101000001" =>
            inv <= conv_std_logic_vector(261504,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4219945,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(199477266,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101000010" =>
            inv <= conv_std_logic_vector(261502,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4285642,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(103593845,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101000011" =>
            inv <= conv_std_logic_vector(261500,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4351339,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(142588522,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101000100" =>
            inv <= conv_std_logic_vector(261498,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4417037,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(48026823,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101000101" =>
            inv <= conv_std_logic_vector(261496,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4482735,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(88347226,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101000110" =>
            inv <= conv_std_logic_vector(261494,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4548433,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(263551224,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101000111" =>
            inv <= conv_std_logic_vector(261492,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4614133,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(36769906,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101001000" =>
            inv <= conv_std_logic_vector(261490,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4679832,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(213312155,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101001001" =>
            inv <= conv_std_logic_vector(261488,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4745532,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(256309059,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101001010" =>
            inv <= conv_std_logic_vector(261486,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4811233,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(165762621,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101001011" =>
            inv <= conv_std_logic_vector(261484,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4876934,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(210109787,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101001100" =>
            inv <= conv_std_logic_vector(261482,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4942636,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(120917613,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101001101" =>
            inv <= conv_std_logic_vector(261480,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5008338,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(166624068,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101001110" =>
            inv <= conv_std_logic_vector(261478,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5074041,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(78795186,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101001111" =>
            inv <= conv_std_logic_vector(261476,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5139744,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(125868425,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101010000" =>
            inv <= conv_std_logic_vector(261474,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5205448,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(39410329,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101010001" =>
            inv <= conv_std_logic_vector(261472,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5271152,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(87859376,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101010010" =>
            inv <= conv_std_logic_vector(261470,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5336857,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(2781090,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101010011" =>
            inv <= conv_std_logic_vector(261468,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5402562,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(52613438,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101010100" =>
            inv <= conv_std_logic_vector(261466,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5468267,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(237358419,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101010101" =>
            inv <= conv_std_logic_vector(261464,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5533974,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(20147124,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101010110" =>
            inv <= conv_std_logic_vector(261462,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5599680,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(206287919,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101010111" =>
            inv <= conv_std_logic_vector(261460,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5665387,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(258912403,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101011000" =>
            inv <= conv_std_logic_vector(261458,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5731095,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(178022066,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101011001" =>
            inv <= conv_std_logic_vector(261456,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5796803,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(232054873,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101011010" =>
            inv <= conv_std_logic_vector(261454,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5862512,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(152577368,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101011011" =>
            inv <= conv_std_logic_vector(261452,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5928221,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(208027007,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101011100" =>
            inv <= conv_std_logic_vector(261450,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5993931,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(129969822,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101011101" =>
            inv <= conv_std_logic_vector(261448,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6059641,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(186844290,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101011110" =>
            inv <= conv_std_logic_vector(261446,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6125352,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(110216442,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101011111" =>
            inv <= conv_std_logic_vector(261444,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6191063,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(168523735,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101100000" =>
            inv <= conv_std_logic_vector(261442,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6256775,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(93333220,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101100001" =>
            inv <= conv_std_logic_vector(261440,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6322487,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(153082353,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101100010" =>
            inv <= conv_std_logic_vector(261438,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6388200,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(79337165,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101100011" =>
            inv <= conv_std_logic_vector(261436,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6453913,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(140535621,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101100100" =>
            inv <= conv_std_logic_vector(261434,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6519627,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(68244774,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101100101" =>
            inv <= conv_std_logic_vector(261432,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6585341,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(130901057,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101100110" =>
            inv <= conv_std_logic_vector(261430,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6651056,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(60072032,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101100111" =>
            inv <= conv_std_logic_vector(261428,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6716771,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(124194644,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101101000" =>
            inv <= conv_std_logic_vector(261426,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6782487,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(54835943,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101101001" =>
            inv <= conv_std_logic_vector(261424,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6848203,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(120433383,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101101010" =>
            inv <= conv_std_logic_vector(261422,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6913920,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(52552996,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101101011" =>
            inv <= conv_std_logic_vector(261421,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6946778,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(203440839,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101101100" =>
            inv <= conv_std_logic_vector(261419,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7012496,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(69566203,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101101101" =>
            inv <= conv_std_logic_vector(261417,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7078214,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(70654699,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101101110" =>
            inv <= conv_std_logic_vector(261415,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7143932,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(206708322,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101101111" =>
            inv <= conv_std_logic_vector(261413,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7209651,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(209294124,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101110000" =>
            inv <= conv_std_logic_vector(261411,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7275371,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(78413591,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101110001" =>
            inv <= conv_std_logic_vector(261409,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7341091,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(82505197,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101110010" =>
            inv <= conv_std_logic_vector(261407,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7406811,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(221569406,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101110011" =>
            inv <= conv_std_logic_vector(261405,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7472532,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(227174289,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101110100" =>
            inv <= conv_std_logic_vector(261403,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7538254,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(99321843,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101110101" =>
            inv <= conv_std_logic_vector(261401,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7603976,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(106448498,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101110110" =>
            inv <= conv_std_logic_vector(261399,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7669698,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(248557271,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101110111" =>
            inv <= conv_std_logic_vector(261397,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7735421,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(257214192,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101111000" =>
            inv <= conv_std_logic_vector(261395,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7801145,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(132421765,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101111001" =>
            inv <= conv_std_logic_vector(261393,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7866869,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(142616931,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101111010" =>
            inv <= conv_std_logic_vector(261391,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7932594,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(19367251,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101111011" =>
            inv <= conv_std_logic_vector(261389,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7998319,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(31109665,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101111100" =>
            inv <= conv_std_logic_vector(261387,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8064044,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(177846168,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101111101" =>
            inv <= conv_std_logic_vector(261385,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8129770,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(191143299,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101111110" =>
            inv <= conv_std_logic_vector(261383,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8195497,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(71003562,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "101111111" =>
            inv <= conv_std_logic_vector(261381,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8261224,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(85863897,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110000000" =>
            inv <= conv_std_logic_vector(261379,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8326951,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(235726809,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110000001" =>
            inv <= conv_std_logic_vector(261377,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8392679,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(252159347,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110000010" =>
            inv <= conv_std_logic_vector(261375,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8458408,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(135162483,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110000011" =>
            inv <= conv_std_logic_vector(261373,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8524137,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(153174178,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110000100" =>
            inv <= conv_std_logic_vector(261371,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8589867,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(37761480,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110000101" =>
            inv <= conv_std_logic_vector(261369,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8655597,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(57361328,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110000110" =>
            inv <= conv_std_logic_vector(261367,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8721327,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(211976226,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110000111" =>
            inv <= conv_std_logic_vector(261365,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8787058,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(233172711,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110001000" =>
            inv <= conv_std_logic_vector(261363,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8852790,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(120952266,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110001001" =>
            inv <= conv_std_logic_vector(261361,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8918522,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(143753360,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110001010" =>
            inv <= conv_std_logic_vector(261359,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8984255,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(33142020,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110001011" =>
            inv <= conv_std_logic_vector(261357,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9049988,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(57555694,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110001100" =>
            inv <= conv_std_logic_vector(261355,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9115721,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(216996886,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110001101" =>
            inv <= conv_std_logic_vector(261353,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9181455,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(243031622,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110001110" =>
            inv <= conv_std_logic_vector(261351,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9247190,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(135662403,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110001111" =>
            inv <= conv_std_logic_vector(261349,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9312925,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(163326679,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110010000" =>
            inv <= conv_std_logic_vector(261347,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9378661,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(57590984,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110010001" =>
            inv <= conv_std_logic_vector(261345,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9444397,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(86893278,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110010010" =>
            inv <= conv_std_logic_vector(261343,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9510133,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(251234532,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110010011" =>
            inv <= conv_std_logic_vector(261341,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9575871,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(13747355,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110010100" =>
            inv <= conv_std_logic_vector(261339,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9641608,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(179738576,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110010101" =>
            inv <= conv_std_logic_vector(261337,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9707346,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(212340806,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110010110" =>
            inv <= conv_std_logic_vector(261335,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9773085,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(111555525,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110010111" =>
            inv <= conv_std_logic_vector(261333,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9838824,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(145820180,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110011000" =>
            inv <= conv_std_logic_vector(261331,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9904564,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(46701306,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110011001" =>
            inv <= conv_std_logic_vector(261329,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9970304,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(82636350,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110011010" =>
            inv <= conv_std_logic_vector(261327,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10036044,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(253627813,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110011011" =>
            inv <= conv_std_logic_vector(261325,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10101786,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(22806772,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110011100" =>
            inv <= conv_std_logic_vector(261323,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10167527,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(195481587,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110011101" =>
            inv <= conv_std_logic_vector(261321,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10233269,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(234782825,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110011110" =>
            inv <= conv_std_logic_vector(261319,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10299012,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(140713496,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110011111" =>
            inv <= conv_std_logic_vector(261317,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10364755,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(181710537,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110100000" =>
            inv <= conv_std_logic_vector(261315,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10430499,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(89340991,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110100001" =>
            inv <= conv_std_logic_vector(261313,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10496243,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(132041793,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110100010" =>
            inv <= conv_std_logic_vector(261311,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10561988,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(41379987,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110100011" =>
            inv <= conv_std_logic_vector(261309,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10627733,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(85793018,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110100100" =>
            inv <= conv_std_logic_vector(261307,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10693478,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(265282876,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110100101" =>
            inv <= conv_std_logic_vector(261305,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10759225,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(42980638,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110100110" =>
            inv <= conv_std_logic_vector(261303,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10824971,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(224195170,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110100111" =>
            inv <= conv_std_logic_vector(261301,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10890719,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(3621583,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110101000" =>
            inv <= conv_std_logic_vector(261299,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10956466,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(186568744,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110101001" =>
            inv <= conv_std_logic_vector(261297,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11022214,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(236167729,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110101010" =>
            inv <= conv_std_logic_vector(261295,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11087963,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(152420527,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110101011" =>
            inv <= conv_std_logic_vector(261293,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11153712,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(203764581,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110101100" =>
            inv <= conv_std_logic_vector(261291,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11219462,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(121766424,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110101101" =>
            inv <= conv_std_logic_vector(261289,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11285212,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(174864010,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110101110" =>
            inv <= conv_std_logic_vector(261287,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11350963,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(94623359,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110101111" =>
            inv <= conv_std_logic_vector(261285,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11416714,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(149482427,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110110000" =>
            inv <= conv_std_logic_vector(261283,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11482466,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(71008255,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110110001" =>
            inv <= conv_std_logic_vector(261281,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11548218,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(127637265,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110110010" =>
            inv <= conv_std_logic_vector(261279,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11613971,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(50936498,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110110011" =>
            inv <= conv_std_logic_vector(261277,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11679724,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(109344419,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110110100" =>
            inv <= conv_std_logic_vector(261275,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11745478,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(34426028,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110110101" =>
            inv <= conv_std_logic_vector(261273,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11811232,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(94620297,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110110110" =>
            inv <= conv_std_logic_vector(261271,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11876987,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(21492737,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110110111" =>
            inv <= conv_std_logic_vector(261269,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11942742,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(83481301,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110111000" =>
            inv <= conv_std_logic_vector(261267,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12008498,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(12153029,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110111001" =>
            inv <= conv_std_logic_vector(261265,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12074254,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(75944853,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110111010" =>
            inv <= conv_std_logic_vector(261263,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12140011,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(6423814,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110111011" =>
            inv <= conv_std_logic_vector(261261,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12205768,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(72026842,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110111100" =>
            inv <= conv_std_logic_vector(261259,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12271526,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(4320978,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110111101" =>
            inv <= conv_std_logic_vector(261258,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12304405,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(21141383,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110111110" =>
            inv <= conv_std_logic_vector(261256,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12370163,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(156129342,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "110111111" =>
            inv <= conv_std_logic_vector(261254,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12435922,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(157813374,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111000000" =>
            inv <= conv_std_logic_vector(261252,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12501682,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(26195972,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111000001" =>
            inv <= conv_std_logic_vector(261250,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12567442,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(29714068,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111000010" =>
            inv <= conv_std_logic_vector(261248,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12633202,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(168370156,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111000011" =>
            inv <= conv_std_logic_vector(261246,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12698963,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(173730767,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111000100" =>
            inv <= conv_std_logic_vector(261244,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12764725,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(45797884,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111000101" =>
            inv <= conv_std_logic_vector(261242,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12830487,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(53009458,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111000110" =>
            inv <= conv_std_logic_vector(261240,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12896249,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(195366963,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111000111" =>
            inv <= conv_std_logic_vector(261238,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12962012,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(204436928,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111001000" =>
            inv <= conv_std_logic_vector(261236,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13027776,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(80222356,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111001001" =>
            inv <= conv_std_logic_vector(261234,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13093540,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(91159668,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111001010" =>
            inv <= conv_std_logic_vector(261232,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13159304,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(237251358,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111001011" =>
            inv <= conv_std_logic_vector(261230,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13225069,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(250064462,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111001100" =>
            inv <= conv_std_logic_vector(261228,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13290835,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(129600456,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111001101" =>
            inv <= conv_std_logic_vector(261226,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13356601,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(144297287,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111001110" =>
            inv <= conv_std_logic_vector(261224,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13422368,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(25721484,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111001111" =>
            inv <= conv_std_logic_vector(261222,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13488135,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(42309975,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111010000" =>
            inv <= conv_std_logic_vector(261220,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13553902,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(194065764,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111010001" =>
            inv <= conv_std_logic_vector(261218,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13619670,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(212554867,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111010010" =>
            inv <= conv_std_logic_vector(261216,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13685439,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(97779777,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111010011" =>
            inv <= conv_std_logic_vector(261214,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13751208,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(118177423,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111010100" =>
            inv <= conv_std_logic_vector(261212,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13816978,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(5314840,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111010101" =>
            inv <= conv_std_logic_vector(261210,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13882748,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(27629467,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111010110" =>
            inv <= conv_std_logic_vector(261208,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13948518,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(185123287,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111010111" =>
            inv <= conv_std_logic_vector(261206,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14014289,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(209363335,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111011000" =>
            inv <= conv_std_logic_vector(261204,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14080061,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(100351083,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111011001" =>
            inv <= conv_std_logic_vector(261202,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14145833,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(126524479,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111011010" =>
            inv <= conv_std_logic_vector(261200,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14211606,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(19449539,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111011011" =>
            inv <= conv_std_logic_vector(261198,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14277379,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(47564719,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111011100" =>
            inv <= conv_std_logic_vector(261196,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14343152,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(210871490,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111011101" =>
            inv <= conv_std_logic_vector(261194,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14408926,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(240936379,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111011110" =>
            inv <= conv_std_logic_vector(261192,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14474701,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(137761877,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111011111" =>
            inv <= conv_std_logic_vector(261190,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14540476,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(169784908,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111100000" =>
            inv <= conv_std_logic_vector(261188,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14606252,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(68573020,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111100001" =>
            inv <= conv_std_logic_vector(261186,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14672028,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(102562628,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111100010" =>
            inv <= conv_std_logic_vector(261184,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14737805,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(3321276,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111100011" =>
            inv <= conv_std_logic_vector(261182,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14803582,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(39285891,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111100100" =>
            inv <= conv_std_logic_vector(261180,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14869359,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(210458963,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111100101" =>
            inv <= conv_std_logic_vector(261178,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14935137,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(248407016,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111100110" =>
            inv <= conv_std_logic_vector(261176,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15000916,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(153132030,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111100111" =>
            inv <= conv_std_logic_vector(261174,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15066695,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(193071440,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111101000" =>
            inv <= conv_std_logic_vector(261172,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15132475,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(99791770,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111101001" =>
            inv <= conv_std_logic_vector(261170,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15198255,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(141730965,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111101010" =>
            inv <= conv_std_logic_vector(261168,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15264036,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(50455039,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111101011" =>
            inv <= conv_std_logic_vector(261166,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15329817,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(94401937,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111101100" =>
            inv <= conv_std_logic_vector(261164,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15395599,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(5138692,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111101101" =>
            inv <= conv_std_logic_vector(261162,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15461381,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(51101718,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111101110" =>
            inv <= conv_std_logic_vector(261160,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15527163,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(232294014,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111101111" =>
            inv <= conv_std_logic_vector(261158,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15592947,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(11846647,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111110000" =>
            inv <= conv_std_logic_vector(261156,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15658730,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(195067454,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111110001" =>
            inv <= conv_std_logic_vector(261154,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15724514,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(245088520,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111110010" =>
            inv <= conv_std_logic_vector(261152,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15790299,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(161910803,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111110011" =>
            inv <= conv_std_logic_vector(261150,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15856084,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(213972758,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111110100" =>
            inv <= conv_std_logic_vector(261148,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15921870,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(132840397,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111110101" =>
            inv <= conv_std_logic_vector(261146,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15987656,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(186951663,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111110110" =>
            inv <= conv_std_logic_vector(261144,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16053443,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(107873077,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111110111" =>
            inv <= conv_std_logic_vector(261142,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16119230,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(164042073,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111111000" =>
            inv <= conv_std_logic_vector(261140,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16185018,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(87025173,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111111001" =>
            inv <= conv_std_logic_vector(261138,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16250806,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(145260319,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111111010" =>
            inv <= conv_std_logic_vector(261136,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16316595,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(70314033,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111111011" =>
            inv <= conv_std_logic_vector(261134,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16382384,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(130623237,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111111100" =>
            inv <= conv_std_logic_vector(261132,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16448174,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(57754962,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111111101" =>
            inv <= conv_std_logic_vector(261130,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16513964,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(120146640,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111111110" =>
            inv <= conv_std_logic_vector(261128,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16579755,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(49365303,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "111111111" =>
            inv <= conv_std_logic_vector(261126,18);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16645546,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(113847871,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN others =>
           inv <= conv_std_logic_vector(0,18);
           logman(52 DOWNTO 29) <= conv_std_logic_vector(0,24);
           logman(28 DOWNTO 1) <= conv_std_logic_vector(0,28);
           logexp <= conv_std_logic_vector(0,11);
    END CASE;
  END PROCESS;

END rtl;
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   DP_LNLUT9.VHD                             ***
--***                                             ***
--***   Function: Look Up Table - LN()            ***
--***                                             ***
--***   Generated by MATLAB Utility               ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_lnlut9 IS
PORT (
      add : IN STD_LOGIC_VECTOR (9 DOWNTO 1);
      inv : OUT STD_LOGIC_VECTOR (12 DOWNTO 1);
      logman : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
      logexp : OUT STD_LOGIC_VECTOR (11 DOWNTO 1)
     );
END dp_lnlut9;

ARCHITECTURE rtl OF dp_lnlut9 IS

BEGIN

  pca: PROCESS (add)
  BEGIN
    CASE add IS
      WHEN "000000000" =>
            inv <= conv_std_logic_vector(2048,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(0,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(0,28);
            logexp <= conv_std_logic_vector(0,11);
      WHEN "000000001" =>
            inv <= conv_std_logic_vector(4089,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12608028,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(166435551,28);
            logexp <= conv_std_logic_vector(1013,11);
      WHEN "000000010" =>
            inv <= conv_std_logic_vector(4081,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14737805,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(3321276,28);
            logexp <= conv_std_logic_vector(1014,11);
      WHEN "000000011" =>
            inv <= conv_std_logic_vector(4073,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7407998,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(148040387,28);
            logexp <= conv_std_logic_vector(1015,11);
      WHEN "000000100" =>
            inv <= conv_std_logic_vector(4065,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15852272,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(51070306,28);
            logexp <= conv_std_logic_vector(1015,11);
      WHEN "000000101" =>
            inv <= conv_std_logic_vector(4057,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3767982,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(94668708,28);
            logexp <= conv_std_logic_vector(1016,11);
      WHEN "000000110" =>
            inv <= conv_std_logic_vector(4049,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8006786,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(237055061,28);
            logexp <= conv_std_logic_vector(1016,11);
      WHEN "000000111" =>
            inv <= conv_std_logic_vector(4041,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12253974,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(192188802,28);
            logexp <= conv_std_logic_vector(1016,11);
      WHEN "000001000" =>
            inv <= conv_std_logic_vector(4033,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16509579,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(20710393,28);
            logexp <= conv_std_logic_vector(1016,11);
      WHEN "000001001" =>
            inv <= conv_std_logic_vector(4026,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1731473,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(180827014,28);
            logexp <= conv_std_logic_vector(1017,11);
      WHEN "000001010" =>
            inv <= conv_std_logic_vector(4018,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3867211,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(126637664,28);
            logexp <= conv_std_logic_vector(1017,11);
      WHEN "000001011" =>
            inv <= conv_std_logic_vector(4010,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6007205,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(228245542,28);
            logexp <= conv_std_logic_vector(1017,11);
      WHEN "000001100" =>
            inv <= conv_std_logic_vector(4003,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7883206,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(5368567,28);
            logexp <= conv_std_logic_vector(1017,11);
      WHEN "000001101" =>
            inv <= conv_std_logic_vector(3995,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10031227,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(104563152,28);
            logexp <= conv_std_logic_vector(1017,11);
      WHEN "000001110" =>
            inv <= conv_std_logic_vector(3987,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12183554,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(132223343,28);
            logexp <= conv_std_logic_vector(1017,11);
      WHEN "000001111" =>
            inv <= conv_std_logic_vector(3980,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14070386,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(93820959,28);
            logexp <= conv_std_logic_vector(1017,11);
      WHEN "000010000" =>
            inv <= conv_std_logic_vector(3972,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16230833,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(108537941,28);
            logexp <= conv_std_logic_vector(1017,11);
      WHEN "000010001" =>
            inv <= conv_std_logic_vector(3965,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(673790,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(140554826,28);
            logexp <= conv_std_logic_vector(1018,11);
      WHEN "000010010" =>
            inv <= conv_std_logic_vector(3957,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1758104,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(208459132,28);
            logexp <= conv_std_logic_vector(1018,11);
      WHEN "000010011" =>
            inv <= conv_std_logic_vector(3950,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2708679,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(147574307,28);
            logexp <= conv_std_logic_vector(1018,11);
      WHEN "000010100" =>
            inv <= conv_std_logic_vector(3943,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3660940,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(102190772,28);
            logexp <= conv_std_logic_vector(1018,11);
      WHEN "000010101" =>
            inv <= conv_std_logic_vector(3935,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4751310,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(193668840,28);
            logexp <= conv_std_logic_vector(1018,11);
      WHEN "000010110" =>
            inv <= conv_std_logic_vector(3928,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5707204,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(201576161,28);
            logexp <= conv_std_logic_vector(1018,11);
      WHEN "000010111" =>
            inv <= conv_std_logic_vector(3920,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6801743,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(47496037,28);
            logexp <= conv_std_logic_vector(1018,11);
      WHEN "000011000" =>
            inv <= conv_std_logic_vector(3913,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7761298,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(63049717,28);
            logexp <= conv_std_logic_vector(1018,11);
      WHEN "000011001" =>
            inv <= conv_std_logic_vector(3906,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8722571,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(103870568,28);
            logexp <= conv_std_logic_vector(1018,11);
      WHEN "000011010" =>
            inv <= conv_std_logic_vector(3899,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9685568,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(213866899,28);
            logexp <= conv_std_logic_vector(1018,11);
      WHEN "000011011" =>
            inv <= conv_std_logic_vector(3891,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10788256,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(148111271,28);
            logexp <= conv_std_logic_vector(1018,11);
      WHEN "000011100" =>
            inv <= conv_std_logic_vector(3884,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11754969,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(190364328,28);
            logexp <= conv_std_logic_vector(1018,11);
      WHEN "000011101" =>
            inv <= conv_std_logic_vector(3877,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12723426,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(191372810,28);
            logexp <= conv_std_logic_vector(1018,11);
      WHEN "000011110" =>
            inv <= conv_std_logic_vector(3870,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13693633,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(232417040,28);
            logexp <= conv_std_logic_vector(1018,11);
      WHEN "000011111" =>
            inv <= conv_std_logic_vector(3863,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14665597,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(135531172,28);
            logexp <= conv_std_logic_vector(1018,11);
      WHEN "000100000" =>
            inv <= conv_std_logic_vector(3856,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15639324,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(440444,28);
            logexp <= conv_std_logic_vector(1018,11);
      WHEN "000100001" =>
            inv <= conv_std_logic_vector(3848,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16754321,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(28021513,28);
            logexp <= conv_std_logic_vector(1018,11);
      WHEN "000100010" =>
            inv <= conv_std_logic_vector(3841,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(477315,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(103375890,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000100011" =>
            inv <= conv_std_logic_vector(3834,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(966969,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(207463933,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000100100" =>
            inv <= conv_std_logic_vector(3827,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1457518,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(261454332,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000100101" =>
            inv <= conv_std_logic_vector(3820,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1948966,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(71112978,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000100110" =>
            inv <= conv_std_logic_vector(3814,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2370924,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(27626077,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000100111" =>
            inv <= conv_std_logic_vector(3807,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2864048,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(7790664,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000101000" =>
            inv <= conv_std_logic_vector(3800,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3358079,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(135806794,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000101001" =>
            inv <= conv_std_logic_vector(3793,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3853021,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(236303861,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000101010" =>
            inv <= conv_std_logic_vector(3786,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4348878,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(138889654,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000101011" =>
            inv <= conv_std_logic_vector(3779,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4845652,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(215058204,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000101100" =>
            inv <= conv_std_logic_vector(3772,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5343348,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(36049681,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000101101" =>
            inv <= conv_std_logic_vector(3766,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5770679,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(216749821,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000101110" =>
            inv <= conv_std_logic_vector(3759,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6270094,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(202231188,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000101111" =>
            inv <= conv_std_logic_vector(3752,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6770440,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(154557048,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000110000" =>
            inv <= conv_std_logic_vector(3745,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7271720,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(201681452,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000110001" =>
            inv <= conv_std_logic_vector(3739,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7702135,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(212518450,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000110010" =>
            inv <= conv_std_logic_vector(3732,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8205160,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(130192328,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000110011" =>
            inv <= conv_std_logic_vector(3725,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8709129,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(153765892,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000110100" =>
            inv <= conv_std_logic_vector(3719,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9141857,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(115454106,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000110101" =>
            inv <= conv_std_logic_vector(3712,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9647589,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(223955336,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000110110" =>
            inv <= conv_std_logic_vector(3706,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10081834,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(106871151,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000110111" =>
            inv <= conv_std_logic_vector(3699,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10589342,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(134545541,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000111000" =>
            inv <= conv_std_logic_vector(3693,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11025114,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(118400992,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000111001" =>
            inv <= conv_std_logic_vector(3686,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11534410,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(203065005,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000111010" =>
            inv <= conv_std_logic_vector(3680,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11971720,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(229464861,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000111011" =>
            inv <= conv_std_logic_vector(3673,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12482818,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(7696520,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000111100" =>
            inv <= conv_std_logic_vector(3667,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12921677,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(49003431,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000111101" =>
            inv <= conv_std_logic_vector(3660,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13434587,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(267260840,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000111110" =>
            inv <= conv_std_logic_vector(3654,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13875007,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(58597277,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "000111111" =>
            inv <= conv_std_logic_vector(3648,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14316150,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(59000478,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "001000000" =>
            inv <= conv_std_logic_vector(3641,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14831735,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(2814011,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "001000001" =>
            inv <= conv_std_logic_vector(3635,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15274454,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(104571506,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "001000010" =>
            inv <= conv_std_logic_vector(3629,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15717905,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(35857837,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "001000011" =>
            inv <= conv_std_logic_vector(3623,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16162089,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(177959810,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "001000100" =>
            inv <= conv_std_logic_vector(3616,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16681235,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(165401956,28);
            logexp <= conv_std_logic_vector(1019,11);
      WHEN "001000101" =>
            inv <= conv_std_logic_vector(3610,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(174901,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(50275830,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001000110" =>
            inv <= conv_std_logic_vector(3604,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(398163,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(88951577,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001000111" =>
            inv <= conv_std_logic_vector(3598,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(621797,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(127737931,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001001000" =>
            inv <= conv_std_logic_vector(3592,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(845804,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(231522955,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001001001" =>
            inv <= conv_std_logic_vector(3585,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1107620,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(57821111,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001001010" =>
            inv <= conv_std_logic_vector(3579,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1332440,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(156464157,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001001011" =>
            inv <= conv_std_logic_vector(3573,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1557638,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(44535294,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001001100" =>
            inv <= conv_std_logic_vector(3567,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1783214,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(62397887,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001001101" =>
            inv <= conv_std_logic_vector(3561,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2009170,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(15263403,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001001110" =>
            inv <= conv_std_logic_vector(3555,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2235506,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(246944822,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001001111" =>
            inv <= conv_std_logic_vector(3549,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2462226,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(29255593,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001010000" =>
            inv <= conv_std_logic_vector(3543,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2689328,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(246376003,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001010001" =>
            inv <= conv_std_logic_vector(3537,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2916816,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(173639564,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001010010" =>
            inv <= conv_std_logic_vector(3531,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3144690,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(161899610,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001010011" =>
            inv <= conv_std_logic_vector(3525,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3372952,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(26928617,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001010100" =>
            inv <= conv_std_logic_vector(3519,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3601602,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(123172243,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001010101" =>
            inv <= conv_std_logic_vector(3513,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3830643,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(1584354,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001010110" =>
            inv <= conv_std_logic_vector(3507,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4060075,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(20252153,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001010111" =>
            inv <= conv_std_logic_vector(3502,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4251568,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(137854980,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001011000" =>
            inv <= conv_std_logic_vector(3496,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4481721,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(231322588,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001011001" =>
            inv <= conv_std_logic_vector(3490,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4712270,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(147480442,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001011010" =>
            inv <= conv_std_logic_vector(3484,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4943215,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(251536037,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001011011" =>
            inv <= conv_std_logic_vector(3478,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5174559,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(105278949,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001011100" =>
            inv <= conv_std_logic_vector(3473,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5367650,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(181375864,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001011101" =>
            inv <= conv_std_logic_vector(3467,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5599727,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(133308340,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001011110" =>
            inv <= conv_std_logic_vector(3461,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5832206,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(80096944,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001011111" =>
            inv <= conv_std_logic_vector(3455,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6065088,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(127763081,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001100000" =>
            inv <= conv_std_logic_vector(3450,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6259466,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(27642512,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001100001" =>
            inv <= conv_std_logic_vector(3444,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6493091,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(120806774,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001100010" =>
            inv <= conv_std_logic_vector(3438,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6727124,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(44281139,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001100011" =>
            inv <= conv_std_logic_vector(3433,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6922463,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(171170237,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001100100" =>
            inv <= conv_std_logic_vector(3427,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7157246,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(240302137,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001100101" =>
            inv <= conv_std_logic_vector(3422,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7353213,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(222094360,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001100110" =>
            inv <= conv_std_logic_vector(3416,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7588752,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(122671437,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001100111" =>
            inv <= conv_std_logic_vector(3411,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7785350,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(239607246,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001101000" =>
            inv <= conv_std_logic_vector(3405,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8021649,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(206841234,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001101001" =>
            inv <= conv_std_logic_vector(3399,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8258365,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(107795018,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001101010" =>
            inv <= conv_std_logic_vector(3394,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8455947,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(226201607,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001101011" =>
            inv <= conv_std_logic_vector(3388,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8693431,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(94327085,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001101100" =>
            inv <= conv_std_logic_vector(3383,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8891655,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(206124156,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001101101" =>
            inv <= conv_std_logic_vector(3378,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9090173,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(99984141,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001101110" =>
            inv <= conv_std_logic_vector(3372,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9328782,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(195833281,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001101111" =>
            inv <= conv_std_logic_vector(3367,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9527948,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(110283065,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001110000" =>
            inv <= conv_std_logic_vector(3361,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9767338,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(282511,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001110001" =>
            inv <= conv_std_logic_vector(3356,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9967156,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(1157748,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001110010" =>
            inv <= conv_std_logic_vector(3351,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10167271,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(250247631,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001110011" =>
            inv <= conv_std_logic_vector(3345,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10407805,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(150148144,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001110100" =>
            inv <= conv_std_logic_vector(3340,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10608580,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(15841264,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001110101" =>
            inv <= conv_std_logic_vector(3335,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10809655,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(92492368,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001110110" =>
            inv <= conv_std_logic_vector(3329,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11051343,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(267282110,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001110111" =>
            inv <= conv_std_logic_vector(3324,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11253084,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(51811246,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001111000" =>
            inv <= conv_std_logic_vector(3319,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11455128,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(21159361,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001111001" =>
            inv <= conv_std_logic_vector(3314,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11657476,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(152694737,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001111010" =>
            inv <= conv_std_logic_vector(3308,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11900698,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(34843865,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001111011" =>
            inv <= conv_std_logic_vector(3303,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12103719,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(266488285,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001111100" =>
            inv <= conv_std_logic_vector(3298,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12307049,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(112230017,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001111101" =>
            inv <= conv_std_logic_vector(3293,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12510687,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(91030082,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001111110" =>
            inv <= conv_std_logic_vector(3288,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12714634,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(186120630,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "001111111" =>
            inv <= conv_std_logic_vector(3282,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12959781,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(79635368,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "010000000" =>
            inv <= conv_std_logic_vector(3277,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13164412,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(194678646,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "010000001" =>
            inv <= conv_std_logic_vector(3272,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13369356,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(165362770,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "010000010" =>
            inv <= conv_std_logic_vector(3267,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13574613,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(248228452,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "010000011" =>
            inv <= conv_std_logic_vector(3262,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13780185,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(164124274,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "010000100" =>
            inv <= conv_std_logic_vector(3257,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13986072,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(171955743,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "010000101" =>
            inv <= conv_std_logic_vector(3252,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14192275,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(263386193,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "010000110" =>
            inv <= conv_std_logic_vector(3247,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14398796,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(162844158,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "010000111" =>
            inv <= conv_std_logic_vector(3242,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14605635,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(132837122,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "010001000" =>
            inv <= conv_std_logic_vector(3237,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14812793,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(168652610,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "010001001" =>
            inv <= conv_std_logic_vector(3232,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15020271,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(266801170,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "010001010" =>
            inv <= conv_std_logic_vector(3227,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15228071,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(156588484,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "010001011" =>
            inv <= conv_std_logic_vector(3222,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15436193,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(105429361,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "010001100" =>
            inv <= conv_std_logic_vector(3217,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15644638,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(113549080,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "010001101" =>
            inv <= conv_std_logic_vector(3212,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15853407,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(182426590,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "010001110" =>
            inv <= conv_std_logic_vector(3207,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16062502,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(46366848,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "010001111" =>
            inv <= conv_std_logic_vector(3202,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16271922,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(246250548,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "010010000" =>
            inv <= conv_std_logic_vector(3197,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16481670,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(250493842,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "010010001" =>
            inv <= conv_std_logic_vector(3193,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16649705,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(179677631,28);
            logexp <= conv_std_logic_vector(1020,11);
      WHEN "010010010" =>
            inv <= conv_std_logic_vector(3188,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(41414,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(182297714,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010010011" =>
            inv <= conv_std_logic_vector(3183,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(146749,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(160926493,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010010100" =>
            inv <= conv_std_logic_vector(3178,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(252250,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(30832263,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010010101" =>
            inv <= conv_std_logic_vector(3173,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(357916,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(200433438,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010010110" =>
            inv <= conv_std_logic_vector(3168,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(463750,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(5068900,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010010111" =>
            inv <= conv_std_logic_vector(3164,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(548536,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(260761497,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010011000" =>
            inv <= conv_std_logic_vector(3159,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(654671,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(140824337,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010011001" =>
            inv <= conv_std_logic_vector(3154,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(760974,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(53287185,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010011010" =>
            inv <= conv_std_logic_vector(3149,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(867445,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(141350373,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010011011" =>
            inv <= conv_std_logic_vector(3145,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(952744,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(102039527,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010011100" =>
            inv <= conv_std_logic_vector(3140,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1059520,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(171297819,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010011101" =>
            inv <= conv_std_logic_vector(3135,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1166467,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(15456691,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010011110" =>
            inv <= conv_std_logic_vector(3131,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1252147,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(19951762,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010011111" =>
            inv <= conv_std_logic_vector(3126,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1359401,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(41610452,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010100000" =>
            inv <= conv_std_logic_vector(3121,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1466826,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(248224675,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010100001" =>
            inv <= conv_std_logic_vector(3117,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1552891,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(141314514,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010100010" =>
            inv <= conv_std_logic_vector(3112,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1660627,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(194757369,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010100011" =>
            inv <= conv_std_logic_vector(3107,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1768537,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(43450957,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010100100" =>
            inv <= conv_std_logic_vector(3103,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1854989,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(219219906,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010100101" =>
            inv <= conv_std_logic_vector(3098,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1963212,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(131015724,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010100110" =>
            inv <= conv_std_logic_vector(3094,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2049916,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(123155162,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010100111" =>
            inv <= conv_std_logic_vector(3089,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2158454,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(50751187,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010101000" =>
            inv <= conv_std_logic_vector(3085,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2245410,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(252626322,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010101001" =>
            inv <= conv_std_logic_vector(3080,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2354265,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(153008713,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010101010" =>
            inv <= conv_std_logic_vector(3076,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2441476,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(156128968,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010101011" =>
            inv <= conv_std_logic_vector(3071,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2550649,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(259057771,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010101100" =>
            inv <= conv_std_logic_vector(3067,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2638116,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(195294519,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010101101" =>
            inv <= conv_std_logic_vector(3062,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2747610,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(198048260,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010101110" =>
            inv <= conv_std_logic_vector(3058,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2835334,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(202805005,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010101111" =>
            inv <= conv_std_logic_vector(3053,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2945151,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(75538772,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010110000" =>
            inv <= conv_std_logic_vector(3049,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3033134,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(19357354,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010110001" =>
            inv <= conv_std_logic_vector(3044,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3143275,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(5155285,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010110010" =>
            inv <= conv_std_logic_vector(3040,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3231518,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(30629091,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010110011" =>
            inv <= conv_std_logic_vector(3035,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3341985,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(108686704,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010110100" =>
            inv <= conv_std_logic_vector(3031,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3430490,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(93632684,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010110101" =>
            inv <= conv_std_logic_vector(3027,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3519112,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(45511961,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010110110" =>
            inv <= conv_std_logic_vector(3022,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3630054,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(73684067,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010110111" =>
            inv <= conv_std_logic_vector(3018,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3718940,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(53706357,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010111000" =>
            inv <= conv_std_logic_vector(3014,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3807944,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(3094116,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010111001" =>
            inv <= conv_std_logic_vector(3009,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3919365,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(8048359,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010111010" =>
            inv <= conv_std_logic_vector(3005,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4008635,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(62108895,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010111011" =>
            inv <= conv_std_logic_vector(3001,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4098024,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(91490091,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010111100" =>
            inv <= conv_std_logic_vector(2996,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4209928,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(114206619,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010111101" =>
            inv <= conv_std_logic_vector(2992,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4299586,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(64350406,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010111110" =>
            inv <= conv_std_logic_vector(2988,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4389363,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(267789889,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "010111111" =>
            inv <= conv_std_logic_vector(2984,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4479262,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(5480265,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011000000" =>
            inv <= conv_std_logic_vector(2979,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4591804,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(43802136,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011000001" =>
            inv <= conv_std_logic_vector(2975,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4681973,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(258711462,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011000010" =>
            inv <= conv_std_logic_vector(2971,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4772265,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(22193356,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011000011" =>
            inv <= conv_std_logic_vector(2967,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4862677,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(227303994,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011000100" =>
            inv <= conv_std_logic_vector(2963,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4953212,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(156841963,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011000101" =>
            inv <= conv_std_logic_vector(2958,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5066553,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(8978848,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011000110" =>
            inv <= conv_std_logic_vector(2954,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5157363,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(112226691,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011000111" =>
            inv <= conv_std_logic_vector(2950,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5248296,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(228718953,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011001000" =>
            inv <= conv_std_logic_vector(2946,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5339353,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(179656048,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011001001" =>
            inv <= conv_std_logic_vector(2942,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5430534,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(55039221,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011001010" =>
            inv <= conv_std_logic_vector(2938,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5521838,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(213672522,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011001011" =>
            inv <= conv_std_logic_vector(2934,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5613267,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(209422987,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011001100" =>
            inv <= conv_std_logic_vector(2929,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5727729,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(122280556,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011001101" =>
            inv <= conv_std_logic_vector(2925,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5819439,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(152340981,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011001110" =>
            inv <= conv_std_logic_vector(2921,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5911275,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(48556746,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011001111" =>
            inv <= conv_std_logic_vector(2917,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6003236,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(171693667,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011010000" =>
            inv <= conv_std_logic_vector(2913,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6095324,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(77591273,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011010001" =>
            inv <= conv_std_logic_vector(2909,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6187538,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(127777649,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011010010" =>
            inv <= conv_std_logic_vector(2905,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6279879,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(147294249,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011010011" =>
            inv <= conv_std_logic_vector(2901,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6372347,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(230004385,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011010100" =>
            inv <= conv_std_logic_vector(2897,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6464943,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(201724446,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011010101" =>
            inv <= conv_std_logic_vector(2893,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6557667,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(157096962,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011010110" =>
            inv <= conv_std_logic_vector(2889,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6650519,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(191157304,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011010111" =>
            inv <= conv_std_logic_vector(2885,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6743500,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(130900404,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011011000" =>
            inv <= conv_std_logic_vector(2881,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6836610,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(72153870,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011011001" =>
            inv <= conv_std_logic_vector(2877,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6929849,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(111144728,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011011010" =>
            inv <= conv_std_logic_vector(2873,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7023218,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(76066192,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011011011" =>
            inv <= conv_std_logic_vector(2869,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7116717,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(63950809,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011011100" =>
            inv <= conv_std_logic_vector(2865,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7210346,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(172237270,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011011101" =>
            inv <= conv_std_logic_vector(2862,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7280654,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(139653305,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011011110" =>
            inv <= conv_std_logic_vector(2858,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7374513,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(23245886,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011011111" =>
            inv <= conv_std_logic_vector(2854,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7468503,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(28873967,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011100000" =>
            inv <= conv_std_logic_vector(2850,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7562624,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(255519588,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011100001" =>
            inv <= conv_std_logic_vector(2846,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7656878,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(265710940,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011100010" =>
            inv <= conv_std_logic_vector(2842,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7751265,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(159266526,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011100011" =>
            inv <= conv_std_logic_vector(2838,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7845785,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(36426622,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011100100" =>
            inv <= conv_std_logic_vector(2834,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7940437,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(266291107,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011100101" =>
            inv <= conv_std_logic_vector(2831,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8011515,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(93413946,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011100110" =>
            inv <= conv_std_logic_vector(2827,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8106402,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(110277380,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011100111" =>
            inv <= conv_std_logic_vector(2823,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8201423,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(222008092,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011101000" =>
            inv <= conv_std_logic_vector(2819,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8296579,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(262447083,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011101001" =>
            inv <= conv_std_logic_vector(2815,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8391871,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(65871042,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011101010" =>
            inv <= conv_std_logic_vector(2812,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8463428,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(160477028,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011101011" =>
            inv <= conv_std_logic_vector(2808,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8558957,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(66030540,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011101100" =>
            inv <= conv_std_logic_vector(2804,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8654622,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(19294193,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011101101" =>
            inv <= conv_std_logic_vector(2800,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8750423,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(124636155,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011101110" =>
            inv <= conv_std_logic_vector(2797,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8822364,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(98044902,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011101111" =>
            inv <= conv_std_logic_vector(2793,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8918405,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(185136678,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011110000" =>
            inv <= conv_std_logic_vector(2789,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9014584,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(176764031,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011110001" =>
            inv <= conv_std_logic_vector(2786,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9086809,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(121288912,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011110010" =>
            inv <= conv_std_logic_vector(2782,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9183230,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(67117648,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011110011" =>
            inv <= conv_std_logic_vector(2778,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9279789,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(210248932,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011110100" =>
            inv <= conv_std_logic_vector(2775,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9352300,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(192854718,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011110101" =>
            inv <= conv_std_logic_vector(2771,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9449104,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(269037,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011110110" =>
            inv <= conv_std_logic_vector(2767,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9546047,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(32810921,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011110111" =>
            inv <= conv_std_logic_vector(2764,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9618846,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(127667797,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011111000" =>
            inv <= conv_std_logic_vector(2760,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9716035,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(77607514,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011111001" =>
            inv <= conv_std_logic_vector(2756,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9813365,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(15613650,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011111010" =>
            inv <= conv_std_logic_vector(2753,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9886455,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(35776871,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011111011" =>
            inv <= conv_std_logic_vector(2749,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9984032,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(150556503,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011111100" =>
            inv <= conv_std_logic_vector(2745,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10081752,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(19947644,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011111101" =>
            inv <= conv_std_logic_vector(2742,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10155135,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(54345836,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011111110" =>
            inv <= conv_std_logic_vector(2738,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10253104,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(97812156,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "011111111" =>
            inv <= conv_std_logic_vector(2735,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10326675,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(55696655,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100000000" =>
            inv <= conv_std_logic_vector(2731,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10424895,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(79654305,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100000001" =>
            inv <= conv_std_logic_vector(2728,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10498654,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(219479460,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100000010" =>
            inv <= conv_std_logic_vector(2724,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10597127,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(32989146,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100000011" =>
            inv <= conv_std_logic_vector(2721,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10671076,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(78331980,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100000100" =>
            inv <= conv_std_logic_vector(2717,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10769802,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(29997091,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100000101" =>
            inv <= conv_std_logic_vector(2714,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10843941,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(243319683,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100000110" =>
            inv <= conv_std_logic_vector(2710,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10942922,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(147572067,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100000111" =>
            inv <= conv_std_logic_vector(2707,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11017253,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(256500550,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100001000" =>
            inv <= conv_std_logic_vector(2703,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11116490,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(198934815,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100001001" =>
            inv <= conv_std_logic_vector(2700,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11191014,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(201586837,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100001010" =>
            inv <= conv_std_logic_vector(2696,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11290509,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(2117744,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100001011" =>
            inv <= conv_std_logic_vector(2693,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11365226,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(167123833,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100001100" =>
            inv <= conv_std_logic_vector(2689,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11464979,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(185321336,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100001101" =>
            inv <= conv_std_logic_vector(2686,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11539891,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(246540176,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100001110" =>
            inv <= conv_std_logic_vector(2682,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11639905,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(39481193,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100001111" =>
            inv <= conv_std_logic_vector(2679,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11715013,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(1327916,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100010000" =>
            inv <= conv_std_logic_vector(2675,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11815287,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(202673946,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100010001" =>
            inv <= conv_std_logic_vector(2672,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11890592,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(71706890,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100010010" =>
            inv <= conv_std_logic_vector(2669,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11965981,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(100723928,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100010011" =>
            inv <= conv_std_logic_vector(2665,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12066632,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(29193386,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100010100" =>
            inv <= conv_std_logic_vector(2662,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12142219,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(93571958,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100010101" =>
            inv <= conv_std_logic_vector(2658,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12243134,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(255701348,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100010110" =>
            inv <= conv_std_logic_vector(2655,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12318921,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(98863551,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100010111" =>
            inv <= conv_std_logic_vector(2652,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12394793,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(125312048,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100011000" =>
            inv <= conv_std_logic_vector(2648,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12496089,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(237443793,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100011001" =>
            inv <= conv_std_logic_vector(2645,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12572162,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(178518688,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100011010" =>
            inv <= conv_std_logic_vector(2642,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12648321,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(208688605,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100011011" =>
            inv <= conv_std_logic_vector(2638,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12750001,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(239940349,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100011100" =>
            inv <= conv_std_logic_vector(2635,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12826363,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(56746753,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100011101" =>
            inv <= conv_std_logic_vector(2632,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12902811,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(138879938,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100011110" =>
            inv <= conv_std_logic_vector(2629,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12979347,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(2730614,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100011111" =>
            inv <= conv_std_logic_vector(2625,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13081530,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(81091197,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100100000" =>
            inv <= conv_std_logic_vector(2622,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13158270,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(1684866,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100100001" =>
            inv <= conv_std_logic_vector(2619,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13235097,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(151292526,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100100010" =>
            inv <= conv_std_logic_vector(2615,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13337671,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(84646293,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100100011" =>
            inv <= conv_std_logic_vector(2612,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13414704,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(173861808,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100100100" =>
            inv <= conv_std_logic_vector(2609,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13491826,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(136139682,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100100101" =>
            inv <= conv_std_logic_vector(2606,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13569037,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(26161775,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100100110" =>
            inv <= conv_std_logic_vector(2602,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13672122,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(249732568,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100100111" =>
            inv <= conv_std_logic_vector(2599,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13749541,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(95394098,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100101000" =>
            inv <= conv_std_logic_vector(2596,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13827049,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(52442312,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100101001" =>
            inv <= conv_std_logic_vector(2593,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13904646,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(176384205,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100101010" =>
            inv <= conv_std_logic_vector(2590,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13982333,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(254484090,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100101011" =>
            inv <= conv_std_logic_vector(2586,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14086057,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(26027470,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100101100" =>
            inv <= conv_std_logic_vector(2583,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14163954,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(214862414,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100101101" =>
            inv <= conv_std_logic_vector(2580,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14241943,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(8054063,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100101110" =>
            inv <= conv_std_logic_vector(2577,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14320021,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(267454282,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100101111" =>
            inv <= conv_std_logic_vector(2574,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14398191,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(244499796,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100110000" =>
            inv <= conv_std_logic_vector(2571,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14476452,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(264567670,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100110001" =>
            inv <= conv_std_logic_vector(2567,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14580943,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(69299566,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100110010" =>
            inv <= conv_std_logic_vector(2564,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14659417,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(233357662,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100110011" =>
            inv <= conv_std_logic_vector(2561,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14737984,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(94818262,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100110100" =>
            inv <= conv_std_logic_vector(2558,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14816642,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(248364916,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100110101" =>
            inv <= conv_std_logic_vector(2555,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14895393,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(215142880,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100110110" =>
            inv <= conv_std_logic_vector(2552,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14974237,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(53372798,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100110111" =>
            inv <= conv_std_logic_vector(2549,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15053173,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(89916221,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100111000" =>
            inv <= conv_std_logic_vector(2546,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15132202,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(114970198,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100111001" =>
            inv <= conv_std_logic_vector(2543,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15211324,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(187374614,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100111010" =>
            inv <= conv_std_logic_vector(2539,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15316966,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(101744986,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100111011" =>
            inv <= conv_std_logic_vector(2536,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15396306,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(246192396,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100111100" =>
            inv <= conv_std_logic_vector(2533,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15475741,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(98762703,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100111101" =>
            inv <= conv_std_logic_vector(2530,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15555269,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(256076770,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100111110" =>
            inv <= conv_std_logic_vector(2527,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15634892,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(241226312,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "100111111" =>
            inv <= conv_std_logic_vector(2524,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15714610,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(114387642,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "101000000" =>
            inv <= conv_std_logic_vector(2521,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15794422,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(204387226,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "101000001" =>
            inv <= conv_std_logic_vector(2518,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15874330,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(34960895,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "101000010" =>
            inv <= conv_std_logic_vector(2515,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15954332,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(203803056,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "101000011" =>
            inv <= conv_std_logic_vector(2512,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16034430,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(235084078,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "101000100" =>
            inv <= conv_std_logic_vector(2509,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16114624,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(190064071,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "101000101" =>
            inv <= conv_std_logic_vector(2506,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16194914,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(130223025,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "101000110" =>
            inv <= conv_std_logic_vector(2503,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16275300,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(117261858,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "101000111" =>
            inv <= conv_std_logic_vector(2500,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16355782,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(213103482,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "101001000" =>
            inv <= conv_std_logic_vector(2497,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16436361,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(211458404,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "101001001" =>
            inv <= conv_std_logic_vector(2494,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16517037,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(174696720,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "101001010" =>
            inv <= conv_std_logic_vector(2491,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16597810,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(165413733,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "101001011" =>
            inv <= conv_std_logic_vector(2488,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16678680,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(246431038,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "101001100" =>
            inv <= conv_std_logic_vector(2485,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16759648,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(212362162,28);
            logexp <= conv_std_logic_vector(1021,11);
      WHEN "101001101" =>
            inv <= conv_std_logic_vector(2482,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(31749,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(63242286,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101001110" =>
            inv <= conv_std_logic_vector(2479,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(72331,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(26152662,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101001111" =>
            inv <= conv_std_logic_vector(2476,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(112962,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(26781090,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101010000" =>
            inv <= conv_std_logic_vector(2474,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(140076,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(213075491,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101010001" =>
            inv <= conv_std_logic_vector(2471,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(180789,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(258223654,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101010010" =>
            inv <= conv_std_logic_vector(2468,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(221552,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(158206290,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101010011" =>
            inv <= conv_std_logic_vector(2465,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(262364,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(213755501,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101010100" =>
            inv <= conv_std_logic_vector(2462,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(303226,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(188850466,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101010101" =>
            inv <= conv_std_logic_vector(2459,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(344138,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(116024386,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101010110" =>
            inv <= conv_std_logic_vector(2456,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(385100,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(27929606,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101010111" =>
            inv <= conv_std_logic_vector(2453,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(426111,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(225773656,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101011000" =>
            inv <= conv_std_logic_vector(2450,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(467173,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(205578013,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101011001" =>
            inv <= conv_std_logic_vector(2448,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(494576,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(87278952,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101011010" =>
            inv <= conv_std_logic_vector(2445,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(535722,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(45542114,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101011011" =>
            inv <= conv_std_logic_vector(2442,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(576918,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(142506767,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101011100" =>
            inv <= conv_std_logic_vector(2439,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(618165,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(143076061,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101011101" =>
            inv <= conv_std_logic_vector(2436,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(659463,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(80711705,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101011110" =>
            inv <= conv_std_logic_vector(2433,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(700811,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(257434563,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101011111" =>
            inv <= conv_std_logic_vector(2431,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(728406,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(17672925,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101100000" =>
            inv <= conv_std_logic_vector(2428,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(769839,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(220454209,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101100001" =>
            inv <= conv_std_logic_vector(2425,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(811324,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(215622313,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101100010" =>
            inv <= conv_std_logic_vector(2422,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(852861,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(37221475,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101100011" =>
            inv <= conv_std_logic_vector(2419,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(894448,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(256293434,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101100100" =>
            inv <= conv_std_logic_vector(2417,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(922202,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(222525409,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101100101" =>
            inv <= conv_std_logic_vector(2414,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(963876,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(196069656,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101100110" =>
            inv <= conv_std_logic_vector(2411,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1005602,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(121961634,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101100111" =>
            inv <= conv_std_logic_vector(2408,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1047380,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(34841718,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101101000" =>
            inv <= conv_std_logic_vector(2405,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1089209,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(237915287,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101101001" =>
            inv <= conv_std_logic_vector(2403,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1117125,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(104353094,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101101010" =>
            inv <= conv_std_logic_vector(2400,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1159042,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(63396520,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101101011" =>
            inv <= conv_std_logic_vector(2397,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1201011,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(137556064,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101101100" =>
            inv <= conv_std_logic_vector(2395,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1229020,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(59568237,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101101101" =>
            inv <= conv_std_logic_vector(2392,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1271077,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(46073956,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101101110" =>
            inv <= conv_std_logic_vector(2389,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1313186,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(241992154,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101101111" =>
            inv <= conv_std_logic_vector(2386,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1355349,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(146057517,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101110000" =>
            inv <= conv_std_logic_vector(2384,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1383487,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(116561426,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101110001" =>
            inv <= conv_std_logic_vector(2381,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1425738,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(150565181,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101110010" =>
            inv <= conv_std_logic_vector(2378,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1468042,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(256758677,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101110011" =>
            inv <= conv_std_logic_vector(2376,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1496275,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(146872826,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101110100" =>
            inv <= conv_std_logic_vector(2373,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1538669,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(6283669,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101110101" =>
            inv <= conv_std_logic_vector(2370,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1581116,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(34459956,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101110110" =>
            inv <= conv_std_logic_vector(2367,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1623616,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(267869958,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101110111" =>
            inv <= conv_std_logic_vector(2365,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1651980,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(227479388,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101111000" =>
            inv <= conv_std_logic_vector(2362,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1694571,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(168535478,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101111001" =>
            inv <= conv_std_logic_vector(2360,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1722995,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(146252604,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101111010" =>
            inv <= conv_std_logic_vector(2357,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1765676,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(165723426,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101111011" =>
            inv <= conv_std_logic_vector(2354,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1808412,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(13198653,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101111100" =>
            inv <= conv_std_logic_vector(2352,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1836932,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(162422791,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101111101" =>
            inv <= conv_std_logic_vector(2349,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1879758,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(253404775,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101111110" =>
            inv <= conv_std_logic_vector(2346,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1922640,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(3516811,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "101111111" =>
            inv <= conv_std_logic_vector(2344,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1951257,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(232810820,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110000000" =>
            inv <= conv_std_logic_vector(2341,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1994230,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(124778707,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110000001" =>
            inv <= conv_std_logic_vector(2338,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2037258,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(44895651,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110000010" =>
            inv <= conv_std_logic_vector(2336,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2065973,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(264640088,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110000011" =>
            inv <= conv_std_logic_vector(2333,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2109093,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(226677719,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110000100" =>
            inv <= conv_std_logic_vector(2331,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2137871,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(62314345,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110000101" =>
            inv <= conv_std_logic_vector(2328,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2181083,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(172467092,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110000110" =>
            inv <= conv_std_logic_vector(2326,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2209922,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(231891008,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110000111" =>
            inv <= conv_std_logic_vector(2323,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2253228,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(60167664,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110001000" =>
            inv <= conv_std_logic_vector(2320,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2296589,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(146717848,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110001001" =>
            inv <= conv_std_logic_vector(2318,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2325528,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(68833327,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110001010" =>
            inv <= conv_std_logic_vector(2315,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2368983,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(45955088,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110001011" =>
            inv <= conv_std_logic_vector(2313,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2397984,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(110242438,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110001100" =>
            inv <= conv_std_logic_vector(2310,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2441533,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(86625006,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110001101" =>
            inv <= conv_std_logic_vector(2308,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2470597,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(97343330,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110001110" =>
            inv <= conv_std_logic_vector(2305,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2514240,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(182382776,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110001111" =>
            inv <= conv_std_logic_vector(2303,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2543367,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(212699904,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110010000" =>
            inv <= conv_std_logic_vector(2300,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2587105,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(248069835,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110010001" =>
            inv <= conv_std_logic_vector(2297,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2630901,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(38353874,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110010010" =>
            inv <= conv_std_logic_vector(2295,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2660129,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(199724201,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110010011" =>
            inv <= conv_std_logic_vector(2292,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2704020,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(118011763,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110010100" =>
            inv <= conv_std_logic_vector(2290,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2733312,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(223026379,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110010101" =>
            inv <= conv_std_logic_vector(2287,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2777299,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(112874067,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110010110" =>
            inv <= conv_std_logic_vector(2285,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2806655,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(236438996,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110010111" =>
            inv <= conv_std_logic_vector(2282,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2850738,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(210574529,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110011000" =>
            inv <= conv_std_logic_vector(2280,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2880159,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(159652923,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110011001" =>
            inv <= conv_std_logic_vector(2278,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2909606,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(60159477,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110011010" =>
            inv <= conv_std_logic_vector(2275,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2953824,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(182033526,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110011011" =>
            inv <= conv_std_logic_vector(2273,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2983336,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(14447396,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110011100" =>
            inv <= conv_std_logic_vector(2270,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3027651,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(225760651,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110011101" =>
            inv <= conv_std_logic_vector(2268,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3057228,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(66680404,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110011110" =>
            inv <= conv_std_logic_vector(2265,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3101641,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(214275106,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110011111" =>
            inv <= conv_std_logic_vector(2263,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3131283,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(140806814,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110100000" =>
            inv <= conv_std_logic_vector(2260,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3175795,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(72289811,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110100001" =>
            inv <= conv_std_logic_vector(2258,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3205502,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(162051533,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110100010" =>
            inv <= conv_std_logic_vector(2256,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3235236,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(70518411,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110100011" =>
            inv <= conv_std_logic_vector(2253,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3279886,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(56927398,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110100100" =>
            inv <= conv_std_logic_vector(2251,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3309685,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(238158383,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110100101" =>
            inv <= conv_std_logic_vector(2248,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3354435,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(21682069,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110100110" =>
            inv <= conv_std_logic_vector(2246,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3384301,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(17671725,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110100111" =>
            inv <= conv_std_logic_vector(2243,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3429149,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(253874147,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110101000" =>
            inv <= conv_std_logic_vector(2241,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3459082,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(144015594,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110101001" =>
            inv <= conv_std_logic_vector(2239,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3489041,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(228915285,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110101010" =>
            inv <= conv_std_logic_vector(2236,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3534031,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(11297232,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110101011" =>
            inv <= conv_std_logic_vector(2234,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3564057,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(102394521,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110101100" =>
            inv <= conv_std_logic_vector(2232,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3594110,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(164843479,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110101101" =>
            inv <= conv_std_logic_vector(2229,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3639240,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(266678657,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110101110" =>
            inv <= conv_std_logic_vector(2227,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3669361,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(179992124,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110101111" =>
            inv <= conv_std_logic_vector(2224,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3714593,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(119109352,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110110000" =>
            inv <= conv_std_logic_vector(2222,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3744781,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(233164434,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110110001" =>
            inv <= conv_std_logic_vector(2220,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3774997,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(128320487,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110110010" =>
            inv <= conv_std_logic_vector(2217,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3820371,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(260492078,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110110011" =>
            inv <= conv_std_logic_vector(2215,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3850655,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(202899023,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110110100" =>
            inv <= conv_std_logic_vector(2213,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3880966,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(241038144,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110110101" =>
            inv <= conv_std_logic_vector(2210,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3926485,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(3486646,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110110110" =>
            inv <= conv_std_logic_vector(2208,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3956864,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(204914613,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110110111" =>
            inv <= conv_std_logic_vector(2206,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3987272,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(11839650,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110111000" =>
            inv <= conv_std_logic_vector(2203,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4032934,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(186275213,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110111001" =>
            inv <= conv_std_logic_vector(2201,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4063411,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(5198727,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110111010" =>
            inv <= conv_std_logic_vector(2199,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4093915,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(13571695,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110111011" =>
            inv <= conv_std_logic_vector(2196,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4139723,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(41866951,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110111100" =>
            inv <= conv_std_logic_vector(2194,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4170296,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(180504741,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110111101" =>
            inv <= conv_std_logic_vector(2192,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4200898,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(19253907,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110111110" =>
            inv <= conv_std_logic_vector(2190,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4231527,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(108649881,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "110111111" =>
            inv <= conv_std_logic_vector(2187,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4277523,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(239373474,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111000000" =>
            inv <= conv_std_logic_vector(2185,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4308223,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(75890782,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111000001" =>
            inv <= conv_std_logic_vector(2183,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4338950,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(211176572,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111000010" =>
            inv <= conv_std_logic_vector(2180,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4385094,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(232816832,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111000011" =>
            inv <= conv_std_logic_vector(2178,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4415892,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(236107455,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111000100" =>
            inv <= conv_std_logic_vector(2176,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4446719,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(49882053,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111000101" =>
            inv <= conv_std_logic_vector(2174,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4477573,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(224979561,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111000110" =>
            inv <= conv_std_logic_vector(2171,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4523909,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(21351166,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111000111" =>
            inv <= conv_std_logic_vector(2169,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4554834,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(221595418,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111001000" =>
            inv <= conv_std_logic_vector(2167,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4585789,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(27048959,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111001001" =>
            inv <= conv_std_logic_vector(2165,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4616771,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(257160862,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111001010" =>
            inv <= conv_std_logic_vector(2163,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4647783,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(120806675,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111001011" =>
            inv <= conv_std_logic_vector(2160,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4694354,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(132686548,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111001100" =>
            inv <= conv_std_logic_vector(2158,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4725437,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(216213494,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111001101" =>
            inv <= conv_std_logic_vector(2156,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4756549,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(251657420,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111001110" =>
            inv <= conv_std_logic_vector(2154,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4787690,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(253378504,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111001111" =>
            inv <= conv_std_logic_vector(2151,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4834456,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(190686783,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111010000" =>
            inv <= conv_std_logic_vector(2149,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4865670,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(36971813,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111010001" =>
            inv <= conv_std_logic_vector(2147,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4896912,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(168546215,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111010010" =>
            inv <= conv_std_logic_vector(2145,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4928184,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(63080520,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111010011" =>
            inv <= conv_std_logic_vector(2143,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4959485,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(3592320,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111010100" =>
            inv <= conv_std_logic_vector(2140,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5006490,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(267447830,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111010101" =>
            inv <= conv_std_logic_vector(2138,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5037864,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(252750919,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111010110" =>
            inv <= conv_std_logic_vector(2136,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5069268,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(66956194,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111010111" =>
            inv <= conv_std_logic_vector(2134,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5100700,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(261701721,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111011000" =>
            inv <= conv_std_logic_vector(2132,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5132163,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(46489821,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111011001" =>
            inv <= conv_std_logic_vector(2130,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5163654,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(241477251,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111011010" =>
            inv <= conv_std_logic_vector(2127,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5210947,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(261928568,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111011011" =>
            inv <= conv_std_logic_vector(2125,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5242513,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(205482523,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111011100" =>
            inv <= conv_std_logic_vector(2123,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5274109,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(74671864,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111011101" =>
            inv <= conv_std_logic_vector(2121,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5305734,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(152972013,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111011110" =>
            inv <= conv_std_logic_vector(2119,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5337389,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(187030043,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111011111" =>
            inv <= conv_std_logic_vector(2117,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5369074,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(191971210,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111100000" =>
            inv <= conv_std_logic_vector(2115,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5400789,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(182963660,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111100001" =>
            inv <= conv_std_logic_vector(2112,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5448418,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(109475927,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111100010" =>
            inv <= conv_std_logic_vector(2110,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5480208,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(132240138,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111100011" =>
            inv <= conv_std_logic_vector(2108,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5512028,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(194484233,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111100100" =>
            inv <= conv_std_logic_vector(2106,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5543879,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(43135919,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111100101" =>
            inv <= conv_std_logic_vector(2104,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5575759,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(230473058,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111100110" =>
            inv <= conv_std_logic_vector(2102,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5607670,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(235075650,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111100111" =>
            inv <= conv_std_logic_vector(2100,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5639612,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(72438727,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111101000" =>
            inv <= conv_std_logic_vector(2098,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5671584,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(26537070,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111101001" =>
            inv <= conv_std_logic_vector(2096,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5703586,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(112954470,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111101010" =>
            inv <= conv_std_logic_vector(2093,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5751647,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(55116163,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111101011" =>
            inv <= conv_std_logic_vector(2091,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5783726,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(3932676,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111101100" =>
            inv <= conv_std_logic_vector(2089,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5815835,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(139964094,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111101101" =>
            inv <= conv_std_logic_vector(2087,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5847975,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(210560941,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111101110" =>
            inv <= conv_std_logic_vector(2085,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5880146,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(231554600,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111101111" =>
            inv <= conv_std_logic_vector(2083,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5912348,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(218822034,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111110000" =>
            inv <= conv_std_logic_vector(2081,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5944581,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(188285963,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111110001" =>
            inv <= conv_std_logic_vector(2079,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5976845,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(155915034,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111110010" =>
            inv <= conv_std_logic_vector(2077,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6009140,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(137724004,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111110011" =>
            inv <= conv_std_logic_vector(2075,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6041466,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(149773915,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111110100" =>
            inv <= conv_std_logic_vector(2073,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6073823,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(208172277,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111110101" =>
            inv <= conv_std_logic_vector(2071,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6106212,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(60637778,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111110110" =>
            inv <= conv_std_logic_vector(2069,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6138631,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(260242308,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111110111" =>
            inv <= conv_std_logic_vector(2067,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6171083,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(17927474,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111111000" =>
            inv <= conv_std_logic_vector(2065,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6203565,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(155294811,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111111001" =>
            inv <= conv_std_logic_vector(2063,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6236079,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(151815941,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111111010" =>
            inv <= conv_std_logic_vector(2061,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6268625,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(23880951,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111111011" =>
            inv <= conv_std_logic_vector(2059,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6301202,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(56363124,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111111100" =>
            inv <= conv_std_logic_vector(2057,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6333810,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(265748209,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111111101" =>
            inv <= conv_std_logic_vector(2055,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6366451,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(131699156,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111111110" =>
            inv <= conv_std_logic_vector(2053,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6399123,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(207669033,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "111111111" =>
            inv <= conv_std_logic_vector(2051,12);
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6431827,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(241853027,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN others =>
           inv <= conv_std_logic_vector(0,12);
           logman(52 DOWNTO 29) <= conv_std_logic_vector(0,24);
           logman(28 DOWNTO 1) <= conv_std_logic_vector(0,28);
           logexp <= conv_std_logic_vector(0,11);
    END CASE;
  END PROCESS;

END rtl;
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   DP_LNLUTPOW.VHD                           ***
--***                                             ***
--***   Function: Look Up Table - LN()            ***
--***                                             ***
--***   Generated by MATLAB Utility               ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_lnlutpow IS
PORT (
      add : IN STD_LOGIC_VECTOR (10 DOWNTO 1);
      logman : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
      logexp : OUT STD_LOGIC_VECTOR (11 DOWNTO 1)
     );
END dp_lnlutpow;

ARCHITECTURE rtl OF dp_lnlutpow IS

BEGIN

  pca: PROCESS (add)
  BEGIN
    CASE add IS
      WHEN "0000000000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(0,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(0,28);
            logexp <= conv_std_logic_vector(0,11);
      WHEN "0000000001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6480943,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(251279855,28);
            logexp <= conv_std_logic_vector(1022,11);
      WHEN "0000000010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6480943,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(251279855,28);
            logexp <= conv_std_logic_vector(1023,11);
      WHEN "0000000011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(666403,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(255568755,28);
            logexp <= conv_std_logic_vector(1024,11);
      WHEN "0000000100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6480943,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(251279855,28);
            logexp <= conv_std_logic_vector(1024,11);
      WHEN "0000000101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12295483,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(246990955,28);
            logexp <= conv_std_logic_vector(1024,11);
      WHEN "0000000110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(666403,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(255568755,28);
            logexp <= conv_std_logic_vector(1025,11);
      WHEN "0000000111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3573673,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(253424305,28);
            logexp <= conv_std_logic_vector(1025,11);
      WHEN "0000001000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6480943,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(251279855,28);
            logexp <= conv_std_logic_vector(1025,11);
      WHEN "0000001001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9388213,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(249135405,28);
            logexp <= conv_std_logic_vector(1025,11);
      WHEN "0000001010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12295483,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(246990955,28);
            logexp <= conv_std_logic_vector(1025,11);
      WHEN "0000001011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15202753,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(244846505,28);
            logexp <= conv_std_logic_vector(1025,11);
      WHEN "0000001100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(666403,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(255568755,28);
            logexp <= conv_std_logic_vector(1026,11);
      WHEN "0000001101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2120038,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(254496530,28);
            logexp <= conv_std_logic_vector(1026,11);
      WHEN "0000001110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3573673,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(253424305,28);
            logexp <= conv_std_logic_vector(1026,11);
      WHEN "0000001111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5027308,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(252352080,28);
            logexp <= conv_std_logic_vector(1026,11);
      WHEN "0000010000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6480943,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(251279855,28);
            logexp <= conv_std_logic_vector(1026,11);
      WHEN "0000010001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7934578,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(250207630,28);
            logexp <= conv_std_logic_vector(1026,11);
      WHEN "0000010010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9388213,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(249135405,28);
            logexp <= conv_std_logic_vector(1026,11);
      WHEN "0000010011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10841848,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(248063180,28);
            logexp <= conv_std_logic_vector(1026,11);
      WHEN "0000010100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12295483,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(246990955,28);
            logexp <= conv_std_logic_vector(1026,11);
      WHEN "0000010101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13749118,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(245918730,28);
            logexp <= conv_std_logic_vector(1026,11);
      WHEN "0000010110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15202753,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(244846505,28);
            logexp <= conv_std_logic_vector(1026,11);
      WHEN "0000010111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16656388,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(243774280,28);
            logexp <= conv_std_logic_vector(1026,11);
      WHEN "0000011000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(666403,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(255568755,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000011001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1393221,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(120814915,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000011010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2120038,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(254496530,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000011011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2846856,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(119742690,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000011100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3573673,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(253424305,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000011101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4300491,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(118670465,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000011110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5027308,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(252352080,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000011111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5754126,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(117598240,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000100000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6480943,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(251279855,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000100001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7207761,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(116526015,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000100010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7934578,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(250207630,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000100011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8661396,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(115453790,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000100100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9388213,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(249135405,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000100101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10115031,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(114381565,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000100110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10841848,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(248063180,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000100111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11568666,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(113309340,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000101000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12295483,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(246990955,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000101001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13022301,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(112237114,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000101010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13749118,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(245918730,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000101011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14475936,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(111164889,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000101100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15202753,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(244846505,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000101101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15929571,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(110092664,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000101110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16656388,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(243774280,28);
            logexp <= conv_std_logic_vector(1027,11);
      WHEN "0000101111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(302995,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(54510220,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0000110000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(666403,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(255568755,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0000110001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1029812,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(188191835,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0000110010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1393221,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(120814915,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0000110011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1756630,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(53437995,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0000110100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2120038,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(254496530,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0000110101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2483447,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(187119610,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0000110110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2846856,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(119742690,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0000110111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3210265,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(52365770,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0000111000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3573673,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(253424305,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0000111001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3937082,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(186047385,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0000111010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4300491,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(118670465,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0000111011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4663900,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(51293545,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0000111100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5027308,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(252352080,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0000111101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5390717,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(184975160,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0000111110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5754126,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(117598240,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0000111111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6117535,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(50221319,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001000000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6480943,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(251279855,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001000001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6844352,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(183902935,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001000010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7207761,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(116526015,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001000011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7571170,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(49149094,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001000100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7934578,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(250207630,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001000101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8297987,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(182830710,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001000110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8661396,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(115453790,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001000111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9024805,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(48076869,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001001000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9388213,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(249135405,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001001001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9751622,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(181758485,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001001010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10115031,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(114381565,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001001011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10478440,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(47004644,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001001100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10841848,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(248063180,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001001101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11205257,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(180686260,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001001110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11568666,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(113309340,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001001111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11932075,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(45932419,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001010000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12295483,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(246990955,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001010001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12658892,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(179614035,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001010010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13022301,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(112237114,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001010011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13385710,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(44860194,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001010100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13749118,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(245918730,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001010101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14112527,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(178541810,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001010110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14475936,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(111164889,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001010111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14839345,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(43787969,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001011000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15202753,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(244846505,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001011001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15566162,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(177469585,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001011010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15929571,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(110092664,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001011011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16292980,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(42715744,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001011100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16656388,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(243774280,28);
            logexp <= conv_std_logic_vector(1028,11);
      WHEN "0001011101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(121290,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(222416408,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001011110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(302995,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(54510220,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001011111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(484699,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(155039488,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001100000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(666403,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(255568755,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001100001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(848108,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(87662567,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001100010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1029812,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(188191835,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001100011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1211517,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(20285647,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001100100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1393221,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(120814915,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001100101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1574925,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(221344183,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001100110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1756630,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(53437995,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001100111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1938334,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(153967262,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001101000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2120038,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(254496530,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001101001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2301743,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(86590342,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001101010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2483447,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(187119610,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001101011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2665152,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(19213422,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001101100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2846856,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(119742690,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001101101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3028560,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(220271958,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001101110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3210265,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(52365770,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001101111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3391969,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(152895037,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001110000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3573673,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(253424305,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001110001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3755378,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(85518117,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001110010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3937082,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(186047385,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001110011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4118787,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(18141197,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001110100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4300491,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(118670465,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001110101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4482195,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(219199733,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001110110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4663900,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(51293545,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001110111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4845604,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(151822812,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001111000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5027308,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(252352080,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001111001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5209013,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(84445892,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001111010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5390717,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(184975160,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001111011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5572422,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(17068972,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001111100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5754126,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(117598240,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001111101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5935830,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(218127508,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001111110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6117535,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(50221319,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0001111111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6299239,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(150750587,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010000000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6480943,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(251279855,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010000001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6662648,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(83373667,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010000010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6844352,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(183902935,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010000011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7026057,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(15996747,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010000100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7207761,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(116526015,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010000101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7389465,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(217055283,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010000110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7571170,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(49149094,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010000111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7752874,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(149678362,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010001000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7934578,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(250207630,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010001001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8116283,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(82301442,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010001010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8297987,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(182830710,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010001011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8479692,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(14924522,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010001100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8661396,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(115453790,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010001101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8843100,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(215983058,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010001110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9024805,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(48076869,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010001111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9206509,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(148606137,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010010000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9388213,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(249135405,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010010001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9569918,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(81229217,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010010010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9751622,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(181758485,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010010011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9933327,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(13852297,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010010100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10115031,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(114381565,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010010101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10296735,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(214910832,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010010110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10478440,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(47004644,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010010111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10660144,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(147533912,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010011000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10841848,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(248063180,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010011001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11023553,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(80156992,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010011010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11205257,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(180686260,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010011011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11386962,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(12780072,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010011100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11568666,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(113309340,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010011101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11750370,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(213838607,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010011110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11932075,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(45932419,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010011111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12113779,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(146461687,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010100000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12295483,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(246990955,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010100001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12477188,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(79084767,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010100010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12658892,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(179614035,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010100011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12840597,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(11707847,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010100100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13022301,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(112237114,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010100101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13204005,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(212766382,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010100110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13385710,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(44860194,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010100111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13567414,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(145389462,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010101000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13749118,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(245918730,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010101001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13930823,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(78012542,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010101010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14112527,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(178541810,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010101011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14294232,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(10635622,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010101100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14475936,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(111164889,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010101101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14657640,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(211694157,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010101110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14839345,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(43787969,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010101111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15021049,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(144317237,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010110000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15202753,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(244846505,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010110001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15384458,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(76940317,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010110010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15566162,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(177469585,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010110011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15747867,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(9563397,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010110100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15929571,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(110092664,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010110101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16111275,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(210621932,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010110110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16292980,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(42715744,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010110111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16474684,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(143245012,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010111000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16656388,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(243774280,28);
            logexp <= conv_std_logic_vector(1029,11);
      WHEN "0010111001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(30438,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(172151774,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0010111010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(121290,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(222416408,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0010111011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(212143,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(4245586,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0010111100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(302995,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(54510220,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0010111101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(393847,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(104774854,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0010111110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(484699,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(155039488,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0010111111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(575551,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(205304121,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011000000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(666403,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(255568755,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011000001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(757256,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(37397933,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011000010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(848108,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(87662567,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011000011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(938960,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(137927201,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011000100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1029812,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(188191835,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011000101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1120664,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(238456469,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011000110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1211517,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(20285647,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011000111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1302369,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(70550281,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011001000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1393221,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(120814915,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011001001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1484073,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(171079549,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011001010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1574925,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(221344183,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011001011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1665778,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(3173361,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011001100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1756630,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(53437995,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011001101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1847482,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(103702629,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011001110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1938334,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(153967262,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011001111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2029186,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(204231896,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011010000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2120038,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(254496530,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011010001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2210891,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(36325708,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011010010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2301743,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(86590342,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011010011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2392595,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(136854976,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011010100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2483447,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(187119610,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011010101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2574299,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(237384244,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011010110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2665152,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(19213422,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011010111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2756004,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(69478056,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011011000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2846856,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(119742690,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011011001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2937708,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(170007324,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011011010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3028560,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(220271958,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011011011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3119413,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(2101136,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011011100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3210265,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(52365770,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011011101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3301117,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(102630404,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011011110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3391969,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(152895037,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011011111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3482821,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(203159671,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011100000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3573673,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(253424305,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011100001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3664526,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(35253483,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011100010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3755378,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(85518117,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011100011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3846230,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(135782751,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011100100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3937082,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(186047385,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011100101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4027934,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(236312019,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011100110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4118787,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(18141197,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011100111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4209639,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(68405831,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011101000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4300491,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(118670465,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011101001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4391343,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(168935099,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011101010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4482195,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(219199733,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011101011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4573048,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(1028911,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011101100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4663900,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(51293545,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011101101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4754752,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(101558178,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011101110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4845604,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(151822812,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011101111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4936456,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(202087446,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011110000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5027308,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(252352080,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011110001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5118161,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(34181258,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011110010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5209013,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(84445892,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011110011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5299865,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(134710526,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011110100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5390717,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(184975160,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011110101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5481569,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(235239794,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011110110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5572422,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(17068972,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011110111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5663274,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(67333606,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011111000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5754126,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(117598240,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011111001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5844978,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(167862874,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011111010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5935830,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(218127508,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011111011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6026682,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(268392142,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011111100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6117535,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(50221319,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011111101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6208387,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(100485953,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011111110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6299239,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(150750587,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0011111111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6390091,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(201015221,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100000000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6480943,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(251279855,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100000001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6571796,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(33109033,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100000010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6662648,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(83373667,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100000011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6753500,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(133638301,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100000100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6844352,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(183902935,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100000101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6935204,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(234167569,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100000110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7026057,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(15996747,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100000111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7116909,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(66261381,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100001000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7207761,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(116526015,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100001001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7298613,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(166790649,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100001010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7389465,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(217055283,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100001011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7480317,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(267319916,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100001100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7571170,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(49149094,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100001101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7662022,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(99413728,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100001110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7752874,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(149678362,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100001111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7843726,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(199942996,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100010000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7934578,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(250207630,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100010001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8025431,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(32036808,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100010010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8116283,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(82301442,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100010011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8207135,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(132566076,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100010100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8297987,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(182830710,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100010101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8388839,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(233095344,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100010110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8479692,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(14924522,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100010111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8570544,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(65189156,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100011000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8661396,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(115453790,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100011001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8752248,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(165718424,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100011010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8843100,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(215983058,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100011011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8933952,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(266247691,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100011100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9024805,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(48076869,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100011101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9115657,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(98341503,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100011110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9206509,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(148606137,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100011111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9297361,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(198870771,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100100000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9388213,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(249135405,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100100001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9479066,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(30964583,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100100010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9569918,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(81229217,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100100011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9660770,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(131493851,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100100100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9751622,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(181758485,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100100101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9842474,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(232023119,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100100110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9933327,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(13852297,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100100111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10024179,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(64116931,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100101000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10115031,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(114381565,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100101001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10205883,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(164646199,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100101010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10296735,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(214910832,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100101011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10387587,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(265175466,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100101100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10478440,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(47004644,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100101101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10569292,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(97269278,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100101110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10660144,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(147533912,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100101111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10750996,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(197798546,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100110000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10841848,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(248063180,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100110001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10932701,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(29892358,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100110010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11023553,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(80156992,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100110011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11114405,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(130421626,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100110100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11205257,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(180686260,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100110101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11296109,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(230950894,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100110110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11386962,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(12780072,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100110111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11477814,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(63044706,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100111000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11568666,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(113309340,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100111001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11659518,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(163573973,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100111010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11750370,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(213838607,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100111011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11841222,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(264103241,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100111100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11932075,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(45932419,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100111101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12022927,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(96197053,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100111110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12113779,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(146461687,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0100111111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12204631,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(196726321,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101000000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12295483,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(246990955,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101000001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12386336,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(28820133,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101000010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12477188,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(79084767,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101000011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12568040,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(129349401,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101000100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12658892,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(179614035,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101000101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12749744,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(229878669,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101000110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12840597,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(11707847,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101000111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12931449,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(61972481,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101001000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13022301,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(112237114,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101001001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13113153,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(162501748,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101001010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13204005,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(212766382,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101001011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13294857,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(263031016,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101001100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13385710,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(44860194,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101001101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13476562,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(95124828,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101001110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13567414,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(145389462,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101001111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13658266,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(195654096,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101010000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13749118,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(245918730,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101010001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13839971,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(27747908,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101010010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13930823,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(78012542,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101010011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14021675,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(128277176,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101010100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14112527,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(178541810,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101010101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14203379,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(228806444,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101010110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14294232,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(10635622,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101010111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14385084,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(60900256,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101011000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14475936,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(111164889,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101011001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14566788,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(161429523,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101011010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14657640,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(211694157,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101011011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14748492,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(261958791,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101011100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14839345,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(43787969,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101011101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14930197,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(94052603,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101011110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15021049,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(144317237,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101011111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15111901,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(194581871,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101100000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15202753,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(244846505,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101100001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15293606,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(26675683,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101100010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15384458,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(76940317,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101100011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15475310,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(127204951,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101100100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15566162,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(177469585,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101100101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15657014,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(227734219,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101100110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15747867,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(9563397,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101100111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15838719,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(59828030,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101101000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15929571,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(110092664,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101101001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16020423,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(160357298,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101101010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16111275,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(210621932,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101101011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16202127,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(260886566,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101101100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16292980,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(42715744,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101101101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16383832,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(92980378,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101101110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16474684,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(143245012,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101101111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16565536,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(193509646,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101110000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16656388,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(243774280,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101110001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16747241,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(25603458,28);
            logexp <= conv_std_logic_vector(1030,11);
      WHEN "0101110010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(30438,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(172151774,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0101110011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(75864,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(197284091,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0101110100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(121290,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(222416408,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0101110101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(166716,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(247548725,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0101110110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(212143,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(4245586,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0101110111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(257569,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(29377903,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0101111000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(302995,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(54510220,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0101111001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(348421,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(79642537,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0101111010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(393847,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(104774854,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0101111011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(439273,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(129907171,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0101111100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(484699,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(155039488,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0101111101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(530125,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(180171805,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0101111110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(575551,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(205304121,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0101111111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(620977,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(230436438,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110000000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(666403,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(255568755,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110000001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(711830,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(12265616,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110000010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(757256,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(37397933,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110000011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(802682,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(62530250,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110000100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(848108,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(87662567,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110000101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(893534,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(112794884,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110000110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(938960,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(137927201,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110000111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(984386,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(163059518,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110001000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1029812,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(188191835,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110001001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1075238,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(213324152,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110001010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1120664,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(238456469,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110001011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1166090,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(263588786,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110001100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1211517,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(20285647,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110001101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1256943,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(45417964,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110001110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1302369,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(70550281,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110001111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1347795,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(95682598,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110010000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1393221,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(120814915,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110010001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1438647,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(145947232,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110010010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1484073,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(171079549,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110010011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1529499,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(196211866,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110010100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1574925,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(221344183,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110010101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1620351,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(246476500,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110010110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1665778,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(3173361,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110010111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1711204,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(28305678,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110011000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1756630,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(53437995,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110011001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1802056,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(78570312,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110011010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1847482,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(103702629,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110011011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1892908,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(128834946,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110011100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1938334,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(153967262,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110011101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1983760,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(179099579,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110011110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2029186,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(204231896,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110011111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2074612,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(229364213,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110100000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2120038,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(254496530,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110100001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2165465,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(11193391,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110100010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2210891,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(36325708,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110100011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2256317,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(61458025,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110100100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2301743,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(86590342,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110100101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2347169,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(111722659,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110100110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2392595,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(136854976,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110100111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2438021,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(161987293,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110101000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2483447,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(187119610,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110101001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2528873,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(212251927,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110101010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2574299,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(237384244,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110101011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2619725,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(262516561,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110101100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2665152,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(19213422,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110101101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2710578,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(44345739,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110101110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2756004,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(69478056,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110101111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2801430,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(94610373,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110110000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2846856,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(119742690,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110110001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2892282,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(144875007,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110110010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2937708,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(170007324,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110110011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2983134,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(195139641,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110110100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3028560,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(220271958,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110110101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3073986,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(245404275,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110110110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3119413,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(2101136,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110110111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3164839,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(27233453,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110111000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3210265,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(52365770,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110111001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3255691,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(77498087,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110111010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3301117,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(102630404,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110111011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3346543,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(127762720,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110111100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3391969,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(152895037,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110111101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3437395,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(178027354,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110111110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3482821,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(203159671,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0110111111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3528247,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(228291988,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111000000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3573673,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(253424305,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111000001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3619100,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(10121166,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111000010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3664526,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(35253483,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111000011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3709952,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(60385800,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111000100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3755378,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(85518117,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111000101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3800804,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(110650434,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111000110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3846230,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(135782751,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111000111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3891656,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(160915068,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111001000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3937082,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(186047385,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111001001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3982508,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(211179702,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111001010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4027934,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(236312019,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111001011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4073360,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(261444336,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111001100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4118787,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(18141197,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111001101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4164213,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(43273514,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111001110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4209639,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(68405831,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111001111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4255065,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(93538148,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111010000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4300491,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(118670465,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111010001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4345917,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(143802782,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111010010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4391343,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(168935099,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111010011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4436769,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(194067416,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111010100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4482195,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(219199733,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111010101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4527621,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(244332050,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111010110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4573048,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(1028911,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111010111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4618474,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(26161228,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111011000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4663900,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(51293545,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111011001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4709326,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(76425861,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111011010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4754752,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(101558178,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111011011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4800178,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(126690495,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111011100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4845604,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(151822812,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111011101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4891030,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(176955129,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111011110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4936456,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(202087446,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111011111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4981882,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(227219763,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111100000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5027308,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(252352080,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111100001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5072735,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(9048941,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111100010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5118161,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(34181258,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111100011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5163587,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(59313575,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111100100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5209013,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(84445892,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111100101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5254439,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(109578209,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111100110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5299865,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(134710526,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111100111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5345291,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(159842843,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111101000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5390717,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(184975160,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111101001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5436143,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(210107477,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111101010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5481569,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(235239794,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111101011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5526995,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(260372111,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111101100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5572422,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(17068972,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111101101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5617848,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(42201289,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111101110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5663274,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(67333606,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111101111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5708700,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(92465923,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111110000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5754126,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(117598240,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111110001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5799552,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(142730557,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111110010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5844978,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(167862874,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111110011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5890404,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(192995191,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111110100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5935830,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(218127508,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111110101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5981256,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(243259825,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111110110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6026682,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(268392142,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111110111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6072109,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(25089003,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111111000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6117535,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(50221319,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111111001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6162961,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(75353636,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111111010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6208387,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(100485953,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111111011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6253813,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(125618270,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111111100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6299239,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(150750587,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111111101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6344665,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(175882904,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111111110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6390091,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(201015221,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "0111111111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6435517,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(226147538,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000000000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6480943,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(251279855,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000000001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6526370,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(7976716,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000000010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6571796,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(33109033,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000000011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6617222,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(58241350,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000000100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6662648,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(83373667,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000000101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6708074,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(108505984,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000000110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6753500,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(133638301,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000000111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6798926,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(158770618,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000001000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6844352,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(183902935,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000001001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6889778,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(209035252,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000001010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6935204,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(234167569,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000001011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6980630,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(259299886,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000001100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7026057,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(15996747,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000001101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7071483,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(41129064,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000001110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7116909,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(66261381,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000001111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7162335,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(91393698,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000010000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7207761,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(116526015,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000010001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7253187,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(141658332,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000010010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7298613,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(166790649,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000010011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7344039,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(191922966,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000010100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7389465,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(217055283,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000010101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7434891,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(242187600,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000010110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7480317,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(267319916,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000010111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7525744,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(24016777,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000011000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7571170,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(49149094,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000011001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7616596,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(74281411,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000011010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7662022,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(99413728,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000011011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7707448,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(124546045,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000011100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7752874,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(149678362,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000011101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7798300,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(174810679,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000011110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7843726,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(199942996,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000011111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7889152,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(225075313,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000100000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7934578,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(250207630,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000100001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7980005,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(6904491,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000100010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8025431,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(32036808,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000100011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8070857,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(57169125,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000100100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8116283,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(82301442,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000100101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8161709,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(107433759,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000100110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8207135,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(132566076,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000100111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8252561,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(157698393,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000101000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8297987,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(182830710,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000101001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8343413,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(207963027,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000101010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8388839,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(233095344,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000101011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8434265,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(258227661,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000101100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8479692,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(14924522,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000101101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8525118,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(40056839,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000101110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8570544,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(65189156,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000101111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8615970,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(90321473,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000110000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8661396,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(115453790,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000110001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8706822,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(140586107,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000110010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8752248,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(165718424,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000110011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8797674,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(190850741,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000110100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8843100,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(215983058,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000110101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8888526,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(241115374,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000110110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8933952,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(266247691,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000110111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(8979379,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(22944552,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000111000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9024805,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(48076869,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000111001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9070231,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(73209186,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000111010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9115657,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(98341503,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000111011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9161083,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(123473820,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000111100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9206509,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(148606137,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000111101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9251935,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(173738454,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000111110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9297361,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(198870771,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1000111111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9342787,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(224003088,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001000000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9388213,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(249135405,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001000001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9433640,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(5832266,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001000010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9479066,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(30964583,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001000011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9524492,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(56096900,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001000100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9569918,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(81229217,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001000101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9615344,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(106361534,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001000110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9660770,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(131493851,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001000111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9706196,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(156626168,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001001000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9751622,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(181758485,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001001001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9797048,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(206890802,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001001010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9842474,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(232023119,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001001011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9887900,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(257155436,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001001100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9933327,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(13852297,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001001101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(9978753,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(38984614,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001001110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10024179,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(64116931,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001001111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10069605,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(89249248,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001010000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10115031,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(114381565,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001010001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10160457,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(139513882,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001010010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10205883,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(164646199,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001010011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10251309,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(189778515,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001010100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10296735,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(214910832,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001010101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10342161,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(240043149,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001010110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10387587,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(265175466,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001010111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10433014,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(21872327,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001011000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10478440,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(47004644,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001011001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10523866,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(72136961,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001011010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10569292,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(97269278,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001011011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10614718,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(122401595,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001011100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10660144,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(147533912,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001011101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10705570,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(172666229,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001011110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10750996,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(197798546,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001011111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10796422,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(222930863,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001100000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10841848,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(248063180,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001100001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10887275,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(4760041,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001100010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10932701,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(29892358,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001100011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(10978127,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(55024675,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001100100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11023553,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(80156992,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001100101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11068979,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(105289309,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001100110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11114405,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(130421626,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001100111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11159831,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(155553943,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001101000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11205257,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(180686260,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001101001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11250683,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(205818577,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001101010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11296109,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(230950894,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001101011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11341535,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(256083211,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001101100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11386962,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(12780072,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001101101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11432388,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(37912389,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001101110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11477814,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(63044706,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001101111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11523240,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(88177023,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001110000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11568666,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(113309340,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001110001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11614092,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(138441657,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001110010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11659518,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(163573973,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001110011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11704944,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(188706290,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001110100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11750370,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(213838607,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001110101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11795796,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(238970924,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001110110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11841222,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(264103241,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001110111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11886649,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(20800102,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001111000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11932075,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(45932419,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001111001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(11977501,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(71064736,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001111010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12022927,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(96197053,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001111011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12068353,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(121329370,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001111100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12113779,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(146461687,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001111101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12159205,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(171594004,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001111110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12204631,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(196726321,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1001111111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12250057,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(221858638,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010000000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12295483,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(246990955,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010000001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12340910,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(3687816,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010000010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12386336,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(28820133,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010000011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12431762,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(53952450,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010000100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12477188,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(79084767,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010000101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12522614,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(104217084,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010000110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12568040,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(129349401,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010000111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12613466,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(154481718,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010001000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12658892,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(179614035,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010001001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12704318,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(204746352,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010001010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12749744,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(229878669,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010001011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12795170,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(255010986,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010001100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12840597,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(11707847,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010001101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12886023,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(36840164,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010001110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12931449,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(61972481,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010001111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(12976875,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(87104798,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010010000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13022301,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(112237114,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010010001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13067727,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(137369431,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010010010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13113153,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(162501748,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010010011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13158579,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(187634065,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010010100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13204005,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(212766382,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010010101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13249431,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(237898699,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010010110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13294857,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(263031016,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010010111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13340284,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(19727877,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010011000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13385710,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(44860194,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010011001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13431136,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(69992511,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010011010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13476562,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(95124828,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010011011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13521988,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(120257145,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010011100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13567414,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(145389462,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010011101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13612840,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(170521779,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010011110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13658266,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(195654096,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010011111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13703692,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(220786413,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010100000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13749118,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(245918730,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010100001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13794545,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(2615591,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010100010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13839971,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(27747908,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010100011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13885397,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(52880225,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010100100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13930823,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(78012542,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010100101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(13976249,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(103144859,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010100110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14021675,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(128277176,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010100111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14067101,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(153409493,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010101000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14112527,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(178541810,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010101001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14157953,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(203674127,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010101010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14203379,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(228806444,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010101011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14248805,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(253938761,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010101100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14294232,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(10635622,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010101101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14339658,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(35767939,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010101110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14385084,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(60900256,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010101111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14430510,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(86032572,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010110000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14475936,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(111164889,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010110001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14521362,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(136297206,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010110010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14566788,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(161429523,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010110011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14612214,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(186561840,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010110100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14657640,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(211694157,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010110101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14703066,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(236826474,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010110110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14748492,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(261958791,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010110111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14793919,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(18655652,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010111000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14839345,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(43787969,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010111001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14884771,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(68920286,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010111010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14930197,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(94052603,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010111011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(14975623,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(119184920,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010111100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15021049,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(144317237,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010111101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15066475,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(169449554,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010111110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15111901,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(194581871,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1010111111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15157327,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(219714188,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011000000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15202753,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(244846505,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011000001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15248180,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(1543366,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011000010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15293606,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(26675683,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011000011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15339032,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(51808000,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011000100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15384458,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(76940317,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011000101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15429884,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(102072634,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011000110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15475310,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(127204951,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011000111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15520736,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(152337268,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011001000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15566162,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(177469585,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011001001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15611588,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(202601902,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011001010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15657014,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(227734219,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011001011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15702440,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(252866536,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011001100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15747867,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(9563397,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011001101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15793293,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(34695713,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011001110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15838719,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(59828030,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011001111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15884145,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(84960347,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011010000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15929571,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(110092664,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011010001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(15974997,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(135224981,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011010010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16020423,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(160357298,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011010011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16065849,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(185489615,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011010100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16111275,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(210621932,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011010101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16156701,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(235754249,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011010110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16202127,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(260886566,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011010111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16247554,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(17583427,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011011000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16292980,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(42715744,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011011001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16338406,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(67848061,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011011010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16383832,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(92980378,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011011011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16429258,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(118112695,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011011100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16474684,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(143245012,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011011101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16520110,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(168377329,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011011110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16565536,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(193509646,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011011111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16610962,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(218641963,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011100000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16656388,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(243774280,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011100001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16701815,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(471141,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011100010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(16747241,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(25603458,28);
            logexp <= conv_std_logic_vector(1031,11);
      WHEN "1011100011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(7725,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(159585615,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011100100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(30438,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(172151774,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011100101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(53151,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(184717932,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011100110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(75864,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(197284091,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011100111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(98577,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(209850249,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011101000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(121290,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(222416408,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011101001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(144003,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(234982566,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011101010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(166716,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(247548725,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011101011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(189429,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(260114883,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011101100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(212143,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(4245586,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011101101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(234856,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(16811744,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011101110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(257569,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(29377903,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011101111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(280282,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(41944061,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011110000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(302995,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(54510220,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011110001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(325708,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(67076378,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011110010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(348421,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(79642537,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011110011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(371134,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(92208695,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011110100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(393847,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(104774854,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011110101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(416560,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(117341012,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011110110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(439273,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(129907171,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011110111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(461986,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(142473329,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011111000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(484699,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(155039488,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011111001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(507412,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(167605646,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011111010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(530125,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(180171805,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011111011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(552838,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(192737963,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011111100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(575551,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(205304121,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011111101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(598264,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(217870280,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011111110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(620977,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(230436438,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1011111111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(643690,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(243002597,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100000000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(666403,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(255568755,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100000001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(689116,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(268134914,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100000010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(711830,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(12265616,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100000011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(734543,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(24831775,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100000100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(757256,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(37397933,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100000101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(779969,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(49964092,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100000110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(802682,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(62530250,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100000111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(825395,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(75096409,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100001000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(848108,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(87662567,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100001001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(870821,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(100228726,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100001010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(893534,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(112794884,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100001011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(916247,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(125361043,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100001100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(938960,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(137927201,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100001101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(961673,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(150493360,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100001110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(984386,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(163059518,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100001111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1007099,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(175625677,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100010000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1029812,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(188191835,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100010001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1052525,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(200757994,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100010010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1075238,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(213324152,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100010011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1097951,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(225890311,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100010100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1120664,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(238456469,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100010101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1143377,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(251022628,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100010110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1166090,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(263588786,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100010111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1188804,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(7719489,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100011000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1211517,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(20285647,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100011001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1234230,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(32851805,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100011010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1256943,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(45417964,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100011011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1279656,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(57984122,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100011100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1302369,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(70550281,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100011101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1325082,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(83116439,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100011110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1347795,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(95682598,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100011111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1370508,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(108248756,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100100000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1393221,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(120814915,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100100001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1415934,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(133381073,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100100010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1438647,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(145947232,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100100011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1461360,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(158513390,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100100100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1484073,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(171079549,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100100101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1506786,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(183645707,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100100110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1529499,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(196211866,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100100111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1552212,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(208778024,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100101000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1574925,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(221344183,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100101001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1597638,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(233910341,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100101010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1620351,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(246476500,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100101011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1643064,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(259042658,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100101100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1665778,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(3173361,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100101101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1688491,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(15739519,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100101110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1711204,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(28305678,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100101111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1733917,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(40871836,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100110000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1756630,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(53437995,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100110001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1779343,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(66004153,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100110010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1802056,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(78570312,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100110011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1824769,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(91136470,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100110100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1847482,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(103702629,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100110101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1870195,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(116268787,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100110110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1892908,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(128834946,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100110111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1915621,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(141401104,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100111000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1938334,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(153967262,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100111001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1961047,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(166533421,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100111010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(1983760,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(179099579,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100111011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2006473,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(191665738,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100111100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2029186,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(204231896,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100111101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2051899,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(216798055,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100111110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2074612,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(229364213,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1100111111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2097325,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(241930372,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101000000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2120038,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(254496530,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101000001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2142751,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(267062689,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101000010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2165465,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(11193391,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101000011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2188178,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(23759550,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101000100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2210891,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(36325708,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101000101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2233604,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(48891867,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101000110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2256317,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(61458025,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101000111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2279030,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(74024184,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101001000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2301743,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(86590342,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101001001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2324456,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(99156501,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101001010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2347169,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(111722659,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101001011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2369882,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(124288818,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101001100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2392595,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(136854976,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101001101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2415308,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(149421135,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101001110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2438021,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(161987293,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101001111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2460734,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(174553452,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101010000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2483447,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(187119610,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101010001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2506160,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(199685769,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101010010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2528873,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(212251927,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101010011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2551586,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(224818086,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101010100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2574299,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(237384244,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101010101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2597012,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(249950403,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101010110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2619725,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(262516561,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101010111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2642439,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(6647263,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101011000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2665152,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(19213422,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101011001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2687865,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(31779580,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101011010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2710578,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(44345739,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101011011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2733291,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(56911897,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101011100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2756004,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(69478056,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101011101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2778717,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(82044214,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101011110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2801430,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(94610373,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101011111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2824143,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(107176531,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101100000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2846856,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(119742690,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101100001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2869569,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(132308848,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101100010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2892282,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(144875007,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101100011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2914995,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(157441165,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101100100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2937708,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(170007324,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101100101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2960421,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(182573482,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101100110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(2983134,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(195139641,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101100111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3005847,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(207705799,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101101000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3028560,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(220271958,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101101001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3051273,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(232838116,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101101010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3073986,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(245404275,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101101011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3096699,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(257970433,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101101100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3119413,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(2101136,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101101101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3142126,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(14667294,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101101110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3164839,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(27233453,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101101111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3187552,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(39799611,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101110000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3210265,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(52365770,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101110001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3232978,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(64931928,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101110010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3255691,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(77498087,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101110011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3278404,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(90064245,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101110100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3301117,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(102630404,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101110101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3323830,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(115196562,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101110110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3346543,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(127762720,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101110111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3369256,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(140328879,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101111000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3391969,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(152895037,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101111001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3414682,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(165461196,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101111010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3437395,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(178027354,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101111011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3460108,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(190593513,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101111100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3482821,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(203159671,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101111101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3505534,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(215725830,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101111110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3528247,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(228291988,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1101111111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3550960,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(240858147,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110000000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3573673,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(253424305,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110000001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3596386,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(265990464,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110000010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3619100,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(10121166,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110000011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3641813,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(22687325,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110000100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3664526,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(35253483,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110000101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3687239,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(47819642,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110000110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3709952,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(60385800,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110000111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3732665,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(72951959,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110001000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3755378,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(85518117,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110001001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3778091,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(98084276,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110001010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3800804,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(110650434,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110001011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3823517,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(123216593,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110001100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3846230,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(135782751,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110001101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3868943,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(148348910,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110001110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3891656,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(160915068,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110001111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3914369,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(173481227,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110010000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3937082,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(186047385,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110010001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3959795,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(198613544,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110010010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(3982508,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(211179702,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110010011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4005221,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(223745860,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110010100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4027934,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(236312019,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110010101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4050647,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(248878177,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110010110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4073360,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(261444336,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110010111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4096074,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(5575038,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110011000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4118787,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(18141197,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110011001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4141500,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(30707355,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110011010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4164213,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(43273514,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110011011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4186926,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(55839672,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110011100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4209639,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(68405831,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110011101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4232352,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(80971989,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110011110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4255065,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(93538148,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110011111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4277778,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(106104306,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110100000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4300491,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(118670465,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110100001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4323204,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(131236623,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110100010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4345917,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(143802782,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110100011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4368630,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(156368940,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110100100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4391343,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(168935099,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110100101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4414056,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(181501257,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110100110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4436769,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(194067416,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110100111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4459482,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(206633574,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110101000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4482195,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(219199733,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110101001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4504908,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(231765891,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110101010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4527621,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(244332050,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110101011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4550334,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(256898208,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110101100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4573048,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(1028911,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110101101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4595761,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(13595069,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110101110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4618474,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(26161228,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110101111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4641187,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(38727386,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110110000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4663900,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(51293545,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110110001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4686613,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(63859703,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110110010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4709326,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(76425861,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110110011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4732039,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(88992020,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110110100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4754752,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(101558178,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110110101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4777465,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(114124337,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110110110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4800178,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(126690495,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110110111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4822891,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(139256654,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110111000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4845604,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(151822812,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110111001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4868317,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(164388971,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110111010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4891030,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(176955129,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110111011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4913743,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(189521288,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110111100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4936456,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(202087446,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110111101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4959169,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(214653605,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110111110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(4981882,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(227219763,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1110111111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5004595,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(239785922,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111000000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5027308,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(252352080,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111000001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5050021,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(264918239,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111000010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5072735,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(9048941,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111000011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5095448,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(21615100,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111000100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5118161,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(34181258,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111000101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5140874,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(46747417,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111000110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5163587,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(59313575,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111000111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5186300,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(71879734,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111001000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5209013,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(84445892,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111001001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5231726,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(97012051,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111001010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5254439,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(109578209,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111001011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5277152,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(122144368,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111001100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5299865,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(134710526,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111001101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5322578,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(147276685,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111001110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5345291,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(159842843,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111001111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5368004,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(172409002,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111010000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5390717,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(184975160,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111010001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5413430,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(197541318,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111010010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5436143,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(210107477,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111010011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5458856,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(222673635,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111010100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5481569,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(235239794,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111010101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5504282,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(247805952,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111010110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5526995,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(260372111,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111010111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5549709,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(4502813,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111011000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5572422,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(17068972,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111011001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5595135,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(29635130,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111011010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5617848,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(42201289,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111011011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5640561,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(54767447,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111011100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5663274,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(67333606,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111011101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5685987,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(79899764,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111011110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5708700,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(92465923,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111011111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5731413,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(105032081,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111100000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5754126,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(117598240,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111100001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5776839,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(130164398,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111100010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5799552,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(142730557,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111100011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5822265,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(155296715,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111100100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5844978,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(167862874,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111100101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5867691,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(180429032,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111100110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5890404,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(192995191,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111100111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5913117,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(205561349,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111101000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5935830,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(218127508,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111101001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5958543,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(230693666,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111101010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(5981256,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(243259825,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111101011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6003969,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(255825983,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111101100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6026682,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(268392142,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111101101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6049396,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(12522844,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111101110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6072109,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(25089003,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111101111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6094822,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(37655161,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111110000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6117535,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(50221319,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111110001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6140248,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(62787478,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111110010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6162961,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(75353636,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111110011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6185674,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(87919795,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111110100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6208387,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(100485953,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111110101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6231100,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(113052112,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111110110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6253813,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(125618270,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111110111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6276526,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(138184429,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111111000" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6299239,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(150750587,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111111001" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6321952,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(163316746,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111111010" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6344665,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(175882904,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111111011" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6367378,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(188449063,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111111100" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6390091,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(201015221,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111111101" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6412804,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(213581380,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111111110" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6435517,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(226147538,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN "1111111111" =>
            logman(52 DOWNTO 29) <= conv_std_logic_vector(6458230,24);
            logman(28 DOWNTO 1) <= conv_std_logic_vector(238713697,28);
            logexp <= conv_std_logic_vector(1032,11);
      WHEN others =>
           logman(52 DOWNTO 29) <= conv_std_logic_vector(0,24);
           logman(28 DOWNTO 1) <= conv_std_logic_vector(0,28);
           logexp <= conv_std_logic_vector(0,11);
    END CASE;
  END PROCESS;

END rtl;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   DP_LNNORM.VHD                             ***
--***                                             ***
--***   Function: Double Precision Normalization  ***
--***   of LN calculation                         ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** Latency = 3 + 2*Speed                       ***
--*************************************************** 

ENTITY dp_lnnorm IS 
GENERIC (
         speed : integer := 1
        ); 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      inman : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
      inexp : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
      
      outman : OUT STD_LOGIC_VECTOR (64 DOWNTO 1);
      outexp : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
      zero : OUT STD_LOGIC
    );
END dp_lnnorm;

ARCHITECTURE rtl OF dp_lnnorm IS

  -- 3+2*speed
  
  signal shift, shiftff : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal zerochk : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal inmanff, outmanff : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal inexpff : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal inmandelbus : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal outmanbus : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal expaddbus, expsubbus : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal expmidbus, expoutbus : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal zeroff : STD_LOGIC_VECTOR (2+2*speed DOWNTO 1);

  component dp_lnclz
  PORT (
        mantissa : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
        leading : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
       );
  end component;
  
  component dp_lnclzpipe
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        mantissa : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
        leading : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
       );
  end component;
     
  component dp_lsft64x6
  PORT (
        inbus : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);
        outbus : OUT STD_LOGIC_VECTOR (64 DOWNTO 1)
      );
  end component;
  
  component dp_lsft64x6pipe
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        inbus : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);
        outbus : OUT STD_LOGIC_VECTOR (64 DOWNTO 1)
      );
  end component;
  
  component fp_del
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
  end component;
             
BEGIN
  
  ppin: PROCESS (sysclk,reset)
  BEGIN
  
    IF (reset = '1') THEN
        
      FOR k IN 1 TO 64 LOOP
        inmanff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 11 LOOP
        inexpff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 2+2*speed LOOP
        zeroff(k) <= '0';
      END LOOP;
      shiftff <= "000000";
      
    ELSIF (rising_edge(sysclk)) THEN
        
      IF (enable = '1') THEN
          
        inmanff <= inman;
        inexpff <= inexp;
      
        zeroff(1) <= zerochk(64);
        FOR k IN 2 TO 2+2*speed LOOP
          zeroff(k) <= zeroff(k-1);
        END LOOP;
      
        shiftff <= shift;
        
      END IF;
  
    END IF;
    
  END PROCESS;
  
  zerochk(1) <= inmanff(1);
  gza: FOR k IN 2 TO 64 GENERATE
    zerochk(k) <= zerochk(k-1) OR inmanff(k);
  END GENERATE;
  
  delma: fp_del
  GENERIC MAP (width=>64,pipes=>1+speed)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>inmanff,cc=>inmandelbus);
  
  gsa: IF (speed = 0) GENERATE
  
    clz: dp_lnclz
    PORT MAP (mantissa=>inmanff,leading=>shift);
  
    sft: dp_lsft64x6
    PORT MAP (inbus=>inmandelbus,shift=>shiftff,
              outbus=>outmanbus);
  
  END GENERATE;

  gsb: IF (speed = 1) GENERATE
  
    clzp: dp_lnclzpipe
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              mantissa=>inmanff,
              leading=>shift);
  
    sftp: dp_lsft64x6pipe
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              inbus=>inmandelbus,shift=>shiftff,
              outbus=>outmanbus);
  
  END GENERATE;
  
  -- add 2 - 1 for right shift to avoid overflow 
  expaddbus <= inexpff + 1;
  
  delxa: fp_del
  GENERIC MAP (width=>11,pipes=>1+speed)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>expaddbus,cc=>expmidbus);
          
  expsubbus <= expmidbus - ("00000" & shiftff);
  
  delxb: fp_del
  GENERIC MAP (width=>11,pipes=>1+speed)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>expsubbus,cc=>expoutbus);

  ppout: PROCESS (sysclk,reset)
  BEGIN
  
    IF (reset = '1') THEN
        
      FOR k IN 1 TO 64 LOOP
        outmanff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
        
      IF (enable = '1') THEN    
        outmanff <= outmanbus;
      END IF;

    END IF;
    
  END PROCESS;
  
  --*** OUTPUTS ***
  outman <= outmanff;
  outexp <= expoutbus;
  zero <= zeroff(2+2*speed);
      
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   DP_LNNORND.VHD                            ***
--***                                             ***
--***   Function: DP LOG Output Block - Simple    ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_lnnornd IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signln : IN STD_LOGIC;
      exponentln : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaln : IN STD_LOGIC_VECTOR (53 DOWNTO 1);
      nanin : IN STD_LOGIC;
      infinityin : IN STD_LOGIC;
      zeroin : IN STD_LOGIC;
        
		signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
      --------------------------------------------------
      nanout : OUT STD_LOGIC;
      overflowout : OUT STD_LOGIC;
      zeroout : OUT STD_LOGIC
		);
END dp_lnnornd;

ARCHITECTURE rtl OF dp_lnnornd IS

  constant expwidth : positive := 11;
  constant manwidth : positive := 52;
  
  signal nanff : STD_LOGIC;
  signal infinityff : STD_LOGIC;
  signal zeroff : STD_LOGIC; 
  signal signff : STD_LOGIC; 
  signal mantissaff : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal exponentff : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  
  signal setmanzero, setexpzero, setmanmax, setexpmax : STD_LOGIC;

BEGIN

  pra: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN
        
      nanff <= '0';
      signff <= '0';
      FOR k IN 1 TO manwidth LOOP
        mantissaff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        exponentff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF(enable = '1') THEN 
      
        signff <= signln;
        nanff <= nanin;
        infinityff <= infinityin;
        zeroff <= zeroin;

        -- nan takes precedence (set max)  
        FOR k IN 1 TO manwidth LOOP
          mantissaff(k) <= (mantissaln(k+1) AND NOT(setmanzero)) OR setmanmax;
        END LOOP;
               
        FOR k IN 1 TO expwidth LOOP
          exponentff(k) <= (exponentln(k) AND NOT(setexpzero)) OR setexpmax;
        END LOOP;
      
      END IF;
             
    END IF;
      
  END PROCESS;
                                                  
--**********************************
--*** CHECK GENERATED CONDITIONS ***   
--**********************************
  
  -- all set to '1' when true
  
  -- set mantissa to 0 when zero or infinity condition
  setmanzero <= NOT(zeroin) OR infinityin;
  -- setmantissa to "11..11" when nan
  setmanmax <= nanin;
  -- set exponent to 0 when zero condition 
  setexpzero <= NOT(zeroin);
  -- set exponent to "11..11" when nan or infinity
  setexpmax <= nanin OR infinityin;
                             
--***************
--*** OUTPUTS ***
--***************

  signout <= signff;   
  mantissaout <= mantissaff;
  exponentout <= exponentff; 
  -----------------------------------------------
  nanout <= nanff;
  overflowout <= infinityff;
  zeroout <= zeroff;

END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   DP_LNRND.VHD                              ***
--***                                             ***
--***   Function: DP LOG Output Block - Rounded   ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_lnrnd IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signln : IN STD_LOGIC;
      exponentln : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaln : IN STD_LOGIC_VECTOR (53 DOWNTO 1);
      nanin : IN STD_LOGIC;
      infinityin : IN STD_LOGIC;
      zeroin : IN STD_LOGIC;
        
		signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
      --------------------------------------------------
      nanout : OUT STD_LOGIC;
      overflowout : OUT STD_LOGIC;
      zeroout : OUT STD_LOGIC
		);
END dp_lnrnd;

ARCHITECTURE rtl OF dp_lnrnd IS

  constant expwidth : positive := 11;
  constant manwidth : positive := 52;
  
  type exponentfftype IS ARRAY (2 DOWNTO 1) OF STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  
  signal zerovec : STD_LOGIC_VECTOR (manwidth-1 DOWNTO 1);
  signal nanff : STD_LOGIC_VECTOR (2 DOWNTO 1);
  signal zeroff : STD_LOGIC_VECTOR (2 DOWNTO 1);
  signal signff : STD_LOGIC_VECTOR (2 DOWNTO 1);
  signal infinityff : STD_LOGIC_VECTOR (2 DOWNTO 1);
  signal manoverflowbitff : STD_LOGIC; 
  signal roundmantissaff, mantissaff : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal exponentnode : STD_LOGIC_VECTOR (expwidth+2 DOWNTO 1);
  signal exponentoneff : STD_LOGIC_VECTOR (expwidth+2 DOWNTO 1);
  signal exponenttwoff : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
    
  signal manoverflow : STD_LOGIC_VECTOR (manwidth+1 DOWNTO 1);
  signal setmanzero, setmanmax : STD_LOGIC;
  signal setexpzero, setexpmax : STD_LOGIC;

BEGIN
    
  gzv: FOR k IN 1 TO manwidth-1 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  pra: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN
        
      nanff <= "00";
      signff <= "00";
      FOR k IN 1 TO manwidth LOOP
        roundmantissaff(k) <= '0';
        mantissaff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth+2 LOOP
        exponentoneff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        exponenttwoff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF(enable = '1') THEN 
      
        nanff(1) <= nanin;
        nanff(2) <= nanff(1);
        infinityff(1) <= infinityin;
        infinityff(2) <= infinityff(1);
        zeroff(1) <= zeroin;
        zeroff(2) <= zeroff(1);
        signff(1) <= signln;
        signff(2) <= signff(1);
       
        manoverflowbitff <= manoverflow(manwidth+1);
        
        roundmantissaff <= mantissaln(manwidth+1 DOWNTO 2) + (zerovec & mantissaln(1));
        
        FOR k IN 1 TO manwidth LOOP
          mantissaff(k) <= (roundmantissaff(k) AND NOT(setmanzero)) OR setmanmax;
        END LOOP;
        
        exponentoneff(expwidth+2 DOWNTO 1) <= "00" & exponentln;                 
        FOR k IN 1 TO expwidth LOOP
          exponenttwoff(k) <= (exponentnode(k) AND NOT(setexpzero)) OR setexpmax;
        END LOOP;
      
      END IF;
             
    END IF;
      
  END PROCESS;
  
  exponentnode <= exponentoneff(expwidth+2 DOWNTO 1) + 
                 (zerovec(expwidth+1 DOWNTO 1) & manoverflowbitff);

--*********************************
--*** PREDICT MANTISSA OVERFLOW ***   
--*********************************
     
  manoverflow(1) <= mantissaln(1);
  gmoa: FOR k IN 2 TO manwidth+1 GENERATE
    manoverflow(k) <= manoverflow(k-1) AND mantissaln(k);
  END GENERATE; 
                                                                 
--**********************************
--*** CHECK GENERATED CONDITIONS ***   
--**********************************
  
  -- all set to '1' when condition true
  
  -- set mantissa to 0 when infinity or zero condition
  setmanzero <= NOT(zeroff(1)) OR infinityff(1);
  -- setmantissa to "11..11" when nan
  setmanmax <= nanff(1);
  -- set exponent to 0 when zero condition 
  setexpzero <= NOT(zeroff(1));
  -- set exponent to "11..11" when nan or infinity
  setexpmax <= nanff(1) OR infinityff(1);
                             
--***************
--*** OUTPUTS ***
--***************
  
  signout <= signff(2);
  mantissaout <= mantissaff;
  exponentout <= exponenttwoff; 
  -----------------------------------------------
  nanout <= nanff(2);
  overflowout <= infinityff(2);
  zeroout <= zeroff(2);

END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   DP_LNRNDPIPE.VHD                          ***
--***                                             ***
--***   Function: DP LOG Output Block - Pipelined ***
--***   Round                                     ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_lnrndpipe IS 
GENERIC (synthesize : integer := 1); 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signln : IN STD_LOGIC;
      exponentln : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaln : IN STD_LOGIC_VECTOR (53 DOWNTO 1);
      nanin : IN STD_LOGIC;
      infinityin : IN STD_LOGIC;
      zeroin : IN STD_LOGIC;
        
		signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
      --------------------------------------------------
      nanout : OUT STD_LOGIC;
      overflowout : OUT STD_LOGIC;
      zeroout : OUT STD_LOGIC
		);
END dp_lnrndpipe;

ARCHITECTURE rtl OF dp_lnrndpipe IS

  constant expwidth : positive := 11;
  constant manwidth : positive := 52;
  
  type exponentfftype IS ARRAY (3 DOWNTO 1) OF STD_LOGIC_VECTOR (expwidth+2 DOWNTO 1);
  
  signal zerovec : STD_LOGIC_VECTOR (manwidth+1 DOWNTO 1);
  signal nanff : STD_LOGIC_VECTOR (3 DOWNTO 1);
  signal zeroff : STD_LOGIC_VECTOR (3 DOWNTO 1);
  signal infinityff : STD_LOGIC_VECTOR (3 DOWNTO 1);
  signal signff : STD_LOGIC_VECTOR (3 DOWNTO 1);
  signal roundmantissanode : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal mantissaff : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal exponentff : exponentfftype;
       
  signal manoverflow : STD_LOGIC_VECTOR (manwidth+1 DOWNTO 1);
  signal manoverflowff : STD_LOGIC;
  signal setmanzero, setmanmax : STD_LOGIC;
  signal setexpzero, setexpmax : STD_LOGIC;

  component dp_fxadd 
  GENERIC (
           width : positive := 64;
           pipes : positive := 1;
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
        carryin : IN STD_LOGIC;
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
  end component;
  
BEGIN
    
  gzv: FOR k IN 1 TO manwidth+1 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  pra: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN

      nanff <= "000";
      signff <= "000";
      infinityff <= "000";
      zeroff <= "000";
      manoverflowff <= '0';
      FOR k IN 1 TO manwidth LOOP
        mantissaff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        exponentff(1)(k) <= '0';
        exponentff(2)(k) <= '0';
        exponentff(3)(k) <= '0';
      END LOOP;
        
    ELSIF (rising_edge(sysclk)) THEN
    
      IF(enable = '1') THEN 
      
        nanff(1) <= nanin;
        nanff(2) <= nanff(1);
        nanff(3) <= nanff(2);
        infinityff(1) <= infinityin;
        infinityff(2) <= infinityff(1);
        infinityff(3) <= infinityff(2);
        zeroff(1) <= zeroin;
        zeroff(2) <= zeroff(1);
        zeroff(3) <= zeroff(2);
        signff(1) <= signln;
        signff(2) <= signff(1);
        signff(3) <= signff(2);
        
        manoverflowff <= manoverflow(53);
        
        -- nan takes precedence (set max)  
        FOR k IN 1 TO manwidth LOOP
          mantissaff(k) <= (roundmantissanode(k) AND NOT(setmanzero)) OR setmanmax;
        END LOOP;
        
        exponentff(1)(expwidth+2 DOWNTO 1) <= "00" & exponentln(expwidth DOWNTO 1);
        exponentff(2)(expwidth+2 DOWNTO 1) <= (exponentff(1)(expwidth+2 DOWNTO 1)) + 
                                              (zerovec(expwidth+1 DOWNTO 1) & manoverflowff);                 
        FOR k IN 1 TO expwidth LOOP
          exponentff(3)(k) <= (exponentff(2)(k) AND NOT(setexpzero)) OR setexpmax;
        END LOOP;
      
      END IF;
             
    END IF;
      
  END PROCESS;
       
  rndadd: dp_fxadd 
  GENERIC MAP(width=>manwidth,pipes=>2,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>mantissaln(manwidth+1 DOWNTO 2),bb=>zerovec(manwidth DOWNTO 1),
            carryin=>mantissaln(1),
            cc=>roundmantissanode);

--*********************************
--*** PREDICT MANTISSA OVERFLOW ***   
--*********************************
     
  manoverflow(1) <= mantissaln(1);
  gmoa: FOR k IN 2 TO 53 GENERATE
    manoverflow(k) <= manoverflow(k-1) AND mantissaln(k);
  END GENERATE;                                           
    
--**********************************
--*** CHECK GENERATED CONDITIONS ***   
--**********************************
                    
  -- all set to '1' when true
  
  -- set mantissa to 0 when infinity or zero condition
  setmanzero <= infinityff(2) OR NOT(zeroff(2));
  -- setmantissa to "11..11" when nan
  setmanmax <= nanff(2);
  -- set exponent to 0 when zero condition 
  setexpzero <= NOT(zeroff(2));
  -- set exponent to "11..11" when nan or infinity
  setexpmax <= nanff(2) OR infinityff(2);
            
--***************
--*** OUTPUTS ***
--***************

  signout <= signff(3);
  mantissaout <= mantissaff;
  exponentout <= exponentff(3)(expwidth DOWNTO 1); 
  -----------------------------------------------
  nanout <= nanff(3);
  overflowout <= infinityff(3);
  zeroout <= zeroff(3);
  
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   DOUBLE PRECISION LOG(LN) - TOP LEVEL      ***
--***                                             ***
--***   DP_LOG.VHD                                ***
--***                                             ***
--***   Function: IEEE754 DP LN()                 ***
--***                                             ***
--***   11/08/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** Latency = 27 + 7*DoubleSpeed +              ***
--***           RoundConvert*(1+DoubleSpeed)      ***
--*** DoubleSpeed = 0, RoundConvert = 0 : 27      ***
--*** DoubleSpeed = 1, RoundConvert = 0 : 34      ***
--*** DoubleSpeed = 0, RoundConvert = 1 : 28      ***
--*** DoubleSpeed = 1, RoundConvert = 1 : 36      ***
--***                                             ***
--***************************************************

ENTITY dp_log IS 
GENERIC (
         roundconvert : integer := 0; -- 0 = no round, 1 = round
         doublespeed : integer := 0; -- 0/1
         device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
         synthesize : integer := 1      -- 0/1    
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (52 DOWNTO 1);

		  signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
      --------------------------------------------------
      nanout : OUT STD_LOGIC;
      overflowout : OUT STD_LOGIC;
      zeroout : OUT STD_LOGIC
		);
END dp_log;

ARCHITECTURE rtl OF dp_log IS
  
  constant expwidth : positive := 11;
  constant manwidth : positive := 52;
  
  constant coredepth : positive := 26 + 7*doublespeed;

  signal signinff : STD_LOGIC_VECTOR (2 DOWNTO 1);
  signal maninff : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal expinff : STD_LOGIC_VECTOR (expwidth DOWNTO 1);   
  signal signnode : STD_LOGIC;
  signal mantissanode : STD_LOGIC_VECTOR (53 DOWNTO 1);
  signal exponentnode : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal zeronode : STD_LOGIC;
              
  -- conditions
  signal zeroman : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal zeroexp : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal maxexp : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal zeromaninff : STD_LOGIC;
  signal zeroexpinff : STD_LOGIC;
  signal maxexpinff : STD_LOGIC;
  signal naninff : STD_LOGIC;
  signal nanff : STD_LOGIC_VECTOR (coredepth-3 DOWNTO 1);
  signal infinityinff : STD_LOGIC;
  signal infinityff : STD_LOGIC_VECTOR (coredepth-3 DOWNTO 1);
      
  component dp_ln_core 
  GENERIC (
           doublespeed : integer := 0; -- 0/1
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 1 -- 0/1       
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aaman : IN STD_LOGIC_VECTOR (52 DOWNTO 1); 
        aaexp : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
      
        ccman : OUT STD_LOGIC_VECTOR (53 DOWNTO 1);
        ccexp : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
        ccsgn : OUT STD_LOGIC;
        zeroout : OUT STD_LOGIC
       );
  end component;
  
  component dp_lnnornd
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        signln : IN STD_LOGIC;
        exponentln : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
        mantissaln : IN STD_LOGIC_VECTOR (53 DOWNTO 1);
        nanin : IN STD_LOGIC;
        infinityin : IN STD_LOGIC;
        zeroin : IN STD_LOGIC;

        signout : OUT STD_LOGIC;
        exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
        mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
        --------------------------------------------------
        nanout : OUT STD_LOGIC;
        overflowout : OUT STD_LOGIC;
        zeroout : OUT STD_LOGIC
		  );
  end component;
                        
  component dp_lnrnd
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        signln : IN STD_LOGIC;
        exponentln : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
        mantissaln : IN STD_LOGIC_VECTOR (53 DOWNTO 1);
        nanin : IN STD_LOGIC;
        infinityin : IN STD_LOGIC;
        zeroin : IN STD_LOGIC;

        signout : OUT STD_LOGIC;
        exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
        mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
        --------------------------------------------------
        nanout : OUT STD_LOGIC;
        overflowout : OUT STD_LOGIC;
        zeroout : OUT STD_LOGIC
		  );
  end component;

  component dp_lnrndpipe
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        signln : IN STD_LOGIC;
        exponentln : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
        mantissaln : IN STD_LOGIC_VECTOR (53 DOWNTO 1);
        nanin : IN STD_LOGIC;
        infinityin : IN STD_LOGIC;
        zeroin : IN STD_LOGIC;

        signout : OUT STD_LOGIC;
        exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
        mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
        --------------------------------------------------
        nanout : OUT STD_LOGIC;
        overflowout : OUT STD_LOGIC;
        zeroout : OUT STD_LOGIC
		  );
  end component;
  
BEGIN

  pma: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN

      FOR k IN 1 TO manwidth LOOP
        maninff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        expinff(k) <= '0';
      END LOOP;
      signinff <= "00";
    
    ELSIF (rising_edge(sysclk)) THEN

      IF (enable = '1') THEN

        maninff <= mantissain;
        expinff <= exponentin;
        signinff(1) <= signin;
        signinff(2) <= signinff(1);
                                                  
      END IF;
  
    END IF;
  
  END PROCESS;

--********************
--*** CHECK INPUTS ***
--********************

  zeroman(1) <= maninff(1);
  gca: FOR k IN 2 TO manwidth GENERATE
    zeroman(k) <= zeroman(k-1) OR maninff(k);
  END GENERATE; 
  zeroexp(1) <= expinff(1);
  gcb: FOR k IN 2 TO expwidth GENERATE
    zeroexp(k) <= zeroexp(k-1) OR expinff(k);
  END GENERATE;
  maxexp(1) <= expinff(1);
  gcc: FOR k IN 2 TO expwidth GENERATE
    maxexp(k) <= maxexp(k-1) AND expinff(k);
  END GENERATE;

  pcc: PROCESS (sysclk,reset)
  BEGIN
    
    IF (reset = '1') THEN
      
      zeromaninff <= '0';
      zeroexpinff <= '0';
      maxexpinff <= '0';  
      naninff <= '0';
      FOR k IN 1 TO coredepth-3 LOOP
        nanff(k) <= '0';
      END LOOP;
     
    ELSIF (rising_edge(sysclk)) THEN
            
      IF (enable = '1') THEN

        zeromaninff <= NOT(zeroman(manwidth));
        zeroexpinff <= NOT(zeroexp(expwidth));
        maxexpinff <= maxexp(expwidth);
    
        -- infinity when exp = zero
        -- nan when man != 0, exp = max
    
        -- all ffs '1' when condition true
        naninff <= (zeromaninff AND maxexpinff) OR signinff(2);
        infinityinff <= zeroexpinff OR maxexpinff;

        -- nan output when nan input
        nanff(1) <= naninff;
        FOR k IN 2 TO coredepth-3 LOOP
          nanff(k) <= nanff(k-1);
        END LOOP;
        
        infinityff(1) <= infinityinff;
        FOR k IN 2 TO coredepth-3 LOOP
          infinityff(k) <= infinityff(k-1);
        END LOOP;
      
      END IF;
   
    END IF;

  END PROCESS;


--***************
--*** LN CORE ***
--***************

  lncore: dp_ln_core
  GENERIC MAP (doublespeed=>doublespeed,device=>device,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aaman=>mantissain,aaexp=>exponentin,
            ccman=>mantissanode,ccexp=>exponentnode,ccsgn=>signnode,
            zeroout=>zeronode);
  
--************************
--*** ROUND AND OUTPUT ***
--************************

  gra: IF (roundconvert = 0) GENERATE

    norndout: dp_lnnornd
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              signln=>signnode,
              exponentln=>exponentnode,
              mantissaln=>mantissanode,
              nanin=>nanff(coredepth-3),
              infinityin=>infinityff(coredepth-3),
              zeroin=>zeronode,

              signout=>signout,
              exponentout=>exponentout,
              mantissaout=>mantissaout,
              nanout=>nanout,overflowout=>overflowout,zeroout=>zeroout);
            
  END GENERATE;
  
  grb: IF (roundconvert = 1 AND doublespeed = 0) GENERATE

    rndout: dp_lnrnd
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              signln=>signnode,
              exponentln=>exponentnode,
              mantissaln=>mantissanode,
              nanin=>nanff(coredepth-3),
              infinityin=>infinityff(coredepth-3),
              zeroin=>zeronode,

              signout=>signout,
              exponentout=>exponentout,
              mantissaout=>mantissaout,
              nanout=>nanout,overflowout=>overflowout,zeroout=>zeroout);
            
  END GENERATE;

  grc: IF (roundconvert = 1 AND doublespeed = 1) GENERATE
    
    rndoutpipe: dp_lnrndpipe
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              signln=>signnode,
              exponentln=>exponentnode,
              mantissaln=>mantissanode,
              nanin=>nanff(coredepth-3),
              infinityin=>infinityff(coredepth-3),
              zeroin=>zeronode,

              signout=>signout,
              exponentout=>exponentout,
              mantissaout=>mantissaout,
              nanout=>nanout,overflowout=>overflowout,zeroout=>zeroout);
            
  END GENERATE;
  
END rtl;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOAT CONVERT - CORE LEVEL                ***
--***                                             ***
--***   DP_LSFT64.VHD                             ***
--***                                             ***
--***   Function: Combinatorial Left Shift 64     ***
--***             Bits                            ***
--***                                             ***
--***   01/12/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_lsft64 IS
PORT (
      inbus : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
      shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);      
        
      outbus : OUT STD_LOGIC_VECTOR (64 DOWNTO 1)    
     );
END dp_lsft64;

ARCHITECTURE rtl of dp_lsft64 IS

  signal levzip, levone, levtwo, levthr : STD_LOGIC_VECTOR (64 DOWNTO 1);
  
BEGIN

  levzip <= inbus;
  
  gla: FOR k IN 4 TO 64 GENERATE
    levone(k) <= (levzip(k)   AND NOT(shift(2)) AND NOT(shift(1))) OR 
                 (levzip(k-1) AND NOT(shift(2)) AND     shift(1)) OR
                 (levzip(k-2) AND     shift(2)  AND NOT(shift(1))) OR
                 (levzip(k-3) AND     shift(2)  AND     shift(1));
  END GENERATE;
  levone(3) <= (levzip(3) AND NOT(shift(2)) AND NOT(shift(1))) OR 
               (levzip(2) AND NOT(shift(2)) AND     shift(1)) OR
               (levzip(1) AND     shift(2)  AND NOT(shift(1)));
  levone(2) <= (levzip(2) AND NOT(shift(2)) AND NOT(shift(1))) OR 
               (levzip(1) AND NOT(shift(2)) AND     shift(1));                
  levone(1) <= (levzip(1) AND NOT(shift(2)) AND NOT(shift(1)));
                               
  glba: FOR k IN 13 TO 64 GENERATE
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR 
                 (levone(k-4)  AND NOT(shift(4)) AND     shift(3)) OR
                 (levone(k-8)  AND     shift(4)  AND NOT(shift(3))) OR
                 (levone(k-12) AND     shift(4)  AND     shift(3));
  END GENERATE;  
  glbb: FOR k IN 9 TO 12 GENERATE            
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR 
                 (levone(k-4)  AND NOT(shift(4)) AND     shift(3)) OR
                 (levone(k-8)  AND     shift(4)  AND NOT(shift(3)));             
  END GENERATE;
  glbc: FOR k IN 5 TO 8 GENERATE            
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR 
                 (levone(k-4)  AND NOT(shift(4)) AND     shift(3));           
  END GENERATE;  
  glbd: FOR k IN 1 TO 4 GENERATE            
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3)));          
  END GENERATE;    

  glca: FOR k IN 49 TO 64 GENERATE
    levthr(k) <= (levtwo(k)    AND NOT(shift(6)) AND NOT(shift(5))) OR 
                 (levtwo(k-16) AND NOT(shift(6)) AND     shift(5)) OR
                 (levtwo(k-32) AND     shift(6)  AND NOT(shift(5))) OR
                 (levtwo(k-48) AND     shift(6)  AND     shift(5));
  END GENERATE;  
  glcb: FOR k IN 33 TO 48 GENERATE
    levthr(k) <= (levtwo(k)    AND NOT(shift(6)) AND NOT(shift(5))) OR 
                 (levtwo(k-16) AND NOT(shift(6)) AND     shift(5)) OR
                 (levtwo(k-32) AND     shift(6)  AND NOT(shift(5)));
  END GENERATE; 
  glcc: FOR k IN 17 TO 32 GENERATE
    levthr(k) <= (levtwo(k)    AND NOT(shift(6)) AND NOT(shift(5))) OR 
                 (levtwo(k-16) AND NOT(shift(6)) AND     shift(5));
  END GENERATE; 
  glcd: FOR k IN 1 TO 16 GENERATE
    levthr(k) <= (levtwo(k)    AND NOT(shift(6)) AND NOT(shift(5)));
  END GENERATE; 
      
  outbus <= levthr;
  
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   DP_LSFT64X6.VHD                           ***
--***                                             ***
--***   Function: Double Precision Left Shift     ***
--***   (Combinatorial)                           ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_lsft64x6 IS 
PORT (
      inbus : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
      shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);
      outbus : OUT STD_LOGIC_VECTOR (64 DOWNTO 1)
    );
END dp_lsft64x6;

ARCHITECTURE rtl OF dp_lsft64x6 IS

  signal leftone, lefttwo, leftthr : STD_LOGIC_VECTOR (64 DOWNTO 1);
            
BEGIN
  
  leftone(1) <=  inbus(1)     AND NOT(shift(2)) AND NOT(shift(1));
  leftone(2) <= (inbus(2)     AND NOT(shift(2)) AND NOT(shift(1))) OR
                (inbus(1)     AND NOT(shift(2)) AND     shift(1)); 
  leftone(3) <= (inbus(3)     AND NOT(shift(2)) AND NOT(shift(1))) OR
                (inbus(2)     AND NOT(shift(2)) AND     shift(1)) OR
                (inbus(1)     AND     shift(2)  AND NOT(shift(1))); 
  gla: FOR k IN 4 TO 64 GENERATE
    leftone(k) <= (inbus(k)   AND NOT(shift(2)) AND NOT(shift(1))) OR
                  (inbus(k-1) AND NOT(shift(2)) AND     shift(1)) OR
                  (inbus(k-2) AND     shift(2)  AND NOT(shift(1))) OR
                  (inbus(k-3) AND     shift(2)  AND     shift(1));
  END GENERATE;
             
  glb: FOR k IN 1 TO 4 GENERATE
    lefttwo(k) <=  leftone(k)    AND NOT(shift(4)) AND NOT(shift(3));
  END GENERATE;
  glc: FOR k IN 5 TO 8 GENERATE
    lefttwo(k) <= (leftone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                  (leftone(k-4)  AND NOT(shift(4)) AND     shift(3)); 
  END GENERATE;
  gld: FOR k IN 9 TO 12 GENERATE
    lefttwo(k) <= (leftone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                  (leftone(k-4)  AND NOT(shift(4)) AND     shift(3)) OR
                  (leftone(k-8)  AND     shift(4)  AND NOT(shift(3))); 
  END GENERATE;
  gle: FOR k IN 13 TO 64 GENERATE
    lefttwo(k) <= (leftone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                  (leftone(k-4)  AND NOT(shift(4)) AND     shift(3)) OR
                  (leftone(k-8)  AND     shift(4)  AND NOT(shift(3)))  OR
                  (leftone(k-12) AND     shift(4)  AND     shift(3)); 
  END GENERATE;
  
  glf: FOR k IN 1 TO 16 GENERATE
    leftthr(k) <=  lefttwo(k)    AND NOT(shift(6)) AND NOT(shift(5));
  END GENERATE;
  glg: FOR k IN 17 TO 32 GENERATE
    leftthr(k) <= (lefttwo(k)    AND NOT(shift(6)) AND NOT(shift(5))) OR
                  (lefttwo(k-16) AND NOT(shift(6)) AND     shift(5)); 
  END GENERATE;
  glh: FOR k IN 33 TO 48 GENERATE
    leftthr(k) <= (lefttwo(k)    AND NOT(shift(6)) AND NOT(shift(5))) OR
                  (lefttwo(k-16) AND NOT(shift(6)) AND     shift(5)) OR
                  (lefttwo(k-32) AND     shift(6)  AND NOT(shift(5))); 
  END GENERATE;
  gli: FOR k IN 49 TO 64 GENERATE
    leftthr(k) <= (lefttwo(k)    AND NOT(shift(6)) AND NOT(shift(5))) OR
                  (lefttwo(k-16) AND NOT(shift(6)) AND     shift(5)) OR
                  (lefttwo(k-32) AND     shift(6)  AND NOT(shift(5)))  OR
                  (lefttwo(k-48) AND     shift(6)  AND     shift(5)); 
  END GENERATE;
    
  outbus <= leftthr;        
            
END rtl;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOAT CONVERT - CORE LEVEL                ***
--***                                             ***
--***   DP_LSFT64X64.VHD                          ***
--***                                             ***
--***   Function: Combinatorial Left Shift        ***
--***             (max 1.52 to 64.0)              ***
--***                                             ***
--***   07/12/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_lsft64x64 IS
PORT (
      inbus : IN STD_LOGIC_VECTOR (116 DOWNTO 1);
      shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);      
        
      outbus : OUT STD_LOGIC_VECTOR (116 DOWNTO 1)    
     );
END dp_lsft64x64;

ARCHITECTURE rtl of dp_lsft64x64 IS

  signal levzip, levone, levtwo, levthr : STD_LOGIC_VECTOR (116 DOWNTO 1);
 
BEGIN
  
  levzip <= inbus;
  
  gla: FOR k IN 4 TO 116 GENERATE
    levone(k) <= (levzip(k)   AND NOT(shift(2)) AND NOT(shift(1))) OR 
                 (levzip(k-1) AND NOT(shift(2)) AND     shift(1)) OR
                 (levzip(k-2) AND     shift(2)  AND NOT(shift(1))) OR
                 (levzip(k-3) AND     shift(2)  AND     shift(1));
  END GENERATE;
  levone(3) <= (levzip(3) AND NOT(shift(2)) AND NOT(shift(1))) OR 
               (levzip(2) AND NOT(shift(2)) AND     shift(1)) OR
               (levzip(1) AND     shift(2)  AND NOT(shift(1)));
  levone(2) <= (levzip(2) AND NOT(shift(2)) AND NOT(shift(1))) OR 
               (levzip(1) AND NOT(shift(2)) AND     shift(1));                
  levone(1) <= (levzip(1) AND NOT(shift(2)) AND NOT(shift(1)));
                               
  glba: FOR k IN 13 TO 116 GENERATE
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR 
                 (levone(k-4)  AND NOT(shift(4)) AND     shift(3)) OR
                 (levone(k-8)  AND     shift(4)  AND NOT(shift(3))) OR
                 (levone(k-12) AND     shift(4)  AND     shift(3));
  END GENERATE;  
  glbb: FOR k IN 9 TO 12 GENERATE            
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR 
                 (levone(k-4)  AND NOT(shift(4)) AND     shift(3)) OR
                 (levone(k-8)  AND     shift(4)  AND NOT(shift(3)));             
  END GENERATE;
  glbc: FOR k IN 5 TO 8 GENERATE            
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR 
                 (levone(k-4)  AND NOT(shift(4)) AND     shift(3));           
  END GENERATE;  
  glbd: FOR k IN 1 TO 4 GENERATE            
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3)));          
  END GENERATE;    

  glca: FOR k IN 49 TO 116 GENERATE
    levthr(k) <= (levtwo(k)    AND NOT(shift(6)) AND NOT(shift(5))) OR 
                 (levtwo(k-16) AND NOT(shift(6)) AND     shift(5)) OR
                 (levtwo(k-32) AND     shift(6)  AND NOT(shift(5))) OR
                 (levtwo(k-48) AND     shift(6)  AND     shift(5));
  END GENERATE;  
  glcb: FOR k IN 33 TO 48 GENERATE
    levthr(k) <= (levtwo(k)    AND NOT(shift(6)) AND NOT(shift(5))) OR 
                 (levtwo(k-16) AND NOT(shift(6)) AND     shift(5)) OR
                 (levtwo(k-32) AND     shift(6)  AND NOT(shift(5)));
  END GENERATE; 
  glcc: FOR k IN 17 TO 32 GENERATE
    levthr(k) <= (levtwo(k)    AND NOT(shift(6)) AND NOT(shift(5))) OR 
                 (levtwo(k-16) AND NOT(shift(6)) AND     shift(5));
  END GENERATE; 
  glcd: FOR k IN 1 TO 16 GENERATE
    levthr(k) <= (levtwo(k)    AND NOT(shift(6)) AND NOT(shift(5)));
  END GENERATE; 
      
  outbus <= levthr;
  
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   DP_LSFT64X6PIPE.VHD                       ***
--***                                             ***
--***   Function: Double Precision Left Shift     ***
--***   (Pipelined)                               ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_lsft64x6pipe IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      inbus : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
      shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);
      outbus : OUT STD_LOGIC_VECTOR (64 DOWNTO 1)
    );
END dp_lsft64x6pipe;

ARCHITECTURE rtl OF dp_lsft64x6pipe IS

  signal leftone, lefttwo, leftthr : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal lefttwoff : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal shiftff : STD_LOGIC_VECTOR (6 DOWNTO 5);
            
BEGIN
  
  leftone(1) <=  inbus(1)     AND NOT(shift(2)) AND NOT(shift(1));
  leftone(2) <= (inbus(2)     AND NOT(shift(2)) AND NOT(shift(1))) OR
                (inbus(1)     AND NOT(shift(2)) AND     shift(1)); 
  leftone(3) <= (inbus(3)     AND NOT(shift(2)) AND NOT(shift(1))) OR
                (inbus(2)     AND NOT(shift(2)) AND     shift(1)) OR
                (inbus(1)     AND     shift(2)  AND NOT(shift(1))); 
  gla: FOR k IN 4 TO 64 GENERATE
    leftone(k) <= (inbus(k)   AND NOT(shift(2)) AND NOT(shift(1))) OR
                  (inbus(k-1) AND NOT(shift(2)) AND     shift(1)) OR
                  (inbus(k-2) AND     shift(2)  AND NOT(shift(1))) OR
                  (inbus(k-3) AND     shift(2)  AND     shift(1));
  END GENERATE;
             
  glb: FOR k IN 1 TO 4 GENERATE
    lefttwo(k) <=  leftone(k)    AND NOT(shift(4)) AND NOT(shift(3));
  END GENERATE;
  glc: FOR k IN 5 TO 8 GENERATE
    lefttwo(k) <= (leftone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                  (leftone(k-4)  AND NOT(shift(4)) AND     shift(3)); 
  END GENERATE;
  gld: FOR k IN 9 TO 12 GENERATE
    lefttwo(k) <= (leftone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                  (leftone(k-4)  AND NOT(shift(4)) AND     shift(3)) OR
                  (leftone(k-8)  AND     shift(4)  AND NOT(shift(3))); 
  END GENERATE;
  gle: FOR k IN 13 TO 64 GENERATE
    lefttwo(k) <= (leftone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                  (leftone(k-4)  AND NOT(shift(4)) AND     shift(3)) OR
                  (leftone(k-8)  AND     shift(4)  AND NOT(shift(3)))  OR
                  (leftone(k-12) AND     shift(4)  AND     shift(3)); 
  END GENERATE;
  
  ppa: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN
        
      FOR k IN 1 TO 64 LOOP
        lefttwoff(k) <= '0';
      END LOOP;
      shiftff <= "00";
      
    ELSIF (rising_edge(sysclk)) THEN
    
      lefttwoff <= lefttwo;
      shiftff <= shift(6 DOWNTO 5);
              
    END IF;
      
  END PROCESS;
  
  glf: FOR k IN 1 TO 16 GENERATE
    leftthr(k) <=  lefttwoff(k)    AND NOT(shiftff(6)) AND NOT(shiftff(5));
  END GENERATE;
  glg: FOR k IN 17 TO 32 GENERATE
    leftthr(k) <= (lefttwoff(k)    AND NOT(shiftff(6)) AND NOT(shiftff(5))) OR
                  (lefttwoff(k-16) AND NOT(shiftff(6)) AND     shiftff(5)); 
  END GENERATE;
  glh: FOR k IN 33 TO 48 GENERATE
    leftthr(k) <= (lefttwoff(k)    AND NOT(shiftff(6)) AND NOT(shiftff(5))) OR
                  (lefttwoff(k-16) AND NOT(shiftff(6)) AND     shiftff(5)) OR
                  (lefttwoff(k-32) AND     shiftff(6)  AND NOT(shiftff(5))); 
  END GENERATE;
  gli: FOR k IN 49 TO 64 GENERATE
    leftthr(k) <= (lefttwoff(k)    AND NOT(shiftff(6)) AND NOT(shiftff(5))) OR
                  (lefttwoff(k-16) AND NOT(shiftff(6)) AND     shiftff(5)) OR
                  (lefttwoff(k-32) AND     shiftff(6)  AND NOT(shiftff(5)))  OR
                  (lefttwoff(k-48) AND     shiftff(6)  AND     shiftff(5)); 
  END GENERATE;
    
  outbus <= leftthr;        
            
END rtl;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOAT CONVERT - CORE LEVEL                **
--***                                             ***
--***   DP_LSFTPIPE64.VHD                         ***
--***                                             ***
--***   Function: Pipelined Left Shift 64 Bits    ***
--***                                             ***
--***   01/12/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_lsftpipe64 IS
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      inbus : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
      shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);      
        
      outbus : OUT STD_LOGIC_VECTOR (64 DOWNTO 1)    
     );
END dp_lsftpipe64;

ARCHITECTURE rtl of dp_lsftpipe64 IS

  signal levzip, levone, levtwo, levtwoff, levthr : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal shiftff : STD_LOGIC_VECTOR (6 DOWNTO 5);
  
BEGIN

  levzip <= inbus;
  
  gla: FOR k IN 4 TO 64 GENERATE
    levone(k) <= (levzip(k)   AND NOT(shift(2)) AND NOT(shift(1))) OR 
                 (levzip(k-1) AND NOT(shift(2)) AND     shift(1)) OR
                 (levzip(k-2) AND     shift(2)  AND NOT(shift(1))) OR
                 (levzip(k-3) AND     shift(2)  AND     shift(1));
  END GENERATE;
  levone(3) <= (levzip(3) AND NOT(shift(2)) AND NOT(shift(1))) OR 
               (levzip(2) AND NOT(shift(2)) AND     shift(1)) OR
               (levzip(1) AND     shift(2)  AND NOT(shift(1)));
  levone(2) <= (levzip(2) AND NOT(shift(2)) AND NOT(shift(1))) OR 
               (levzip(1) AND NOT(shift(2)) AND     shift(1));                
  levone(1) <= (levzip(1) AND NOT(shift(2)) AND NOT(shift(1)));
                               
  glba: FOR k IN 13 TO 64 GENERATE
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR 
                 (levone(k-4)  AND NOT(shift(4)) AND     shift(3)) OR
                 (levone(k-8)  AND     shift(4)  AND NOT(shift(3))) OR
                 (levone(k-12) AND     shift(4)  AND     shift(3));
  END GENERATE;  
  glbb: FOR k IN 9 TO 12 GENERATE            
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR 
                 (levone(k-4)  AND NOT(shift(4)) AND     shift(3)) OR
                 (levone(k-8)  AND     shift(4)  AND NOT(shift(3)));             
  END GENERATE;
  glbc: FOR k IN 5 TO 8 GENERATE            
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR 
                 (levone(k-4)  AND NOT(shift(4)) AND     shift(3));           
  END GENERATE;  
  glbd: FOR k IN 1 TO 4 GENERATE            
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3)));          
  END GENERATE;    
  
  pp: PROCESS (sysclk,reset)
  BEGIN
    
    IF (reset = '1') THEN
        
      FOR k IN 1 TO 64 LOOP
        levtwoff(k) <= '0';
      END LOOP;
      shiftff <= "00";
      
    ELSIF (rising_edge(sysclk)) THEN
        
      IF (enable = '1') THEN
          
        levtwoff <= levtwo;
        shiftff <= shift(6 DOWNTO 5);
        
      END IF;
  
    END IF;
    
  END PROCESS;
  
  glca: FOR k IN 49 TO 64 GENERATE
    levthr(k) <= (levtwoff(k)    AND NOT(shiftff(6)) AND NOT(shiftff(5))) OR 
                 (levtwoff(k-16) AND NOT(shiftff(6)) AND     shiftff(5)) OR
                 (levtwoff(k-32) AND     shiftff(6)  AND NOT(shiftff(5))) OR
                 (levtwoff(k-48) AND     shiftff(6)  AND     shiftff(5));
  END GENERATE;  
  glcb: FOR k IN 33 TO 48 GENERATE
    levthr(k) <= (levtwoff(k)    AND NOT(shiftff(6)) AND NOT(shiftff(5))) OR 
                 (levtwoff(k-16) AND NOT(shiftff(6)) AND     shiftff(5)) OR
                 (levtwoff(k-32) AND     shiftff(6)  AND NOT(shiftff(5)));
  END GENERATE; 
  glcc: FOR k IN 17 TO 32 GENERATE
    levthr(k) <= (levtwoff(k)    AND NOT(shiftff(6)) AND NOT(shiftff(5))) OR 
                 (levtwoff(k-16) AND NOT(shiftff(6)) AND     shiftff(5));
  END GENERATE; 
  glcd: FOR k IN 1 TO 16 GENERATE
    levthr(k) <= (levtwoff(k)    AND NOT(shiftff(6)) AND NOT(shiftff(5)));
  END GENERATE; 
      
  outbus <= levthr;
  
END rtl;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOAT CONVERT - CORE LEVEL                ***
--***                                             ***
--***   DP_LSFTPIPE64X64.VHD                      ***
--***                                             ***
--***   Function: Pipelined Left Shift            ***
--***             (max 1.52 to 64.0)              ***
--***                                             ***
--***   07/12/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_lsftpipe64x64 IS
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      inbus : IN STD_LOGIC_VECTOR (116 DOWNTO 1);
      shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);      
        
      outbus : OUT STD_LOGIC_VECTOR (116 DOWNTO 1)    
     );
END dp_lsftpipe64x64;

ARCHITECTURE rtl of dp_lsftpipe64x64 IS

  signal levzip, levone, levtwo, levthr : STD_LOGIC_VECTOR (116 DOWNTO 1);
  signal levtwoff : STD_LOGIC_VECTOR (116 DOWNTO 1);
  signal shiftff : STD_LOGIC_VECTOR (6 DOWNTO 5);
 
BEGIN
  
  levzip <= inbus;
  
  gla: FOR k IN 4 TO 116 GENERATE
    levone(k) <= (levzip(k)   AND NOT(shift(2)) AND NOT(shift(1))) OR 
                 (levzip(k-1) AND NOT(shift(2)) AND     shift(1)) OR
                 (levzip(k-2) AND     shift(2)  AND NOT(shift(1))) OR
                 (levzip(k-3) AND     shift(2)  AND     shift(1));
  END GENERATE;
  levone(3) <= (levzip(3) AND NOT(shift(2)) AND NOT(shift(1))) OR 
               (levzip(2) AND NOT(shift(2)) AND     shift(1)) OR
               (levzip(1) AND     shift(2)  AND NOT(shift(1)));
  levone(2) <= (levzip(2) AND NOT(shift(2)) AND NOT(shift(1))) OR 
               (levzip(1) AND NOT(shift(2)) AND     shift(1));                
  levone(1) <= (levzip(1) AND NOT(shift(2)) AND NOT(shift(1)));
                               
  glba: FOR k IN 13 TO 116 GENERATE
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR 
                 (levone(k-4)  AND NOT(shift(4)) AND     shift(3)) OR
                 (levone(k-8)  AND     shift(4)  AND NOT(shift(3))) OR
                 (levone(k-12) AND     shift(4)  AND     shift(3));
  END GENERATE;  
  glbb: FOR k IN 9 TO 12 GENERATE            
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR 
                 (levone(k-4)  AND NOT(shift(4)) AND     shift(3)) OR
                 (levone(k-8)  AND     shift(4)  AND NOT(shift(3)));             
  END GENERATE;
  glbc: FOR k IN 5 TO 8 GENERATE            
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR 
                 (levone(k-4)  AND NOT(shift(4)) AND     shift(3));           
  END GENERATE;  
  glbd: FOR k IN 1 TO 4 GENERATE            
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3)));          
  END GENERATE;    

  pp: PROCESS (sysclk,reset)
  BEGIN
    
    IF (reset = '1') THEN
        
      FOR k IN 1 TO 116 LOOP
        levtwoff(k) <= '0';
      END LOOP;
      shiftff <= "00";
      
    ELSIF (rising_edge(sysclk)) THEN
        
      IF (enable = '1') THEN
          
        levtwoff <= levtwo;
        shiftff <= shift(6 DOWNTO 5);
        
      END IF;
  
    END IF;
    
  END PROCESS;
  
  glca: FOR k IN 49 TO 116 GENERATE
    levthr(k) <= (levtwoff(k)    AND NOT(shiftff(6)) AND NOT(shiftff(5))) OR 
                 (levtwoff(k-16) AND NOT(shiftff(6)) AND     shiftff(5)) OR
                 (levtwoff(k-32) AND     shiftff(6)  AND NOT(shiftff(5))) OR
                 (levtwoff(k-48) AND     shiftff(6)  AND     shiftff(5));
  END GENERATE;  
  glcb: FOR k IN 33 TO 48 GENERATE
    levthr(k) <= (levtwoff(k)    AND NOT(shiftff(6)) AND NOT(shiftff(5))) OR 
                 (levtwoff(k-16) AND NOT(shiftff(6)) AND     shiftff(5)) OR
                 (levtwoff(k-32) AND     shiftff(6)  AND NOT(shiftff(5)));
  END GENERATE; 
  glcc: FOR k IN 17 TO 32 GENERATE
    levthr(k) <= (levtwoff(k)    AND NOT(shiftff(6)) AND NOT(shiftff(5))) OR 
                 (levtwoff(k-16) AND NOT(shiftff(6)) AND     shiftff(5));
  END GENERATE; 
  glcd: FOR k IN 1 TO 16 GENERATE
    levthr(k) <= (levtwoff(k)    AND NOT(shiftff(6)) AND NOT(shiftff(5)));
  END GENERATE; 
      
  outbus <= levthr;
  
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   ALTERA FLOATING POINT DATAPATH COMPILER   ***
--***                                             ***
--***   DP_NEG.VHD                                ***
--***                                             ***
--***   Function: Single Precision Negative Value ***
--***                                             ***
--***   Created 12/09/09                          ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_neg IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (52 DOWNTO 1);

		  signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
		  satout, zeroout, nanout : OUT STD_LOGIC
		);
END dp_neg;

ARCHITECTURE rtl OF dp_neg IS
 
  signal signff : STD_LOGIC;
  signal exponentff : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal mantissaff : STD_LOGIC_VECTOR (52 DOWNTO 1);
  signal expnode : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal expzerochk, expmaxchk : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal expzero, expmax : STD_LOGIC;
  signal manzerochk : STD_LOGIC_VECTOR (52 DOWNTO 1);
  signal manzero, mannonzero : STD_LOGIC; 

BEGIN
    
  pin: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
    
      signff <= '0';
      FOR k IN 1 TO 11 LOOP
        exponentff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 52 LOOP
        mantissaff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF (enable = '1') THEN
          
        signff <= NOT(signin);
        exponentff <= exponentin;
        mantissaff <= mantissain;
        
      END IF;
    
    END IF;  
      
  END PROCESS;

  expzerochk(1) <= exponentff(1);
  expmaxchk(1) <= exponentff(1);
  gxa: FOR k IN 2 TO 11 GENERATE
    expzerochk(k) <= expzerochk(k-1) OR exponentff(k);
    expmaxchk(k) <= expmaxchk(k-1) AND exponentff(k);
  END GENERATE;
  expzero <= NOT(expzerochk(11));
  expmax <= expmaxchk(11);
  
  manzerochk(1) <= mantissaff(1);
  gma: FOR k IN 2 TO 52 GENERATE
    manzerochk(k) <= manzerochk(k-1) OR mantissaff(k);
  END GENERATE;
  manzero <= NOT(manzerochk(52));
  mannonzero <= manzerochk(52);
  
  signout <= signff;
  exponentout <= exponentff;
  mantissaout <= mantissaff;
  satout <= expmax AND manzero;
  zeroout <= expzero;
  nanout <= expmax AND mannonzero;

END rtl;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   DOUBLE PRECISION MULTIPLIER - CORE LEVEL  ***
--***                                             ***
--***   DP_POS.VHD                                ***
--***                                             ***
--***   Function: Local Count Leading Zeroes      ***
--***                                             ***
--***   14/07/07 ML                               ***
--***                                             ***
--***   (c) 2007 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_pos IS
GENERIC (start : integer := 10);
PORT (
      ingroup : IN STD_LOGIC_VECTOR (6 DOWNTO 1);
      
      position : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)   
     );
END dp_pos;

ARCHITECTURE rtl of dp_pos IS
  
BEGIN

ptab: PROCESS (ingroup)
BEGIN

  CASE ingroup IS
      
      WHEN "000000" => position <= conv_std_logic_vector(0,6);
          
      WHEN "000001" => position <= conv_std_logic_vector(start+5,6);
          
      WHEN "000010" => position <= conv_std_logic_vector(start+4,6);
      WHEN "000011" => position <= conv_std_logic_vector(start+4,6); 
          
      WHEN "000100" => position <= conv_std_logic_vector(start+3,6);
      WHEN "000101" => position <= conv_std_logic_vector(start+3,6);
      WHEN "000110" => position <= conv_std_logic_vector(start+3,6);
      WHEN "000111" => position <= conv_std_logic_vector(start+3,6);
       
      WHEN "001000" => position <= conv_std_logic_vector(start+2,6); 
      WHEN "001001" => position <= conv_std_logic_vector(start+2,6);
      WHEN "001010" => position <= conv_std_logic_vector(start+2,6);
      WHEN "001011" => position <= conv_std_logic_vector(start+2,6);
      WHEN "001100" => position <= conv_std_logic_vector(start+2,6);
      WHEN "001101" => position <= conv_std_logic_vector(start+2,6);
      WHEN "001110" => position <= conv_std_logic_vector(start+2,6);
      WHEN "001111" => position <= conv_std_logic_vector(start+2,6); 
              
      WHEN "010000" => position <= conv_std_logic_vector(start+1,6);
      WHEN "010001" => position <= conv_std_logic_vector(start+1,6);
      WHEN "010010" => position <= conv_std_logic_vector(start+1,6);
      WHEN "010011" => position <= conv_std_logic_vector(start+1,6);
      WHEN "010100" => position <= conv_std_logic_vector(start+1,6);
      WHEN "010101" => position <= conv_std_logic_vector(start+1,6);
      WHEN "010110" => position <= conv_std_logic_vector(start+1,6);
      WHEN "010111" => position <= conv_std_logic_vector(start+1,6);
      WHEN "011000" => position <= conv_std_logic_vector(start+1,6);
      WHEN "011001" => position <= conv_std_logic_vector(start+1,6);
      WHEN "011010" => position <= conv_std_logic_vector(start+1,6);
      WHEN "011011" => position <= conv_std_logic_vector(start+1,6);
      WHEN "011100" => position <= conv_std_logic_vector(start+1,6);
      WHEN "011101" => position <= conv_std_logic_vector(start+1,6);
      WHEN "011110" => position <= conv_std_logic_vector(start+1,6); 
      WHEN "011111" => position <= conv_std_logic_vector(start+1,6);  
 
      WHEN "100000" => position <= conv_std_logic_vector(start,6);
      WHEN "100001" => position <= conv_std_logic_vector(start,6);
      WHEN "100010" => position <= conv_std_logic_vector(start,6);
      WHEN "100011" => position <= conv_std_logic_vector(start,6);
      WHEN "100100" => position <= conv_std_logic_vector(start,6);
      WHEN "100101" => position <= conv_std_logic_vector(start,6);
      WHEN "100110" => position <= conv_std_logic_vector(start,6);
      WHEN "100111" => position <= conv_std_logic_vector(start,6);
      WHEN "101000" => position <= conv_std_logic_vector(start,6);
      WHEN "101001" => position <= conv_std_logic_vector(start,6);
      WHEN "101010" => position <= conv_std_logic_vector(start,6);
      WHEN "101011" => position <= conv_std_logic_vector(start,6);
      WHEN "101100" => position <= conv_std_logic_vector(start,6);
      WHEN "101101" => position <= conv_std_logic_vector(start,6);
      WHEN "101110" => position <= conv_std_logic_vector(start,6); 
      WHEN "101111" => position <= conv_std_logic_vector(start,6);      
      WHEN "110000" => position <= conv_std_logic_vector(start,6);
      WHEN "110001" => position <= conv_std_logic_vector(start,6);
      WHEN "110010" => position <= conv_std_logic_vector(start,6);
      WHEN "110011" => position <= conv_std_logic_vector(start,6);
      WHEN "110100" => position <= conv_std_logic_vector(start,6);
      WHEN "110101" => position <= conv_std_logic_vector(start,6);
      WHEN "110110" => position <= conv_std_logic_vector(start,6);
      WHEN "110111" => position <= conv_std_logic_vector(start,6);
      WHEN "111000" => position <= conv_std_logic_vector(start,6);
      WHEN "111001" => position <= conv_std_logic_vector(start,6);
      WHEN "111010" => position <= conv_std_logic_vector(start,6);
      WHEN "111011" => position <= conv_std_logic_vector(start,6);
      WHEN "111100" => position <= conv_std_logic_vector(start,6);
      WHEN "111101" => position <= conv_std_logic_vector(start,6);
      WHEN "111110" => position <= conv_std_logic_vector(start,6); 
      WHEN "111111" => position <= conv_std_logic_vector(start,6);
          
      WHEN others => position <= conv_std_logic_vector(0,6);
          
  END CASE;
               
END PROCESS;    
    
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   DP_RSFT64X6.VHD                           ***
--***                                             ***
--***   Function: Double Precision Right Shift    ***
--***   (Combinatorial)                           ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_rsft64x5 IS 
PORT (
      inbus : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
      shift : IN STD_LOGIC_VECTOR (5 DOWNTO 1);
      outbus : OUT STD_LOGIC_VECTOR (64 DOWNTO 1)
    );
END dp_rsft64x5;

ARCHITECTURE rtl OF dp_rsft64x5 IS

  signal rightone, righttwo, rightthr : STD_LOGIC_VECTOR (64 DOWNTO 1);
            
BEGIN

  gra: FOR k IN 1 TO 61 GENERATE
    rightone(k) <= (inbus(k)   AND NOT(shift(2)) AND NOT(shift(1))) OR
                   (inbus(k+1) AND NOT(shift(2)) AND     shift(1)) OR
                   (inbus(k+2) AND     shift(2)  AND NOT(shift(1))) OR
                   (inbus(k+3) AND     shift(2)  AND     shift(1));
  END GENERATE;
  rightone(62) <= (inbus(62) AND NOT(shift(2)) AND NOT(shift(1))) OR
                  (inbus(63) AND NOT(shift(2)) AND     shift(1)) OR
                  (inbus(64) AND     shift(2)  AND NOT(shift(1))); 
  rightone(63) <= (inbus(63) AND NOT(shift(2)) AND NOT(shift(1))) OR
                  (inbus(64) AND NOT(shift(2)) AND     shift(1));
  rightone(64) <=  inbus(64) AND NOT(shift(2)) AND NOT(shift(1));
  
  grb: FOR k IN 1 TO 52 GENERATE
    righttwo(k) <= (rightone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                   (rightone(k+4)  AND NOT(shift(4)) AND     shift(3)) OR
                   (rightone(k+8)  AND     shift(4)  AND NOT(shift(3))) OR
                   (rightone(k+12) AND     shift(4)  AND     shift(3)); 
  END GENERATE;
  grc: FOR k IN 53 TO 56 GENERATE
    righttwo(k) <= (rightone(k)   AND NOT(shift(4)) AND NOT(shift(3))) OR
                   (rightone(k+4) AND NOT(shift(4)) AND     shift(3)) OR
                   (rightone(k+8) AND     shift(4)  AND NOT(shift(3))); 
  END GENERATE; 
  grd: FOR k IN 57 TO 60 GENERATE
    righttwo(k) <= (rightone(k)   AND NOT(shift(4)) AND NOT(shift(3))) OR
                   (rightone(k+4) AND NOT(shift(4)) AND     shift(3));
  END GENERATE; 
  gre: FOR k IN 61 TO 64 GENERATE
    righttwo(k) <= (rightone(k)   AND NOT(shift(4)) AND NOT(shift(3)));
  END GENERATE;  
  
  grf: FOR k IN 1 TO 48 GENERATE
    rightthr(k) <= (righttwo(k)    AND NOT(shift(5))) OR 
                   (righttwo(k+16) AND shift(5));
  END GENERATE;
  grg: FOR k IN 49 TO 64 GENERATE
    rightthr(k) <= (righttwo(k)    AND NOT(shift(5)));
  END GENERATE;
  
  outbus <= rightthr;        
            
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   DP_LSFT64X6.VHD                           ***
--***                                             ***
--***   Function: Double Precision Left Shift     ***
--***   (Combinatorial)                           ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_rsft64x5pipe IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      inbus : IN STD_LOGIC_VECTOR (64 DOWNTO 1);
      shift : IN STD_LOGIC_VECTOR (5 DOWNTO 1);
      outbus : OUT STD_LOGIC_VECTOR (64 DOWNTO 1)
    );
END dp_rsft64x5pipe;

ARCHITECTURE rtl OF dp_rsft64x5pipe IS

  signal rightone, righttwo, rightthr : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal righttwoff : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal shiftff : STD_LOGIC;
            
BEGIN

  gra: FOR k IN 1 TO 61 GENERATE
    rightone(k) <= (inbus(k)   AND NOT(shift(2)) AND NOT(shift(1))) OR
                   (inbus(k+1) AND NOT(shift(2)) AND     shift(1)) OR
                   (inbus(k+2) AND     shift(2)  AND NOT(shift(1))) OR
                   (inbus(k+3) AND     shift(2)  AND     shift(1));
  END GENERATE;
  rightone(62) <= (inbus(62) AND NOT(shift(2)) AND NOT(shift(1))) OR
                  (inbus(63) AND NOT(shift(2)) AND     shift(1)) OR
                  (inbus(64) AND     shift(2)  AND NOT(shift(1))); 
  rightone(63) <= (inbus(63) AND NOT(shift(2)) AND NOT(shift(1))) OR
                  (inbus(64) AND NOT(shift(2)) AND     shift(1));
  rightone(64) <=  inbus(64) AND NOT(shift(2)) AND NOT(shift(1));
  
  grb: FOR k IN 1 TO 52 GENERATE
    righttwo(k) <= (rightone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                   (rightone(k+4)  AND NOT(shift(4)) AND     shift(3)) OR
                   (rightone(k+8)  AND     shift(4)  AND NOT(shift(3))) OR
                   (rightone(k+12) AND     shift(4)  AND     shift(3)); 
  END GENERATE;
  grc: FOR k IN 53 TO 56 GENERATE
    righttwo(k) <= (rightone(k)   AND NOT(shift(4)) AND NOT(shift(3))) OR
                   (rightone(k+4) AND NOT(shift(4)) AND     shift(3)) OR
                   (rightone(k+8) AND     shift(4)  AND NOT(shift(3))); 
  END GENERATE; 
  grd: FOR k IN 57 TO 60 GENERATE
    righttwo(k) <= (rightone(k)   AND NOT(shift(4)) AND NOT(shift(3))) OR
                   (rightone(k+4) AND NOT(shift(4)) AND     shift(3));
  END GENERATE; 
  gre: FOR k IN 61 TO 64 GENERATE
    righttwo(k) <= (rightone(k)   AND NOT(shift(4)) AND NOT(shift(3)));
  END GENERATE;  
  
  ppa: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN
        
      FOR k IN 1 TO 64 LOOP
        righttwoff(k) <= '0';
      END LOOP;
      shiftff <= '0';
      
    ELSIF (rising_edge(sysclk)) THEN
    
      righttwoff <= righttwo;
      shiftff <= shift(5);
              
    END IF;
      
  END PROCESS;
  
  grf: FOR k IN 1 TO 48 GENERATE
    rightthr(k) <= (righttwoff(k)    AND NOT(shiftff)) OR 
                   (righttwoff(k+16) AND     shiftff);
  END GENERATE;
  grg: FOR k IN 49 TO 64 GENERATE
    rightthr(k) <= (righttwoff(k)    AND NOT(shiftff));
  END GENERATE;
  
  outbus <= rightthr;        
            
END rtl;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOAT CONVERT - CORE LEVEL                ***
--***                                             ***
--***   DP_RSFT64X64.VHD                          ***
--***                                             ***
--***   Function: Combinatorial Right Shift       ***
--***             (max 64.0 to 1.52)              ***
--***                                             ***
--***   07/12/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***   29/07/09 - signed number problem fixed    ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_rsft64x64 IS
PORT (
      inbus : IN STD_LOGIC_VECTOR (116 DOWNTO 1);
      shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);      
        
      outbus : OUT STD_LOGIC_VECTOR (116 DOWNTO 1)    
     );
END dp_rsft64x64;

ARCHITECTURE rtl of dp_rsft64x64 IS

  signal levzip, levone, levtwo, levthr : STD_LOGIC_VECTOR (116 DOWNTO 1);
 
BEGIN
  
  levzip <= inbus;
  
  -- unsigned input
  
  gla: FOR k IN 1 TO 113 GENERATE
    levone(k) <= (levzip(k)   AND NOT(shift(2)) AND NOT(shift(1))) OR 
                 (levzip(k+1) AND NOT(shift(2)) AND     shift(1)) OR
                 (levzip(k+2) AND     shift(2)  AND NOT(shift(1))) OR
                 (levzip(k+3) AND     shift(2)  AND     shift(1));
  END GENERATE;
  -- 29/07/65 always shift 116, else will fill with zeros
  -- fixed here and other lines
  levone(114) <= (levzip(114) AND NOT(shift(2)) AND NOT(shift(1))) OR 
                 (levzip(115) AND NOT(shift(2)) AND     shift(1)) OR
                 (levzip(116) AND     shift(2)  AND NOT(shift(1))) OR
                 (levzip(116) AND     shift(2)  AND     shift(1));
  levone(115) <= (levzip(115) AND NOT(shift(2)) AND NOT(shift(1))) OR 
                 (levzip(116) AND NOT(shift(2)) AND     shift(1)) OR 
                 (levzip(116) AND     shift(2)  AND NOT(shift(1))) OR 
                 (levzip(116) AND     shift(2)  AND     shift(1));                
  levone(116) <= levzip(116);
                               
  glba: FOR k IN 1 TO 104 GENERATE
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR 
                 (levone(k+4)  AND NOT(shift(4)) AND     shift(3)) OR
                 (levone(k+8)  AND     shift(4)  AND NOT(shift(3))) OR
                 (levone(k+12) AND     shift(4)  AND     shift(3));
  END GENERATE;  
  glbb: FOR k IN 105 TO 108 GENERATE            
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR 
                 (levone(k+4)  AND NOT(shift(4)) AND     shift(3)) OR
                 (levone(k+8)  AND     shift(4)  AND NOT(shift(3))) OR
                 (levone(116)  AND     shift(4)  AND     shift(3));             
  END GENERATE;
  glbc: FOR k IN 109 TO 112 GENERATE            
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR 
                 (levone(k+4)  AND NOT(shift(4)) AND     shift(3)) OR
                 (levone(116)  AND     shift(4)  AND NOT(shift(3))) OR
                 (levone(116)  AND     shift(4)  AND     shift(3));           
  END GENERATE;  
  glbd: FOR k IN 113 TO 116 GENERATE            
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
				 (levone(116)  AND (shift(4) OR shift(3)));
  END GENERATE;    

  glca: FOR k IN 1 TO 66 GENERATE
    levthr(k) <= (levtwo(k)    AND NOT(shift(6)) AND NOT(shift(5))) OR 
                 (levtwo(k+16) AND NOT(shift(6)) AND     shift(5)) OR
                 (levtwo(k+32) AND     shift(6)  AND NOT(shift(5))) OR
                 (levtwo(k+48) AND     shift(6)  AND     shift(5));
  END GENERATE;  
  glcb: FOR k IN 67 TO 84 GENERATE
    levthr(k) <= (levtwo(k)    AND NOT(shift(6)) AND NOT(shift(5))) OR 
                 (levtwo(k+16) AND NOT(shift(6)) AND     shift(5)) OR
                 (levtwo(k+32) AND     shift(6)  AND NOT(shift(5))) OR
                 (levtwo(116)  AND     shift(6)  AND     shift(5));
  END GENERATE; 
  glcc: FOR k IN 85 TO 100 GENERATE
    levthr(k) <= (levtwo(k)    AND NOT(shift(6)) AND NOT(shift(5))) OR 
                 (levtwo(k+16) AND NOT(shift(6)) AND     shift(5)) OR
                 (levtwo(116)  AND     shift(6)  AND NOT(shift(5))) OR
                 (levtwo(116)  AND     shift(6)  AND     shift(5));
  END GENERATE; 
  glcd: FOR k IN 101 TO 116 GENERATE
    levthr(k) <= (levtwo(k)    AND NOT(shift(6)) AND NOT(shift(5))) OR
	             (levtwo(116)  AND (shift(6) OR shift(5)));
  END GENERATE; 
      
  outbus <= levthr;
  
END rtl;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOAT CONVERT - CORE LEVEL                ***
--***                                             ***
--***   DP_RSFTPIPE64X64.VHD                      ***
--***                                             ***
--***   Function: Pipelined Right Shift           ***
--***             (max 64.0 to 1.52)              ***
--***                                             ***
--***   07/12/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***   29/07/09 - signed number problem fixed    ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_rsftpipe64x64 IS
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      inbus : IN STD_LOGIC_VECTOR (116 DOWNTO 1);
      shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);      
        
      outbus : OUT STD_LOGIC_VECTOR (116 DOWNTO 1)    
     );
END dp_rsftpipe64x64;

ARCHITECTURE rtl of dp_rsftpipe64x64 IS

  signal levzip, levone, levtwo, levthr : STD_LOGIC_VECTOR (116 DOWNTO 1);
  signal levtwoff : STD_LOGIC_VECTOR (116 DOWNTO 1);
  signal shiftff : STD_LOGIC_VECTOR (6 DOWNTO 5);
 
BEGIN
  
  levzip <= inbus;
  
  -- unsigned input
  
  gla: FOR k IN 1 TO 113 GENERATE
    levone(k) <= (levzip(k)   AND NOT(shift(2)) AND NOT(shift(1))) OR 
                 (levzip(k+1) AND NOT(shift(2)) AND     shift(1)) OR
                 (levzip(k+2) AND     shift(2)  AND NOT(shift(1))) OR
                 (levzip(k+3) AND     shift(2)  AND     shift(1));
  END GENERATE;
  -- 29/07/65 always shift 116, else will fill with zeros
  -- fixed here and other lines
  levone(114) <= (levzip(114) AND NOT(shift(2)) AND NOT(shift(1))) OR 
                 (levzip(115) AND NOT(shift(2)) AND     shift(1)) OR
                 (levzip(116) AND     shift(2)  AND NOT(shift(1))) OR
                 (levzip(116) AND     shift(2)  AND     shift(1));
  levone(115) <= (levzip(115) AND NOT(shift(2)) AND NOT(shift(1))) OR 
                 (levzip(116) AND NOT(shift(2)) AND     shift(1)) OR 
                 (levzip(116) AND     shift(2)  AND NOT(shift(1))) OR 
                 (levzip(116) AND     shift(2)  AND     shift(1));                
  levone(116) <= levzip(116);
                               
  glba: FOR k IN 1 TO 104 GENERATE
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR 
                 (levone(k+4)  AND NOT(shift(4)) AND     shift(3)) OR
                 (levone(k+8)  AND     shift(4)  AND NOT(shift(3))) OR
                 (levone(k+12) AND     shift(4)  AND     shift(3));
  END GENERATE;  
  glbb: FOR k IN 105 TO 108 GENERATE            
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR 
                 (levone(k+4)  AND NOT(shift(4)) AND     shift(3)) OR
                 (levone(k+8)  AND     shift(4)  AND NOT(shift(3))) OR
                 (levone(116)  AND     shift(4)  AND     shift(3));             
  END GENERATE;
  glbc: FOR k IN 109 TO 112 GENERATE            
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR 
                 (levone(k+4)  AND NOT(shift(4)) AND     shift(3)) OR
                 (levone(116)  AND     shift(4)  AND NOT(shift(3))) OR
                 (levone(116)  AND     shift(4)  AND     shift(3));           
  END GENERATE;  
  glbd: FOR k IN 113 TO 116 GENERATE            
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
				 (levone(116)  AND (shift(4) OR shift(3)));
  END GENERATE; 
   
  pp: PROCESS (sysclk,reset)
  BEGIN
    
    IF (reset = '1') THEN
        
      FOR k IN 1 TO 116 LOOP
        levtwoff(k) <= '0';
      END LOOP;
      shiftff <= "00";
      
    ELSIF (rising_edge(sysclk)) THEN
        
      IF (enable = '1') THEN
          
        levtwoff <= levtwo;
        shiftff <= shift(6 DOWNTO 5);
        
      END IF;
  
    END IF;
    
  END PROCESS;

  glca: FOR k IN 1 TO 66 GENERATE
    levthr(k) <= (levtwoff(k)    AND NOT(shiftff(6)) AND NOT(shiftff(5))) OR 
                 (levtwoff(k+16) AND NOT(shiftff(6)) AND     shiftff(5)) OR
                 (levtwoff(k+32) AND     shiftff(6)  AND NOT(shiftff(5))) OR
                 (levtwoff(k+48) AND     shiftff(6)  AND     shiftff(5));
  END GENERATE;  
  glcb: FOR k IN 67 TO 84 GENERATE
    levthr(k) <= (levtwoff(k)    AND NOT(shiftff(6)) AND NOT(shift(5))) OR 
                 (levtwoff(k+16) AND NOT(shiftff(6)) AND     shift(5)) OR
                 (levtwoff(k+32) AND     shiftff(6)  AND NOT(shift(5))) OR
                 (levtwoff(116)  AND     shiftff(6)  AND     shift(5));
  END GENERATE; 
  glcc: FOR k IN 85 TO 100 GENERATE
    levthr(k) <= (levtwoff(k)    AND NOT(shiftff(6)) AND NOT(shiftff(5))) OR 
                 (levtwoff(k+16) AND NOT(shiftff(6)) AND     shiftff(5)) OR
                 (levtwoff(116)  AND     shiftff(6)  AND NOT(shiftff(5))) OR
                 (levtwoff(116)  AND     shiftff(6)  AND     shiftff(5));
  END GENERATE; 
  glcd: FOR k IN 101 TO 116 GENERATE
    levthr(k) <= (levtwoff(k)    AND NOT(shiftff(6)) AND NOT(shiftff(5))) OR
	             (levtwoff(116)  AND (shiftff(6) OR shiftff(5)));
  END GENERATE; 
      
  outbus <= levthr;
  
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   DOUBLE PRECISION SQUARE ROOT - TOP LEVEL  ***
--***                                             ***
--***   DP_SQR.VHD                                ***
--***                                             ***
--***   Function: IEEE754 DP Square Root          ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** Latency = 57                                ***
--*** Based on FPROOT1.VHD (12/06)                ***
--***************************************************

ENTITY dp_sqr IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (52 DOWNTO 1);

		  signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1);
      --------------------------------------------------
      nanout : OUT STD_LOGIC;
      invalidout : OUT STD_LOGIC
		);
END dp_sqr;

ARCHITECTURE rtl OF dp_sqr IS
  
  constant manwidth : positive := 52;
  constant expwidth : positive := 11;
  
  type expfftype IS ARRAY (manwidth+4 DOWNTO 1) OF STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  
  signal signinff : STD_LOGIC;
  signal maninff : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal expinff : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal signff : STD_LOGIC_VECTOR (manwidth+4 DOWNTO 1);
  signal expnode, expdiv : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal expff : expfftype;
  signal radicand : STD_LOGIC_VECTOR (manwidth+3 DOWNTO 1);
  signal squareroot : STD_LOGIC_VECTOR (manwidth+2 DOWNTO 1);
  signal roundff, manff : STD_LOGIC_VECTOR (manwidth DOWNTO 1); 
  signal roundbit : STD_LOGIC;
  signal preadjust : STD_LOGIC;
  signal zerovec : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal offset : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
    
  -- conditions
  signal nanmanff, nanexpff : STD_LOGIC_VECTOR (manwidth+4 DOWNTO 1);
  signal zeroexpff, zeromanff : STD_LOGIC_VECTOR (manwidth+3 DOWNTO 1); 
  signal expinzero, expinmax : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal maninzero : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal expzero, expmax, manzero : STD_LOGIC;
  signal infinitycondition, nancondition : STD_LOGIC;

  component fp_sqrroot IS 
  GENERIC (width : positive := 52);
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        rad : IN STD_LOGIC_VECTOR (width+1 DOWNTO 1);

		  root : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
		  );
	end component;
		
BEGIN
    
  gzva: FOR k IN 1 TO manwidth GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  gxoa: FOR k IN 1 TO expwidth-1 GENERATE
    offset(k) <= '1';
  END GENERATE;
  offset(expwidth) <= '0';

  pma: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
      
      signinff <= '0';
      FOR k IN 1 TO manwidth LOOP
        maninff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        expinff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO manwidth+4 LOOP
        signff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO manwidth+4 LOOP
        FOR j IN 1 TO expwidth LOOP
          expff(k)(j) <= '0';
        END LOOP;
      END LOOP;
      FOR k IN 1 TO manwidth LOOP
        roundff(k) <= '0';
        manff(k) <= '0';
      END LOOP;
  
    ELSIF (rising_edge(sysclk)) THEN

      signinff <= signin;
      maninff <= mantissain;
      expinff <= exponentin;
    
      signff(1) <= signinff;
      FOR k IN 2 TO manwidth+4 LOOP
        signff(k) <= signff(k-1);
      END LOOP;
      
      expff(1)(expwidth DOWNTO 1) <= expdiv;
      expff(2)(expwidth DOWNTO 1) <= expff(1)(expwidth DOWNTO 1) + offset;
      FOR k IN 3 TO manwidth+3 LOOP
        expff(k)(expwidth DOWNTO 1) <= expff(k-1)(expwidth DOWNTO 1);
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        expff(manwidth+4)(k) <= (expff(manwidth+3)(k) AND zeroexpff(manwidth+3)) OR nanexpff(manwidth+3);
      END LOOP;
    
      roundff <= squareroot(manwidth+1 DOWNTO 2) + (zerovec(manwidth-1 DOWNTO 1) & roundbit);
    
      FOR k IN 1 TO manwidth LOOP
        manff(k) <= (roundff(k) AND zeromanff(manwidth+3)) OR nanmanff(manwidth+3);
      END LOOP;
  
    END IF;
  
  END PROCESS;

--*******************
--*** CONDITIONS ***
--*******************

  pcc: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
      
      FOR k IN 1 TO manwidth+4 LOOP
        nanmanff(k) <= '0';
        nanexpff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO manwidth+3 LOOP
        zeroexpff(k) <= '0';
        zeromanff(k) <= '0';
      END LOOP;
    
    ELSIF (rising_edge(sysclk)) THEN
      
      nanmanff(1) <= nancondition; -- level 1
      nanexpff(1) <= nancondition OR infinitycondition; -- also max exp when infinity
      FOR k IN 2 TO manwidth+4 LOOP
        nanmanff(k) <= nanmanff(k-1);
        nanexpff(k) <= nanexpff(k-1);
      END LOOP;

      zeromanff(1) <= expzero AND NOT(infinitycondition); -- level 1
      zeroexpff(1) <= expzero; -- level 1
      FOR k IN 2 TO manwidth+3 LOOP
        zeromanff(k) <= zeromanff(k-1);
        zeroexpff(k) <= zeroexpff(k-1);
      END LOOP;
    
    END IF;
  
  END PROCESS;

--*******************
--*** SQUARE ROOT ***
--*******************

  -- if exponent is odd, double mantissa and adjust exponent
  -- core latency manwidth+2 = 54
  -- top latency = core + 1 (input) + 2 (output) = 57
  sqr: fp_sqrroot 
  GENERIC MAP (width=>manwidth+2)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            rad=>radicand,
            root=>squareroot);

  radicand(1) <= '0';
  radicand(2) <= maninff(1) AND NOT(preadjust);
  gra: FOR k IN 3 TO manwidth+1 GENERATE
    radicand(k) <= (maninff(k-1) AND NOT(preadjust)) OR (maninff(k-2) AND preadjust);
  END GENERATE; 
  radicand(manwidth+2) <= NOT(preadjust) OR (maninff(manwidth) AND preadjust);
  radicand(manwidth+3) <= preadjust;   

--****************
--*** EXPONENT ***
--****************

  -- subtract 1023, divide result/2, if odd - preadjust
  -- if zero input, zero exponent and mantissa
  expnode <= expinff - offset;

  preadjust <= expnode(1);

  expdiv <= expnode(expwidth) & expnode(expwidth DOWNTO 2);

--*************
--*** ROUND ***
--*************

  -- only need to round up, round to nearest not possible out of root
  roundbit <= squareroot(1);

--*********************
--*** SPECIAL CASES ***
--*********************
-- 1. if negative input, invalid operation, NAN  (unless -0)
-- 2. -0 in -0 out
-- 3. infinity in, invalid operation, infinity out
-- 4. NAN in, invalid operation, NAN

  -- '0' if 0 
  expinzero(1) <= expinff(1);
  gxza: FOR k IN 2 TO expwidth GENERATE
    expinzero(k) <= expinzero(k-1) OR expinff(k);
  END GENERATE;
  expzero <= expinzero(expwidth); -- '0' when zero
                 
  -- '1' if nan or infinity
  expinmax(1) <= expinff(1);
  gxia: FOR k IN 2 TO expwidth GENERATE
    expinmax(k) <= expinmax(k-1) AND expinff(k);
  END GENERATE;
  expmax <= expinmax(expwidth); -- '1' when true
          
  -- '1' if not zero or infinity
  maninzero(1) <= maninff(1);
  gmza: FOR k IN 2 TO manwidth GENERATE
    maninzero(k) <= maninzero(k-1) OR maninff(k);
  END GENERATE;
  manzero <= maninzero(manwidth); 
    
  infinitycondition <= NOT(manzero) AND expmax; 

  nancondition <= (signinff AND expzero) OR (expmax AND manzero);
                
--***************
--*** OUTPUTS ***
--***************

  signout <= signff(manwidth+4);
  exponentout <= expff(manwidth+4)(expwidth DOWNTO 1);   
  mantissaout <= manff;
  -----------------------------------------------
  nanout <= nanmanff(manwidth+4);
  invalidout <= nanmanff(manwidth+4);

END rtl;



LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   DOUBLE PRECISION CORE LIBRARY             ***
--***                                             ***
--***   DP_SUBB.VHD                               ***
--***                                             ***
--***   Function: Behavioral Fixed Point Subtract ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_subb IS 
GENERIC (
         width : positive := 64;
         pipes : positive := 1
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      borrowin : IN STD_LOGIC;
      
      cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
     );
END dp_subb;

ARCHITECTURE rtl OF dp_subb IS

  type pipefftype IS ARRAY (pipes DOWNTO 1) OF STD_LOGIC_VECTOR (width DOWNTO 1);
  
  signal bbinv : STD_LOGIC_VECTOR (width DOWNTO 1);
  signal delff : STD_LOGIC_VECTOR (width DOWNTO 1);
  signal pipeff : pipefftype;
  signal ccnode : STD_LOGIC_VECTOR (width DOWNTO 1);
  signal zerovec : STD_LOGIC_VECTOR (width-1 DOWNTO 1);
    
BEGIN
  
  gza: FOR k IN 1 TO width-1 GENERATE
    zerovec(k) <= '0';
  END GENERATE;

  gia: FOR k IN 1 TO width GENERATE
    bbinv(k) <= NOT(bb(k));
  END GENERATE;
  
  -- lpm_add_sub subs 1's complement of bb
  ccnode <= aa + bbinv + (zerovec & borrowin);
  
  gda: IF (pipes = 1) GENERATE
  
    pda: PROCESS (sysclk,reset)
    BEGIN

      IF (reset = '1') THEN
    
        FOR k IN 1 TO width LOOP
          delff(k) <= '0';
        END LOOP;
     
      ELSIF (rising_edge(sysclk)) THEN

        IF (enable = '1') THEN   
          delff <= ccnode;
        END IF;

      END IF;

    END PROCESS;
    
    cc <= delff;
    
  END GENERATE;
  
  gpa: IF (pipes > 1) GENERATE
  
    ppa: PROCESS (sysclk,reset)
    BEGIN

      IF (reset = '1') THEN
        
        FOR k IN 1 TO pipes LOOP 
          FOR j IN 1 TO width LOOP
            pipeff(k)(j) <= '0';
          END LOOP;
        END LOOP;
   
      ELSIF (rising_edge(sysclk)) THEN

        IF (enable = '1') THEN   
          pipeff(1)(width DOWNTO 1) <= ccnode;
          FOR k IN 2 TO pipes LOOP
            pipeff(k)(width DOWNTO 1) <= pipeff(k-1)(width DOWNTO 1);
          END LOOP;
        END IF;

      END IF;

    END PROCESS;

    cc <= pipeff(pipes)(width DOWNTO 1);
          
  END GENERATE;
       
END rtl;


LIBRARY ieee;
LIBRARY work;
LIBRARY lpm;
USE lpm.all;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   DOUBLE PRECISION CORE LIBRARY             ***
--***                                             ***
--***   DP_ADDS.VHD                               ***
--***                                             ***
--***   Function: Synthesizable Fixed Point       ***
--***   Subtractor                                ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY dp_subs IS
GENERIC (
         width : positive := 64;
         pipes : positive := 1
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      borrowin : IN STD_LOGIC;
      
      cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
     );
END dp_subs;

ARCHITECTURE syn of dp_subs IS

  component lpm_add_sub
  GENERIC (
		     lpm_direction		: STRING;
		     lpm_hint		: STRING;
		     lpm_pipeline		: NATURAL;
		     lpm_type		: STRING;
		     lpm_width		: NATURAL
	       );
	PORT (
			dataa	: IN STD_LOGIC_VECTOR (lpm_width-1 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (lpm_width-1 DOWNTO 0);
			cin	: IN STD_LOGIC ;
			clken	: IN STD_LOGIC ;
			aclr	: IN STD_LOGIC ;
			clock	: IN STD_LOGIC ;
			result	: OUT STD_LOGIC_VECTOR (lpm_width-1 DOWNTO 0)
	     );
  end component;

BEGIN
  
  addtwo: lpm_add_sub
  GENERIC MAP (
		       lpm_direction => "SUB",
		       lpm_hint => "ONE_INPUT_IS_CONSTANT=NO,CIN_USED=YES",
		       lpm_pipeline => pipes,
		       lpm_type => "LPM_ADD_SUB",
		       lpm_width => width
	           )
  PORT MAP (
  		    dataa => aa,
		    datab => bb,
		    cin => borrowin,
		    clken => enable,
		    aclr => reset,
		    clock => sysclk,
		    result => cc
	       );  
  
END syn;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--*** Notes: Latency = 53                         ***
--***************************************************
-- input -1 to 1, output 0 to pi
ENTITY fp_acos IS 
GENERIC (synthesize : integer := 1); 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (23 DOWNTO 1);

      signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (23 DOWNTO 1)
		);
END fp_acos ;

ARCHITECTURE rtl OF fp_acos  IS

  type term_exponentfftype IS ARRAY (3 DOWNTO 1) OF STD_LOGIC_VECTOR (9 DOWNTO 1);
  type acos_sumfftype IS ARRAY (2 DOWNTO 1) OF STD_LOGIC_VECTOR (36 DOWNTO 1);
  
  signal pi : STD_LOGIC_VECTOR (36 DOWNTO 1);
  
  signal prep_signout : STD_LOGIC;
  signal numerator_exponent : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal numerator_mantissa : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal denominator_exponent : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal denominator_mantissa : STD_LOGIC_VECTOR (36 DOWNTO 1);
  
  signal signff : STD_LOGIC_VECTOR (43 DOWNTO 1);
  
  signal invsqr_exponent : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal invsqr_mantissa : STD_LOGIC_VECTOR (36 DOWNTO 1);
  
  signal del_numerator_exponent : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal del_numerator_mantissa : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal term_mantissa : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal pi_term, acos_term, acos_sum : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal acos_fixedpoint : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal term_exponentff : term_exponentfftype;

  signal acos_sumff : acos_sumfftype;
  signal acos_shift, acos_shiftff : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal shiftzeroout : STD_LOGIC;
  signal acos_mantissabus : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal acos_mantissaff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal mantissaoutff : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal zeroexponentff : STD_LOGIC;
  signal exponentadjustff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal exponentoutff : STD_LOGIC_VECTOR (8 DOWNTO 1);

  -- latency = 8
	component fp_acos_prep1
	GENERIC (synthesize : integer := 0);
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        signin : IN STD_LOGIC;
        exponentin: IN STD_LOGIC_VECTOR (8 DOWNTO 1);
        mantissain : IN STD_LOGIC_VECTOR (23 DOWNTO 1);

        signout : OUT STD_LOGIC;
		    numerator_exponent : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
		    numerator_mantissa : OUT STD_LOGIC_VECTOR (36 DOWNTO 1);
		    denominator_exponent : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
		    denominator_mantissa : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
		  );
	 end component;
	 
	-- latency = 17
	component fp_invsqr_trig1
  GENERIC (synthesize : integer := 1); 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        exponentin: IN STD_LOGIC_VECTOR (8 DOWNTO 1);
        mantissain : IN STD_LOGIC_VECTOR (36 DOWNTO 1);

        exponentout : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
        mantissaout : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
		  );
	end component;
		
	-- latency = 22
  component fp_atan_core1 IS 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        exponentin : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
        mantissain : IN STD_LOGIC_VECTOR (36 DOWNTO 1);

        atan : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
		  );
	end component;
		
  component fp_fxmul
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36;
           pipes : positive := 1;
           accuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1); 
      
        result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
       );
  end component;
  
  component fp_del 
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
   end component;	

  component fp_clz36 
  PORT (
        mantissa : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
      
        leading : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
     );
  end component;

	component fp_lsft36
  PORT (
        inbus : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);

	     outbus : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
	    );
	 end component;
	    			
BEGIN
  
  pi <= x"C90FDAA22";
  
  -- latency 8: input level 0, output level 8
  cprep: fp_acos_prep1
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            signin=>signin,exponentin=>exponentin,mantissain=>mantissain,
            signout=>prep_signout,
            numerator_exponent=>numerator_exponent,
            numerator_mantissa=>numerator_mantissa,
            denominator_exponent=>denominator_exponent,
            denominator_mantissa=>denominator_mantissa);
  
  -- latency 17: input level 8, output level 25 
  cisqr: fp_invsqr_trig1
  GENERIC MAP (synthesize=>0)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            exponentin=>denominator_exponent,
            mantissain=>denominator_mantissa,
            exponentout=>invsqr_exponent,
            mantissaout=>invsqr_mantissa);

  -- input level 8, output level 25
  cdnx: fp_del 
  GENERIC MAP (width=>8,pipes=>17)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>numerator_exponent,
            cc=>del_numerator_exponent);
  -- input level 8, output level 25                       
  cdnm: fp_del 
  GENERIC MAP (width=>36,pipes=>17)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>numerator_mantissa,
            cc=>del_numerator_mantissa);
  
  -- input level 25, output level 28
  cma: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>36,widthcc=>36,pipes=>3,
               synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>del_numerator_mantissa,
            databb=>invsqr_mantissa,
            result=>term_mantissa);
            
  pxa: PROCESS (sysclk,reset)
  BEGIN
    
    IF (reset = '1') THEN
      FOR k IN 1 TO 3 LOOP
        FOR j IN 1 TO 9 LOOP
          term_exponentff(1)(k) <= '0';
          term_exponentff(2)(k) <= '0';
          term_exponentff(3)(k) <= '0';
        END LOOP;
      END LOOP;
    ELSIF (rising_edge(sysclk)) THEN
      IF (enable = '1') THEN
        term_exponentff(1)(9 DOWNTO 1) <= ('0' & del_numerator_exponent) + ('0' & invsqr_exponent) - 126;
        term_exponentff(2)(9 DOWNTO 1) <= term_exponentff(1)(9 DOWNTO 1);
        term_exponentff(3)(9 DOWNTO 1) <= term_exponentff(2)(9 DOWNTO 1);
      END IF;
    END IF;
    
  END PROCESS;

  -- input level 28, output level 49
  cat: fp_atan_core1
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            exponentin=>term_exponentff(3)(8 DOWNTO 1),
            mantissain=>term_mantissa,
            atan=>acos_fixedpoint);
  
  gpa: FOR k IN 1 TO 36 GENERATE
    pi_term(k) <= pi(k) AND signff(41);
    acos_term(k) <= acos_fixedpoint(k) XOR signff(41);
  END GENERATE;
  acos_sum <= pi_term + acos_term + signff(41);
  
  poa: PROCESS (sysclk,reset)
  BEGIN
    
    IF (reset = '1') THEN
      
      FOR k IN 1 TO 43 LOOP
        signff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 6 LOOP
        acos_shiftff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 36 LOOP
        acos_sumff(1)(k) <= '0';
        acos_sumff(2)(k) <= '0';
        acos_mantissaff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 23 LOOP
        mantissaoutff(k) <= '0';
      END LOOP;
      zeroexponentff <= '0';
      FOR k IN 1 TO 8 LOOP
        exponentadjustff(k) <= '0';
        exponentoutff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN
        
        signff(1) <= prep_signout;
        FOR k IN 2 TO 43 LOOP
          signff(k) <= signff(k-1);
        END LOOP;
        
        acos_sumff(1)(36 DOWNTO 1) <= acos_sum;  -- level 50
        acos_sumff(2)(36 DOWNTO 1) <= acos_sumff(1)(36 DOWNTO 1);  -- level 51

        acos_shiftff <= acos_shift;  -- level 51
        
        acos_mantissaff <= acos_mantissabus;  -- level 52
        -- check for overflow not needed?
        mantissaoutff <= acos_mantissaff(35 DOWNTO 13) + acos_mantissaff(12);  -- level 52
        
        -- if CLZ output = 0 and positive input, output = 0
        zeroexponentff <= NOT(signff(43)) AND shiftzeroout;
        
        exponentadjustff <= 128 - ("00" & acos_shiftff);  -- level 52
        FOR k IN 1 TO 8 LOOP
          exponentoutff(k) <= exponentadjustff(k) AND NOT(zeroexponentff);  -- level 53
        END LOOP;
        
      END IF;
      
    END IF;
    
  END PROCESS; 
   
  czo: fp_clz36 
  PORT MAP (mantissa=>acos_sumff(1)(36 DOWNTO 1),
            leading=>acos_shift);
            
  clso: fp_lsft36
  PORT MAP (inbus=>acos_sumff(2)(36 DOWNTO 1),
            shift=>acos_shiftff,
            outbus=>acos_mantissabus);
            
  shiftzeroout <= NOT(acos_shiftff(6) OR acos_shiftff(5) OR acos_shiftff(4) OR 
                      acos_shiftff(3) OR acos_shiftff(2) OR acos_shiftff(1));
    
  --*** OUTPUTS *** 
  signout <= '0';
  exponentout <= exponentoutff;
  mantissaout <= mantissaoutff;
   
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_ACOS_PREP1.VHD                         ***
--***                                             ***
--***   Function: Single Precision Floating Point ***
--***   ACOS/ASIN Setup - generate 1-x, 1-x*x     ***
--***                                             ***
--***   23/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes: Latency = 8                          ***
--***************************************************

ENTITY fp_acos_prep1 IS 
GENERIC (synthesize : integer := 0);
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin: IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (23 DOWNTO 1);

      signout : OUT STD_LOGIC;
		  numerator_exponent : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
		  numerator_mantissa : OUT STD_LOGIC_VECTOR (36 DOWNTO 1);
		  denominator_exponent : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
		  denominator_mantissa : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
		);
END fp_acos_prep1 ;

ARCHITECTURE rtl OF fp_acos_prep1  IS

  type denominator_shiftfftype IS ARRAY (3 DOWNTO 1) OF STD_LOGIC_VECTOR (8 DOWNTO 1);
  type numerator_fixedpointfftype IS ARRAY (4 DOWNTO 1) OF STD_LOGIC_VECTOR (36 DOWNTO 1);
  type denominator_fixedpointfftype IS ARRAY (2 DOWNTO 1) OF STD_LOGIC_VECTOR (36 DOWNTO 1);
  
  signal zerovec : STD_LOGIC_VECTOR (36 DOWNTO 1);
  
  signal signff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal mantissainff : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal exponentinff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal mantissaextendff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal numerator_shiftff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal denominator_shiftff : denominator_shiftfftype;
  signal x_fixedpointff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal x_squared_fixedpointff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal numerator_fixedpointff : numerator_fixedpointfftype;
  signal denominator_fixedpointff : denominator_fixedpointfftype;
  signal numerator_leadingff, denominator_leadingff : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal numerator_mantissaff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal denominator_mantissaff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal numerator_exponentff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal denominator_exponentff : STD_LOGIC_VECTOR (8 DOWNTO 1);

  signal mantissaextend : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal x_fixedpoint : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal x_squared : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal numerator_mantissanode : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal numerator_exponentnode : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal x_squared_fixedpoint : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal denominator_mantissanode : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal denominator_exponentnode : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal numerator_leading : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal denominator_leading : STD_LOGIC_VECTOR (6 DOWNTO 1);

  component fp_fxmul
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36;
           pipes : positive := 1;
           accuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1); 
      
        result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
       );
  end component;
    
	component fp_rsft36
  PORT (
        inbus : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);

	     outbus : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
	    );
	 end component;

  component fp_clz36 
  PORT (
        mantissa : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
      
        leading : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
     );
  end component;

	component fp_lsft36
  PORT (
        inbus : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);

	     outbus : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
	    );
	 end component;
	   	 	
BEGIN
    
  gzva: FOR k IN 1 TO 36 GENERATE
    zerovec(k) <= '0';
  END GENERATE;

  pinx: PROCESS (sysclk,reset)
  BEGIN
    
    IF  (reset = '1') THEN
      
      FOR k IN 1 TO 8 LOOP
        signff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 23 LOOP
        mantissainff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 36 LOOP
        mantissaextendff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 8 LOOP
        exponentinff(k) <= '0';
        numerator_shiftff(k) <= '0';
        denominator_shiftff(1)(k) <= '0';
        denominator_shiftff(2)(k) <= '0';
        denominator_shiftff(3)(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 36 LOOP
        x_fixedpointff(k) <= '0';
        x_squared_fixedpointff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 4 LOOP
        FOR j IN 1 TO 36 LOOP
          numerator_fixedpointff(k)(j) <= '0';
        END LOOP;
      END LOOP;
      FOR k IN 1 TO 2 LOOP
        FOR j IN 1 TO 36 LOOP
          denominator_fixedpointff(k)(j) <= '0';
        END LOOP;
      END LOOP;
      FOR k IN 1 TO 6 LOOP
        numerator_leadingff(k) <= '0';
        denominator_leadingff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 36 LOOP
        numerator_mantissaff(k) <= '0';
        denominator_mantissaff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 8 LOOP
        numerator_exponentff(k) <= '0';
        denominator_exponentff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN
        
        signff(1) <= signin;
        FOR k IN 2 TO 8 LOOP
          signff(k) <= signff(k-1);
        END LOOP;
        
        mantissainff <= mantissain;  -- level 1
        exponentinff <= exponentin;  -- level 1
        
        mantissaextendff <= mantissaextend;  -- level 2
        
        numerator_shiftff <= 127 - exponentinff; -- exponent will always be 127 or less, level 2
        
        denominator_shiftff(1)(8 DOWNTO 1) <= 253 - (exponentinff(7 DOWNTO 1) & '0');  -- level 2
        denominator_shiftff(2)(8 DOWNTO 1) <= denominator_shiftff(1)(8 DOWNTO 1);  -- level 3
        denominator_shiftff(3)(8 DOWNTO 1) <= denominator_shiftff(2)(8 DOWNTO 1);  -- level 4
        
        x_fixedpointff <= x_fixedpoint;  -- level 3
        
        numerator_fixedpointff(1)(36 DOWNTO 1) <= ('1' & zerovec(35 DOWNTO 1)) - x_fixedpointff;  -- level 4
        numerator_fixedpointff(2)(36 DOWNTO 1) <= numerator_fixedpointff(1)(36 DOWNTO 1);  -- level 5
        numerator_fixedpointff(3)(36 DOWNTO 1) <= numerator_fixedpointff(2)(36 DOWNTO 1);  -- level 6
        numerator_fixedpointff(4)(36 DOWNTO 1) <= numerator_fixedpointff(3)(36 DOWNTO 1);  -- level 7
        
        x_squared_fixedpointff <= x_squared_fixedpoint; -- level 5
        
        denominator_fixedpointff(1)(36 DOWNTO 1) <= ('1' & zerovec(35 DOWNTO 1)) - x_squared_fixedpointff;  -- level 6
        denominator_fixedpointff(2)(36 DOWNTO 1) <= denominator_fixedpointff(1)(36 DOWNTO 1);  -- level 7
        
        numerator_leadingff <= numerator_leading;  -- level 7
        denominator_leadingff <= denominator_leading;  -- level 7
        
        numerator_mantissaff <= numerator_mantissanode;
        numerator_exponentff <= numerator_exponentnode;
        denominator_mantissaff <= denominator_mantissanode;
        denominator_exponentff <= denominator_exponentnode;
         
      END IF;
    
    END IF;
  
  END PROCESS;
 
  mantissaextend <= '1' & mantissainff & zerovec(12 DOWNTO 1);
  
  numsr: fp_rsft36
  PORT MAP (inbus=>mantissaextendff,shift=>numerator_shiftff(6 DOWNTO 1),
            outbus=>x_fixedpoint);
             
  mulxx: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>36,widthcc=>36,pipes=>3,
               synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>mantissaextend,databb=>mantissaextend,
            result=>x_squared);
        
  -- if x^2 <0.5, 1 bit normalization shift, output exp = 126
  densr: fp_rsft36
  PORT MAP (inbus=>x_squared,shift=>denominator_shiftff(3)(6 DOWNTO 1),
            outbus=>x_squared_fixedpoint);            

  ccznum: fp_clz36 
  PORT MAP (mantissa=>numerator_fixedpointff(3)(36 DOWNTO 1),
            leading=>numerator_leading);
            
  csftnum: fp_lsft36
  PORT MAP (inbus=>numerator_fixedpointff(4)(36 DOWNTO 1),shift=>numerator_leadingff,
            outbus=>numerator_mantissanode);
            
  numerator_exponentnode <= 127 - ("00" & numerator_leadingff); 

  cczd: fp_clz36 
  PORT MAP (mantissa=>denominator_fixedpointff(1)(36 DOWNTO 1),
            leading=>denominator_leading); 
            
  cnd: fp_lsft36
  PORT MAP (inbus=>denominator_fixedpointff(2)(36 DOWNTO 1),shift=>denominator_leadingff,
            outbus=>denominator_mantissanode);
            
  denominator_exponentnode <= 127 - ("00" & denominator_leadingff); 
  
  --*** OUTPUTS ***
  signout <= signff(8);
  numerator_mantissa <= numerator_mantissaff;
  numerator_exponent <= numerator_exponentff;
  denominator_mantissa <= denominator_mantissaff;
  denominator_exponent <= denominator_exponentff;        

END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--*** Notes: Latency = 53                         ***
--***************************************************
-- input -1 to 1, output -pi/2 to pi/2
ENTITY fp_asin IS 
GENERIC (synthesize : integer := 1); 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (23 DOWNTO 1);

      signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (23 DOWNTO 1)
		);
END fp_asin;

ARCHITECTURE rtl OF fp_asin  IS

  type term_exponentfftype IS ARRAY (3 DOWNTO 1) OF STD_LOGIC_VECTOR (9 DOWNTO 1);
  type asin_sumfftype IS ARRAY (2 DOWNTO 1) OF STD_LOGIC_VECTOR (36 DOWNTO 1);
  
  signal piovertwo : STD_LOGIC_VECTOR (36 DOWNTO 1);
  
  signal prep_signout : STD_LOGIC;
  signal numerator_exponent : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal numerator_mantissa : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal denominator_exponent : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal denominator_mantissa : STD_LOGIC_VECTOR (36 DOWNTO 1);
  
  signal signff : STD_LOGIC_VECTOR (45 DOWNTO 1);
  
  signal invsqr_exponent : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal invsqr_mantissa : STD_LOGIC_VECTOR (36 DOWNTO 1);
  
  signal del_numerator_exponent : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal del_numerator_mantissa : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal term_mantissa : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal asin_sum : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal acos_fixedpoint : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal term_exponentff : term_exponentfftype;

  signal small_mantissa : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal small_exponent : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal exponentinff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal exponentcheck : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal small_inputff : STD_LOGIC_VECTOR (50 DOWNTO 1);
      
  signal asin_sumff : asin_sumfftype;
  signal asin_shift, asin_shiftff : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal asin_mantissabus : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal asin_mantissaff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal mantissaoutff : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal exponentadjustff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal exponentadjustnode : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal exponentoutff : STD_LOGIC_VECTOR (8 DOWNTO 1);

  -- latency = 8
	component fp_acos_prep1
	GENERIC (synthesize : integer := 0);
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        signin : IN STD_LOGIC;
        exponentin: IN STD_LOGIC_VECTOR (8 DOWNTO 1);
        mantissain : IN STD_LOGIC_VECTOR (23 DOWNTO 1);

        signout : OUT STD_LOGIC;
		    numerator_exponent : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
		    numerator_mantissa : OUT STD_LOGIC_VECTOR (36 DOWNTO 1);
		    denominator_exponent : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
		    denominator_mantissa : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
		  );
	 end component;
	 
	-- latency = 17
	component fp_invsqr_trig1
  GENERIC (synthesize : integer := 1); 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        exponentin: IN STD_LOGIC_VECTOR (8 DOWNTO 1);
        mantissain : IN STD_LOGIC_VECTOR (36 DOWNTO 1);

        exponentout : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
        mantissaout : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
		  );
	end component;
		
	-- latency = 22
  component fp_atan_core1 IS 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        exponentin : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
        mantissain : IN STD_LOGIC_VECTOR (36 DOWNTO 1);

        atan : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
		  );
	end component;
		
  component fp_fxmul
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36;
           pipes : positive := 1;
           accuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1); 
      
        result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
       );
  end component;
  
  component fp_del 
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
   end component;	

  component fp_clz36 
  PORT (
        mantissa : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
      
        leading : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
     );
  end component;

	component fp_lsft36
  PORT (
        inbus : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);

	     outbus : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
	    );
	 end component;
	    			
BEGIN

  piovertwo <= x"6487ED511";
  
  -- latency 8: input level 0, output level 8
  cprep: fp_acos_prep1
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            signin=>signin,exponentin=>exponentin,mantissain=>mantissain,
            signout=>prep_signout,
            numerator_exponent=>numerator_exponent,
            numerator_mantissa=>numerator_mantissa,
            denominator_exponent=>denominator_exponent,
            denominator_mantissa=>denominator_mantissa);
  
  -- latency 17: input level 8, output level 25 
  cisqr: fp_invsqr_trig1
  GENERIC MAP (synthesize=>0)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            exponentin=>denominator_exponent,
            mantissain=>denominator_mantissa,
            exponentout=>invsqr_exponent,
            mantissaout=>invsqr_mantissa);

  -- input level 8, output level 25
  cdnx: fp_del 
  GENERIC MAP (width=>8,pipes=>17)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>numerator_exponent,
            cc=>del_numerator_exponent);
  -- input level 8, output level 25                       
  cdnm: fp_del 
  GENERIC MAP (width=>36,pipes=>17)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>numerator_mantissa,
            cc=>del_numerator_mantissa);
  
  -- input level 25, output level 28
  cma: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>36,widthcc=>36,pipes=>3,
               synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>del_numerator_mantissa,
            databb=>invsqr_mantissa,
            result=>term_mantissa);
            
  pxa: PROCESS (sysclk,reset)
  BEGIN
    
    IF (reset = '1') THEN
      FOR k IN 1 TO 3 LOOP
        FOR j IN 1 TO 9 LOOP
          term_exponentff(1)(k) <= '0';
          term_exponentff(2)(k) <= '0';
          term_exponentff(3)(k) <= '0';
        END LOOP;
      END LOOP;
    ELSIF (rising_edge(sysclk)) THEN
      IF (enable = '1') THEN
        term_exponentff(1)(9 DOWNTO 1) <= ('0' & del_numerator_exponent) + ('0' & invsqr_exponent) - 126;
        term_exponentff(2)(9 DOWNTO 1) <= term_exponentff(1)(9 DOWNTO 1);
        term_exponentff(3)(9 DOWNTO 1) <= term_exponentff(2)(9 DOWNTO 1);
      END IF;
    END IF;
    
  END PROCESS;

  -- input level 28, output level 49
  cat: fp_atan_core1
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            exponentin=>term_exponentff(3)(8 DOWNTO 1),
            mantissain=>term_mantissa,
            atan=>acos_fixedpoint);

  asin_sum <= piovertwo - acos_fixedpoint;
  
  --*** handle small inputs ****
  dsma: fp_del
  GENERIC MAP (width=>23,pipes=>51)
  PORT MAP (sysclk=>sysclk,reset=>'0',enable=>enable, -- no resets for memory
            aa=>mantissain,
            cc=>small_mantissa); 
  dsxa: fp_del
  GENERIC MAP (width=>8,pipes=>51)
  PORT MAP (sysclk=>sysclk,reset=>'0',enable=>enable, -- no resets for memory
            aa=>exponentin,
            cc=>small_exponent); 
        
  exponentcheck <= exponentinff - 115;
                
  psa: PROCESS (sysclk,reset)
  BEGIN
  
    IF (reset = '1') THEN

      exponentinff <= "00000000";
      FOR k IN 1 TO 50 LOOP
        small_inputff(k) <= '0';
      END LOOP;
    
    ELSIF(rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN

        exponentinff <= exponentin;
        small_inputff(1) <= exponentcheck(8);
        FOR k IN 2 TO 50 LOOP
          small_inputff(k) <= small_inputff(k-1);
        END LOOP;
        
      END IF;
    
    END IF;
  
  END PROCESS;
  
  poa: PROCESS (sysclk,reset)
  BEGIN
    
    IF (reset = '1') THEN
      
      FOR k IN 1 TO 45 LOOP
        signff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 6 LOOP
        asin_shiftff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 36 LOOP
        asin_sumff(1)(k) <= '0';
        asin_sumff(2)(k) <= '0';
        asin_mantissaff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 23 LOOP
        mantissaoutff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 8 LOOP
        exponentadjustff(k) <= '0';
        exponentoutff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN
        
        signff(1) <= prep_signout;
        FOR k IN 2 TO 45 LOOP
          signff(k) <= signff(k-1);
        END LOOP;
        
        asin_sumff(1)(36 DOWNTO 1) <= asin_sum;  -- level 50
        asin_sumff(2)(36 DOWNTO 1) <= asin_sumff(1)(36 DOWNTO 1);  -- level 51

        asin_shiftff <= asin_shift;  -- level 51

        FOR k IN 1 TO 12 LOOP
          asin_mantissaff(k) <= asin_mantissabus(k) AND NOT(small_inputff(50));  -- level 52
        END LOOP;
        FOR k IN 1 TO 23 LOOP
          asin_mantissaff(k+12) <= (asin_mantissabus(k+12) AND NOT(small_inputff(50))) OR
                                   (small_mantissa(k) AND small_inputff(50));
        END LOOP;
        asin_mantissaff(36) <= asin_mantissabus (36);
        
        -- check for overflow not needed?
        mantissaoutff <= asin_mantissaff(35 DOWNTO 13) + asin_mantissaff(12);  -- level 52
    
        FOR k IN 1 TO 8 LOOP
          exponentadjustff(k) <= (exponentadjustnode(k) AND NOT(small_inputff(50))) OR
                                 (small_exponent(k) AND small_inputff(50));  -- level 52
        END LOOP;
        FOR k IN 1 TO 8 LOOP
          exponentoutff(k) <= exponentadjustff(k);  -- level 53
        END LOOP;
        
      END IF;
      
    END IF;
    
  END PROCESS; 
   
  exponentadjustnode <= 128 - ("00" & asin_shiftff);
  
  czo: fp_clz36 
  PORT MAP (mantissa=>asin_sumff(1)(36 DOWNTO 1),
            leading=>asin_shift);
            
  clso: fp_lsft36
  PORT MAP (inbus=>asin_sumff(2)(36 DOWNTO 1),
            shift=>asin_shiftff,
            outbus=>asin_mantissabus);
    
  --*** OUTPUTS *** 
  signout <= signff(45);
  exponentout <= exponentoutff;
  mantissaout <= mantissaoutff;
   
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_ATAN.VHD                              ***
--***                                             ***
--***   Function: Single Precision Floating Point ***
--***   ArcTangent                                ***
--***                                             ***
--***   23/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** NOTES                                       ***
--***************************************************
-- slight improvement when "roundbit" is used i.e. round up from
-- X.4999 - exact number of bits to be used needs to be tweaked

ENTITY fp_atan IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (23 DOWNTO 1);

      signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (23 DOWNTO 1)
		);
END fp_atan;

ARCHITECTURE rtl OF fp_atan IS
  
  constant coredepth : positive := 12;
  
  constant b_precision : positive := 10;
  
  type exponentinfftype IS ARRAY (coredepth-2 DOWNTO 1) OF STD_LOGIC_VECTOR (10 DOWNTO 1);
  type exponenttopfftype IS ARRAY (coredepth-3 DOWNTO 1) OF STD_LOGIC_VECTOR (10 DOWNTO 1);
  type mantissabpfftype IS ARRAY (2*coredepth+10 DOWNTO 1) OF STD_LOGIC_VECTOR (23 DOWNTO 1); -- SPR: 380600
  type termfftype IS ARRAY (2 DOWNTO 1) OF STD_LOGIC_VECTOR (36 DOWNTO 1);
  
  signal zerovec : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal pi_over_two : STD_LOGIC_VECTOR (36 DOWNTO 1);
  
  signal inputnumber : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal delinputnumber : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal topquotient : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal topquotientnumber : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal exponentoffset : STD_LOGIC_VECTOR (10 DOWNTO 1);
  
  signal exponentinff : exponentinfftype;
  signal idselectff : STD_LOGIC_VECTOR (2*coredepth+10 DOWNTO 1); -- SPR: 380600
  signal pathselectff : STD_LOGIC_VECTOR (2*coredepth+9 DOWNTO 1);
  signal exponenttopff : exponenttopfftype;
  signal forward_shiftff, inverse_shiftff : STD_LOGIC_VECTOR (10 DOWNTO 1);
  signal a_shiftff : STD_LOGIC_VECTOR (10 DOWNTO 1);
  signal a_fixedpointff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal a_fixedpointbus : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal a_mantissanode : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal pathcheck : STD_LOGIC_VECTOR (9 DOWNTO 1);

  signal a_fixedpoint : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal b_fixedpoint : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal c_fixedpoint : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal ab_fixedpoint : STD_LOGIC_VECTOR (37 DOWNTO 1);
  signal ab_plusone : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal numerator, denominator : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal addterm : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal b_address : STD_LOGIC_VECTOR (10 DOWNTO 1);
  signal lutterm : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal dellutterm : STD_LOGIC_VECTOR (36 DOWNTO 1);
  
  signal signff : STD_LOGIC_VECTOR (2*coredepth+11 DOWNTO 1);
  signal mantissabpff : mantissabpfftype; -- SPR: 380600
  signal atantermff : termfftype;
  signal large_atanff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal small_mantissa, small_mantissaff : STD_LOGIC_VECTOR (36 DOWNTO 1); 
  signal large_mantissa, large_mantissaff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal mux_mantissa : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal small_count, small_countff : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal small_overflowbus, large_overflowbus : STD_LOGIC_VECTOR (24 DOWNTO 1);
  signal small_overflowff, large_overflowff : STD_LOGIC;
  signal mux_overflow : STD_LOGIC;
  signal roundbit : STD_LOGIC;
  signal mantissa_roundff : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal mantissa_bypass : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal exponent_outff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal small_exponent_adjust, large_exponent_adjust : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal exponent_adjust, exponent_adjustff : STD_LOGIC_VECTOR (8 DOWNTO 1);

  -- SPR: 380600
  signal expinzero : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal expzero : STD_LOGIC;
  
	component fp_inv_core
  GENERIC (synthesize : integer := 1); 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        divisor : IN STD_LOGIC_VECTOR (36 DOWNTO 1);

		    quotient : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
		    );
  end component;

	component fp_rsft36
  PORT (
        inbus : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);

	     outbus : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
	    );
	 end component;

  component fp_del 
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
   end component;	
   
  component fp_fxmul
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36;
           pipes : positive := 1;
           accuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1); 
      
        result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
       );
  end component;
  
  component fp_atanlut
  PORT (
        add : IN STD_LOGIC_VECTOR (10 DOWNTO 1);
        data : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
       );
  end component;

  component fp_clz36
  PORT (
        mantissa : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
       
        leading : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
       );
  end component;

  component fp_lsft36 IS 
  PORT (
        inbus : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);

	     outbus : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
	    );
	end component;
	       	    
BEGIN
        
  gza: FOR k IN 1 TO 36 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  pi_over_two <= x"C90FDAA22"; -- 1.57...
  
  --*** Invert Input ***
  inputnumber <= '1' & mantissain & "000000000000";

  -- will give output between 0.5 and 0.99999...
  -- will always need to be normalized
  invcore: fp_inv_core
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            divisor=>inputnumber,
            quotient=>topquotient);
      
  exponentoffset <= conv_std_logic_vector (127,10);
  
  pinx: PROCESS (sysclk,reset)
  BEGIN
    
    IF  (reset = '1') THEN
      
      FOR k IN 1 TO coredepth-2 LOOP
        FOR j IN 1 TO 8 LOOP
          exponentinff(k)(j) <= '0';
        END LOOP;
      END LOOP;
      FOR k IN 1 TO 2*coredepth+9 LOOP
        pathselectff(k) <= '0';
      END LOOP;
	  -- SPR: 380600
      FOR k IN 1 TO 2*coredepth+10 LOOP
        idselectff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO coredepth-3 LOOP
        FOR j IN 1 TO 10 LOOP
          exponenttopff(k)(j) <= '0';
        END LOOP;
      END LOOP;
      FOR k IN 1 TO 10 LOOP
        forward_shiftff(k) <= '0';
        inverse_shiftff(k) <= '0';
        a_shiftff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 36 LOOP
        a_fixedpointff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN
      
        exponentinff(1)(8 DOWNTO 1) <= exponentin;
        FOR k IN 2 TO coredepth-2 LOOP
          exponentinff(k)(8 DOWNTO 1) <= exponentinff(k-1)(8 DOWNTO 1);
        END LOOP;
        
        pathselectff(1) <= pathcheck(9);
        FOR k IN 2 TO 2*coredepth+9 LOOP
          pathselectff(k) <= pathselectff(k-1); 
        END LOOP;
		
		-- SPR: 380600
		idselectff(1) <= expzero;
        FOR k IN 2 TO 2*coredepth+10 LOOP
          idselectff(k) <= idselectff(k-1); 
        END LOOP;
        
        -- exponent for inverse, used when exponent > 126
        exponenttopff(1)(10 DOWNTO 1) <= exponentoffset - ("00" & exponentinff(1)(8 DOWNTO 1));
        exponenttopff(2)(10 DOWNTO 1) <= exponenttopff(1)(10 DOWNTO 1) + exponentoffset;
        exponenttopff(3)(10 DOWNTO 1) <= exponenttopff(2)(10 DOWNTO 1) - 1;
        -- inverse always less than 1, decrement exponent
        FOR k IN 4 TO coredepth-3 LOOP
          exponenttopff(k)(10 DOWNTO 1) <= exponenttopff(k-1)(10 DOWNTO 1);
        END LOOP;
        
        forward_shiftff <= "0001111111" - ("00" & exponentinff(coredepth-2)(8 DOWNTO 1));
        inverse_shiftff <= "0001111111" - exponenttopff(coredepth-3)(10 DOWNTO 1);
        
        FOR k IN 1 TO 6 LOOP
          a_shiftff(k) <= (forward_shiftff(k) AND NOT(pathselectff(coredepth-2))) OR 
                          (inverse_shiftff(k) AND     pathselectff(coredepth-2)); 
        END LOOP;
        
        a_fixedpointff <= a_fixedpointbus;
   
      END IF;
      
    END IF;
    
  END PROCESS;    

  -- if <=126 (<= 0.999999), use atan(x) path, else use (pi/2-atan(1/x)) path
  pathcheck <= "001111110" - ('0' & exponentinff(1)(8 DOWNTO 1));
  
  cdma: fp_del 
  GENERIC MAP (width=>36,pipes=>coredepth)  -- 12 for inv_core
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>inputnumber,
            cc=>delinputnumber);
            
  topquotientnumber <= topquotient(35 DOWNTO 1) & '0';
  gma: FOR k IN 1 TO 36 GENERATE
    a_mantissanode(k) <= (delinputnumber(k)    AND NOT(pathselectff(coredepth-1))) OR
                         (topquotientnumber(k) AND     pathselectff(coredepth-1));
  END GENERATE;

  casr: fp_rsft36
  PORT MAP (inbus=>a_mantissanode,shift=>a_shiftff(6 DOWNTO 1),
            outbus=>a_fixedpointbus);
      
  a_fixedpoint <= a_fixedpointff;    
  b_fixedpoint <= a_fixedpointff(36 DOWNTO 37-b_precision) & zerovec(36-b_precision DOWNTO 1);
  c_fixedpoint <= a_fixedpointff(36-b_precision DOWNTO 1) & zerovec(b_precision DOWNTO 1); 
  
  cmone: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>36,widthcc=>37,
               pipes=>3)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>a_fixedpoint,databb=>b_fixedpoint,
            result=>ab_fixedpoint);
            
  ab_plusone <= '1' & ab_fixedpoint(35 DOWNTO 1); -- ab_fixedpoint always 1/4 true value
            
  invtwo: fp_inv_core
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            divisor=>ab_plusone,
            quotient=>denominator);
  
  cdc: fp_del 
  GENERIC MAP (width=>36,pipes=>coredepth+3)  -- inv_core and 3 for 36*36 mult
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>c_fixedpoint,
            cc=>numerator);
                      
  cmtwo: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>36,widthcc=>36,
               pipes=>3)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>numerator,databb=>denominator,
            result=>addterm);         

  b_address <= a_fixedpoint(36 DOWNTO 37-b_precision);
 
  clut: fp_atanlut
  PORT MAP (add=>b_address,
            data=>lutterm);
            
  cdlut: fp_del 
  GENERIC MAP (width=>36,pipes=>18)  -- 12 for inv_core and 3 for 36*36 mult
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>lutterm,
            cc=>dellutterm);
  
  pimo: PROCESS (sysclk,reset)
  BEGIN
    
    IF  (reset = '1') THEN
      
      FOR k IN 1 TO 2*coredepth+11 LOOP
        signff(k) <= '0';
      END LOOP;
	  
	  -- SPR: 380600
      FOR k IN 1 TO 2*coredepth+10 LOOP
		FOR j IN 1 TO 23 LOOP
		  mantissabpff(k)(j) <= '0';
		END LOOP;
      END LOOP;
	  
      FOR k IN 1 TO 36 LOOP
        atantermff(1)(k) <= '0';
        atantermff(2)(k) <= '0';
        large_atanff(k) <= '0';
        small_mantissaff(k) <= '0';
        large_mantissaff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 6 LOOP
        small_countff(k) <= '0';
      END LOOP;
      small_overflowff <= '0';
      large_overflowff <= '0';
      FOR k IN 1 TO 23 LOOP
        mantissa_roundff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 8 LOOP
        exponent_outff(k) <= '0';
      END LOOP;

    ELSIF (rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN
      
        signff(1) <= signin;
		mantissabpff(1)(23 DOWNTO 1) <= mantissain(23 DOWNTO 1);
        FOR k IN 2 TO 2*coredepth+11 LOOP
          signff(k) <= signff(k-1);
        END LOOP;
		
		-- SPR: 380600
        FOR k IN 2 TO 2*coredepth+10 LOOP
		  mantissabpff(k)(23 DOWNTO 1) <= mantissabpff(k-1)(23 DOWNTO 1);
        END LOOP;
        
        atantermff(1)(36 DOWNTO 1) <= dellutterm + (zerovec(9 DOWNTO 1) & addterm(36 DOWNTO 10));
        atantermff(2)(36 DOWNTO 1) <= atantermff(1)(36 DOWNTO 1);
        
        -- always in the range 0.78 to pi/2
        large_atanff(36 DOWNTO 1) <= pi_over_two - atantermff(1)(36 DOWNTO 1);
            
        small_countff <= small_count;

        large_mantissaff <= large_mantissa;
        small_mantissaff <= small_mantissa;
        
        small_overflowff <= small_overflowbus(24);
        large_overflowff <= large_overflowbus(24);
        
        exponent_adjustff <= exponent_adjust;
        
        --mantissa_roundff <= mux_mantissa(35 DOWNTO 13) + mux_mantissa(12);
        mantissa_roundff <= mux_mantissa(35 DOWNTO 13) + roundbit;
        exponent_outff <= "01111111" - exponent_adjustff + mux_overflow;
        
      END IF;
      
    END IF;
    
  END PROCESS;  
  
  roundbit <= mux_mantissa(12) OR 
             (mux_mantissa(11) AND mux_mantissa(10) AND mux_mantissa(9) AND mux_mantissa(8) AND 
              mux_mantissa(7)  AND mux_mantissa(6)  AND mux_mantissa(5) AND mux_mantissa(4) AND 
              mux_mantissa(3)  AND mux_mantissa(2));

  ccsat: fp_clz36
  PORT MAP (mantissa=>atantermff(1)(36 DOWNTO 1),
            leading=>small_count);
  
  cssat: fp_lsft36
  PORT MAP (inbus=>atantermff(2)(36 DOWNTO 1),shift=>small_countff,
            outbus=>small_mantissa);
            
  small_overflowbus(1) <= small_mantissa(12);
  gova: FOR k IN 2 TO 24 GENERATE
    small_overflowbus(k) <= small_overflowbus(k-1) AND small_mantissa(k+11);
  END GENERATE;
            
  glma: FOR k IN 1 TO 35 GENERATE
    large_mantissa(k+1) <= (large_atanff(k)   AND NOT(large_atanff(36))) OR
                           (large_atanff(k+1) AND     large_atanff(36));
  END GENERATE;
  large_mantissa(1) <= '0';

  large_overflowbus(1) <= large_mantissa(12);
  govb: FOR k IN 2 TO 24 GENERATE
    large_overflowbus(k) <= large_overflowbus(k-1) AND large_mantissa(k+11);
  END GENERATE;
  
  gmma: FOR k IN 1 TO 36 GENERATE
    mux_mantissa(k) <= (small_mantissaff(k) AND NOT(pathselectff(2*coredepth+9))) OR
                       (large_mantissaff(k) AND     pathselectff(2*coredepth+9));
  END GENERATE;
  
  mux_overflow <= (small_overflowff AND NOT(pathselectff(2*coredepth+9))) OR
                  (large_overflowff AND     pathselectff(2*coredepth+9));
  
  large_exponent_adjust <= "0000000" & NOT(large_atanff(36));
  small_exponent_adjust <= "00" & small_countff;
  gxa: FOR k IN 1 TO 8 GENERATE
    exponent_adjust(k) <= (small_exponent_adjust(k) AND NOT(pathselectff(2*coredepth+8))) OR
                          (large_exponent_adjust(k) AND     pathselectff(2*coredepth+8));
  END GENERATE;
  
  -- SPR: 380600
  bypass: FOR k IN 1 TO 23 GENERATE
    mantissa_bypass(k) <= (mantissa_roundff(k) AND NOT(idselectff(2*coredepth+10))) OR
							(mantissabpff(2*coredepth+10)(k) AND idselectff(2*coredepth+10));
  END GENERATE;

  -- SPR: 380600
  expinzero(1) <= exponentinff(1)(1);
  gxza: FOR k IN 2 TO 8 GENERATE
    expinzero(k) <= expinzero(k-1) OR exponentinff(1)(k);
  END GENERATE;
  expzero <= NOT(expinzero(8)); -- '0' when zero

  --*** OUTPUTS ***
  signout <= signff(2*coredepth+11);
  exponentout <= (others => '0') when idselectff(2*coredepth+10) = '1' else exponent_outff; -- SPR: 380600
  mantissaout <= mantissa_bypass;

end rtl;

		    
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_ATAN_CORE1.VHD                         ***
--***                                             ***
--***   Function: Single Precision Floating Point ***
--***   ATAN Core for ACOS/ASIN Function          ***
--***                                             ***
--***   23/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** 1. Latency = 21                             ***
--*** 2. Valid for inputs < 1                     ***
--***************************************************

ENTITY fp_atan_core1 IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (36 DOWNTO 1);

      atan : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
		);
END fp_atan_core1;

ARCHITECTURE rtl OF fp_atan_core1 IS
  
  constant b_precision : positive := 10;
  
  signal zerovec : STD_LOGIC_VECTOR (36 DOWNTO 1);

  signal mantissainff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal exponentinff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal a_fixedpointff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal luttermff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal ab_plusoneff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal atan_sumff : STD_LOGIC_VECTOR (36 DOWNTO 1);

  signal a_shift : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal a_fixedpoint : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal b_fixedpoint : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal c_fixedpoint : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal b_address : STD_LOGIC_VECTOR (10 DOWNTO 1);
  signal lutterm : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal dellutterm : STD_LOGIC_VECTOR (36 DOWNTO 1); 
  signal ab_fixedpoint : STD_LOGIC_VECTOR (37 DOWNTO 1);
  signal numerator, denominator : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal addterm : STD_LOGIC_VECTOR (36 DOWNTO 1);
         
	component fp_inv_core
  GENERIC (synthesize : integer := 1); 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        divisor : IN STD_LOGIC_VECTOR (36 DOWNTO 1);

		    quotient : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
		    );
  end component;

	component fp_rsft36
  PORT (
        inbus : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);

	     outbus : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
	    );
	 end component;

  component fp_del 
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
   end component;	
   
  component fp_fxmul
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36;
           pipes : positive := 1;
           accuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1); 
      
        result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
       );
  end component;
  
  component fp_atanlut
  PORT (
        add : IN STD_LOGIC_VECTOR (10 DOWNTO 1);
        data : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
       );
  end component;
	    
BEGIN
        
  gza: FOR k IN 1 TO 36 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  pinx: PROCESS (sysclk,reset)
  BEGIN
    
    IF  (reset = '1') THEN

      FOR k IN 1 TO 36 LOOP
        mantissainff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 8 LOOP
        exponentinff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 36 LOOP
        a_fixedpointff(k) <= '0';
        luttermff(k) <= '0';
        ab_plusoneff(k) <= '0';
        atan_sumff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN
        
        mantissainff <= mantissain;  -- level 1
        exponentinff <= exponentin;  -- level 1
        
        a_fixedpointff <= a_fixedpoint; -- level 2
        
        luttermff <= lutterm; -- level 4
        
        ab_plusoneff <= '1' & ab_fixedpoint(35 DOWNTO 1); -- ab_fixedpoint always 1/4 true value, level 6
        
        atan_sumff <= dellutterm + (zerovec(9 DOWNTO 1) & addterm(36 DOWNTO 10));
         
      END IF;
    
    END IF;
  
  END PROCESS;
  
  a_shift <= 127 - exponentinff; -- a_exponent will always be 126 or less
  
  asr: fp_rsft36
  PORT MAP (inbus=>mantissainff,shift=>a_shift(6 DOWNTO 1),
            outbus=>a_fixedpoint);
            
  b_fixedpoint <= a_fixedpoint(36 DOWNTO 37-b_precision) & zerovec(36-b_precision DOWNTO 1);
  c_fixedpoint <= a_fixedpoint(36-b_precision DOWNTO 1) & zerovec(b_precision DOWNTO 1); 
  
  b_address <= a_fixedpointff(36 DOWNTO 37-b_precision);
 
  -- level 3
  clut: fp_atanlut
  PORT MAP (add=>b_address,
            data=>lutterm);
  
  -- level 3 in, level 20 out
  cdlut: fp_del 
  GENERIC MAP (width=>36,pipes=>17) 
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>luttermff,
            cc=>dellutterm);

  -- level 1 in, level 17 out
  cdnum: fp_del 
  GENERIC MAP (width=>36,pipes=>16)  
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>c_fixedpoint,
            cc=>numerator);
            
  -- level 2 in, level 5 out             
  cmab: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>36,widthcc=>37,
               pipes=>3,synthesize=>0)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>a_fixedpoint,databb=>b_fixedpoint,
            result=>ab_fixedpoint);
                
  -- level 5 in, level 17 out
  cinv: fp_inv_core
  GENERIC MAP (synthesize=>0) 
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            divisor=>ab_plusoneff,
            quotient=>denominator);
         
  -- level 17 in, level 20 out   
  cmo: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>36,widthcc=>36,
               pipes=>3,synthesize=>0)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>numerator,databb=>denominator,
            result=>addterm);         
            
  --*** OUTPUTS ***
  atan <= atan_sumff;

end rtl;

		    LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_ATANLUT.VHD                            ***
--***                                             ***
--***   Function: ArcTangent Look Up Table        ***
--***   (Generated by MATLAB Utility)             ***
--***                                             ***
--***   22/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_atanlut IS
PORT (
      add : IN STD_LOGIC_VECTOR (10 DOWNTO 1);
      data : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
     );
END fp_atanlut;

ARCHITECTURE rtl OF fp_atanlut IS

BEGIN

  pca: PROCESS (add)
  BEGIN
    CASE add IS
      WHEN "0000000000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(0,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(0,18);
      WHEN "0000000001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(255,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(262058,18);
      WHEN "0000000010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(511,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(261461,18);
      WHEN "0000000011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(767,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(259840,18);
      WHEN "0000000100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(1023,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(256682,18);
      WHEN "0000000101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(1279,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(251477,18);
      WHEN "0000000110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(1535,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(243713,18);
      WHEN "0000000111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(1791,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(232877,18);
      WHEN "0000001000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(2047,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(218459,18);
      WHEN "0000001001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(2303,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(199947,18);
      WHEN "0000001010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(2559,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(176830,18);
      WHEN "0000001011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(2815,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(148596,18);
      WHEN "0000001100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(3071,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(114736,18);
      WHEN "0000001101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(3327,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(74739,18);
      WHEN "0000001110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(3583,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(28094,18);
      WHEN "0000001111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(3838,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(236436,18);
      WHEN "0000010000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(4094,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(174967,18);
      WHEN "0000010001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(4350,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(105322,18);
      WHEN "0000010010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(4606,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(26992,18);
      WHEN "0000010011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(4861,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(201613,18);
      WHEN "0000010100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(5117,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(104389,18);
      WHEN "0000010101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(5372,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(259100,18);
      WHEN "0000010110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(5628,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(140951,18);
      WHEN "0000010111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(5884,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(11580,18);
      WHEN "0000011000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(6139,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(132624,18);
      WHEN "0000011001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(6394,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(241434,18);
      WHEN "0000011010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(6650,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(75361,18);
      WHEN "0000011011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(6905,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(158188,18);
      WHEN "0000011100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(7160,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(227268,18);
      WHEN "0000011101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(7416,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(19954,18);
      WHEN "0000011110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(7671,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(60030,18);
      WHEN "0000011111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(7926,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(84851,18);
      WHEN "0000100000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(8181,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(93916,18);
      WHEN "0000100001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(8436,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(86725,18);
      WHEN "0000100010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(8691,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(62776,18);
      WHEN "0000100011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(8946,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(21573,18);
      WHEN "0000100100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(9200,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(224760,18);
      WHEN "0000100101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(9455,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(147552,18);
      WHEN "0000100110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(9710,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(51596,18);
      WHEN "0000100111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(9964,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(198541,18);
      WHEN "0000101000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(10219,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(63603,18);
      WHEN "0000101001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(10473,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(170578,18);
      WHEN "0000101010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(10727,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(256827,18);
      WHEN "0000101011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(10982,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(59715,18);
      WHEN "0000101100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(11236,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(103038,18);
      WHEN "0000101101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(11490,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(124162,18);
      WHEN "0000101110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(11744,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(122599,18);
      WHEN "0000101111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(11998,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(97859,18);
      WHEN "0000110000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(12252,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(49456,18);
      WHEN "0000110001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(12505,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(239047,18);
      WHEN "0000110010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(12759,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(141859,18);
      WHEN "0000110011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(13013,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(19553,18);
      WHEN "0000110100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(13266,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(133790,18);
      WHEN "0000110101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(13519,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(221944,18);
      WHEN "0000110110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(13773,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(21390,18);
      WHEN "0000110111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(14026,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(55937,18);
      WHEN "0000111000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(14279,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(62963,18);
      WHEN "0000111001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(14532,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(41991,18);
      WHEN "0000111010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(14784,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(254689,18);
      WHEN "0000111011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(15037,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(176296,18);
      WHEN "0000111100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(15290,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(68480,18);
      WHEN "0000111101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(15542,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(192916,18);
      WHEN "0000111110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(15795,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(24844,18);
      WHEN "0000111111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(16047,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(88083,18);
      WHEN "0001000000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(16299,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(120021,18);
      WHEN "0001000001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(16551,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(120191,18);
      WHEN "0001000010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(16803,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(88130,18);
      WHEN "0001000011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(17055,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(23371,18);
      WHEN "0001000100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(17306,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(187599,18);
      WHEN "0001000101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(17558,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(56063,18);
      WHEN "0001000110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(17809,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(152592,18);
      WHEN "0001000111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(18060,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(214584,18);
      WHEN "0001001000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(18311,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(241584,18);
      WHEN "0001001001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(18562,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(233135,18);
      WHEN "0001001010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(18813,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(188785,18);
      WHEN "0001001011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(19064,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(108082,18);
      WHEN "0001001100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(19314,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(252719,18);
      WHEN "0001001101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(19565,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(97960,18);
      WHEN "0001001110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(19815,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(167646,18);
      WHEN "0001001111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(20065,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(199187,18);
      WHEN "0001010000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(20315,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(192140,18);
      WHEN "0001010001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(20565,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(146062,18);
      WHEN "0001010010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(20815,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(60512,18);
      WHEN "0001010011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(21064,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(197196,18);
      WHEN "0001010100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(21314,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(31389,18);
      WHEN "0001010101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(21563,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(86943,18);
      WHEN "0001010110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(21812,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(101281,18);
      WHEN "0001010111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(22061,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(73969,18);
      WHEN "0001011000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(22310,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(4579,18);
      WHEN "0001011001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(22558,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(154826,18);
      WHEN "0001011010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(22806,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(262139,18);
      WHEN "0001011011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(23055,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(63948,18);
      WHEN "0001011100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(23303,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(84120,18);
      WHEN "0001011101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(23551,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(60088,18);
      WHEN "0001011110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(23798,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(253578,18);
      WHEN "0001011111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(24046,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(139883,18);
      WHEN "0001100000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(24293,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(242876,18);
      WHEN "0001100001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(24541,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(37856,18);
      WHEN "0001100010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(24788,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(48697,18);
      WHEN "0001100011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(25035,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(12847,18);
      WHEN "0001100100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(25281,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(192040,18);
      WHEN "0001100101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(25528,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(61583,18);
      WHEN "0001100110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(25774,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(145360,18);
      WHEN "0001100111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(26020,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(180824,18);
      WHEN "0001101000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(26266,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(167574,18);
      WHEN "0001101001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(26512,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(105213,18);
      WHEN "0001101010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(26757,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(255489,18);
      WHEN "0001101011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(27003,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(93717,18);
      WHEN "0001101100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(27248,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(143796,18);
      WHEN "0001101101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(27493,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(143189,18);
      WHEN "0001101110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(27738,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(91508,18);
      WHEN "0001101111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(27982,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(250512,18);
      WHEN "0001110000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(28227,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(95529,18);
      WHEN "0001110001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(28471,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(150463,18);
      WHEN "0001110010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(28715,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(152791,18);
      WHEN "0001110011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(28959,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(102135,18);
      WHEN "0001110100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(29202,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(260263,18);
      WHEN "0001110101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(29446,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(102513,18);
      WHEN "0001110110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(29689,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(152801,18);
      WHEN "0001110111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(29932,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(148615,18);
      WHEN "0001111000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(30175,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(89586,18);
      WHEN "0001111001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(30417,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(237492,18);
      WHEN "0001111010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(30660,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(67684,18);
      WHEN "0001111011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(30902,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(104088,18);
      WHEN "0001111100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(31144,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(84201,18);
      WHEN "0001111101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(31386,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(7666,18);
      WHEN "0001111110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(31627,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(136273,18);
      WHEN "0001111111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(31868,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(207526,18);
      WHEN "0010000000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(32109,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(221074,18);
      WHEN "0010000001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(32350,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(176570,18);
      WHEN "0010000010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(32591,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(73668,18);
      WHEN "0010000011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(32831,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(174167,18);
      WHEN "0010000100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(33071,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(215584,18);
      WHEN "0010000101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(33311,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(197579,18);
      WHEN "0010000110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(33551,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(119815,18);
      WHEN "0010000111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(33790,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(244102,18);
      WHEN "0010001000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(34030,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(45819,18);
      WHEN "0010001001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(34269,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(48923,18);
      WHEN "0010001010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(34507,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(253089,18);
      WHEN "0010001011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(34746,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(133701,18);
      WHEN "0010001100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(34984,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(214724,18);
      WHEN "0010001101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(35222,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(233694,18);
      WHEN "0010001110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(35460,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(190291,18);
      WHEN "0010001111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(35698,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(84200,18);
      WHEN "0010010000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(35935,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(177249,18);
      WHEN "0010010001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(36172,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(206983,18);
      WHEN "0010010010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(36409,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(173093,18);
      WHEN "0010010011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(36646,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(75271,18);
      WHEN "0010010100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(36882,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(175356,18);
      WHEN "0010010101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(37118,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(210901,18);
      WHEN "0010010110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(37354,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(181607,18);
      WHEN "0010010111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(37590,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(87173,18);
      WHEN "0010011000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(37825,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(189450,18);
      WHEN "0010011001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(38060,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(226000,18);
      WHEN "0010011010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(38295,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(196531,18);
      WHEN "0010011011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(38530,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(100754,18);
      WHEN "0010011100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(38764,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(200528,18);
      WHEN "0010011101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(38998,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(233423,18);
      WHEN "0010011110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(39232,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(199158,18);
      WHEN "0010011111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(39466,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(97454,18);
      WHEN "0010100000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(39699,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(190176,18);
      WHEN "0010100001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(39932,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(214908,18);
      WHEN "0010100010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(40165,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(171374,18);
      WHEN "0010100011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(40398,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(59307,18);
      WHEN "0010100100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(40630,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(140580,18);
      WHEN "0010100101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(40862,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(152786,18);
      WHEN "0010100110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(41094,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(95661,18);
      WHEN "0010100111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(41325,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(231088,18);
      WHEN "0010101000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(41557,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(34520,18);
      WHEN "0010101001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(41788,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(29989,18);
      WHEN "0010101010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(42018,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(217242,18);
      WHEN "0010101011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(42249,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(71738,18);
      WHEN "0010101100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(42479,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(117517,18);
      WHEN "0010101101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(42709,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(92187,18);
      WHEN "0010101110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(42938,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(257648,18);
      WHEN "0010101111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(43168,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(89371,18);
      WHEN "0010110000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(43397,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(111402,18);
      WHEN "0010110001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(43626,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(61360,18);
      WHEN "0010110010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(43854,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(201155,18);
      WHEN "0010110011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(44083,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(6265,18);
      WHEN "0010110100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(44311,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(747,18);
      WHEN "0010110101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(44538,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(184374,18);
      WHEN "0010110110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(44766,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(32631,18);
      WHEN "0010110111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(44993,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(69583,18);
      WHEN "0010111000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(45220,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(32865,18);
      WHEN "0010111001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(45446,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(184401,18);
      WHEN "0010111010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(45672,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(261830,18);
      WHEN "0010111011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(45899,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(2795,18);
      WHEN "0010111100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(46124,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(193515,18);
      WHEN "0010111101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(46350,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(47349,18);
      WHEN "0010111110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(46575,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(88377,18);
      WHEN "0010111111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(46800,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(54250,18);
      WHEN "0011000000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(47024,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(206908,18);
      WHEN "0011000001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(47249,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(21864,18);
      WHEN "0011000010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(47473,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(23207,18);
      WHEN "0011000011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(47696,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(210741,18);
      WHEN "0011000100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(47920,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(59984,18);
      WHEN "0011000101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(48143,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(95032,18);
      WHEN "0011000110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(48366,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(53554,18);
      WHEN "0011000111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(48588,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(197504,18);
      WHEN "0011001000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(48811,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(2412,18);
      WHEN "0011001001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(49032,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(254526,18);
      WHEN "0011001010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(49254,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(167234,18);
      WHEN "0011001011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(49476,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(2502,18);
      WHEN "0011001100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(49697,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(22299,18);
      WHEN "0011001101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(49917,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(226451,18);
      WHEN "0011001110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(50138,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(90499,18);
      WHEN "0011001111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(50358,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(138562,18);
      WHEN "0011010000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(50578,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(108329,18);
      WHEN "0011010001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(50797,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(261779,18);
      WHEN "0011010010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(51017,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(74462,18);
      WHEN "0011010011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(51236,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(70506,18);
      WHEN "0011010100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(51454,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(249754,18);
      WHEN "0011010101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(51673,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(87760,18);
      WHEN "0011010110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(51891,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(108660,18);
      WHEN "0011010111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(52109,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(50158,18);
      WHEN "0011011000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(52326,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(174249,18);
      WHEN "0011011001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(52543,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(218642,18);
      WHEN "0011011010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(52760,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(183192,18);
      WHEN "0011011011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(52977,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(67756,18);
      WHEN "0011011100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(53193,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(134338,18);
      WHEN "0011011101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(53409,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(120655,18);
      WHEN "0011011110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(53625,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(26571,18);
      WHEN "0011011111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(53840,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(114096,18);
      WHEN "0011100000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(54055,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(120953,18);
      WHEN "0011100001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(54270,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(47013,18);
      WHEN "0011100010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(54484,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(154291,18);
      WHEN "0011100011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(54698,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(180519,18);
      WHEN "0011100100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(54912,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(125572,18);
      WHEN "0011100101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(55125,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(251472,18);
      WHEN "0011100110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(55339,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(33813,18);
      WHEN "0011100111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(55551,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(258909,18);
      WHEN "0011101000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(55764,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(140212,18);
      WHEN "0011101001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(55976,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(201898,18);
      WHEN "0011101010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(56188,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(181710,18);
      WHEN "0011101011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(56400,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(79540,18);
      WHEN "0011101100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(56611,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(157424,18);
      WHEN "0011101101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(56822,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(153114,18);
      WHEN "0011101110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(57033,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(66506,18);
      WHEN "0011101111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(57243,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(159643,18);
      WHEN "0011110000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(57453,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(170281,18);
      WHEN "0011110001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(57663,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(98325,18);
      WHEN "0011110010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(57872,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(205822,18);
      WHEN "0011110011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(58081,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(230535,18);
      WHEN "0011110100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(58290,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(172373,18);
      WHEN "0011110101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(58499,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(31247,18);
      WHEN "0011110110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(58707,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(69214,18);
      WHEN "0011110111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(58915,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(24044,18);
      WHEN "0011111000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(59122,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(157797,18);
      WHEN "0011111001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(59329,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(208248,18);
      WHEN "0011111010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(59536,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(175318,18);
      WHEN "0011111011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(59743,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(58929,18);
      WHEN "0011111100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(59949,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(121149,18);
      WHEN "0011111101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(60155,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(99760,18);
      WHEN "0011111110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(60360,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(256834,18);
      WHEN "0011111111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(60566,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(68012,18);
      WHEN "0100000000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(60771,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(57516,18);
      WHEN "0100000001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(60975,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(225277,18);
      WHEN "0100000010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(61180,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(46944,18);
      WHEN "0100000011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(61384,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(46741,18);
      WHEN "0100000100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(61587,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(224608,18);
      WHEN "0100000101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(61791,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(56198,18);
      WHEN "0100000110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(61994,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(65741,18);
      WHEN "0100000111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(62196,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(253182,18);
      WHEN "0100001000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(62399,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(94178,18);
      WHEN "0100001001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(62601,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(112967,18);
      WHEN "0100001010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(62803,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(47353,18);
      WHEN "0100001011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(63004,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(159433,18);
      WHEN "0100001100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(63205,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(187015,18);
      WHEN "0100001101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(63406,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(130055,18);
      WHEN "0100001110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(63606,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(250654,18);
      WHEN "0100001111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(63807,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(24481,18);
      WHEN "0100010000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(64006,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(237930,18);
      WHEN "0100010001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(64206,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(104530,18);
      WHEN "0100010010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(64405,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(148532,18);
      WHEN "0100010011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(64604,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(107758,18);
      WHEN "0100010100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(64802,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(244320,18);
      WHEN "0100010101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(65001,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(33897,18);
      WHEN "0100010110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(65199,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(747,18);
      WHEN "0100010111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(65396,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(144844,18);
      WHEN "0100011000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(65593,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(204016,18);
      WHEN "0100011001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(65790,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(178238,18);
      WHEN "0100011010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(65987,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(67488,18);
      WHEN "0100011011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(66183,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(133888,18);
      WHEN "0100011100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(66379,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(115273,18);
      WHEN "0100011101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(66575,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(11625,18);
      WHEN "0100011110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(66770,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(85072,18);
      WHEN "0100011111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(66965,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(73455,18);
      WHEN "0100100000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(67159,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(238902,18);
      WHEN "0100100001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(67354,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(57115,18);
      WHEN "0100100010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(67548,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(52371,18);
      WHEN "0100100011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(67741,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(224661,18);
      WHEN "0100100100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(67935,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(49688,18);
      WHEN "0100100101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(68128,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(51735,18);
      WHEN "0100100110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(68320,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(230798,18);
      WHEN "0100100111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(68513,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(62585,18);
      WHEN "0100101000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(68705,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(71382,18);
      WHEN "0100101001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(68896,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(257190,18);
      WHEN "0100101010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(69088,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(95722,18);
      WHEN "0100101011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(69279,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(111268,18);
      WHEN "0100101100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(69470,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(41689,18);
      WHEN "0100101101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(69660,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(149135,18);
      WHEN "0100101110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(69850,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(171468,18);
      WHEN "0100101111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(70040,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(108696,18);
      WHEN "0100110000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(70229,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(222974,18);
      WHEN "0100110001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(70418,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(252170,18);
      WHEN "0100110010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(70607,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(196294,18);
      WHEN "0100110011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(70796,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(55362,18);
      WHEN "0100110100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(70984,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(91533,18);
      WHEN "0100110101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(71172,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(42680,18);
      WHEN "0100110110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(71359,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(170964,18);
      WHEN "0100110111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(71546,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(214261,18);
      WHEN "0100111000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(71733,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(172591,18);
      WHEN "0100111001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(71920,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(45977,18);
      WHEN "0100111010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(72106,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(96586,18);
      WHEN "0100111011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(72292,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(62298,18);
      WHEN "0100111100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(72477,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(205284,18);
      WHEN "0100111101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(72663,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(1281,18);
      WHEN "0100111110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(72847,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(236752,18);
      WHEN "0100111111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(73032,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(125293,18);
      WHEN "0101000000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(73216,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(191223,18);
      WHEN "0101000001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(73400,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(172431,18);
      WHEN "0101000010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(73584,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(68949,18);
      WHEN "0101000011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(73767,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(142957,18);
      WHEN "0101000100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(73950,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(132346,18);
      WHEN "0101000101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(74133,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(37152,18);
      WHEN "0101000110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(74315,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(119559,18);
      WHEN "0101000111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(74497,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(117461,18);
      WHEN "0101001000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(74679,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(30899,18);
      WHEN "0101001001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(74860,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(122058,18);
      WHEN "0101001010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(75041,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(128837,18);
      WHEN "0101001011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(75222,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(51281,18);
      WHEN "0101001100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(75402,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(151578,18);
      WHEN "0101001101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(75582,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(167630,18);
      WHEN "0101001110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(75762,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(99484,18);
      WHEN "0101001111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(75941,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(209334,18);
      WHEN "0101010000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(76120,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(235084,18);
      WHEN "0101010001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(76299,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(176784,18);
      WHEN "0101010010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(76478,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(34487,18);
      WHEN "0101010011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(76656,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(70389,18);
      WHEN "0101010100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(76834,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(22400,18);
      WHEN "0101010101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(77011,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(152718,18);
      WHEN "0101010110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(77188,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(199256,18);
      WHEN "0101010111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(77365,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(162070,18);
      WHEN "0101011000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(77542,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(41217,18);
      WHEN "0101011001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(77718,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(98901,18);
      WHEN "0101011010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(77894,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(73038,18);
      WHEN "0101011011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(78069,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(225832,18);
      WHEN "0101011100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(78245,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(33058,18);
      WHEN "0101011101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(78420,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(19065,18);
      WHEN "0101011110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(78594,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(183917,18);
      WHEN "0101011111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(78769,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(3392,18);
      WHEN "0101100000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(78943,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(1843,18);
      WHEN "0101100001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(79116,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(179336,18);
      WHEN "0101100010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(79290,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(11651,18);
      WHEN "0101100011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(79463,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(23144,18);
      WHEN "0101100100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(79635,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(213885,18);
      WHEN "0101100101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(79808,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(59656,18);
      WHEN "0101100110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(79980,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(84815,18);
      WHEN "0101100111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(80152,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(27291,18);
      WHEN "0101101000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(80323,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(149301,18);
      WHEN "0101101001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(80494,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(188773,18);
      WHEN "0101101010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(80665,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(145784,18);
      WHEN "0101101011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(80836,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(20408,18);
      WHEN "0101101100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(81006,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(74865,18);
      WHEN "0101101101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(81176,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(47089,18);
      WHEN "0101101110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(81345,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(199302,18);
      WHEN "0101101111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(81515,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(7293,18);
      WHEN "0101110000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(81683,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(257575,18);
      WHEN "0101110001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(81852,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(163796,18);
      WHEN "0101110010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(82020,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(250325,18);
      WHEN "0101110011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(82188,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(255100,18);
      WHEN "0101110100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(82356,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(178203,18);
      WHEN "0101110101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(82524,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(19719,18);
      WHEN "0101110110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(82691,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(41874,18);
      WHEN "0101110111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(82857,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(244755,18);
      WHEN "0101111000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(83024,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(104158,18);
      WHEN "0101111001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(83190,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(144458,18);
      WHEN "0101111010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(83356,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(103598,18);
      WHEN "0101111011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(83521,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(243810,18);
      WHEN "0101111100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(83687,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(40895,18);
      WHEN "0101111101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(83852,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(19229,18);
      WHEN "0101111110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(84016,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(178903,18);
      WHEN "0101111111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(84180,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(257864,18);
      WHEN "0110000000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(84344,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(256201,18);
      WHEN "0110000001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(84508,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(174008,18);
      WHEN "0110000010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(84672,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(11377,18);
      WHEN "0110000011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(84835,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(30546,18);
      WHEN "0110000100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(84997,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(231607,18);
      WHEN "0110000101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(85160,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(90368,18);
      WHEN "0110000110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(85322,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(131213,18);
      WHEN "0110000111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(85484,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(92091,18);
      WHEN "0110001000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(85645,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(235245,18);
      WHEN "0110001001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(85807,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(36483,18);
      WHEN "0110001010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(85968,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(20191,18);
      WHEN "0110001011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(86128,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(186467,18);
      WHEN "0110001100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(86289,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(11121,18);
      WHEN "0110001101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(86449,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(18541,18);
      WHEN "0110001110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(86608,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(208828,18);
      WHEN "0110001111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(86768,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(57793,18);
      WHEN "0110010000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(86927,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(89826,18);
      WHEN "0110010001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(87086,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(42884,18);
      WHEN "0110010010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(87244,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(179213,18);
      WHEN "0110010011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(87402,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(236772,18);
      WHEN "0110010100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(87560,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(215665,18);
      WHEN "0110010101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(87718,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(115995,18);
      WHEN "0110010110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(87875,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(200010,18);
      WHEN "0110010111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(88032,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(205672,18);
      WHEN "0110011000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(88189,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(133084,18);
      WHEN "0110011001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(88345,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(244498,18);
      WHEN "0110011010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(88502,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(15731,18);
      WHEN "0110011011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(88657,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(233323,18);
      WHEN "0110011100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(88813,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(110948,18);
      WHEN "0110011101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(88968,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(173002,18);
      WHEN "0110011110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(89123,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(157449,18);
      WHEN "0110011111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(89278,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(64397,18);
      WHEN "0110100000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(89432,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(156101,18);
      WHEN "0110100001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(89586,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(170525,18);
      WHEN "0110100010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(89740,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(107780,18);
      WHEN "0110100011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(89893,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(230119,18);
      WHEN "0110100100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(90047,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(13365,18);
      WHEN "0110100101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(90199,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(244062,18);
      WHEN "0110100110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(90352,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(135889,18);
      WHEN "0110100111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(90504,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(213247,18);
      WHEN "0110101000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(90656,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(214103,18);
      WHEN "0110101001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(90808,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(138570,18);
      WHEN "0110101010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(90959,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(248907,18);
      WHEN "0110101011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(91111,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(20937,18);
      WHEN "0110101100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(91261,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(241208,18);
      WHEN "0110101101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(91412,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(123401,18);
      WHEN "0110101110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(91562,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(191920,18);
      WHEN "0110101111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(91712,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(184734,18);
      WHEN "0110110000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(91862,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(101960,18);
      WHEN "0110110001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(92011,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(205858,18);
      WHEN "0110110010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(92160,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(234399,18);
      WHEN "0110110011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(92309,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(187700,18);
      WHEN "0110110100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(92458,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(65877,18);
      WHEN "0110110101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(92606,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(131192,18);
      WHEN "0110110110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(92754,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(121618,18);
      WHEN "0110110111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(92902,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(37273,18);
      WHEN "0110111000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(93049,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(140418,18);
      WHEN "0110111001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(93196,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(169029,18);
      WHEN "0110111010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(93343,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(123223,18);
      WHEN "0110111011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(93490,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(3119,18);
      WHEN "0110111100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(93636,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(70981,18);
      WHEN "0110111101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(93782,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(64784,18);
      WHEN "0110111110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(93927,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(246792,18);
      WHEN "0110111111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(94073,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(92836,18);
      WHEN "0111000000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(94218,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(127326,18);
      WHEN "0111000001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(94363,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(88237,18);
      WHEN "0111000010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(94507,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(237834,18);
      WHEN "0111000011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(94652,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(51950,18);
      WHEN "0111000100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(94796,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(54995,18);
      WHEN "0111000101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(94939,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(247090,18);
      WHEN "0111000110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(95083,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(104069,18);
      WHEN "0111000111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(95226,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(150342,18);
      WHEN "0111001000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(95369,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(123886,18);
      WHEN "0111001001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(95512,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(24825,18);
      WHEN "0111001010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(95654,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(115424,18);
      WHEN "0111001011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(95796,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(133663,18);
      WHEN "0111001100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(95938,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(79665,18);
      WHEN "0111001101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(96079,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(215697,18);
      WHEN "0111001110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(96221,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(17594,18);
      WHEN "0111001111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(96362,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(9768,18);
      WHEN "0111010000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(96502,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(192343,18);
      WHEN "0111010001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(96643,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(41154,18);
      WHEN "0111010010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(96783,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(80615,18);
      WHEN "0111010011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(96923,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(48704,18);
      WHEN "0111010100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(97062,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(207691,18);
      WHEN "0111010101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(97202,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(33412,18);
      WHEN "0111010110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(97341,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(50281,18);
      WHEN "0111010111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(97479,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(258422,18);
      WHEN "0111011000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(97618,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(133671,18);
      WHEN "0111011001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(97756,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(200444,18);
      WHEN "0111011010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(97894,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(196720,18);
      WHEN "0111011011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(98032,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(122625,18);
      WHEN "0111011100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(98169,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(240430,18);
      WHEN "0111011101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(98307,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(25971,18);
      WHEN "0111011110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(98444,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(3664,18);
      WHEN "0111011111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(98580,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(173633,18);
      WHEN "0111100000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(98717,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(11717,18);
      WHEN "0111100001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(98853,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(42330,18);
      WHEN "0111100010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(98989,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(3456,18);
      WHEN "0111100011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(99124,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(157363,18);
      WHEN "0111100100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(99259,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(242035,18);
      WHEN "0111100101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(99394,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(257599,18);
      WHEN "0111100110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(99529,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(204180,18);
      WHEN "0111100111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(99664,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(81908,18);
      WHEN "0111101000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(99798,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(153051,18);
      WHEN "0111101001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(99932,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(155593,18);
      WHEN "0111101010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(100066,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(89662,18);
      WHEN "0111101011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(100199,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(217528,18);
      WHEN "0111101100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(100333,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(15031,18);
      WHEN "0111101101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(100466,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(6586,18);
      WHEN "0111101110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(100598,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(192320,18);
      WHEN "0111101111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(100731,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(48074,18);
      WHEN "0111110000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(100863,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(98261,18);
      WHEN "0111110001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(100995,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(80868,18);
      WHEN "0111110010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(101126,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(258163,18);
      WHEN "0111110011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(101258,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(105988,18);
      WHEN "0111110100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(101389,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(148759,18);
      WHEN "0111110101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(101520,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(124458,18);
      WHEN "0111110110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(101651,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(33214,18);
      WHEN "0111110111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(101781,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(137298,18);
      WHEN "0111111000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(101911,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(174695,18);
      WHEN "0111111001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(102041,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(145532,18);
      WHEN "0111111010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(102171,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(49937,18);
      WHEN "0111111011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(102300,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(150182,18);
      WHEN "0111111100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(102429,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(184251,18);
      WHEN "0111111101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(102558,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(152273,18);
      WHEN "0111111110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(102687,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(54374,18);
      WHEN "0111111111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(102815,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(152827,18);
      WHEN "1000000000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(102943,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(185617,18);
      WHEN "1000000001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(103071,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(152870,18);
      WHEN "1000000010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(103199,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(54715,18);
      WHEN "1000000011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(103326,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(153425,18);
      WHEN "1000000100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(103453,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(186982,18);
      WHEN "1000000101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(103580,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(155515,18);
      WHEN "1000000110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(103707,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(59152,18);
      WHEN "1000000111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(103833,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(160165,18);
      WHEN "1000001000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(103959,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(196538,18);
      WHEN "1000001001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(104085,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(168399,18);
      WHEN "1000001010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(104211,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(75875,18);
      WHEN "1000001011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(104336,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(181239,18);
      WHEN "1000001100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(104461,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(222475,18);
      WHEN "1000001101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(104586,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(199709,18);
      WHEN "1000001110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(104711,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(113070,18);
      WHEN "1000001111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(104835,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(224830,18);
      WHEN "1000010000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(104960,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(10829,18);
      WHEN "1000010001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(105083,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(257625,18);
      WHEN "1000010010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(105207,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(178916,18);
      WHEN "1000010011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(105331,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(36971,18);
      WHEN "1000010100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(105454,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(94064,18);
      WHEN "1000010101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(105577,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(88176,18);
      WHEN "1000010110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(105700,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(19436,18);
      WHEN "1000010111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(105822,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(150116,18);
      WHEN "1000011000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(105944,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(218198,18);
      WHEN "1000011001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(106066,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(223809,18);
      WHEN "1000011010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(106188,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(167077,18);
      WHEN "1000011011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(106310,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(48129,18);
      WHEN "1000011100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(106431,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(129236,18);
      WHEN "1000011101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(106552,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(148382,18);
      WHEN "1000011110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(106673,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(105692,18);
      WHEN "1000011111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(106794,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(1293,18);
      WHEN "1000100000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(106914,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(97458,18);
      WHEN "1000100001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(107034,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(132167,18);
      WHEN "1000100010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(107154,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(105548,18);
      WHEN "1000100011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(107274,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(17728,18);
      WHEN "1000100100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(107393,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(130976,18);
      WHEN "1000100101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(107512,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(183276,18);
      WHEN "1000100110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(107631,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(174753,18);
      WHEN "1000100111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(107750,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(105533,18);
      WHEN "1000101000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(107868,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(237887,18);
      WHEN "1000101001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(107987,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(47653,18);
      WHEN "1000101010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(108105,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(59244,18);
      WHEN "1000101011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(108223,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(10643,18);
      WHEN "1000101100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(108340,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(164119,18);
      WHEN "1000101101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(108457,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(257653,18);
      WHEN "1000101110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(108575,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(29228,18);
      WHEN "1000101111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(108692,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(3255,18);
      WHEN "1000110000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(108808,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(179862,18);
      WHEN "1000110001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(108925,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(34885,18);
      WHEN "1000110010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(109041,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(92737,18);
      WHEN "1000110011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(109157,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(91399,18);
      WHEN "1000110100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(109273,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(30995,18);
      WHEN "1000110101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(109388,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(173795,18);
      WHEN "1000110110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(109503,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(257779,18);
      WHEN "1000110111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(109619,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(20928,18);
      WHEN "1000111000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(109733,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(249798,18);
      WHEN "1000111001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(109848,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(158081,18);
      WHEN "1000111010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(109963,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(8045,18);
      WHEN "1000111011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(110077,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(61959,18);
      WHEN "1000111100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(110191,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(57801,18);
      WHEN "1000111101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(110304,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(257841,18);
      WHEN "1000111110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(110418,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(137913,18);
      WHEN "1000111111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(110531,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(222429,18);
      WHEN "1001000000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(110644,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(249369,18);
      WHEN "1001000001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(110757,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(218855,18);
      WHEN "1001000010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(110870,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(131010,18);
      WHEN "1001000011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(110982,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(248102,18);
      WHEN "1001000100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(111095,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(45965,18);
      WHEN "1001000101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(111207,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(49010,18);
      WHEN "1001000110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(111318,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(257360,18);
      WHEN "1001000111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(111430,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(146848,18);
      WHEN "1001001000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(111541,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(241886,18);
      WHEN "1001001001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(111653,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(18306,18);
      WHEN "1001001010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(111764,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(520,18);
      WHEN "1001001011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(111874,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(188648,18);
      WHEN "1001001100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(111985,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(58525,18);
      WHEN "1001001101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(112095,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(134560,18);
      WHEN "1001001110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(112205,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(154730,18);
      WHEN "1001001111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(112315,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(119156,18);
      WHEN "1001010000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(112425,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(27960,18);
      WHEN "1001010001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(112534,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(143406,18);
      WHEN "1001010010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(112643,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(203471,18);
      WHEN "1001010011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(112752,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(208276,18);
      WHEN "1001010100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(112861,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(157941,18);
      WHEN "1001010101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(112970,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(52586,18);
      WHEN "1001010110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(113078,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(154475,18);
      WHEN "1001010111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(113186,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(201584,18);
      WHEN "1001011000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(113294,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(194033,18);
      WHEN "1001011001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(113402,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(131941,18);
      WHEN "1001011010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(113510,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(15429,18);
      WHEN "1001011011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(113617,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(106759,18);
      WHEN "1001011100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(113724,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(143905,18);
      WHEN "1001011101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(113831,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(126988,18);
      WHEN "1001011110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(113938,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(56126,18);
      WHEN "1001011111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(114044,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(193581,18);
      WHEN "1001100000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(114151,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(15184,18);
      WHEN "1001100001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(114257,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(45342,18);
      WHEN "1001100010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(114363,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(22027,18);
      WHEN "1001100011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(114468,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(207502,18);
      WHEN "1001100100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(114574,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(77597,18);
      WHEN "1001100101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(114679,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(156717,18);
      WHEN "1001100110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(114784,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(182836,18);
      WHEN "1001100111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(114889,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(156070,18);
      WHEN "1001101000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(114994,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(76538,18);
      WHEN "1001101001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(115098,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(206498,18);
      WHEN "1001101010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(115203,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(21782,18);
      WHEN "1001101011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(115307,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(46791,18);
      WHEN "1001101100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(115411,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(19500,18);
      WHEN "1001101101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(115514,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(202167,18);
      WHEN "1001101110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(115618,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(70622,18);
      WHEN "1001101111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(115721,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(149267,18);
      WHEN "1001110000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(115824,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(176075,18);
      WHEN "1001110001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(115927,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(151160,18);
      WHEN "1001110010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(116030,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(74638,18);
      WHEN "1001110011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(116132,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(208767,18);
      WHEN "1001110100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(116235,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(29375,18);
      WHEN "1001110101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(116337,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(60864,18);
      WHEN "1001110110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(116439,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(41205,18);
      WHEN "1001110111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(116540,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(232655,18);
      WHEN "1001111000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(116642,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(111041,18);
      WHEN "1001111001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(116743,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(200765,18);
      WHEN "1001111010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(116844,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(239796,18);
      WHEN "1001111011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(116945,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(228248,18);
      WHEN "1001111100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(117046,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(166234,18);
      WHEN "1001111101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(117147,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(53867,18);
      WHEN "1001111110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(117247,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(153404,18);
      WHEN "1001111111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(117347,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(202814,18);
      WHEN "1010000000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(117447,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(202209,18);
      WHEN "1010000001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(117547,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(151701,18);
      WHEN "1010000010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(117647,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(51403,18);
      WHEN "1010000011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(117746,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(163571,18);
      WHEN "1010000100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(117845,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(226171,18);
      WHEN "1010000101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(117944,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(239317,18);
      WHEN "1010000110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(118043,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(203118,18);
      WHEN "1010000111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(118142,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(117687,18);
      WHEN "1010001000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(118240,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(245278,18);
      WHEN "1010001001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(118339,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(61714,18);
      WHEN "1010001010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(118437,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(91393,18);
      WHEN "1010001011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(118535,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(72282,18);
      WHEN "1010001100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(118633,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(4490,18);
      WHEN "1010001101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(118730,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(150272,18);
      WHEN "1010001110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(118827,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(247594,18);
      WHEN "1010001111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(118925,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(34421,18);
      WHEN "1010010000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(119022,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(35150,18);
      WHEN "1010010001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(119118,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(249890,18);
      WHEN "1010010010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(119215,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(154463,18);
      WHEN "1010010011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(119312,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(11120,18);
      WHEN "1010010100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(119408,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(82116,18);
      WHEN "1010010101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(119504,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(105413,18);
      WHEN "1010010110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(119600,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(81120,18);
      WHEN "1010010111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(119696,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(9344,18);
      WHEN "1010011000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(119791,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(152339,18);
      WHEN "1010011001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(119886,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(248066,18);
      WHEN "1010011010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(119982,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(34490,18);
      WHEN "1010011011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(120077,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(36005,18);
      WHEN "1010011100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(120171,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(252718,18);
      WHEN "1010011101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(120266,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(160448,18);
      WHEN "1010011110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(120361,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(21445,18);
      WHEN "1010011111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(120455,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(97961,18);
      WHEN "1010100000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(120549,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(127955,18);
      WHEN "1010100001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(120643,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(111535,18);
      WHEN "1010100010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(120737,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(48807,18);
      WHEN "1010100011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(120830,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(202019,18);
      WHEN "1010100100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(120924,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(46988,18);
      WHEN "1010100101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(121017,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(108109,18);
      WHEN "1010100110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(121110,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(123341,18);
      WHEN "1010100111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(121203,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(92789,18);
      WHEN "1010101000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(121296,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(16558,18);
      WHEN "1010101001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(121388,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(156895,18);
      WHEN "1010101010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(121480,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(251761,18);
      WHEN "1010101011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(121573,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(39116,18);
      WHEN "1010101100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(121665,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(43350,18);
      WHEN "1010101101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(121757,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(2424,18);
      WHEN "1010101110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(121848,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(178584,18);
      WHEN "1010101111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(121940,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(47646,18);
      WHEN "1010110000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(122031,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(134000,18);
      WHEN "1010110001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(122122,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(175604,18);
      WHEN "1010110010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(122213,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(172562,18);
      WHEN "1010110011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(122304,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(124974,18);
      WHEN "1010110100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(122395,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(32943,18);
      WHEN "1010110101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(122485,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(158715,18);
      WHEN "1010110110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(122575,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(240246,18);
      WHEN "1010110111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(122666,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(15495,18);
      WHEN "1010111000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(122756,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(8850,18);
      WHEN "1010111001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(122845,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(220412,18);
      WHEN "1010111010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(122935,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(125994,18);
      WHEN "1010111011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(123024,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(249984,18);
      WHEN "1010111100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(123114,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(68194,18);
      WHEN "1010111101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(123203,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(105012,18);
      WHEN "1010111110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(123292,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(98395,18);
      WHEN "1010111111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(123381,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(48441,18);
      WHEN "1011000000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(123469,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(217394,18);
      WHEN "1011000001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(123558,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(81065,18);
      WHEN "1011000010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(123646,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(163841,18);
      WHEN "1011000011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(123734,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(203676,18);
      WHEN "1011000100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(123822,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(200670,18);
      WHEN "1011000101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(123910,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(154921,18);
      WHEN "1011000110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(123998,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(66526,18);
      WHEN "1011000111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(124085,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(197727,18);
      WHEN "1011001000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(124173,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(24335,18);
      WHEN "1011001001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(124260,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(70734,18);
      WHEN "1011001010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(124347,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(74878,18);
      WHEN "1011001011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(124434,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(36865,18);
      WHEN "1011001100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(124520,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(218933,18);
      WHEN "1011001101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(124607,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(96893,18);
      WHEN "1011001110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(124693,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(195129,18);
      WHEN "1011001111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(124779,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(251593,18);
      WHEN "1011010000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(124866,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(4237,18);
      WHEN "1011010001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(124951,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(239588,18);
      WHEN "1011010010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(125037,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(171311,18);
      WHEN "1011010011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(125123,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(61644,18);
      WHEN "1011010100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(125208,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(172827,18);
      WHEN "1011010101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(125293,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(242811,18);
      WHEN "1011010110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(125379,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(9546,18);
      WHEN "1011010111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(125463,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(259559,18);
      WHEN "1011011000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(125548,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(206512,18);
      WHEN "1011011001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(125633,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(112644,18);
      WHEN "1011011010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(125717,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(240192,18);
      WHEN "1011011011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(125802,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(64962,18);
      WHEN "1011011100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(125886,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(111335,18);
      WHEN "1011011101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(125970,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(117261,18);
      WHEN "1011011110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(126054,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(82832,18);
      WHEN "1011011111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(126138,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(8142,18);
      WHEN "1011100000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(126221,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(155428,18);
      WHEN "1011100001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(126305,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(492,18);
      WHEN "1011100010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(126388,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(67717,18);
      WHEN "1011100011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(126471,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(95050,18);
      WHEN "1011100100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(126554,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(82582,18);
      WHEN "1011100101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(126637,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(30405,18);
      WHEN "1011100110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(126719,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(200755,18);
      WHEN "1011100111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(126802,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(69435,18);
      WHEN "1011101000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(126884,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(160824,18);
      WHEN "1011101001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(126966,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(212868,18);
      WHEN "1011101010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(127048,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(225659,18);
      WHEN "1011101011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(127130,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(199286,18);
      WHEN "1011101100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(127212,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(133839,18);
      WHEN "1011101101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(127294,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(29409,18);
      WHEN "1011101110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(127375,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(148230,18);
      WHEN "1011101111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(127456,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(228246,18);
      WHEN "1011110000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(127538,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(7403,18);
      WHEN "1011110001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(127619,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(10079,18);
      WHEN "1011110010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(127699,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(236362,18);
      WHEN "1011110011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(127780,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(162053,18);
      WHEN "1011110100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(127861,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(49384,18);
      WHEN "1011110101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(127941,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(160588,18);
      WHEN "1011110110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(128021,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(233609,18);
      WHEN "1011110111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(128102,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(6390,18);
      WHEN "1011111000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(128182,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(3308,18);
      WHEN "1011111001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(128261,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(224450,18);
      WHEN "1011111010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(128341,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(145614,18);
      WHEN "1011111011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(128421,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(29034,18);
      WHEN "1011111100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(128500,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(136938,18);
      WHEN "1011111101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(128579,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(207270,18);
      WHEN "1011111110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(128658,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(240116,18);
      WHEN "1011111111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(128737,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(235563,18);
      WHEN "1100000000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(128816,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(193696,18);
      WHEN "1100000001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(128895,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(114602,18);
      WHEN "1100000010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(128973,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(260510,18);
      WHEN "1100000011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(129052,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(107217,18);
      WHEN "1100000100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(129130,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(179097,18);
      WHEN "1100000101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(129208,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(214091,18);
      WHEN "1100000110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(129286,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(212284,18);
      WHEN "1100000111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(129364,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(173760,18);
      WHEN "1100001000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(129442,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(98604,18);
      WHEN "1100001001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(129519,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(249044,18);
      WHEN "1100001010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(129597,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(100876,18);
      WHEN "1100001011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(129674,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(178473,18);
      WHEN "1100001100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(129751,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(219772,18);
      WHEN "1100001101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(129828,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(224859,18);
      WHEN "1100001110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(129905,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(193817,18);
      WHEN "1100001111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(129982,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(126728,18);
      WHEN "1100010000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(130059,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(23675,18);
      WHEN "1100010001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(130135,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(146885,18);
      WHEN "1100010010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(130211,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(234296,18);
      WHEN "1100010011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(130288,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(23847,18);
      WHEN "1100010100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(130364,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(39908,18);
      WHEN "1100010101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(130440,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(20417,18);
      WHEN "1100010110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(130515,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(227599,18);
      WHEN "1100010111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(130591,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(137248,18);
      WHEN "1100011000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(130667,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(11588,18);
      WHEN "1100011001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(130742,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(112847,18);
      WHEN "1100011010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(130817,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(178959,18);
      WHEN "1100011011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(130892,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(210006,18);
      WHEN "1100011100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(130967,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(206068,18);
      WHEN "1100011101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(131042,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(167226,18);
      WHEN "1100011110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(131117,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(93560,18);
      WHEN "1100011111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(131191,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(247293,18);
      WHEN "1100100000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(131266,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(104218,18);
      WHEN "1100100001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(131340,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(188702,18);
      WHEN "1100100010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(131414,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(238680,18);
      WHEN "1100100011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(131488,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(254231,18);
      WHEN "1100100100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(131562,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(235435,18);
      WHEN "1100100101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(131636,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(182370,18);
      WHEN "1100100110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(131710,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(95115,18);
      WHEN "1100100111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(131783,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(235893,18);
      WHEN "1100101000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(131857,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(80492,18);
      WHEN "1100101001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(131930,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(153280,18);
      WHEN "1100101010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(132003,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(192190,18);
      WHEN "1100101011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(132076,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(197300,18);
      WHEN "1100101100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(132149,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(168687,18);
      WHEN "1100101101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(132222,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(106429,18);
      WHEN "1100101110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(132295,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(10602,18);
      WHEN "1100101111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(132367,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(143428,18);
      WHEN "1100110000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(132439,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(242839,18);
      WHEN "1100110001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(132512,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(46768,18);
      WHEN "1100110010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(132584,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(79578,18);
      WHEN "1100110011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(132656,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(79203,18);
      WHEN "1100110100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(132728,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(45718,18);
      WHEN "1100110101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(132799,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(241342,18);
      WHEN "1100110110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(132871,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(141864,18);
      WHEN "1100110111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(132943,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(9502,18);
      WHEN "1100111000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(133014,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(106476,18);
      WHEN "1100111001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(133085,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(170717,18);
      WHEN "1100111010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(133156,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(202300,18);
      WHEN "1100111011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(133227,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(201300,18);
      WHEN "1100111100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(133298,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(167790,18);
      WHEN "1100111101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(133369,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(101845,18);
      WHEN "1100111110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(133440,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(3539,18);
      WHEN "1100111111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(133510,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(135090,18);
      WHEN "1101000000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(133580,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(234429,18);
      WHEN "1101000001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(133651,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(39483,18);
      WHEN "1101000010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(133721,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(74615,18);
      WHEN "1101000011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(133791,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(77754,18);
      WHEN "1101000100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(133861,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(48973,18);
      WHEN "1101000101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(133930,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(250488,18);
      WHEN "1101000110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(134000,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(158085,18);
      WHEN "1101000111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(134070,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(33979,18);
      WHEN "1101001000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(134139,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(140388,18);
      WHEN "1101001001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(134208,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(215238,18);
      WHEN "1101001010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(134277,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(258603,18);
      WHEN "1101001011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(134347,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(8409,18);
      WHEN "1101001100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(134415,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(251160,18);
      WHEN "1101001101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(134484,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(200497,18);
      WHEN "1101001110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(134553,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(118633,18);
      WHEN "1101001111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(134622,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(5640,18);
      WHEN "1101010000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(134690,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(123732,18);
      WHEN "1101010001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(134758,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(210837,18);
      WHEN "1101010010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(134827,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(4881,18);
      WHEN "1101010011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(134895,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(30222,18);
      WHEN "1101010100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(134963,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(24786,18);
      WHEN "1101010101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(135030,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(250788,18);
      WHEN "1101010110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(135098,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(184008,18);
      WHEN "1101010111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(135166,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(86662,18);
      WHEN "1101011000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(135233,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(220961,18);
      WHEN "1101011001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(135301,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(62688,18);
      WHEN "1101011010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(135368,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(136199,18);
      WHEN "1101011011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(135435,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(179420,18);
      WHEN "1101011100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(135502,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(192419,18);
      WHEN "1101011101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(135569,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(175264,18);
      WHEN "1101011110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(135636,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(128025,18);
      WHEN "1101011111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(135703,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(50768,18);
      WHEN "1101100000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(135769,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(205708,18);
      WHEN "1101100001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(135836,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(68622,18);
      WHEN "1101100010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(135902,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(163868,18);
      WHEN "1101100011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(135968,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(229368,18);
      WHEN "1101100100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(136035,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(3045,18);
      WHEN "1101100101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(136101,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(9256,18);
      WHEN "1101100110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(136166,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(248067,18);
      WHEN "1101100111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(136232,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(195258,18);
      WHEN "1101101000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(136298,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(113037,18);
      WHEN "1101101001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(136364,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(1473,18);
      WHEN "1101101010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(136429,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(122776,18);
      WHEN "1101101011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(136494,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(214867,18);
      WHEN "1101101100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(136560,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(15669,18);
      WHEN "1101101101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(136625,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(49536,18);
      WHEN "1101101110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(136690,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(54389,18);
      WHEN "1101101111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(136755,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(30294,18);
      WHEN "1101110000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(136819,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(239461,18);
      WHEN "1101110001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(136884,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(157665,18);
      WHEN "1101110010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(136949,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(47117,18);
      WHEN "1101110011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(137013,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(170026,18);
      WHEN "1101110100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(137078,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(2168,18);
      WHEN "1101110101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(137142,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(67895,18);
      WHEN "1101110110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(137206,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(105128,18);
      WHEN "1101110111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(137270,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(113931,18);
      WHEN "1101111000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(137334,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(94369,18);
      WHEN "1101111001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(137398,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(46504,18);
      WHEN "1101111010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(137461,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(232546,18);
      WHEN "1101111011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(137525,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(128269,18);
      WHEN "1101111100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(137588,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(258024,18);
      WHEN "1101111101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(137652,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(97588,18);
      WHEN "1101111110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(137715,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(171311,18);
      WHEN "1101111111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(137778,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(217112,18);
      WHEN "1110000000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(137841,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(235053,18);
      WHEN "1110000001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(137904,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(225198,18);
      WHEN "1110000010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(137967,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(187609,18);
      WHEN "1110000011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(138030,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(122349,18);
      WHEN "1110000100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(138093,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(29478,18);
      WHEN "1110000101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(138155,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(171204,18);
      WHEN "1110000110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(138218,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(23299,18);
      WHEN "1110000111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(138280,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(110115,18);
      WHEN "1110001000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(138342,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(169567,18);
      WHEN "1110001001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(138404,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(201718,18);
      WHEN "1110001010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(138466,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(206629,18);
      WHEN "1110001011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(138528,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(184361,18);
      WHEN "1110001100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(138590,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(134974,18);
      WHEN "1110001101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(138652,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(58530,18);
      WHEN "1110001110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(138713,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(217232,18);
      WHEN "1110001111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(138775,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(86854,18);
      WHEN "1110010000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(138836,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(191743,18);
      WHEN "1110010001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(138898,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(7673,18);
      WHEN "1110010010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(138959,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(58989,18);
      WHEN "1110010011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(139020,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(83609,18);
      WHEN "1110010100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(139081,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(81593,18);
      WHEN "1110010101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(139142,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(52999,18);
      WHEN "1110010110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(139202,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(260030,18);
      WHEN "1110010111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(139263,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(178459,18);
      WHEN "1110011000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(139324,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(70488,18);
      WHEN "1110011001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(139384,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(198320,18);
      WHEN "1110011010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(139445,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(37726,18);
      WHEN "1110011011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(139505,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(113052,18);
      WHEN "1110011100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(139565,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(162212,18);
      WHEN "1110011101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(139625,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(185266,18);
      WHEN "1110011110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(139685,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(182271,18);
      WHEN "1110011111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(139745,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(153286,18);
      WHEN "1110100000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(139805,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(98367,18);
      WHEN "1110100001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(139865,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(17573,18);
      WHEN "1110100010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(139924,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(173106,18);
      WHEN "1110100011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(139984,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(40734,18);
      WHEN "1110100100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(140043,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(144803,18);
      WHEN "1110100101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(140102,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(223226,18);
      WHEN "1110100110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(140162,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(13916,18);
      WHEN "1110100111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(140221,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(41217,18);
      WHEN "1110101000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(140280,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(43044,18);
      WHEN "1110101001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(140339,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(19451,18);
      WHEN "1110101010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(140397,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(232640,18);
      WHEN "1110101011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(140456,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(158378,18);
      WHEN "1110101100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(140515,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(58866,18);
      WHEN "1110101101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(140573,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(196304,18);
      WHEN "1110101110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(140632,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(46459,18);
      WHEN "1110101111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(140690,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(133676,18);
      WHEN "1110110000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(140748,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(195865,18);
      WHEN "1110110001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(140806,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(233082,18);
      WHEN "1110110010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(140864,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(245382,18);
      WHEN "1110110011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(140922,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(232821,18);
      WHEN "1110110100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(140980,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(195453,18);
      WHEN "1110110101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(141038,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(133334,18);
      WHEN "1110110110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(141096,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(46517,18);
      WHEN "1110110111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(141153,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(197201,18);
      WHEN "1110111000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(141211,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(61153,18);
      WHEN "1110111001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(141268,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(162716,18);
      WHEN "1110111010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(141325,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(239798,18);
      WHEN "1110111011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(141383,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(30311,18);
      WHEN "1110111100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(141440,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(58595,18);
      WHEN "1110111101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(141497,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(62561,18);
      WHEN "1110111110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(141554,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(42262,18);
      WHEN "1110111111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(141610,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(259896,18);
      WHEN "1111000000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(141667,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(191228,18);
      WHEN "1111000001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(141724,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(98455,18);
      WHEN "1111000010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(141780,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(243774,18);
      WHEN "1111000011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(141837,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(102950,18);
      WHEN "1111000100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(141893,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(200324,18);
      WHEN "1111000101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(141950,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(11660,18);
      WHEN "1111000110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(142006,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(61299,18);
      WHEN "1111000111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(142062,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(87149,18);
      WHEN "1111001000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(142118,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(89262,18);
      WHEN "1111001001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(142174,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(67691,18);
      WHEN "1111001010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(142230,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(22487,18);
      WHEN "1111001011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(142285,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(215847,18);
      WHEN "1111001100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(142341,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(123533,18);
      WHEN "1111001101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(142397,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(7742,18);
      WHEN "1111001110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(142452,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(130668,18);
      WHEN "1111001111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(142507,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(230220,18);
      WHEN "1111010000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(142563,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(44304,18);
      WHEN "1111010001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(142618,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(97259,18);
      WHEN "1111010010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(142673,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(126992,18);
      WHEN "1111010011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(142728,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(133554,18);
      WHEN "1111010100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(142783,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(116996,18);
      WHEN "1111010101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(142838,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(77368,18);
      WHEN "1111010110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(142893,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(14720,18);
      WHEN "1111010111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(142947,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(191247,18);
      WHEN "1111011000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(143002,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(82710,18);
      WHEN "1111011001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(143056,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(213448,18);
      WHEN "1111011010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(143111,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(59223,18);
      WHEN "1111011011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(143165,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(144372,18);
      WHEN "1111011100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(143219,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(206801,18);
      WHEN "1111011101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(143273,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(246559,18);
      WHEN "1111011110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(143328,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(1553,18);
      WHEN "1111011111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(143381,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(258262,18);
      WHEN "1111100000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(143435,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(230304,18);
      WHEN "1111100001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(143489,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(179872,18);
      WHEN "1111100010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(143543,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(107014,18);
      WHEN "1111100011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(143597,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(11781,18);
      WHEN "1111100100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(143650,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(156363,18);
      WHEN "1111100101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(143704,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(16522,18);
      WHEN "1111100110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(143757,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(116595,18);
      WHEN "1111100111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(143810,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(194484,18);
      WHEN "1111101000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(143863,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(250238,18);
      WHEN "1111101001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(143917,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(21762,18);
      WHEN "1111101010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(143970,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(33391,18);
      WHEN "1111101011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(144023,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(23028,18);
      WHEN "1111101100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(144075,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(252866,18);
      WHEN "1111101101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(144128,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(198664,18);
      WHEN "1111101110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(144181,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(122614,18);
      WHEN "1111101111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(144234,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(24761,18);
      WHEN "1111110000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(144286,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(167299,18);
      WHEN "1111110001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(144339,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(25984,18);
      WHEN "1111110010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(144391,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(125154,18);
      WHEN "1111110011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(144443,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(202709,18);
      WHEN "1111110100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(144495,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(258698,18);
      WHEN "1111110101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(144548,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(31022,18);
      WHEN "1111110110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(144600,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(44016,18);
      WHEN "1111110111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(144652,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(35582,18);
      WHEN "1111111000" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(144704,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(5766,18);
      WHEN "1111111001" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(144755,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(216758,18);
      WHEN "1111111010" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(144807,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(144317,18);
      WHEN "1111111011" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(144859,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(50632,18);
      WHEN "1111111100" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(144910,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(197892,18);
      WHEN "1111111101" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(144962,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(61856,18);
      WHEN "1111111110" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(145013,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(166857,18);
      WHEN "1111111111" =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(145064,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(250795,18);
      WHEN others =>
           data(36 DOWNTO 19) <= conv_std_logic_vector(0,18);
           data(18 DOWNTO 1) <= conv_std_logic_vector(0,18);
    END CASE;
  END PROCESS;

END rtl;

LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_CLZ23.VHD                              ***
--***                                             ***
--***   Function: 23 bit Count Leading Zeros      ***
--***                                             ***
--***   22/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_clz23 IS
PORT (
      mantissa : IN STD_LOGIC_VECTOR (23 DOWNTO 1);
      
      leading : OUT STD_LOGIC_VECTOR (5 DOWNTO 1)    
     );
END fp_clz23;

ARCHITECTURE zzz of fp_clz23 IS

  type positiontype IS ARRAY (4 DOWNTO 1) OF STD_LOGIC_VECTOR (5 DOWNTO 1);
  
  signal position, positionmux : positiontype;
  signal zerogroup, firstzero : STD_LOGIC_VECTOR (4 DOWNTO 1);
  signal mannode : STD_LOGIC_VECTOR (6 DOWNTO 1);
  
  component fp_pos51
  GENERIC (start: integer := 0);
  PORT 
       (
        ingroup : IN STD_LOGIC_VECTOR (6 DOWNTO 1); 
        
        position : OUT STD_LOGIC_VECTOR (5 DOWNTO 1)    
       );
  end component;
  
BEGIN

zerogroup(1) <= mantissa(23) OR mantissa(22) OR mantissa(21) OR mantissa(20) OR mantissa(19) OR mantissa(18);
zerogroup(2) <= mantissa(17) OR mantissa(16) OR mantissa(15) OR mantissa(14) OR mantissa(13) OR mantissa(12);
zerogroup(3) <= mantissa(11) OR mantissa(10) OR mantissa(9) OR mantissa(8) OR mantissa(7) OR mantissa(6);
zerogroup(4) <= mantissa(5) OR mantissa(4) OR mantissa(3) OR mantissa(2) OR mantissa(1);

firstzero(1) <= zerogroup(1);
firstzero(2) <= NOT(zerogroup(1)) AND zerogroup(2);
firstzero(3) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND zerogroup(3);
firstzero(4) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND zerogroup(4);
                
pone: fp_pos51 
GENERIC MAP (start=>0) 
PORT MAP (ingroup=>mantissa(23 DOWNTO 18),position=>position(1)(5 DOWNTO 1));
ptwo: fp_pos51 
GENERIC MAP (start=>6) 
PORT MAP (ingroup=>mantissa(17 DOWNTO 12),position=>position(2)(5 DOWNTO 1));
pthr: fp_pos51 
GENERIC MAP (start=>12) 
PORT MAP (ingroup=>mantissa(11 DOWNTO 6),position=>position(3)(5 DOWNTO 1));    
pfiv: fp_pos51 
GENERIC MAP (start=>18) 
PORT MAP (ingroup=>mannode,position=>position(4)(5 DOWNTO 1));    
    
mannode <= mantissa(5 DOWNTO 1) & '0';
                
gma: FOR k IN 1 TO 5 GENERATE
  positionmux(1)(k) <= position(1)(k) AND firstzero(1);
  gmb: FOR j IN 2 TO 4 GENERATE
    positionmux(j)(k) <= positionmux(j-1)(k) OR (position(j)(k) AND firstzero(j));
  END GENERATE;
END GENERATE;
  
leading <= positionmux(4)(5 DOWNTO 1);
                                               
END zzz;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_CLZ36.VHD                              ***
--***                                             ***
--***   Function: 36 bit Count Leading Zeros      ***
--***                                             ***
--***   22/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_clz36 IS
PORT (
      mantissa : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
      
      leading : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
     );
END fp_clz36;

ARCHITECTURE zzz of fp_clz36 IS

  type positiontype IS ARRAY (6 DOWNTO 1) OF STD_LOGIC_VECTOR (6 DOWNTO 1);
  
  signal position, positionmux : positiontype;
  signal zerogroup, firstzero : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal mannode : STD_LOGIC_VECTOR (6 DOWNTO 1);
  
  component fp_pos52
  GENERIC (start: integer := 0);
  PORT 
       (
        ingroup : IN STD_LOGIC_VECTOR (6 DOWNTO 1); 
        
        position : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
       );
  end component;
  
BEGIN

zerogroup(1) <= mantissa(36) OR mantissa(35) OR mantissa(34) OR mantissa(33) OR mantissa(32) OR mantissa(31);
zerogroup(2) <= mantissa(30) OR mantissa(29) OR mantissa(28) OR mantissa(27) OR mantissa(26) OR mantissa(25);
zerogroup(3) <= mantissa(24) OR mantissa(23) OR mantissa(22) OR mantissa(21) OR mantissa(20) OR mantissa(19);
zerogroup(4) <= mantissa(18) OR mantissa(17) OR mantissa(16) OR mantissa(15) OR mantissa(14) OR mantissa(13);
zerogroup(5) <= mantissa(12) OR mantissa(11) OR mantissa(10) OR mantissa(9) OR mantissa(8) OR mantissa(7);
zerogroup(6) <= mantissa(6) OR mantissa(5) OR mantissa(4) OR mantissa(3) OR mantissa(2) OR mantissa(1);

firstzero(1) <= zerogroup(1);
firstzero(2) <= NOT(zerogroup(1)) AND zerogroup(2);
firstzero(3) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND zerogroup(3);
firstzero(4) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND zerogroup(4);
firstzero(5) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND NOT(zerogroup(4)) 
                AND zerogroup(5);
firstzero(6) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND NOT(zerogroup(4)) AND NOT(zerogroup(5)) 
                AND zerogroup(6);
                
pone: fp_pos52 
GENERIC MAP (start=>0) 
PORT MAP (ingroup=>mantissa(36 DOWNTO 31),position=>position(1)(6 DOWNTO 1));
ptwo: fp_pos52 
GENERIC MAP (start=>6) 
PORT MAP (ingroup=>mantissa(30 DOWNTO 25),position=>position(2)(6 DOWNTO 1));
pthr: fp_pos52 
GENERIC MAP (start=>12) 
PORT MAP (ingroup=>mantissa(24 DOWNTO 19),position=>position(3)(6 DOWNTO 1));    
pfor: fp_pos52 
GENERIC MAP (start=>18) 
PORT MAP (ingroup=>mantissa(18 DOWNTO 13),position=>position(4)(6 DOWNTO 1));
pfiv: fp_pos52 
GENERIC MAP (start=>24) 
PORT MAP (ingroup=>mantissa(12 DOWNTO 7),position=>position(5)(6 DOWNTO 1));
psix: fp_pos52 
GENERIC MAP (start=>30) 
PORT MAP (ingroup=>mantissa(6 DOWNTO 1),position=>position(6)(6 DOWNTO 1));
                
gma: FOR k IN 1 TO 6 GENERATE
  positionmux(1)(k) <= position(1)(k) AND firstzero(1);
  gmb: FOR j IN 2 TO 6 GENERATE
    positionmux(j)(k) <= positionmux(j-1)(k) OR (position(j)(k) AND firstzero(j));
  END GENERATE;
END GENERATE;
  
leading <= positionmux(6)(6 DOWNTO 1);
                                               
END zzz;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_CLZ36X6.VHD                            ***
--***                                             ***
--***   Function: 6 bit Count Leading Zeros in a  ***
--***   36 bit number                             ***
--***                                             ***
--***   22/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_clz36x6 IS
PORT (
      mantissa : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
      
      leading : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
     );
END fp_clz36x6;

ARCHITECTURE rtl of fp_clz36x6 IS

  type positiontype IS ARRAY (6 DOWNTO 1) OF STD_LOGIC_VECTOR (6 DOWNTO 1);
  
  signal position, positionmux : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal zerogroup : STD_LOGIC;
  
  component fp_pos52
  GENERIC (start: integer := 0);
  PORT 
       (
        ingroup : IN STD_LOGIC_VECTOR (6 DOWNTO 1); 
        
        position : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
       );
  end component;
  
BEGIN

  zerogroup <= mantissa(36) OR mantissa(35) OR mantissa(34) OR mantissa(33) OR mantissa(32) OR mantissa(31);
                
  pone: fp_pos52 
  GENERIC MAP (start=>0) 
  PORT MAP (ingroup=>mantissa(36 DOWNTO 31),position=>position(6 DOWNTO 1));
                
  gma: FOR k IN 1 TO 6 GENERATE
    positionmux(k) <= position(k) AND zerogroup;
  END GENERATE;
  
  leading <= positionmux;
                                               
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_CORDIC_ATAN1.VHD                       ***
--***                                             ***
--***   Function: ATAN Values Table for SIN and   ***
--***   COS CORDIC Core                           ***
--***                                             ***
--***   22/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_cordic_atan1 IS 
GENERIC (start : positive := 32;
         width : positive := 32;
         indexpoint : positive := 1);
PORT (
      indexbit : IN STD_LOGIC;

	    arctan : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
	  );
END fp_cordic_atan1;

ARCHITECTURE sft OF fp_cordic_atan1 IS
  
  type atantype IS ARRAY (48 DOWNTO 1) OF STD_LOGIC_VECTOR (48 DOWNTO 1); 
  
  signal atannum : atantype;
  
BEGIN
   
  -- "00" + 46 bits
  atannum(1)(48 DOWNTO 1) <= x"3243F6A8885A";
  atannum(2)(48 DOWNTO 1) <= x"1DAC670561BB";
  atannum(3)(48 DOWNTO 1) <= x"0FADBAFC9640";
  atannum(4)(48 DOWNTO 1) <= x"07F56EA6AB0C";
  atannum(5)(48 DOWNTO 1) <= x"03FEAB76E5A0";
  atannum(6)(48 DOWNTO 1) <= x"01FFD55BBA97"; 
  atannum(7)(48 DOWNTO 1) <= x"00FFFAAADDDC";
  atannum(8)(48 DOWNTO 1) <= x"007FFF5556EF";
  atannum(9)(48 DOWNTO 1) <= x"003FFFEAAAB7";
  
  atannum(10)(48 DOWNTO 1) <= x"001FFFFD5556";
  atannum(11)(48 DOWNTO 1) <= x"000FFFFFAAAB"; 
  atannum(12)(48 DOWNTO 1) <= x"0007FFFFF555";
  atannum(13)(48 DOWNTO 1) <= x"0003FFFFFEAB";
  atannum(14)(48 DOWNTO 1) <= x"0001FFFFFFD5";
  atannum(15)(48 DOWNTO 1) <= x"0000FFFFFFFB";
  atannum(16)(48 DOWNTO 1) <= x"00007FFFFFFF"; 
  atannum(17)(48 DOWNTO 1) <= x"000040000000";
  atannum(18)(48 DOWNTO 1) <= x"000020000000";
  atannum(19)(48 DOWNTO 1) <= x"000010000000";
  
  atannum(20)(48 DOWNTO 1) <= x"000008000000";
  atannum(21)(48 DOWNTO 1) <= x"000004000000"; 
  atannum(22)(48 DOWNTO 1) <= x"000002000000";
  atannum(23)(48 DOWNTO 1) <= x"000001000000";
  atannum(24)(48 DOWNTO 1) <= x"000000800000";
  atannum(25)(48 DOWNTO 1) <= x"000000400000";
  atannum(26)(48 DOWNTO 1) <= x"000000200000";  
  atannum(27)(48 DOWNTO 1) <= x"000000100000";
  atannum(28)(48 DOWNTO 1) <= x"000000080000";
  atannum(29)(48 DOWNTO 1) <= x"000000040000";
  
  atannum(30)(48 DOWNTO 1) <= x"000000020000";
  atannum(31)(48 DOWNTO 1) <= x"000000010000"; 
  atannum(32)(48 DOWNTO 1) <= x"000000008000";
  atannum(33)(48 DOWNTO 1) <= x"000000004000";
  atannum(34)(48 DOWNTO 1) <= x"000000002000";
  atannum(35)(48 DOWNTO 1) <= x"000000001000";
  atannum(36)(48 DOWNTO 1) <= x"000000000800";  
  atannum(37)(48 DOWNTO 1) <= x"000000000400";
  atannum(38)(48 DOWNTO 1) <= x"000000000200";
  atannum(39)(48 DOWNTO 1) <= x"000000000100";
  
  atannum(40)(48 DOWNTO 1) <= x"000000000080";
  atannum(41)(48 DOWNTO 1) <= x"000000000040"; 
  atannum(42)(48 DOWNTO 1) <= x"000000000020";
  atannum(43)(48 DOWNTO 1) <= x"000000000010";
  atannum(44)(48 DOWNTO 1) <= x"000000000008";
  atannum(45)(48 DOWNTO 1) <= x"000000000004";
  atannum(46)(48 DOWNTO 1) <= x"000000000002";  
  atannum(47)(48 DOWNTO 1) <= x"000000000001";
  atannum(48)(48 DOWNTO 1) <= x"000000000000";
    
  pca: PROCESS (indexbit)
  BEGIN
  
    CASE indexbit IS
      WHEN '0' => arctan <= atannum(start)(48 DOWNTO 49-width);
      WHEN '1' => arctan <= atannum(start+indexpoint)(48-indexpoint DOWNTO 49-indexpoint-width);
      WHEN others => arctan <= atannum(48)(width DOWNTO 1);
    END CASE;
  
  END PROCESS;
  
END sft;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_CORDIC_M1.VHD                          ***
--***                                             ***
--***   Function: SIN and COS CORDIC with early   ***
--***   Termination Algorithm (Multiplier)        ***
--***                                             ***
--***   22/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** 1. estimates lower iterations of cordic     ***
--*** using Z value and multiplier                ***
--*** 2. multiplier at level (depth-4) for best   ***
--*** results try depth = width/2+4               ***
--***************************************************
 
ENTITY fp_cordic_m1 IS
GENERIC (
         width : positive := 36;
         depth : positive := 20;
         indexpoint : positive := 2
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      radians : IN STD_LOGIC_VECTOR (width DOWNTO 1); --'0'&[width-1:1]   
      indexbit : IN STD_LOGIC;   
      sincosbit : IN STD_LOGIC; -- 0 = cos, 1 = sin

      sincos : OUT STD_LOGIC_VECTOR (width DOWNTO 1)     
     );
END fp_cordic_m1;

ARCHITECTURE rtl of fp_cordic_m1 IS
  
  constant cordic_depth : positive := depth - 4;
  
  type datapathtype IS ARRAY (cordic_depth DOWNTO 1) OF STD_LOGIC_VECTOR (width DOWNTO 1);
  type atantype IS ARRAY (cordic_depth DOWNTO 1) OF STD_LOGIC_VECTOR (width DOWNTO 1);

  signal zerovec : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal indexpointnum, startindex : STD_LOGIC_VECTOR (4 DOWNTO 1);
  signal indexbitff : STD_LOGIC_VECTOR (cordic_depth+3 DOWNTO 1);
  signal sincosbitff : STD_LOGIC_VECTOR (cordic_depth+3 DOWNTO 1);
  signal x_start_node : STD_LOGIC_VECTOR (width DOWNTO 1);
  signal radians_load_node : STD_LOGIC_VECTOR (width DOWNTO 1);
  signal x_pipeff : datapathtype;
  signal y_pipeff : datapathtype;
  signal z_pipeff : datapathtype;
  signal x_prenode, x_prenodeone, x_prenodetwo : datapathtype;
  signal x_subnode, x_pipenode : datapathtype;
  signal y_prenode, y_prenodeone, y_prenodetwo  : datapathtype;
  signal y_subnode, y_pipenode : datapathtype;
  signal z_subnode, z_pipenode : datapathtype;
  signal atannode : atantype;

  signal multiplier_input : STD_LOGIC_VECTOR (width DOWNTO 1);
  signal multipliernode : STD_LOGIC_VECTOR (2*width DOWNTO 1);
  signal sincosff : STD_LOGIC_VECTOR (width DOWNTO 1);
  signal delay_input : STD_LOGIC_VECTOR (width DOWNTO 1);
  signal delay_pipe : STD_LOGIC_VECTOR (width DOWNTO 1);
  signal pre_estimate : STD_LOGIC_VECTOR (width DOWNTO 1);
  signal estimate : STD_LOGIC_VECTOR (width DOWNTO 1);
  signal post_estimate : STD_LOGIC_VECTOR (width DOWNTO 1);
  
  component fp_cordic_start1
  GENERIC (width : positive := 36);
  PORT (
        index : IN STD_LOGIC_VECTOR (4 DOWNTO 1);    

        value : OUT STD_LOGIC_VECTOR (width DOWNTO 1)     
       );
  end component;
   
  component fp_cordic_atan1
  GENERIC (start : positive := 32;
           width : positive := 32;
           indexpoint : positive := 1);
  PORT (
        indexbit : IN STD_LOGIC;

	      arctan : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
	    );
	end component;
	  
  component fp_sgn_mul3s
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1);

	      result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
	     );
	end component;
	
  component fp_del 
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
   end component;
    
BEGIN
 
  -- maximum width supported = 36 (width of start table)
  -- depth <= width
  -- maximum indexpoint = 10 (atan_table width - 10 > maximum width)
  gprma: IF (width > 36) GENERATE
    assert false report "maximum width is 36" severity error;
  END GENERATE;
  gprmb: IF (depth > width) GENERATE
    assert false report "depth cannot exceed (width-6)" severity error;
  END GENERATE;
  gprmc: IF (indexpoint > 10) GENERATE
    assert false report "maximum indexpoint is 10" severity error;
  END GENERATE;
     
  -- max radians = 1.57 = 01100100....
  -- max atan(2^-0)= 0.785 = 00110010.....
  -- x start (0.607) = 0010011011....

  indexpointnum <= conv_std_logic_vector (indexpoint,4);

  gipa: FOR k IN 1 TO 4 GENERATE
    startindex(k) <= indexpointnum(k) AND indexbit;
  END GENERATE;
  
  cxs: fp_cordic_start1
  GENERIC MAP (width=>width)
  PORT MAP (index=>startindex,value=>x_start_node);
  
  gra: FOR k IN 1 TO indexpoint GENERATE
    radians_load_node(k) <= (radians(k) AND NOT(indexbit));
  END GENERATE;
  grb: FOR k IN indexpoint+1 TO width GENERATE
    radians_load_node(k) <= (radians(k) AND NOT(indexbit)) OR 
                            (radians(k-indexpoint) AND indexbit);
  END GENERATE;
       
  zerovec <= x"000000000";
  
  ppa: PROCESS (sysclk,reset)
  BEGIN
  
    IF (reset = '1') THEN
        
      FOR k IN 1 TO cordic_depth+3 LOOP
        indexbitff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO cordic_depth+3 LOOP
        sincosbitff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO cordic_depth LOOP
        FOR j IN 1 TO width LOOP
          x_pipeff(k)(j) <= '0';
          y_pipeff(k)(j) <= '0';
          z_pipeff(k)(j) <= '0';
        END LOOP;
      END LOOP;
    
    ELSIF(rising_edge(sysclk)) THEN
            
      IF (enable = '1') THEN
          
        indexbitff(1) <= indexbit;
        FOR k IN 2 TO cordic_depth+3 LOOP
          indexbitff(k) <= indexbitff(k-1);
        END LOOP;
        
        sincosbitff(1) <= sincosbit;
        FOR k IN 2 TO cordic_depth+3 LOOP
          sincosbitff(k) <= sincosbitff(k-1);
        END LOOP;
        
        x_pipeff(1)(width DOWNTO 1) <= x_start_node;
        y_pipeff(1)(width DOWNTO 1) <= conv_std_logic_vector(0,width);
        z_pipeff(1)(width DOWNTO 1) <= radians_load_node;   
      
        -- z(1) always positive
        x_pipeff(2)(width DOWNTO 1) <= x_pipeff(1)(width DOWNTO 1); -- subtraction value always 0 here anyway
        y_pipeff(2)(width DOWNTO 1) <= y_pipeff(1)(width DOWNTO 1) + y_subnode(2)(width DOWNTO 1);
        z_pipeff(2)(width DOWNTO 1) <= z_pipeff(1)(width DOWNTO 1) - atannode(1)(width DOWNTO 1);
        
        FOR k IN 3 TO cordic_depth LOOP
          x_pipeff(k)(width DOWNTO 1) <= x_pipenode(k)(width DOWNTO 1);
          y_pipeff(k)(width DOWNTO 1) <= y_pipenode(k)(width DOWNTO 1);
          z_pipeff(k)(width DOWNTO 1) <= z_pipenode(k)(width DOWNTO 1);
        END LOOP;
        
      END IF;
      
    END IF;
  
  END PROCESS;
  
  gya: FOR k IN 1 TO width-indexpoint GENERATE
    y_subnode(2)(k) <= (x_pipeff(1)(k) AND NOT indexbitff(1)) OR (x_pipeff(1)(k+indexpoint) AND indexbitff(1));
  END GENERATE;
  gyb: FOR k IN (width-(indexpoint-1)) TO width GENERATE
    y_subnode(2)(k) <= (x_pipeff(1)(k) AND NOT indexbitff(1));
  END GENERATE;
  
  gpa: FOR k IN 3 TO cordic_depth GENERATE
    gpb: FOR j IN width+3-k TO width GENERATE
      x_prenodeone(k)(j) <= NOT(y_pipeff(k-1)(width));
      y_prenodeone(k)(j) <= x_pipeff(k-1)(width);
    END GENERATE;
    gpc: FOR j IN width+3-indexpoint-k TO width GENERATE
      x_prenodetwo(k)(j) <= NOT(y_pipeff(k-1)(width));
      y_prenodetwo(k)(j) <= x_pipeff(k-1)(width);
    END GENERATE;
    gpd: FOR j IN 1 TO width+2-k GENERATE
      x_prenodeone(k)(j) <= NOT(y_pipeff(k-1)(j+k-2));
      y_prenodeone(k)(j) <= x_pipeff(k-1)(j+k-2);
    END GENERATE;
    gpe: FOR j IN 1 TO width+2-indexpoint-k GENERATE
      x_prenodetwo(k)(j) <= NOT(y_pipeff(k-1)(j+k-2+indexpoint));
      y_prenodetwo(k)(j) <= x_pipeff(k-1)(j+k-2+indexpoint);
    END GENERATE;
    
    gpf: FOR j IN 1 TO width GENERATE
      x_prenode(k)(j) <= (x_prenodeone(k)(j) AND NOT(indexbitff(k-1))) OR 
                         (x_prenodetwo(k)(j) AND indexbitff(k-1));
      y_prenode(k)(j) <= (y_prenodeone(k)(j) AND NOT(indexbitff(k-1))) OR 
                         (y_prenodetwo(k)(j) AND indexbitff(k-1));
    END GENERATE;
    
    gpg: FOR j IN 1 TO width GENERATE
      x_subnode(k)(j) <= x_prenode(k)(j) XOR z_pipeff(k-1)(width);
      y_subnode(k)(j) <= y_prenode(k)(j) XOR z_pipeff(k-1)(width);
      z_subnode(k)(j) <= NOT(atannode(k-1)(j)) XOR z_pipeff(k-1)(width);
    END GENERATE;

    x_pipenode(k)(width DOWNTO 1) <= x_pipeff(k-1)(width DOWNTO 1) + 
                                     x_subnode(k)(width DOWNTO 1) + z_pipeff(k-1)(width);
                                     
    y_pipenode(k)(width DOWNTO 1) <= y_pipeff(k-1)(width DOWNTO 1) + 
                                     y_subnode(k)(width DOWNTO 1) + z_pipeff(k-1)(width);
                                     
    z_pipenode(k)(width DOWNTO 1) <= z_pipeff(k-1)(width DOWNTO 1) + 
                                     z_subnode(k)(width DOWNTO 1) + z_pipeff(k-1)(width);

  END GENERATE;
  
  gata: FOR k IN 1 TO cordic_depth GENERATE
    cata: fp_cordic_atan1
    GENERIC MAP (start=>k,width=>width,indexpoint=>indexpoint)
    PORT MAP (indexbit=>indexbitff(k),arctan=>atannode(k)(width DOWNTO 1));
  END GENERATE;
	
	gma: FOR k IN 1 TO width GENERATE
	  multiplier_input(k) <= (x_pipeff(cordic_depth)(k) AND sincosbitff(cordic_depth)) OR
	                         (y_pipeff(cordic_depth)(k) AND NOT(sincosbitff(cordic_depth)));
	  delay_input(k) <= (x_pipeff(cordic_depth)(k) AND NOT(sincosbitff(cordic_depth))) OR
	                    (y_pipeff(cordic_depth)(k) AND sincosbitff(cordic_depth));
	END GENERATE;
  
  cmx: fp_sgn_mul3s
  GENERIC MAP (widthaa=>width,widthbb=>width,widthcc=>2*width)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>multiplier_input,
            databb=>z_pipeff(cordic_depth)(width DOWNTO 1),
            result=>multipliernode);
	
  pma: PROCESS (sysclk,reset)
  BEGIN
    IF (reset = '1') THEN
      FOR k IN 1 TO width LOOP
        sincosff(k) <= '0';
      END LOOP;
    ELSIF(rising_edge(sysclk)) THEN
      IF (enable = '1') THEN     
        sincosff <= delay_pipe + post_estimate + NOT(sincosbitff(cordic_depth+3));
      END IF; 
    END IF;  
  END PROCESS;
  
  pre_estimate <= multipliernode(2*width-2 DOWNTO width-1);
  gea: FOR k IN 1 TO width-indexpoint GENERATE
    estimate(k) <= (pre_estimate(k) AND NOT(indexbitff(cordic_depth+3))) OR
                   (pre_estimate(k+indexpoint) AND indexbitff(cordic_depth+3));
  END GENERATE;
  geb: FOR k IN width-indexpoint+1 TO width GENERATE
    estimate(k) <= (pre_estimate(k) AND NOT(indexbitff(cordic_depth+3))) OR
                   (pre_estimate(width) AND indexbitff(cordic_depth+3));
  END GENERATE;
  -- add estimate for sin, subtract for cos
  gec: FOR k IN 1 TO width GENERATE
    post_estimate(k) <= estimate(k) XOR NOT(sincosbitff(cordic_depth+3));
  END GENERATE;
  
  cda: fp_del
  GENERIC MAP (width=>width,pipes=>3)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>delay_input,
            cc=>delay_pipe);

  sincos <= sincosff;
      
END rtl;
LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_CORDIC_START1.VHD                      ***
--***                                             ***
--***   Function: Table for Initial Value of X    ***
--***   for SIN and COS CORDIC Core               ***
--***                                             ***
--***   22/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_cordic_start1 IS
GENERIC (width : positive := 36);
PORT (
      index : IN STD_LOGIC_VECTOR (4 DOWNTO 1);    

      value : OUT STD_LOGIC_VECTOR (width DOWNTO 1)     
     );
END fp_cordic_start1;

ARCHITECTURE rtl of fp_cordic_start1 IS

  signal valuenode : STD_LOGIC_VECTOR (36 DOWNTO 1);
  
BEGIN

  pva: PROCESS (index)
  BEGIN
   
    CASE index IS
      WHEN "0000" => valuenode <= x"26DD3B6A1";
      WHEN "0001" => valuenode <= x"36F656C5A";
      WHEN "0010" => valuenode <= x"3D731DFFB";
      WHEN "0011" => valuenode <= x"3F5743B24";
      WHEN "0100" => valuenode <= x"3FD574860";
      WHEN "0101" => valuenode <= x"3FF557499";
      WHEN "0110" => valuenode <= x"3FFD5574A";
      WHEN "0111" => valuenode <= x"3FFF55575";
      WHEN "1000" => valuenode <= x"3FFFD5557";
      WHEN "1001" => valuenode <= x"3FFFF5555";
      WHEN "1010" => valuenode <= x"3FFFFD555";
      WHEN "1011" => valuenode <= x"3FFFFF555";
      WHEN "1101" => valuenode <= x"3FFFFFD55";
      WHEN "1100" => valuenode <= x"3FFFFFF55";
      WHEN "1111" => valuenode <= x"3FFFFFFD5";
      WHEN "1110" => valuenode <= x"3FFFFFFF5";
      WHEN others => valuenode <= x"000000000";
    END CASE;

  END PROCESS;
  
  value <= valuenode (36 DOWNTO 37-width);
  
END rtl;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_COS1.VHD                               ***
--***                                             ***
--***   Function: Single Precision COS Core       ***
--***                                             ***
--***   10/01/10 ML                               ***
--***                                             ***
--***   (c) 2010 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** 1. Input < 0.5 radians, take sin(pi/2-input)***
--*** 2. latency = depth + range_depth (11) + 6   ***
--*** (1 less than sin)                           ***
--***************************************************

ENTITY fp_cos IS
GENERIC (
          device : integer := 0;
          width : positive := 36;
          depth : positive := 20;
          indexpoint : positive := 2
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (8 DOWNTO 1); 
      mantissain : IN STD_LOGIC_VECTOR (23 DOWNTO 1); 

      signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (8 DOWNTO 1); 
      mantissaout : OUT STD_LOGIC_VECTOR (23 DOWNTO 1) 
     );
END fp_cos;

ARCHITECTURE rtl of fp_cos IS

  constant cordic_width : positive := width;
  constant cordic_depth : positive := depth;
  constant range_depth : positive := 11;

  signal piovertwo : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal zerovec : STD_LOGIC_VECTOR (36 DOWNTO 1);

  -- range reduction
  signal circle : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal negcircle : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal quadrantsign, quadrantselect : STD_LOGIC;
  signal positive_quadrant, negative_quadrant : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal fraction_quadrant : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal one_term : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal quadrant : STD_LOGIC_VECTOR (34 DOWNTO 1);
  
  -- circle to radians mult
  signal radiansnode : STD_LOGIC_VECTOR (cordic_width DOWNTO 1);
  signal indexcheck : STD_LOGIC_VECTOR (16 DOWNTO 1);
  signal indexbit : STD_LOGIC;
  
  signal signinff : STD_LOGIC_VECTOR (range_depth DOWNTO 1);
  signal selectoutputff : STD_LOGIC_VECTOR (range_depth+cordic_depth+5 DOWNTO 1);
  signal signcalcff : STD_LOGIC_VECTOR (cordic_depth+6 DOWNTO 1);
  signal quadrant_sumff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal select_sincosff : STD_LOGIC_VECTOR (4 DOWNTO 1);

  signal fixed_sincos : STD_LOGIC_VECTOR (cordic_width DOWNTO 1);
  signal fixed_sincosnode : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal fixed_sincosff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  
  signal countnode : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal countff : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal mantissanormnode : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal mantissanormff : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal exponentnormnode : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal exponentnormff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal overflownode : STD_LOGIC_VECTOR (24 DOWNTO 1);
 
  component fp_range1
  GENERIC (device : integer);
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        signin : IN STD_LOGIC;
        exponentin : IN STD_LOGIC_VECTOR (8 DOWNTO 1); 
        mantissain : IN STD_LOGIC_VECTOR (23 DOWNTO 1); 

        circle : OUT STD_LOGIC_VECTOR (36 DOWNTO 1);
        negcircle : OUT STD_LOGIC_VECTOR (36 DOWNTO 1) 
       );
  end component;
   
  component fp_cordic_m1
  GENERIC (
         width : positive := 36;
         depth : positive := 20;
         indexpoint : positive := 2
        );  
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        radians : IN STD_LOGIC_VECTOR (width DOWNTO 1); --'0'&[width-1:1]   
        indexbit : IN STD_LOGIC;   
        sincosbit : IN STD_LOGIC;

        sincos : OUT STD_LOGIC_VECTOR (width DOWNTO 1)     
       );
  end component;
    
  component fp_clz36 IS
  PORT (
        mantissa : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
      
        leading : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
       );
  end component;

  component fp_lsft36 IS 
  PORT (
        inbus : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);

         outbus : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
        );
    end component;

  component fp_fxmul
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36;
           pipes : positive := 1;
           accuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1); 
      
        result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
       );
  end component;
   
  component fp_del IS
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
   end component;
   
  BEGIN
    
    -- pi/2 = 1.57
    piovertwo <= x"c90fdaa22";
  
    zerovec <= x"000000000";
                  
    --*** RANGE REDUCTION ***
    crr: fp_range1
    GENERIC MAP(device=>device)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              signin=>signin,exponentin=>exponentin,mantissain=>mantissain,
              circle=>circle,negcircle=>negcircle); 

    quadrantsign <= (NOT(circle(36)) AND circle(35)) OR
                    (circle(36) AND NOT(circle(35))); -- cos negative in quadrants 2&3
    
    quadrantselect <= circle(35); -- cos (1-x) in quadants 2&4
    
    gra: FOR k IN 1 TO 34 GENERATE
      quadrant(k) <= (circle(k) AND NOT(quadrantselect)) OR
                     (negcircle(k) AND quadrantselect);
    END GENERATE;   
    
    -- if quadrant >0.5 (when quadrant(34) = 1), use quadrant, else use 1-quadrant, and take sin rather than cos
    -- do this to maximize input value, not output value
    positive_quadrant <= '0' & quadrant & '0';
    gnqa: FOR k IN 1 TO 36 GENERATE
      negative_quadrant(k) <= NOT(positive_quadrant(k));
      fraction_quadrant(k) <= (positive_quadrant(k) AND quadrant(34)) OR
                              (negative_quadrant(k) AND NOT(quadrant(34)));
    END GENERATE;

    one_term <= NOT(quadrant(34)) & zerovec(35 DOWNTO 1); -- 0 if positive quadrant
      
    pfa: PROCESS (sysclk,reset)
    BEGIN        
      IF (reset = '1') THEN
          
        FOR k IN 1 TO range_depth LOOP
          signinff(k) <= '0';
        END LOOP;
        FOR k IN 1 TO cordic_depth+6 LOOP
          signcalcff(k) <= '0';
        END LOOP;
        FOR k IN 1 TO 36 LOOP
          quadrant_sumff(k) <= '0';
        END LOOP;
        FOR k IN 1 TO 4 LOOP
          select_sincosff(k) <= '0';
        END LOOP;
 
      ELSIF (rising_edge(sysclk)) THEN
         
        IF (enable = '1') THEN
        
          signinff(1) <= signin;
          FOR k IN 2 TO range_depth LOOP
            signinff(k) <= signinff(k-1);
          END LOOP;
          -- level range_depth+1 to range_depth+cordic_depth+6
          signcalcff(1) <= quadrantsign; 
          FOR k IN 2 TO cordic_depth+6 LOOP
            signcalcff(k) <= signcalcff(k-1);
          END LOOP;
          
          -- range 0-0.9999
          quadrant_sumff <= one_term + fraction_quadrant + quadrant(34); -- level range_depth+1
          
          -- level range depth+1 to range_depth+4 
          select_sincosff(1) <= NOT(quadrant(34));
          FOR k IN 2 TO 4 LOOP
            select_sincosff(k) <= select_sincosff(k-1);
          END LOOP;
   
        END IF;
         
      END IF;
        
    END PROCESS;

    -- levels range_depth+2,3,4
    cmul: fp_fxmul  
    GENERIC MAP (widthaa=>36,widthbb=>36,widthcc=>cordic_width,
                 pipes=>3,synthesize=>1)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              dataaa=>quadrant_sumff,databb=>piovertwo,
              result=>radiansnode);
                    
    indexcheck(1) <= radiansnode(cordic_width-1);
    gica: FOR k IN 2 TO 16 GENERATE
      indexcheck(k) <= indexcheck(k-1) OR radiansnode(cordic_width-k);
    END GENERATE;
    -- for safety, give an extra bit of space
    indexbit <= NOT(indexcheck(indexpoint+1));
   
    ccc: fp_cordic_m1
    GENERIC MAP (width=>cordic_width,depth=>cordic_depth,indexpoint=>indexpoint)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              radians=>radiansnode,
              indexbit=>indexbit,
              sincosbit=>select_sincosff(4),
              sincos=>fixed_sincos);
   
    gfxa: IF (width < 36) GENERATE
      fixed_sincosnode <= fixed_sincos & zerovec(36-width DOWNTO 1);
    END GENERATE;
    gfxb: IF (width = 36) GENERATE
      fixed_sincosnode <= fixed_sincos;
    END GENERATE;
    
    clz: fp_clz36
    PORT MAP (mantissa=>fixed_sincosnode,leading=>countnode);
        
    sft: fp_lsft36  
    PORT MAP (inbus=>fixed_sincosff,shift=>countff,
              outbus=>mantissanormnode);
    
    -- maximum sin or cos = 1.0 = 1.0e127 single precision
    -- 1e128 - 1 (leading one) gives correct number
    exponentnormnode <= "10000000" - ("00" & countff); 
    
    overflownode(1) <= mantissanormnode(12);
    gova: FOR k IN 2 TO 24 GENERATE
      overflownode(k) <= mantissanormnode(k+11) AND overflownode(k-1);
    END GENERATE;
    
    -- OUTPUT
    poa: PROCESS (sysclk,reset)
    BEGIN
        
      IF (reset = '1') THEN
          
        FOR k IN 1 TO 36 LOOP
          fixed_sincosff(k) <= '0';
        END LOOP;
        countff <= "000000";
        FOR k IN 1 TO 23 LOOP
          mantissanormff(k) <= '0';
        END LOOP;
        FOR k IN 1 TO 8 LOOP
          exponentnormff(k) <= '0';
        END LOOP;

      ELSIF (rising_edge(sysclk)) THEN
          
        IF (enable = '1') THEN
           
          fixed_sincosff <= fixed_sincosnode; -- level range_depth+cordic_depth+5
          countff <= countnode; -- level range_depth+4+cordic_depth+5

          -- level range_depth+cordic_depth+6
          mantissanormff <= mantissanormnode(35 DOWNTO 13) + mantissanormnode(12);
          exponentnormff <= exponentnormnode(8 DOWNTO 1) + overflownode(24);
          
        END IF;
        
      END IF;
      
    END PROCESS;
    
    mantissaout <= mantissanormff; 
    exponentout <= exponentnormff;
    signout <= signcalcff(cordic_depth+6);    
    
  END rtl;
  
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_DEL.VHD                                ***
--***                                             ***
--***   Function: Generic Bus Delay               ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_del IS 
GENERIC (
         width : positive := 64;
         pipes : positive := 1
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      
      cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
     );
END fp_del;

ARCHITECTURE rtl OF fp_del IS

  component fp_del_one IS 
  GENERIC (width : positive := 64);
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
   end component;
   
  component fp_del_var IS 
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
   end component;
 
            
BEGIN

  genone: IF (pipes = 1) GENERATE
  
    delone: fp_del_one
    GENERIC MAP (width=>width)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>aa,cc=>cc);
              
  END GENERATE;
            
  genvar: IF (pipes > 1) GENERATE
  
    delvar: fp_del_var
    GENERIC MAP (width=>width,pipes=>pipes)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>aa,cc=>cc);
              
  END GENERATE;            
            
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_DEL_ONE.VHD                            ***
--***                                             ***
--***   Function: Single Block Bus Delay          ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_del_one IS 
GENERIC (width : positive := 64);
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      
      cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
     );
END fp_del_one ;

ARCHITECTURE rtl OF fp_del_one  IS

  signal delff : STD_LOGIC_VECTOR (width DOWNTO 1);
            
BEGIN

  pda: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN

      FOR k IN 1 TO width LOOP
        delff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN
        delff(width DOWNTO 1) <= aa;
      END IF;
    
    END IF;
      
  END PROCESS;
    
  cc <= delff(width DOWNTO 1);
    
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_DEL.VHD                                ***
--***                                             ***
--***   Function: Multiple Clock Bus Delay        ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_del_var IS 
GENERIC (
         width : positive := 64;
         pipes : positive := 1
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      
      cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
     );
END fp_del_var ;

ARCHITECTURE rtl OF fp_del_var  IS

  type delfftype IS ARRAY (pipes DOWNTO 1) OF STD_LOGIC_VECTOR (width DOWNTO 1);

  signal delff : delfftype;
            
BEGIN

  pda: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN

      FOR k IN 1 TO pipes LOOP
        FOR j IN 1 TO width LOOP
          delff(k)(j) <= '0';
        END LOOP;
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN
        delff(1)(width DOWNTO 1) <= aa;
        FOR k IN 2 TO pipes LOOP
          delff(k)(width DOWNTO 1) <= delff(k-1)(width DOWNTO 1);
        END LOOP;
      END IF;
    
    END IF;
      
  END PROCESS;
    
  cc <= delff(pipes)(width DOWNTO 1);
    
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_DELBIT.VHD                             ***
--***                                             ***
--***   Function: Generic Bit Delay               ***
--***                                             ***
--***   01/12/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_delbit IS 
GENERIC (
         pipes : positive := 1
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      aa : IN STD_LOGIC; 
      
      cc : OUT STD_LOGIC
     );
END fp_delbit;

ARCHITECTURE rtl OF fp_delbit IS

  component fp_delbit_one IS 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC; 
      
        cc : OUT STD_LOGIC
       );
   end component;
   
  component fp_delbit_var IS 
  GENERIC (
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC; 
      
        cc : OUT STD_LOGIC
       );
   end component;
 
            
BEGIN

  genone: IF (pipes = 1) GENERATE
  
    delone: fp_delbit_one
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>aa,cc=>cc);
              
  END GENERATE;
            
  genvar: IF (pipes > 1) GENERATE
  
    delvar: fp_delbit_var
    GENERIC MAP (pipes=>pipes)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>aa,cc=>cc);
              
  END GENERATE;            
            
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_DELBIT_ONE.VHD                         ***
--***                                             ***
--***   Function: Single Bit Delay                ***
--***                                             ***
--***   01/12/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_delbit_one IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      aa : IN STD_LOGIC; 
      
      cc : OUT STD_LOGIC
     );
END fp_delbit_one ;

ARCHITECTURE rtl OF fp_delbit_one  IS

  signal delff : STD_LOGIC;
            
BEGIN

  pda: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN

      delff <= '0';
      
    ELSIF (rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN
        delff <= aa;
      END IF;
    
    END IF;
      
  END PROCESS;
    
  cc <= delff;
    
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_DELBIT_VAR.VHD                         ***
--***                                             ***
--***   Function: Multiple Bit Delay              ***
--***                                             ***
--***   01/12/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_delbit_var IS 
GENERIC (
         pipes : positive := 1
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      aa : IN STD_LOGIC; 
      
      cc : OUT STD_LOGIC
     );
END fp_delbit_var ;

ARCHITECTURE rtl OF fp_delbit_var  IS

  signal delff : STD_LOGIC_VECTOR (pipes DOWNTO 1);
            
BEGIN

  pda: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN

      FOR k IN 1 TO pipes LOOP
        delff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN
        delff(1) <= aa;
        FOR k IN 2 TO pipes LOOP
          delff(k) <= delff(k-1);
        END LOOP;
      END IF;
    
    END IF;
      
  END PROCESS;
    
  cc <= delff(pipes);
    
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   SINGLE PRECISION DIVIDER - CORE           ***
--***                                             ***
--***   FP_DIV_CORE.VHD                           ***
--***                                             ***
--***   Function: Fixed Point 36 Bit Divider      ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** Latency = 13                                ***
--***************************************************

ENTITY fp_div_core IS 
GENERIC (synthesize : integer := 1);
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      dividend : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
      divisor : IN STD_LOGIC_VECTOR (36 DOWNTO 1);

		quotient : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
		);
END fp_div_core;

ARCHITECTURE rtl OF fp_div_core IS

  signal zerovec : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal guess : STD_LOGIC_VECTOR (18 DOWNTO 1);         
  signal dividenddel : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal divisordel : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal scaledivisor : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal scaledividend : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal nextguessnode : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal nextguessff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal scaledividendff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal quotientnode : STD_LOGIC_VECTOR (72 DOWNTO 1);
  
  signal leadone, leadzip, leader : STD_LOGIC;
  
  component fp_div_est IS 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        divisor : IN STD_LOGIC_VECTOR (19 DOWNTO 1);

		  invdivisor : OUT STD_LOGIC_VECTOR (18 DOWNTO 1)
		  );
  end component;
  
  component fp_del
  GENERIC (
           width : positive := 64;
           pipes : positive := 2
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
       
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
   end component;  
   
  component fp_fxmul 
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36;
           pipes : positive := 1;
           accuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1); 
      
        result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
       );
  end component;
   
BEGIN
  
  gza: FOR k IN 1 TO 36 GENERATE
    zerovec(k) <= '0';
  END GENERATE;

  estcore: fp_div_est
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            divisor=>divisor(36 DOWNTO 18),invdivisor=>guess);

  deltop: fp_del
  GENERIC MAP (width=>36,pipes=>5)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>dividend,cc=>dividenddel);
            
  delbot: fp_del
  GENERIC MAP (width=>36,pipes=>5)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>divisor,cc=>divisordel);
   
  ppa: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN
        
      FOR k IN 1 TO 36 LOOP
        nextguessff(k) <= '0';
        scaledividendff(k) <= '0';
      END LOOP;
         
    ELSIF (rising_edge(sysclk)) THEN
    
      IF (enable = '1') THEN
          
        nextguessff <= nextguessnode;
        scaledividendff <= scaledividend;
 
      END IF;
         
    END IF;
  
  END PROCESS;
  
  leadone <= nextguessff(35) AND nextguessff(34) AND nextguessff(33) AND 
             nextguessff(32) AND nextguessff(31) AND nextguessff(30) AND nextguessff(29) AND 
             nextguessff(28) AND nextguessff(27) AND nextguessff(26) AND nextguessff(25) AND 
             nextguessff(24) AND nextguessff(23) AND nextguessff(22) AND nextguessff(21) AND 
             nextguessff(20) AND nextguessff(19);-- AND nextguessff(18);
  
  leadzip <= NOT(nextguessff(35) OR nextguessff(34) OR nextguessff(33) OR 
                 nextguessff(32) OR nextguessff(31) OR nextguessff(30) OR nextguessff(29) OR 
                 nextguessff(28) OR nextguessff(27) OR nextguessff(26) OR nextguessff(25) OR 
                 nextguessff(24) OR nextguessff(23) OR nextguessff(22) OR nextguessff(21) OR 
                 nextguessff(20) OR nextguessff(19));-- OR nextguessff(18));
                 
  leader <= leadone XOR leadzip;
            
  -- 36 * 18, magnitude will be very close to 1 (1.00..00XXX or 0.11..11XXX)
  mulone: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>18,widthcc=>36,pipes=>3,
               synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>divisordel,databb=>guess,
            result=>scaledivisor);            
        
  -- 36 * 18, as 1<divisor<2 and 1<dividend<1 and 0.5<guess<1, 0.5<scaledividend<2
  multwo: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>18,widthcc=>36,pipes=>3,
               synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>dividenddel,databb=>guess,
            result=>scaledividend); 

  -- 2.0 - about 1 = about 1 (1.00..00XXX or 0.11..11XXX)
  --nextguessnode <= ("10" & zerovec(35 DOWNTO 1)) - ('0' & scaledivisor);
  
  nextguessnode(20 DOWNTO 1) <= zerovec(20 DOWNTO 1) - scaledivisor(20 DOWNTO 1);
  gng: FOR k IN 21 TO 35 GENERATE
    nextguessnode(k) <= scaledivisor(36);
  END GENERATE;
  nextguessnode(36) <= scaledivisor(35);

  multthr: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>36,widthcc=>72,pipes=>3,
               synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>scaledividendff,databb=>nextguessff,
            result=>quotientnode); 
         
  quotient <= quotientnode(71 DOWNTO 36);

END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_DIV_EST.VHD                            ***
--***                                             ***
--***   Function: Estimates 18 Bit Inverse        ***
--***                                             ***
--***   Used by both single and double dividers   ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** 1. Inverse of 18 bit header                 ***
--*** (not including leading '1')                 ***
--*** 2. Uses 20 bit precision tables - 18 bits   ***
--*** drops a bit occasionally                    ***
--***************************************************

ENTITY fp_div_est IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      divisor : IN STD_LOGIC_VECTOR (19 DOWNTO 1);

		invdivisor : OUT STD_LOGIC_VECTOR (18 DOWNTO 1)
		);
END fp_div_est;

ARCHITECTURE rtl OF fp_div_est IS

  type twodelfftype IS ARRAY (2 DOWNTO 1) OF STD_LOGIC_VECTOR (9 DOWNTO 1);
  type ziplutdelfftype IS ARRAY (2 DOWNTO 1) OF STD_LOGIC_VECTOR (20 DOWNTO 1);
  
  signal zerovec : STD_LOGIC_VECTOR (17 DOWNTO 1);
  signal one, two : STD_LOGIC_VECTOR (9 DOWNTO 1);
  signal oneaddff, zipaddff : STD_LOGIC_VECTOR (9 DOWNTO 1);
  signal onelut, onelutff : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal ziplut, ziplutff : STD_LOGIC_VECTOR (20 DOWNTO 1);
  signal onetwo : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal twodelff : twodelfftype;
  signal ziplutdelff : ziplutdelfftype;
  signal invdivisorff : STD_LOGIC_VECTOR (20 DOWNTO 1);
         
  component fp_div_lut1 IS
  PORT (
        add : IN STD_LOGIC_VECTOR (9 DOWNTO 1);
		  data : OUT STD_LOGIC_VECTOR (11 DOWNTO 1)
       );
  end component;
    
  component fp_div_lut0 IS
  PORT (
        add : IN STD_LOGIC_VECTOR (9 DOWNTO 1);
		  data : OUT STD_LOGIC_VECTOR (20 DOWNTO 1)
       );
  end component;
  
  component fp_fxmul  
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36;
           pipes : positive := 1;
           accuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1); 
      
        result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
       );
  end component; 
    
BEGIN
  
  gza: FOR k IN 1 TO 17 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  one <= divisor(18 DOWNTO 10);
  two <= divisor(9 DOWNTO 1);
  
  -- these register seperate to make the LUTs into memories
  pma: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN

      FOR k IN 1 TO 9 LOOP
        oneaddff(k) <= '0';
        zipaddff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 11 LOOP
        onelutff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 20 LOOP
        ziplutff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN
        oneaddff <= one;
        zipaddff <= one;
        onelutff <= onelut;
        ziplutff <= ziplut;
      END IF;
    
    END IF;
      
  END PROCESS;
    
  upper: fp_div_lut1 PORT MAP (add=>oneaddff,data=>onelut);
  
  lower: fp_div_lut0 PORT MAP (add=>zipaddff,data=>ziplut);
  
  pra: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN

      FOR k IN 1 TO 2 LOOP
        FOR j IN 1 TO 9 LOOP
          twodelff(k)(j) <= '0';
        END LOOP;
      END LOOP;
      FOR k IN 1 TO 2 LOOP
        FOR j IN 1 TO 9 LOOP
          ziplutdelff(k)(j) <= '0';
        END LOOP;
      END LOOP;
      FOR k IN 1 TO 20 LOOP
        invdivisorff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN
          
        twodelff(1)(9 DOWNTO 1) <= two;
        twodelff(2)(9 DOWNTO 1) <= twodelff(1)(9 DOWNTO 1);
        
        ziplutdelff(1)(20 DOWNTO 1) <= ziplutff;
        ziplutdelff(2)(20 DOWNTO 1) <= ziplutdelff(1)(20 DOWNTO 1);
        
        invdivisorff <= ziplutdelff(2)(20 DOWNTO 1) - 
                       (zerovec(9 DOWNTO 1) & onetwo);
        
      END IF;
    
    END IF;
      
  END PROCESS;
 
  mulcore: fp_fxmul
  GENERIC MAP (widthaa=>11,widthbb=>9,widthcc=>11,pipes=>2)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>onelutff,databb=>twodelff(2)(9 DOWNTO 1),
            result=>onetwo);
  
  invdivisor <= invdivisorff(20 DOWNTO 3);
    
END rtl;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_DIV_LUT0.VHD                           ***
--***                                             ***
--***   Function: Look Up Table - Inverse         ***
--***                                             ***
--***   Generated by MATLAB Utility               ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_div_lut0 IS
PORT (
      add : IN STD_LOGIC_VECTOR (9 DOWNTO 1);
		data : OUT STD_LOGIC_VECTOR (20 DOWNTO 1)
);
END fp_div_lut0;

ARCHITECTURE rtl OF fp_div_lut0 IS

BEGIN

  pca: PROCESS (add)
  BEGIN
    CASE add IS
      WHEN "000000000" => data <= conv_std_logic_vector(1048575,20);
      WHEN "000000001" => data <= conv_std_logic_vector(1046531,20);
      WHEN "000000010" => data <= conv_std_logic_vector(1044495,20);
      WHEN "000000011" => data <= conv_std_logic_vector(1042467,20);
      WHEN "000000100" => data <= conv_std_logic_vector(1040447,20);
      WHEN "000000101" => data <= conv_std_logic_vector(1038434,20);
      WHEN "000000110" => data <= conv_std_logic_vector(1036429,20);
      WHEN "000000111" => data <= conv_std_logic_vector(1034432,20);
      WHEN "000001000" => data <= conv_std_logic_vector(1032443,20);
      WHEN "000001001" => data <= conv_std_logic_vector(1030461,20);
      WHEN "000001010" => data <= conv_std_logic_vector(1028487,20);
      WHEN "000001011" => data <= conv_std_logic_vector(1026521,20);
      WHEN "000001100" => data <= conv_std_logic_vector(1024562,20);
      WHEN "000001101" => data <= conv_std_logic_vector(1022610,20);
      WHEN "000001110" => data <= conv_std_logic_vector(1020666,20);
      WHEN "000001111" => data <= conv_std_logic_vector(1018729,20);
      WHEN "000010000" => data <= conv_std_logic_vector(1016800,20);
      WHEN "000010001" => data <= conv_std_logic_vector(1014878,20);
      WHEN "000010010" => data <= conv_std_logic_vector(1012963,20);
      WHEN "000010011" => data <= conv_std_logic_vector(1011055,20);
      WHEN "000010100" => data <= conv_std_logic_vector(1009155,20);
      WHEN "000010101" => data <= conv_std_logic_vector(1007262,20);
      WHEN "000010110" => data <= conv_std_logic_vector(1005375,20);
      WHEN "000010111" => data <= conv_std_logic_vector(1003496,20);
      WHEN "000011000" => data <= conv_std_logic_vector(1001624,20);
      WHEN "000011001" => data <= conv_std_logic_vector(999759,20);
      WHEN "000011010" => data <= conv_std_logic_vector(997900,20);
      WHEN "000011011" => data <= conv_std_logic_vector(996049,20);
      WHEN "000011100" => data <= conv_std_logic_vector(994205,20);
      WHEN "000011101" => data <= conv_std_logic_vector(992367,20);
      WHEN "000011110" => data <= conv_std_logic_vector(990536,20);
      WHEN "000011111" => data <= conv_std_logic_vector(988712,20);
      WHEN "000100000" => data <= conv_std_logic_vector(986894,20);
      WHEN "000100001" => data <= conv_std_logic_vector(985083,20);
      WHEN "000100010" => data <= conv_std_logic_vector(983279,20);
      WHEN "000100011" => data <= conv_std_logic_vector(981482,20);
      WHEN "000100100" => data <= conv_std_logic_vector(979691,20);
      WHEN "000100101" => data <= conv_std_logic_vector(977906,20);
      WHEN "000100110" => data <= conv_std_logic_vector(976128,20);
      WHEN "000100111" => data <= conv_std_logic_vector(974357,20);
      WHEN "000101000" => data <= conv_std_logic_vector(972591,20);
      WHEN "000101001" => data <= conv_std_logic_vector(970833,20);
      WHEN "000101010" => data <= conv_std_logic_vector(969080,20);
      WHEN "000101011" => data <= conv_std_logic_vector(967334,20);
      WHEN "000101100" => data <= conv_std_logic_vector(965594,20);
      WHEN "000101101" => data <= conv_std_logic_vector(963861,20);
      WHEN "000101110" => data <= conv_std_logic_vector(962133,20);
      WHEN "000101111" => data <= conv_std_logic_vector(960412,20);
      WHEN "000110000" => data <= conv_std_logic_vector(958697,20);
      WHEN "000110001" => data <= conv_std_logic_vector(956988,20);
      WHEN "000110010" => data <= conv_std_logic_vector(955286,20);
      WHEN "000110011" => data <= conv_std_logic_vector(953589,20);
      WHEN "000110100" => data <= conv_std_logic_vector(951898,20);
      WHEN "000110101" => data <= conv_std_logic_vector(950213,20);
      WHEN "000110110" => data <= conv_std_logic_vector(948534,20);
      WHEN "000110111" => data <= conv_std_logic_vector(946862,20);
      WHEN "000111000" => data <= conv_std_logic_vector(945195,20);
      WHEN "000111001" => data <= conv_std_logic_vector(943533,20);
      WHEN "000111010" => data <= conv_std_logic_vector(941878,20);
      WHEN "000111011" => data <= conv_std_logic_vector(940229,20);
      WHEN "000111100" => data <= conv_std_logic_vector(938585,20);
      WHEN "000111101" => data <= conv_std_logic_vector(936947,20);
      WHEN "000111110" => data <= conv_std_logic_vector(935314,20);
      WHEN "000111111" => data <= conv_std_logic_vector(933688,20);
      WHEN "001000000" => data <= conv_std_logic_vector(932067,20);
      WHEN "001000001" => data <= conv_std_logic_vector(930451,20);
      WHEN "001000010" => data <= conv_std_logic_vector(928842,20);
      WHEN "001000011" => data <= conv_std_logic_vector(927237,20);
      WHEN "001000100" => data <= conv_std_logic_vector(925639,20);
      WHEN "001000101" => data <= conv_std_logic_vector(924046,20);
      WHEN "001000110" => data <= conv_std_logic_vector(922458,20);
      WHEN "001000111" => data <= conv_std_logic_vector(920876,20);
      WHEN "001001000" => data <= conv_std_logic_vector(919299,20);
      WHEN "001001001" => data <= conv_std_logic_vector(917727,20);
      WHEN "001001010" => data <= conv_std_logic_vector(916161,20);
      WHEN "001001011" => data <= conv_std_logic_vector(914601,20);
      WHEN "001001100" => data <= conv_std_logic_vector(913045,20);
      WHEN "001001101" => data <= conv_std_logic_vector(911495,20);
      WHEN "001001110" => data <= conv_std_logic_vector(909950,20);
      WHEN "001001111" => data <= conv_std_logic_vector(908410,20);
      WHEN "001010000" => data <= conv_std_logic_vector(906876,20);
      WHEN "001010001" => data <= conv_std_logic_vector(905347,20);
      WHEN "001010010" => data <= conv_std_logic_vector(903822,20);
      WHEN "001010011" => data <= conv_std_logic_vector(902303,20);
      WHEN "001010100" => data <= conv_std_logic_vector(900789,20);
      WHEN "001010101" => data <= conv_std_logic_vector(899281,20);
      WHEN "001010110" => data <= conv_std_logic_vector(897777,20);
      WHEN "001010111" => data <= conv_std_logic_vector(896278,20);
      WHEN "001011000" => data <= conv_std_logic_vector(894784,20);
      WHEN "001011001" => data <= conv_std_logic_vector(893295,20);
      WHEN "001011010" => data <= conv_std_logic_vector(891812,20);
      WHEN "001011011" => data <= conv_std_logic_vector(890333,20);
      WHEN "001011100" => data <= conv_std_logic_vector(888859,20);
      WHEN "001011101" => data <= conv_std_logic_vector(887389,20);
      WHEN "001011110" => data <= conv_std_logic_vector(885925,20);
      WHEN "001011111" => data <= conv_std_logic_vector(884465,20);
      WHEN "001100000" => data <= conv_std_logic_vector(883011,20);
      WHEN "001100001" => data <= conv_std_logic_vector(881561,20);
      WHEN "001100010" => data <= conv_std_logic_vector(880116,20);
      WHEN "001100011" => data <= conv_std_logic_vector(878675,20);
      WHEN "001100100" => data <= conv_std_logic_vector(877239,20);
      WHEN "001100101" => data <= conv_std_logic_vector(875808,20);
      WHEN "001100110" => data <= conv_std_logic_vector(874382,20);
      WHEN "001100111" => data <= conv_std_logic_vector(872960,20);
      WHEN "001101000" => data <= conv_std_logic_vector(871543,20);
      WHEN "001101001" => data <= conv_std_logic_vector(870131,20);
      WHEN "001101010" => data <= conv_std_logic_vector(868723,20);
      WHEN "001101011" => data <= conv_std_logic_vector(867319,20);
      WHEN "001101100" => data <= conv_std_logic_vector(865920,20);
      WHEN "001101101" => data <= conv_std_logic_vector(864526,20);
      WHEN "001101110" => data <= conv_std_logic_vector(863136,20);
      WHEN "001101111" => data <= conv_std_logic_vector(861751,20);
      WHEN "001110000" => data <= conv_std_logic_vector(860369,20);
      WHEN "001110001" => data <= conv_std_logic_vector(858993,20);
      WHEN "001110010" => data <= conv_std_logic_vector(857621,20);
      WHEN "001110011" => data <= conv_std_logic_vector(856253,20);
      WHEN "001110100" => data <= conv_std_logic_vector(854889,20);
      WHEN "001110101" => data <= conv_std_logic_vector(853530,20);
      WHEN "001110110" => data <= conv_std_logic_vector(852176,20);
      WHEN "001110111" => data <= conv_std_logic_vector(850825,20);
      WHEN "001111000" => data <= conv_std_logic_vector(849479,20);
      WHEN "001111001" => data <= conv_std_logic_vector(848137,20);
      WHEN "001111010" => data <= conv_std_logic_vector(846799,20);
      WHEN "001111011" => data <= conv_std_logic_vector(845465,20);
      WHEN "001111100" => data <= conv_std_logic_vector(844136,20);
      WHEN "001111101" => data <= conv_std_logic_vector(842811,20);
      WHEN "001111110" => data <= conv_std_logic_vector(841490,20);
      WHEN "001111111" => data <= conv_std_logic_vector(840173,20);
      WHEN "010000000" => data <= conv_std_logic_vector(838860,20);
      WHEN "010000001" => data <= conv_std_logic_vector(837552,20);
      WHEN "010000010" => data <= conv_std_logic_vector(836247,20);
      WHEN "010000011" => data <= conv_std_logic_vector(834946,20);
      WHEN "010000100" => data <= conv_std_logic_vector(833650,20);
      WHEN "010000101" => data <= conv_std_logic_vector(832358,20);
      WHEN "010000110" => data <= conv_std_logic_vector(831069,20);
      WHEN "010000111" => data <= conv_std_logic_vector(829785,20);
      WHEN "010001000" => data <= conv_std_logic_vector(828504,20);
      WHEN "010001001" => data <= conv_std_logic_vector(827227,20);
      WHEN "010001010" => data <= conv_std_logic_vector(825955,20);
      WHEN "010001011" => data <= conv_std_logic_vector(824686,20);
      WHEN "010001100" => data <= conv_std_logic_vector(823421,20);
      WHEN "010001101" => data <= conv_std_logic_vector(822160,20);
      WHEN "010001110" => data <= conv_std_logic_vector(820903,20);
      WHEN "010001111" => data <= conv_std_logic_vector(819650,20);
      WHEN "010010000" => data <= conv_std_logic_vector(818400,20);
      WHEN "010010001" => data <= conv_std_logic_vector(817155,20);
      WHEN "010010010" => data <= conv_std_logic_vector(815913,20);
      WHEN "010010011" => data <= conv_std_logic_vector(814675,20);
      WHEN "010010100" => data <= conv_std_logic_vector(813440,20);
      WHEN "010010101" => data <= conv_std_logic_vector(812210,20);
      WHEN "010010110" => data <= conv_std_logic_vector(810983,20);
      WHEN "010010111" => data <= conv_std_logic_vector(809760,20);
      WHEN "010011000" => data <= conv_std_logic_vector(808540,20);
      WHEN "010011001" => data <= conv_std_logic_vector(807324,20);
      WHEN "010011010" => data <= conv_std_logic_vector(806112,20);
      WHEN "010011011" => data <= conv_std_logic_vector(804903,20);
      WHEN "010011100" => data <= conv_std_logic_vector(803699,20);
      WHEN "010011101" => data <= conv_std_logic_vector(802497,20);
      WHEN "010011110" => data <= conv_std_logic_vector(801299,20);
      WHEN "010011111" => data <= conv_std_logic_vector(800105,20);
      WHEN "010100000" => data <= conv_std_logic_vector(798915,20);
      WHEN "010100001" => data <= conv_std_logic_vector(797728,20);
      WHEN "010100010" => data <= conv_std_logic_vector(796544,20);
      WHEN "010100011" => data <= conv_std_logic_vector(795364,20);
      WHEN "010100100" => data <= conv_std_logic_vector(794187,20);
      WHEN "010100101" => data <= conv_std_logic_vector(793014,20);
      WHEN "010100110" => data <= conv_std_logic_vector(791845,20);
      WHEN "010100111" => data <= conv_std_logic_vector(790678,20);
      WHEN "010101000" => data <= conv_std_logic_vector(789516,20);
      WHEN "010101001" => data <= conv_std_logic_vector(788356,20);
      WHEN "010101010" => data <= conv_std_logic_vector(787200,20);
      WHEN "010101011" => data <= conv_std_logic_vector(786048,20);
      WHEN "010101100" => data <= conv_std_logic_vector(784899,20);
      WHEN "010101101" => data <= conv_std_logic_vector(783753,20);
      WHEN "010101110" => data <= conv_std_logic_vector(782610,20);
      WHEN "010101111" => data <= conv_std_logic_vector(781471,20);
      WHEN "010110000" => data <= conv_std_logic_vector(780335,20);
      WHEN "010110001" => data <= conv_std_logic_vector(779203,20);
      WHEN "010110010" => data <= conv_std_logic_vector(778073,20);
      WHEN "010110011" => data <= conv_std_logic_vector(776947,20);
      WHEN "010110100" => data <= conv_std_logic_vector(775825,20);
      WHEN "010110101" => data <= conv_std_logic_vector(774705,20);
      WHEN "010110110" => data <= conv_std_logic_vector(773589,20);
      WHEN "010110111" => data <= conv_std_logic_vector(772476,20);
      WHEN "010111000" => data <= conv_std_logic_vector(771366,20);
      WHEN "010111001" => data <= conv_std_logic_vector(770259,20);
      WHEN "010111010" => data <= conv_std_logic_vector(769156,20);
      WHEN "010111011" => data <= conv_std_logic_vector(768055,20);
      WHEN "010111100" => data <= conv_std_logic_vector(766958,20);
      WHEN "010111101" => data <= conv_std_logic_vector(765864,20);
      WHEN "010111110" => data <= conv_std_logic_vector(764773,20);
      WHEN "010111111" => data <= conv_std_logic_vector(763685,20);
      WHEN "011000000" => data <= conv_std_logic_vector(762600,20);
      WHEN "011000001" => data <= conv_std_logic_vector(761519,20);
      WHEN "011000010" => data <= conv_std_logic_vector(760440,20);
      WHEN "011000011" => data <= conv_std_logic_vector(759364,20);
      WHEN "011000100" => data <= conv_std_logic_vector(758292,20);
      WHEN "011000101" => data <= conv_std_logic_vector(757222,20);
      WHEN "011000110" => data <= conv_std_logic_vector(756156,20);
      WHEN "011000111" => data <= conv_std_logic_vector(755092,20);
      WHEN "011001000" => data <= conv_std_logic_vector(754032,20);
      WHEN "011001001" => data <= conv_std_logic_vector(752974,20);
      WHEN "011001010" => data <= conv_std_logic_vector(751920,20);
      WHEN "011001011" => data <= conv_std_logic_vector(750868,20);
      WHEN "011001100" => data <= conv_std_logic_vector(749819,20);
      WHEN "011001101" => data <= conv_std_logic_vector(748774,20);
      WHEN "011001110" => data <= conv_std_logic_vector(747731,20);
      WHEN "011001111" => data <= conv_std_logic_vector(746691,20);
      WHEN "011010000" => data <= conv_std_logic_vector(745654,20);
      WHEN "011010001" => data <= conv_std_logic_vector(744619,20);
      WHEN "011010010" => data <= conv_std_logic_vector(743588,20);
      WHEN "011010011" => data <= conv_std_logic_vector(742560,20);
      WHEN "011010100" => data <= conv_std_logic_vector(741534,20);
      WHEN "011010101" => data <= conv_std_logic_vector(740511,20);
      WHEN "011010110" => data <= conv_std_logic_vector(739491,20);
      WHEN "011010111" => data <= conv_std_logic_vector(738474,20);
      WHEN "011011000" => data <= conv_std_logic_vector(737460,20);
      WHEN "011011001" => data <= conv_std_logic_vector(736448,20);
      WHEN "011011010" => data <= conv_std_logic_vector(735439,20);
      WHEN "011011011" => data <= conv_std_logic_vector(734433,20);
      WHEN "011011100" => data <= conv_std_logic_vector(733430,20);
      WHEN "011011101" => data <= conv_std_logic_vector(732429,20);
      WHEN "011011110" => data <= conv_std_logic_vector(731431,20);
      WHEN "011011111" => data <= conv_std_logic_vector(730436,20);
      WHEN "011100000" => data <= conv_std_logic_vector(729444,20);
      WHEN "011100001" => data <= conv_std_logic_vector(728454,20);
      WHEN "011100010" => data <= conv_std_logic_vector(727467,20);
      WHEN "011100011" => data <= conv_std_logic_vector(726483,20);
      WHEN "011100100" => data <= conv_std_logic_vector(725501,20);
      WHEN "011100101" => data <= conv_std_logic_vector(724522,20);
      WHEN "011100110" => data <= conv_std_logic_vector(723545,20);
      WHEN "011100111" => data <= conv_std_logic_vector(722572,20);
      WHEN "011101000" => data <= conv_std_logic_vector(721600,20);
      WHEN "011101001" => data <= conv_std_logic_vector(720632,20);
      WHEN "011101010" => data <= conv_std_logic_vector(719666,20);
      WHEN "011101011" => data <= conv_std_logic_vector(718702,20);
      WHEN "011101100" => data <= conv_std_logic_vector(717742,20);
      WHEN "011101101" => data <= conv_std_logic_vector(716783,20);
      WHEN "011101110" => data <= conv_std_logic_vector(715828,20);
      WHEN "011101111" => data <= conv_std_logic_vector(714874,20);
      WHEN "011110000" => data <= conv_std_logic_vector(713924,20);
      WHEN "011110001" => data <= conv_std_logic_vector(712976,20);
      WHEN "011110010" => data <= conv_std_logic_vector(712030,20);
      WHEN "011110011" => data <= conv_std_logic_vector(711087,20);
      WHEN "011110100" => data <= conv_std_logic_vector(710146,20);
      WHEN "011110101" => data <= conv_std_logic_vector(709208,20);
      WHEN "011110110" => data <= conv_std_logic_vector(708273,20);
      WHEN "011110111" => data <= conv_std_logic_vector(707339,20);
      WHEN "011111000" => data <= conv_std_logic_vector(706409,20);
      WHEN "011111001" => data <= conv_std_logic_vector(705481,20);
      WHEN "011111010" => data <= conv_std_logic_vector(704555,20);
      WHEN "011111011" => data <= conv_std_logic_vector(703631,20);
      WHEN "011111100" => data <= conv_std_logic_vector(702710,20);
      WHEN "011111101" => data <= conv_std_logic_vector(701792,20);
      WHEN "011111110" => data <= conv_std_logic_vector(700876,20);
      WHEN "011111111" => data <= conv_std_logic_vector(699962,20);
      WHEN "100000000" => data <= conv_std_logic_vector(699050,20);
      WHEN "100000001" => data <= conv_std_logic_vector(698141,20);
      WHEN "100000010" => data <= conv_std_logic_vector(697235,20);
      WHEN "100000011" => data <= conv_std_logic_vector(696330,20);
      WHEN "100000100" => data <= conv_std_logic_vector(695428,20);
      WHEN "100000101" => data <= conv_std_logic_vector(694529,20);
      WHEN "100000110" => data <= conv_std_logic_vector(693631,20);
      WHEN "100000111" => data <= conv_std_logic_vector(692736,20);
      WHEN "100001000" => data <= conv_std_logic_vector(691844,20);
      WHEN "100001001" => data <= conv_std_logic_vector(690953,20);
      WHEN "100001010" => data <= conv_std_logic_vector(690065,20);
      WHEN "100001011" => data <= conv_std_logic_vector(689179,20);
      WHEN "100001100" => data <= conv_std_logic_vector(688296,20);
      WHEN "100001101" => data <= conv_std_logic_vector(687414,20);
      WHEN "100001110" => data <= conv_std_logic_vector(686535,20);
      WHEN "100001111" => data <= conv_std_logic_vector(685659,20);
      WHEN "100010000" => data <= conv_std_logic_vector(684784,20);
      WHEN "100010001" => data <= conv_std_logic_vector(683912,20);
      WHEN "100010010" => data <= conv_std_logic_vector(683042,20);
      WHEN "100010011" => data <= conv_std_logic_vector(682174,20);
      WHEN "100010100" => data <= conv_std_logic_vector(681308,20);
      WHEN "100010101" => data <= conv_std_logic_vector(680444,20);
      WHEN "100010110" => data <= conv_std_logic_vector(679583,20);
      WHEN "100010111" => data <= conv_std_logic_vector(678724,20);
      WHEN "100011000" => data <= conv_std_logic_vector(677867,20);
      WHEN "100011001" => data <= conv_std_logic_vector(677012,20);
      WHEN "100011010" => data <= conv_std_logic_vector(676160,20);
      WHEN "100011011" => data <= conv_std_logic_vector(675309,20);
      WHEN "100011100" => data <= conv_std_logic_vector(674461,20);
      WHEN "100011101" => data <= conv_std_logic_vector(673614,20);
      WHEN "100011110" => data <= conv_std_logic_vector(672770,20);
      WHEN "100011111" => data <= conv_std_logic_vector(671928,20);
      WHEN "100100000" => data <= conv_std_logic_vector(671088,20);
      WHEN "100100001" => data <= conv_std_logic_vector(670251,20);
      WHEN "100100010" => data <= conv_std_logic_vector(669415,20);
      WHEN "100100011" => data <= conv_std_logic_vector(668581,20);
      WHEN "100100100" => data <= conv_std_logic_vector(667750,20);
      WHEN "100100101" => data <= conv_std_logic_vector(666920,20);
      WHEN "100100110" => data <= conv_std_logic_vector(666093,20);
      WHEN "100100111" => data <= conv_std_logic_vector(665267,20);
      WHEN "100101000" => data <= conv_std_logic_vector(664444,20);
      WHEN "100101001" => data <= conv_std_logic_vector(663623,20);
      WHEN "100101010" => data <= conv_std_logic_vector(662803,20);
      WHEN "100101011" => data <= conv_std_logic_vector(661986,20);
      WHEN "100101100" => data <= conv_std_logic_vector(661171,20);
      WHEN "100101101" => data <= conv_std_logic_vector(660358,20);
      WHEN "100101110" => data <= conv_std_logic_vector(659546,20);
      WHEN "100101111" => data <= conv_std_logic_vector(658737,20);
      WHEN "100110000" => data <= conv_std_logic_vector(657930,20);
      WHEN "100110001" => data <= conv_std_logic_vector(657124,20);
      WHEN "100110010" => data <= conv_std_logic_vector(656321,20);
      WHEN "100110011" => data <= conv_std_logic_vector(655520,20);
      WHEN "100110100" => data <= conv_std_logic_vector(654720,20);
      WHEN "100110101" => data <= conv_std_logic_vector(653923,20);
      WHEN "100110110" => data <= conv_std_logic_vector(653127,20);
      WHEN "100110111" => data <= conv_std_logic_vector(652334,20);
      WHEN "100111000" => data <= conv_std_logic_vector(651542,20);
      WHEN "100111001" => data <= conv_std_logic_vector(650752,20);
      WHEN "100111010" => data <= conv_std_logic_vector(649965,20);
      WHEN "100111011" => data <= conv_std_logic_vector(649179,20);
      WHEN "100111100" => data <= conv_std_logic_vector(648395,20);
      WHEN "100111101" => data <= conv_std_logic_vector(647612,20);
      WHEN "100111110" => data <= conv_std_logic_vector(646832,20);
      WHEN "100111111" => data <= conv_std_logic_vector(646054,20);
      WHEN "101000000" => data <= conv_std_logic_vector(645277,20);
      WHEN "101000001" => data <= conv_std_logic_vector(644503,20);
      WHEN "101000010" => data <= conv_std_logic_vector(643730,20);
      WHEN "101000011" => data <= conv_std_logic_vector(642959,20);
      WHEN "101000100" => data <= conv_std_logic_vector(642190,20);
      WHEN "101000101" => data <= conv_std_logic_vector(641423,20);
      WHEN "101000110" => data <= conv_std_logic_vector(640657,20);
      WHEN "101000111" => data <= conv_std_logic_vector(639894,20);
      WHEN "101001000" => data <= conv_std_logic_vector(639132,20);
      WHEN "101001001" => data <= conv_std_logic_vector(638372,20);
      WHEN "101001010" => data <= conv_std_logic_vector(637614,20);
      WHEN "101001011" => data <= conv_std_logic_vector(636857,20);
      WHEN "101001100" => data <= conv_std_logic_vector(636103,20);
      WHEN "101001101" => data <= conv_std_logic_vector(635350,20);
      WHEN "101001110" => data <= conv_std_logic_vector(634599,20);
      WHEN "101001111" => data <= conv_std_logic_vector(633850,20);
      WHEN "101010000" => data <= conv_std_logic_vector(633102,20);
      WHEN "101010001" => data <= conv_std_logic_vector(632357,20);
      WHEN "101010010" => data <= conv_std_logic_vector(631613,20);
      WHEN "101010011" => data <= conv_std_logic_vector(630870,20);
      WHEN "101010100" => data <= conv_std_logic_vector(630130,20);
      WHEN "101010101" => data <= conv_std_logic_vector(629391,20);
      WHEN "101010110" => data <= conv_std_logic_vector(628654,20);
      WHEN "101010111" => data <= conv_std_logic_vector(627919,20);
      WHEN "101011000" => data <= conv_std_logic_vector(627185,20);
      WHEN "101011001" => data <= conv_std_logic_vector(626454,20);
      WHEN "101011010" => data <= conv_std_logic_vector(625723,20);
      WHEN "101011011" => data <= conv_std_logic_vector(624995,20);
      WHEN "101011100" => data <= conv_std_logic_vector(624268,20);
      WHEN "101011101" => data <= conv_std_logic_vector(623543,20);
      WHEN "101011110" => data <= conv_std_logic_vector(622820,20);
      WHEN "101011111" => data <= conv_std_logic_vector(622098,20);
      WHEN "101100000" => data <= conv_std_logic_vector(621378,20);
      WHEN "101100001" => data <= conv_std_logic_vector(620660,20);
      WHEN "101100010" => data <= conv_std_logic_vector(619943,20);
      WHEN "101100011" => data <= conv_std_logic_vector(619228,20);
      WHEN "101100100" => data <= conv_std_logic_vector(618515,20);
      WHEN "101100101" => data <= conv_std_logic_vector(617803,20);
      WHEN "101100110" => data <= conv_std_logic_vector(617093,20);
      WHEN "101100111" => data <= conv_std_logic_vector(616384,20);
      WHEN "101101000" => data <= conv_std_logic_vector(615677,20);
      WHEN "101101001" => data <= conv_std_logic_vector(614972,20);
      WHEN "101101010" => data <= conv_std_logic_vector(614269,20);
      WHEN "101101011" => data <= conv_std_logic_vector(613567,20);
      WHEN "101101100" => data <= conv_std_logic_vector(612866,20);
      WHEN "101101101" => data <= conv_std_logic_vector(612167,20);
      WHEN "101101110" => data <= conv_std_logic_vector(611470,20);
      WHEN "101101111" => data <= conv_std_logic_vector(610774,20);
      WHEN "101110000" => data <= conv_std_logic_vector(610080,20);
      WHEN "101110001" => data <= conv_std_logic_vector(609388,20);
      WHEN "101110010" => data <= conv_std_logic_vector(608697,20);
      WHEN "101110011" => data <= conv_std_logic_vector(608008,20);
      WHEN "101110100" => data <= conv_std_logic_vector(607320,20);
      WHEN "101110101" => data <= conv_std_logic_vector(606634,20);
      WHEN "101110110" => data <= conv_std_logic_vector(605949,20);
      WHEN "101110111" => data <= conv_std_logic_vector(605266,20);
      WHEN "101111000" => data <= conv_std_logic_vector(604584,20);
      WHEN "101111001" => data <= conv_std_logic_vector(603904,20);
      WHEN "101111010" => data <= conv_std_logic_vector(603226,20);
      WHEN "101111011" => data <= conv_std_logic_vector(602549,20);
      WHEN "101111100" => data <= conv_std_logic_vector(601873,20);
      WHEN "101111101" => data <= conv_std_logic_vector(601199,20);
      WHEN "101111110" => data <= conv_std_logic_vector(600527,20);
      WHEN "101111111" => data <= conv_std_logic_vector(599856,20);
      WHEN "110000000" => data <= conv_std_logic_vector(599186,20);
      WHEN "110000001" => data <= conv_std_logic_vector(598518,20);
      WHEN "110000010" => data <= conv_std_logic_vector(597852,20);
      WHEN "110000011" => data <= conv_std_logic_vector(597187,20);
      WHEN "110000100" => data <= conv_std_logic_vector(596523,20);
      WHEN "110000101" => data <= conv_std_logic_vector(595861,20);
      WHEN "110000110" => data <= conv_std_logic_vector(595200,20);
      WHEN "110000111" => data <= conv_std_logic_vector(594541,20);
      WHEN "110001000" => data <= conv_std_logic_vector(593884,20);
      WHEN "110001001" => data <= conv_std_logic_vector(593227,20);
      WHEN "110001010" => data <= conv_std_logic_vector(592573,20);
      WHEN "110001011" => data <= conv_std_logic_vector(591919,20);
      WHEN "110001100" => data <= conv_std_logic_vector(591267,20);
      WHEN "110001101" => data <= conv_std_logic_vector(590617,20);
      WHEN "110001110" => data <= conv_std_logic_vector(589968,20);
      WHEN "110001111" => data <= conv_std_logic_vector(589320,20);
      WHEN "110010000" => data <= conv_std_logic_vector(588674,20);
      WHEN "110010001" => data <= conv_std_logic_vector(588029,20);
      WHEN "110010010" => data <= conv_std_logic_vector(587386,20);
      WHEN "110010011" => data <= conv_std_logic_vector(586744,20);
      WHEN "110010100" => data <= conv_std_logic_vector(586103,20);
      WHEN "110010101" => data <= conv_std_logic_vector(585464,20);
      WHEN "110010110" => data <= conv_std_logic_vector(584827,20);
      WHEN "110010111" => data <= conv_std_logic_vector(584190,20);
      WHEN "110011000" => data <= conv_std_logic_vector(583555,20);
      WHEN "110011001" => data <= conv_std_logic_vector(582922,20);
      WHEN "110011010" => data <= conv_std_logic_vector(582289,20);
      WHEN "110011011" => data <= conv_std_logic_vector(581658,20);
      WHEN "110011100" => data <= conv_std_logic_vector(581029,20);
      WHEN "110011101" => data <= conv_std_logic_vector(580401,20);
      WHEN "110011110" => data <= conv_std_logic_vector(579774,20);
      WHEN "110011111" => data <= conv_std_logic_vector(579149,20);
      WHEN "110100000" => data <= conv_std_logic_vector(578525,20);
      WHEN "110100001" => data <= conv_std_logic_vector(577902,20);
      WHEN "110100010" => data <= conv_std_logic_vector(577280,20);
      WHEN "110100011" => data <= conv_std_logic_vector(576660,20);
      WHEN "110100100" => data <= conv_std_logic_vector(576042,20);
      WHEN "110100101" => data <= conv_std_logic_vector(575424,20);
      WHEN "110100110" => data <= conv_std_logic_vector(574808,20);
      WHEN "110100111" => data <= conv_std_logic_vector(574193,20);
      WHEN "110101000" => data <= conv_std_logic_vector(573580,20);
      WHEN "110101001" => data <= conv_std_logic_vector(572968,20);
      WHEN "110101010" => data <= conv_std_logic_vector(572357,20);
      WHEN "110101011" => data <= conv_std_logic_vector(571747,20);
      WHEN "110101100" => data <= conv_std_logic_vector(571139,20);
      WHEN "110101101" => data <= conv_std_logic_vector(570532,20);
      WHEN "110101110" => data <= conv_std_logic_vector(569926,20);
      WHEN "110101111" => data <= conv_std_logic_vector(569322,20);
      WHEN "110110000" => data <= conv_std_logic_vector(568719,20);
      WHEN "110110001" => data <= conv_std_logic_vector(568117,20);
      WHEN "110110010" => data <= conv_std_logic_vector(567517,20);
      WHEN "110110011" => data <= conv_std_logic_vector(566917,20);
      WHEN "110110100" => data <= conv_std_logic_vector(566319,20);
      WHEN "110110101" => data <= conv_std_logic_vector(565723,20);
      WHEN "110110110" => data <= conv_std_logic_vector(565127,20);
      WHEN "110110111" => data <= conv_std_logic_vector(564533,20);
      WHEN "110111000" => data <= conv_std_logic_vector(563940,20);
      WHEN "110111001" => data <= conv_std_logic_vector(563348,20);
      WHEN "110111010" => data <= conv_std_logic_vector(562758,20);
      WHEN "110111011" => data <= conv_std_logic_vector(562168,20);
      WHEN "110111100" => data <= conv_std_logic_vector(561580,20);
      WHEN "110111101" => data <= conv_std_logic_vector(560993,20);
      WHEN "110111110" => data <= conv_std_logic_vector(560408,20);
      WHEN "110111111" => data <= conv_std_logic_vector(559824,20);
      WHEN "111000000" => data <= conv_std_logic_vector(559240,20);
      WHEN "111000001" => data <= conv_std_logic_vector(558658,20);
      WHEN "111000010" => data <= conv_std_logic_vector(558078,20);
      WHEN "111000011" => data <= conv_std_logic_vector(557498,20);
      WHEN "111000100" => data <= conv_std_logic_vector(556920,20);
      WHEN "111000101" => data <= conv_std_logic_vector(556343,20);
      WHEN "111000110" => data <= conv_std_logic_vector(555767,20);
      WHEN "111000111" => data <= conv_std_logic_vector(555192,20);
      WHEN "111001000" => data <= conv_std_logic_vector(554619,20);
      WHEN "111001001" => data <= conv_std_logic_vector(554046,20);
      WHEN "111001010" => data <= conv_std_logic_vector(553475,20);
      WHEN "111001011" => data <= conv_std_logic_vector(552905,20);
      WHEN "111001100" => data <= conv_std_logic_vector(552336,20);
      WHEN "111001101" => data <= conv_std_logic_vector(551769,20);
      WHEN "111001110" => data <= conv_std_logic_vector(551202,20);
      WHEN "111001111" => data <= conv_std_logic_vector(550637,20);
      WHEN "111010000" => data <= conv_std_logic_vector(550073,20);
      WHEN "111010001" => data <= conv_std_logic_vector(549509,20);
      WHEN "111010010" => data <= conv_std_logic_vector(548948,20);
      WHEN "111010011" => data <= conv_std_logic_vector(548387,20);
      WHEN "111010100" => data <= conv_std_logic_vector(547827,20);
      WHEN "111010101" => data <= conv_std_logic_vector(547269,20);
      WHEN "111010110" => data <= conv_std_logic_vector(546712,20);
      WHEN "111010111" => data <= conv_std_logic_vector(546155,20);
      WHEN "111011000" => data <= conv_std_logic_vector(545600,20);
      WHEN "111011001" => data <= conv_std_logic_vector(545046,20);
      WHEN "111011010" => data <= conv_std_logic_vector(544494,20);
      WHEN "111011011" => data <= conv_std_logic_vector(543942,20);
      WHEN "111011100" => data <= conv_std_logic_vector(543391,20);
      WHEN "111011101" => data <= conv_std_logic_vector(542842,20);
      WHEN "111011110" => data <= conv_std_logic_vector(542294,20);
      WHEN "111011111" => data <= conv_std_logic_vector(541746,20);
      WHEN "111100000" => data <= conv_std_logic_vector(541200,20);
      WHEN "111100001" => data <= conv_std_logic_vector(540655,20);
      WHEN "111100010" => data <= conv_std_logic_vector(540111,20);
      WHEN "111100011" => data <= conv_std_logic_vector(539569,20);
      WHEN "111100100" => data <= conv_std_logic_vector(539027,20);
      WHEN "111100101" => data <= conv_std_logic_vector(538486,20);
      WHEN "111100110" => data <= conv_std_logic_vector(537947,20);
      WHEN "111100111" => data <= conv_std_logic_vector(537408,20);
      WHEN "111101000" => data <= conv_std_logic_vector(536871,20);
      WHEN "111101001" => data <= conv_std_logic_vector(536334,20);
      WHEN "111101010" => data <= conv_std_logic_vector(535799,20);
      WHEN "111101011" => data <= conv_std_logic_vector(535265,20);
      WHEN "111101100" => data <= conv_std_logic_vector(534732,20);
      WHEN "111101101" => data <= conv_std_logic_vector(534200,20);
      WHEN "111101110" => data <= conv_std_logic_vector(533669,20);
      WHEN "111101111" => data <= conv_std_logic_vector(533139,20);
      WHEN "111110000" => data <= conv_std_logic_vector(532610,20);
      WHEN "111110001" => data <= conv_std_logic_vector(532082,20);
      WHEN "111110010" => data <= conv_std_logic_vector(531555,20);
      WHEN "111110011" => data <= conv_std_logic_vector(531029,20);
      WHEN "111110100" => data <= conv_std_logic_vector(530505,20);
      WHEN "111110101" => data <= conv_std_logic_vector(529981,20);
      WHEN "111110110" => data <= conv_std_logic_vector(529458,20);
      WHEN "111110111" => data <= conv_std_logic_vector(528937,20);
      WHEN "111111000" => data <= conv_std_logic_vector(528416,20);
      WHEN "111111001" => data <= conv_std_logic_vector(527897,20);
      WHEN "111111010" => data <= conv_std_logic_vector(527378,20);
      WHEN "111111011" => data <= conv_std_logic_vector(526860,20);
      WHEN "111111100" => data <= conv_std_logic_vector(526344,20);
      WHEN "111111101" => data <= conv_std_logic_vector(525828,20);
      WHEN "111111110" => data <= conv_std_logic_vector(525314,20);
      WHEN "111111111" => data <= conv_std_logic_vector(524800,20);
      WHEN others => data <= conv_std_logic_vector(0,20);
    END CASE;
  END PROCESS;

END rtl;
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_DIV_LUT1.VHD                           ***
--***                                             ***
--***   Function: Look Up Table - Inverse         ***
--***                                             ***
--***   Generated by MATLAB Utility               ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_div_lut1 IS
PORT (
      add : IN STD_LOGIC_VECTOR (9 DOWNTO 1);
		data : OUT STD_LOGIC_VECTOR (11 DOWNTO 1)
);
END fp_div_lut1;

ARCHITECTURE rtl OF fp_div_lut1 IS

BEGIN

  pca: PROCESS (add)
  BEGIN
    CASE add IS
      WHEN "000000000" => data <= conv_std_logic_vector(2044,11);
      WHEN "000000001" => data <= conv_std_logic_vector(2036,11);
      WHEN "000000010" => data <= conv_std_logic_vector(2028,11);
      WHEN "000000011" => data <= conv_std_logic_vector(2020,11);
      WHEN "000000100" => data <= conv_std_logic_vector(2012,11);
      WHEN "000000101" => data <= conv_std_logic_vector(2005,11);
      WHEN "000000110" => data <= conv_std_logic_vector(1997,11);
      WHEN "000000111" => data <= conv_std_logic_vector(1989,11);
      WHEN "000001000" => data <= conv_std_logic_vector(1982,11);
      WHEN "000001001" => data <= conv_std_logic_vector(1974,11);
      WHEN "000001010" => data <= conv_std_logic_vector(1967,11);
      WHEN "000001011" => data <= conv_std_logic_vector(1959,11);
      WHEN "000001100" => data <= conv_std_logic_vector(1952,11);
      WHEN "000001101" => data <= conv_std_logic_vector(1944,11);
      WHEN "000001110" => data <= conv_std_logic_vector(1937,11);
      WHEN "000001111" => data <= conv_std_logic_vector(1929,11);
      WHEN "000010000" => data <= conv_std_logic_vector(1922,11);
      WHEN "000010001" => data <= conv_std_logic_vector(1915,11);
      WHEN "000010010" => data <= conv_std_logic_vector(1908,11);
      WHEN "000010011" => data <= conv_std_logic_vector(1900,11);
      WHEN "000010100" => data <= conv_std_logic_vector(1893,11);
      WHEN "000010101" => data <= conv_std_logic_vector(1886,11);
      WHEN "000010110" => data <= conv_std_logic_vector(1879,11);
      WHEN "000010111" => data <= conv_std_logic_vector(1872,11);
      WHEN "000011000" => data <= conv_std_logic_vector(1865,11);
      WHEN "000011001" => data <= conv_std_logic_vector(1858,11);
      WHEN "000011010" => data <= conv_std_logic_vector(1851,11);
      WHEN "000011011" => data <= conv_std_logic_vector(1845,11);
      WHEN "000011100" => data <= conv_std_logic_vector(1838,11);
      WHEN "000011101" => data <= conv_std_logic_vector(1831,11);
      WHEN "000011110" => data <= conv_std_logic_vector(1824,11);
      WHEN "000011111" => data <= conv_std_logic_vector(1817,11);
      WHEN "000100000" => data <= conv_std_logic_vector(1811,11);
      WHEN "000100001" => data <= conv_std_logic_vector(1804,11);
      WHEN "000100010" => data <= conv_std_logic_vector(1798,11);
      WHEN "000100011" => data <= conv_std_logic_vector(1791,11);
      WHEN "000100100" => data <= conv_std_logic_vector(1785,11);
      WHEN "000100101" => data <= conv_std_logic_vector(1778,11);
      WHEN "000100110" => data <= conv_std_logic_vector(1772,11);
      WHEN "000100111" => data <= conv_std_logic_vector(1765,11);
      WHEN "000101000" => data <= conv_std_logic_vector(1759,11);
      WHEN "000101001" => data <= conv_std_logic_vector(1752,11);
      WHEN "000101010" => data <= conv_std_logic_vector(1746,11);
      WHEN "000101011" => data <= conv_std_logic_vector(1740,11);
      WHEN "000101100" => data <= conv_std_logic_vector(1734,11);
      WHEN "000101101" => data <= conv_std_logic_vector(1727,11);
      WHEN "000101110" => data <= conv_std_logic_vector(1721,11);
      WHEN "000101111" => data <= conv_std_logic_vector(1715,11);
      WHEN "000110000" => data <= conv_std_logic_vector(1709,11);
      WHEN "000110001" => data <= conv_std_logic_vector(1703,11);
      WHEN "000110010" => data <= conv_std_logic_vector(1697,11);
      WHEN "000110011" => data <= conv_std_logic_vector(1691,11);
      WHEN "000110100" => data <= conv_std_logic_vector(1685,11);
      WHEN "000110101" => data <= conv_std_logic_vector(1679,11);
      WHEN "000110110" => data <= conv_std_logic_vector(1673,11);
      WHEN "000110111" => data <= conv_std_logic_vector(1667,11);
      WHEN "000111000" => data <= conv_std_logic_vector(1661,11);
      WHEN "000111001" => data <= conv_std_logic_vector(1655,11);
      WHEN "000111010" => data <= conv_std_logic_vector(1650,11);
      WHEN "000111011" => data <= conv_std_logic_vector(1644,11);
      WHEN "000111100" => data <= conv_std_logic_vector(1638,11);
      WHEN "000111101" => data <= conv_std_logic_vector(1632,11);
      WHEN "000111110" => data <= conv_std_logic_vector(1627,11);
      WHEN "000111111" => data <= conv_std_logic_vector(1621,11);
      WHEN "001000000" => data <= conv_std_logic_vector(1615,11);
      WHEN "001000001" => data <= conv_std_logic_vector(1610,11);
      WHEN "001000010" => data <= conv_std_logic_vector(1604,11);
      WHEN "001000011" => data <= conv_std_logic_vector(1599,11);
      WHEN "001000100" => data <= conv_std_logic_vector(1593,11);
      WHEN "001000101" => data <= conv_std_logic_vector(1588,11);
      WHEN "001000110" => data <= conv_std_logic_vector(1582,11);
      WHEN "001000111" => data <= conv_std_logic_vector(1577,11);
      WHEN "001001000" => data <= conv_std_logic_vector(1571,11);
      WHEN "001001001" => data <= conv_std_logic_vector(1566,11);
      WHEN "001001010" => data <= conv_std_logic_vector(1561,11);
      WHEN "001001011" => data <= conv_std_logic_vector(1555,11);
      WHEN "001001100" => data <= conv_std_logic_vector(1550,11);
      WHEN "001001101" => data <= conv_std_logic_vector(1545,11);
      WHEN "001001110" => data <= conv_std_logic_vector(1540,11);
      WHEN "001001111" => data <= conv_std_logic_vector(1534,11);
      WHEN "001010000" => data <= conv_std_logic_vector(1529,11);
      WHEN "001010001" => data <= conv_std_logic_vector(1524,11);
      WHEN "001010010" => data <= conv_std_logic_vector(1519,11);
      WHEN "001010011" => data <= conv_std_logic_vector(1514,11);
      WHEN "001010100" => data <= conv_std_logic_vector(1509,11);
      WHEN "001010101" => data <= conv_std_logic_vector(1504,11);
      WHEN "001010110" => data <= conv_std_logic_vector(1499,11);
      WHEN "001010111" => data <= conv_std_logic_vector(1494,11);
      WHEN "001011000" => data <= conv_std_logic_vector(1489,11);
      WHEN "001011001" => data <= conv_std_logic_vector(1484,11);
      WHEN "001011010" => data <= conv_std_logic_vector(1479,11);
      WHEN "001011011" => data <= conv_std_logic_vector(1474,11);
      WHEN "001011100" => data <= conv_std_logic_vector(1469,11);
      WHEN "001011101" => data <= conv_std_logic_vector(1464,11);
      WHEN "001011110" => data <= conv_std_logic_vector(1460,11);
      WHEN "001011111" => data <= conv_std_logic_vector(1455,11);
      WHEN "001100000" => data <= conv_std_logic_vector(1450,11);
      WHEN "001100001" => data <= conv_std_logic_vector(1445,11);
      WHEN "001100010" => data <= conv_std_logic_vector(1440,11);
      WHEN "001100011" => data <= conv_std_logic_vector(1436,11);
      WHEN "001100100" => data <= conv_std_logic_vector(1431,11);
      WHEN "001100101" => data <= conv_std_logic_vector(1426,11);
      WHEN "001100110" => data <= conv_std_logic_vector(1422,11);
      WHEN "001100111" => data <= conv_std_logic_vector(1417,11);
      WHEN "001101000" => data <= conv_std_logic_vector(1413,11);
      WHEN "001101001" => data <= conv_std_logic_vector(1408,11);
      WHEN "001101010" => data <= conv_std_logic_vector(1403,11);
      WHEN "001101011" => data <= conv_std_logic_vector(1399,11);
      WHEN "001101100" => data <= conv_std_logic_vector(1394,11);
      WHEN "001101101" => data <= conv_std_logic_vector(1390,11);
      WHEN "001101110" => data <= conv_std_logic_vector(1385,11);
      WHEN "001101111" => data <= conv_std_logic_vector(1381,11);
      WHEN "001110000" => data <= conv_std_logic_vector(1377,11);
      WHEN "001110001" => data <= conv_std_logic_vector(1372,11);
      WHEN "001110010" => data <= conv_std_logic_vector(1368,11);
      WHEN "001110011" => data <= conv_std_logic_vector(1363,11);
      WHEN "001110100" => data <= conv_std_logic_vector(1359,11);
      WHEN "001110101" => data <= conv_std_logic_vector(1355,11);
      WHEN "001110110" => data <= conv_std_logic_vector(1351,11);
      WHEN "001110111" => data <= conv_std_logic_vector(1346,11);
      WHEN "001111000" => data <= conv_std_logic_vector(1342,11);
      WHEN "001111001" => data <= conv_std_logic_vector(1338,11);
      WHEN "001111010" => data <= conv_std_logic_vector(1334,11);
      WHEN "001111011" => data <= conv_std_logic_vector(1329,11);
      WHEN "001111100" => data <= conv_std_logic_vector(1325,11);
      WHEN "001111101" => data <= conv_std_logic_vector(1321,11);
      WHEN "001111110" => data <= conv_std_logic_vector(1317,11);
      WHEN "001111111" => data <= conv_std_logic_vector(1313,11);
      WHEN "010000000" => data <= conv_std_logic_vector(1309,11);
      WHEN "010000001" => data <= conv_std_logic_vector(1305,11);
      WHEN "010000010" => data <= conv_std_logic_vector(1301,11);
      WHEN "010000011" => data <= conv_std_logic_vector(1297,11);
      WHEN "010000100" => data <= conv_std_logic_vector(1292,11);
      WHEN "010000101" => data <= conv_std_logic_vector(1288,11);
      WHEN "010000110" => data <= conv_std_logic_vector(1284,11);
      WHEN "010000111" => data <= conv_std_logic_vector(1281,11);
      WHEN "010001000" => data <= conv_std_logic_vector(1277,11);
      WHEN "010001001" => data <= conv_std_logic_vector(1273,11);
      WHEN "010001010" => data <= conv_std_logic_vector(1269,11);
      WHEN "010001011" => data <= conv_std_logic_vector(1265,11);
      WHEN "010001100" => data <= conv_std_logic_vector(1261,11);
      WHEN "010001101" => data <= conv_std_logic_vector(1257,11);
      WHEN "010001110" => data <= conv_std_logic_vector(1253,11);
      WHEN "010001111" => data <= conv_std_logic_vector(1249,11);
      WHEN "010010000" => data <= conv_std_logic_vector(1246,11);
      WHEN "010010001" => data <= conv_std_logic_vector(1242,11);
      WHEN "010010010" => data <= conv_std_logic_vector(1238,11);
      WHEN "010010011" => data <= conv_std_logic_vector(1234,11);
      WHEN "010010100" => data <= conv_std_logic_vector(1231,11);
      WHEN "010010101" => data <= conv_std_logic_vector(1227,11);
      WHEN "010010110" => data <= conv_std_logic_vector(1223,11);
      WHEN "010010111" => data <= conv_std_logic_vector(1220,11);
      WHEN "010011000" => data <= conv_std_logic_vector(1216,11);
      WHEN "010011001" => data <= conv_std_logic_vector(1212,11);
      WHEN "010011010" => data <= conv_std_logic_vector(1209,11);
      WHEN "010011011" => data <= conv_std_logic_vector(1205,11);
      WHEN "010011100" => data <= conv_std_logic_vector(1201,11);
      WHEN "010011101" => data <= conv_std_logic_vector(1198,11);
      WHEN "010011110" => data <= conv_std_logic_vector(1194,11);
      WHEN "010011111" => data <= conv_std_logic_vector(1191,11);
      WHEN "010100000" => data <= conv_std_logic_vector(1187,11);
      WHEN "010100001" => data <= conv_std_logic_vector(1184,11);
      WHEN "010100010" => data <= conv_std_logic_vector(1180,11);
      WHEN "010100011" => data <= conv_std_logic_vector(1177,11);
      WHEN "010100100" => data <= conv_std_logic_vector(1173,11);
      WHEN "010100101" => data <= conv_std_logic_vector(1170,11);
      WHEN "010100110" => data <= conv_std_logic_vector(1166,11);
      WHEN "010100111" => data <= conv_std_logic_vector(1163,11);
      WHEN "010101000" => data <= conv_std_logic_vector(1159,11);
      WHEN "010101001" => data <= conv_std_logic_vector(1156,11);
      WHEN "010101010" => data <= conv_std_logic_vector(1153,11);
      WHEN "010101011" => data <= conv_std_logic_vector(1149,11);
      WHEN "010101100" => data <= conv_std_logic_vector(1146,11);
      WHEN "010101101" => data <= conv_std_logic_vector(1142,11);
      WHEN "010101110" => data <= conv_std_logic_vector(1139,11);
      WHEN "010101111" => data <= conv_std_logic_vector(1136,11);
      WHEN "010110000" => data <= conv_std_logic_vector(1133,11);
      WHEN "010110001" => data <= conv_std_logic_vector(1129,11);
      WHEN "010110010" => data <= conv_std_logic_vector(1126,11);
      WHEN "010110011" => data <= conv_std_logic_vector(1123,11);
      WHEN "010110100" => data <= conv_std_logic_vector(1120,11);
      WHEN "010110101" => data <= conv_std_logic_vector(1116,11);
      WHEN "010110110" => data <= conv_std_logic_vector(1113,11);
      WHEN "010110111" => data <= conv_std_logic_vector(1110,11);
      WHEN "010111000" => data <= conv_std_logic_vector(1107,11);
      WHEN "010111001" => data <= conv_std_logic_vector(1104,11);
      WHEN "010111010" => data <= conv_std_logic_vector(1100,11);
      WHEN "010111011" => data <= conv_std_logic_vector(1097,11);
      WHEN "010111100" => data <= conv_std_logic_vector(1094,11);
      WHEN "010111101" => data <= conv_std_logic_vector(1091,11);
      WHEN "010111110" => data <= conv_std_logic_vector(1088,11);
      WHEN "010111111" => data <= conv_std_logic_vector(1085,11);
      WHEN "011000000" => data <= conv_std_logic_vector(1082,11);
      WHEN "011000001" => data <= conv_std_logic_vector(1079,11);
      WHEN "011000010" => data <= conv_std_logic_vector(1076,11);
      WHEN "011000011" => data <= conv_std_logic_vector(1073,11);
      WHEN "011000100" => data <= conv_std_logic_vector(1070,11);
      WHEN "011000101" => data <= conv_std_logic_vector(1067,11);
      WHEN "011000110" => data <= conv_std_logic_vector(1064,11);
      WHEN "011000111" => data <= conv_std_logic_vector(1061,11);
      WHEN "011001000" => data <= conv_std_logic_vector(1058,11);
      WHEN "011001001" => data <= conv_std_logic_vector(1055,11);
      WHEN "011001010" => data <= conv_std_logic_vector(1052,11);
      WHEN "011001011" => data <= conv_std_logic_vector(1049,11);
      WHEN "011001100" => data <= conv_std_logic_vector(1046,11);
      WHEN "011001101" => data <= conv_std_logic_vector(1043,11);
      WHEN "011001110" => data <= conv_std_logic_vector(1040,11);
      WHEN "011001111" => data <= conv_std_logic_vector(1037,11);
      WHEN "011010000" => data <= conv_std_logic_vector(1034,11);
      WHEN "011010001" => data <= conv_std_logic_vector(1031,11);
      WHEN "011010010" => data <= conv_std_logic_vector(1028,11);
      WHEN "011010011" => data <= conv_std_logic_vector(1026,11);
      WHEN "011010100" => data <= conv_std_logic_vector(1023,11);
      WHEN "011010101" => data <= conv_std_logic_vector(1020,11);
      WHEN "011010110" => data <= conv_std_logic_vector(1017,11);
      WHEN "011010111" => data <= conv_std_logic_vector(1014,11);
      WHEN "011011000" => data <= conv_std_logic_vector(1012,11);
      WHEN "011011001" => data <= conv_std_logic_vector(1009,11);
      WHEN "011011010" => data <= conv_std_logic_vector(1006,11);
      WHEN "011011011" => data <= conv_std_logic_vector(1003,11);
      WHEN "011011100" => data <= conv_std_logic_vector(1001,11);
      WHEN "011011101" => data <= conv_std_logic_vector(998,11);
      WHEN "011011110" => data <= conv_std_logic_vector(995,11);
      WHEN "011011111" => data <= conv_std_logic_vector(992,11);
      WHEN "011100000" => data <= conv_std_logic_vector(990,11);
      WHEN "011100001" => data <= conv_std_logic_vector(987,11);
      WHEN "011100010" => data <= conv_std_logic_vector(984,11);
      WHEN "011100011" => data <= conv_std_logic_vector(982,11);
      WHEN "011100100" => data <= conv_std_logic_vector(979,11);
      WHEN "011100101" => data <= conv_std_logic_vector(976,11);
      WHEN "011100110" => data <= conv_std_logic_vector(974,11);
      WHEN "011100111" => data <= conv_std_logic_vector(971,11);
      WHEN "011101000" => data <= conv_std_logic_vector(969,11);
      WHEN "011101001" => data <= conv_std_logic_vector(966,11);
      WHEN "011101010" => data <= conv_std_logic_vector(963,11);
      WHEN "011101011" => data <= conv_std_logic_vector(961,11);
      WHEN "011101100" => data <= conv_std_logic_vector(958,11);
      WHEN "011101101" => data <= conv_std_logic_vector(956,11);
      WHEN "011101110" => data <= conv_std_logic_vector(953,11);
      WHEN "011101111" => data <= conv_std_logic_vector(951,11);
      WHEN "011110000" => data <= conv_std_logic_vector(948,11);
      WHEN "011110001" => data <= conv_std_logic_vector(946,11);
      WHEN "011110010" => data <= conv_std_logic_vector(943,11);
      WHEN "011110011" => data <= conv_std_logic_vector(941,11);
      WHEN "011110100" => data <= conv_std_logic_vector(938,11);
      WHEN "011110101" => data <= conv_std_logic_vector(936,11);
      WHEN "011110110" => data <= conv_std_logic_vector(933,11);
      WHEN "011110111" => data <= conv_std_logic_vector(931,11);
      WHEN "011111000" => data <= conv_std_logic_vector(928,11);
      WHEN "011111001" => data <= conv_std_logic_vector(926,11);
      WHEN "011111010" => data <= conv_std_logic_vector(923,11);
      WHEN "011111011" => data <= conv_std_logic_vector(921,11);
      WHEN "011111100" => data <= conv_std_logic_vector(919,11);
      WHEN "011111101" => data <= conv_std_logic_vector(916,11);
      WHEN "011111110" => data <= conv_std_logic_vector(914,11);
      WHEN "011111111" => data <= conv_std_logic_vector(911,11);
      WHEN "100000000" => data <= conv_std_logic_vector(909,11);
      WHEN "100000001" => data <= conv_std_logic_vector(907,11);
      WHEN "100000010" => data <= conv_std_logic_vector(904,11);
      WHEN "100000011" => data <= conv_std_logic_vector(902,11);
      WHEN "100000100" => data <= conv_std_logic_vector(900,11);
      WHEN "100000101" => data <= conv_std_logic_vector(897,11);
      WHEN "100000110" => data <= conv_std_logic_vector(895,11);
      WHEN "100000111" => data <= conv_std_logic_vector(893,11);
      WHEN "100001000" => data <= conv_std_logic_vector(890,11);
      WHEN "100001001" => data <= conv_std_logic_vector(888,11);
      WHEN "100001010" => data <= conv_std_logic_vector(886,11);
      WHEN "100001011" => data <= conv_std_logic_vector(884,11);
      WHEN "100001100" => data <= conv_std_logic_vector(881,11);
      WHEN "100001101" => data <= conv_std_logic_vector(879,11);
      WHEN "100001110" => data <= conv_std_logic_vector(877,11);
      WHEN "100001111" => data <= conv_std_logic_vector(875,11);
      WHEN "100010000" => data <= conv_std_logic_vector(872,11);
      WHEN "100010001" => data <= conv_std_logic_vector(870,11);
      WHEN "100010010" => data <= conv_std_logic_vector(868,11);
      WHEN "100010011" => data <= conv_std_logic_vector(866,11);
      WHEN "100010100" => data <= conv_std_logic_vector(864,11);
      WHEN "100010101" => data <= conv_std_logic_vector(861,11);
      WHEN "100010110" => data <= conv_std_logic_vector(859,11);
      WHEN "100010111" => data <= conv_std_logic_vector(857,11);
      WHEN "100011000" => data <= conv_std_logic_vector(855,11);
      WHEN "100011001" => data <= conv_std_logic_vector(853,11);
      WHEN "100011010" => data <= conv_std_logic_vector(851,11);
      WHEN "100011011" => data <= conv_std_logic_vector(848,11);
      WHEN "100011100" => data <= conv_std_logic_vector(846,11);
      WHEN "100011101" => data <= conv_std_logic_vector(844,11);
      WHEN "100011110" => data <= conv_std_logic_vector(842,11);
      WHEN "100011111" => data <= conv_std_logic_vector(840,11);
      WHEN "100100000" => data <= conv_std_logic_vector(838,11);
      WHEN "100100001" => data <= conv_std_logic_vector(836,11);
      WHEN "100100010" => data <= conv_std_logic_vector(834,11);
      WHEN "100100011" => data <= conv_std_logic_vector(832,11);
      WHEN "100100100" => data <= conv_std_logic_vector(830,11);
      WHEN "100100101" => data <= conv_std_logic_vector(827,11);
      WHEN "100100110" => data <= conv_std_logic_vector(825,11);
      WHEN "100100111" => data <= conv_std_logic_vector(823,11);
      WHEN "100101000" => data <= conv_std_logic_vector(821,11);
      WHEN "100101001" => data <= conv_std_logic_vector(819,11);
      WHEN "100101010" => data <= conv_std_logic_vector(817,11);
      WHEN "100101011" => data <= conv_std_logic_vector(815,11);
      WHEN "100101100" => data <= conv_std_logic_vector(813,11);
      WHEN "100101101" => data <= conv_std_logic_vector(811,11);
      WHEN "100101110" => data <= conv_std_logic_vector(809,11);
      WHEN "100101111" => data <= conv_std_logic_vector(807,11);
      WHEN "100110000" => data <= conv_std_logic_vector(805,11);
      WHEN "100110001" => data <= conv_std_logic_vector(803,11);
      WHEN "100110010" => data <= conv_std_logic_vector(801,11);
      WHEN "100110011" => data <= conv_std_logic_vector(799,11);
      WHEN "100110100" => data <= conv_std_logic_vector(797,11);
      WHEN "100110101" => data <= conv_std_logic_vector(796,11);
      WHEN "100110110" => data <= conv_std_logic_vector(794,11);
      WHEN "100110111" => data <= conv_std_logic_vector(792,11);
      WHEN "100111000" => data <= conv_std_logic_vector(790,11);
      WHEN "100111001" => data <= conv_std_logic_vector(788,11);
      WHEN "100111010" => data <= conv_std_logic_vector(786,11);
      WHEN "100111011" => data <= conv_std_logic_vector(784,11);
      WHEN "100111100" => data <= conv_std_logic_vector(782,11);
      WHEN "100111101" => data <= conv_std_logic_vector(780,11);
      WHEN "100111110" => data <= conv_std_logic_vector(778,11);
      WHEN "100111111" => data <= conv_std_logic_vector(777,11);
      WHEN "101000000" => data <= conv_std_logic_vector(775,11);
      WHEN "101000001" => data <= conv_std_logic_vector(773,11);
      WHEN "101000010" => data <= conv_std_logic_vector(771,11);
      WHEN "101000011" => data <= conv_std_logic_vector(769,11);
      WHEN "101000100" => data <= conv_std_logic_vector(767,11);
      WHEN "101000101" => data <= conv_std_logic_vector(765,11);
      WHEN "101000110" => data <= conv_std_logic_vector(764,11);
      WHEN "101000111" => data <= conv_std_logic_vector(762,11);
      WHEN "101001000" => data <= conv_std_logic_vector(760,11);
      WHEN "101001001" => data <= conv_std_logic_vector(758,11);
      WHEN "101001010" => data <= conv_std_logic_vector(756,11);
      WHEN "101001011" => data <= conv_std_logic_vector(755,11);
      WHEN "101001100" => data <= conv_std_logic_vector(753,11);
      WHEN "101001101" => data <= conv_std_logic_vector(751,11);
      WHEN "101001110" => data <= conv_std_logic_vector(749,11);
      WHEN "101001111" => data <= conv_std_logic_vector(747,11);
      WHEN "101010000" => data <= conv_std_logic_vector(746,11);
      WHEN "101010001" => data <= conv_std_logic_vector(744,11);
      WHEN "101010010" => data <= conv_std_logic_vector(742,11);
      WHEN "101010011" => data <= conv_std_logic_vector(740,11);
      WHEN "101010100" => data <= conv_std_logic_vector(739,11);
      WHEN "101010101" => data <= conv_std_logic_vector(737,11);
      WHEN "101010110" => data <= conv_std_logic_vector(735,11);
      WHEN "101010111" => data <= conv_std_logic_vector(734,11);
      WHEN "101011000" => data <= conv_std_logic_vector(732,11);
      WHEN "101011001" => data <= conv_std_logic_vector(730,11);
      WHEN "101011010" => data <= conv_std_logic_vector(728,11);
      WHEN "101011011" => data <= conv_std_logic_vector(727,11);
      WHEN "101011100" => data <= conv_std_logic_vector(725,11);
      WHEN "101011101" => data <= conv_std_logic_vector(723,11);
      WHEN "101011110" => data <= conv_std_logic_vector(722,11);
      WHEN "101011111" => data <= conv_std_logic_vector(720,11);
      WHEN "101100000" => data <= conv_std_logic_vector(718,11);
      WHEN "101100001" => data <= conv_std_logic_vector(717,11);
      WHEN "101100010" => data <= conv_std_logic_vector(715,11);
      WHEN "101100011" => data <= conv_std_logic_vector(713,11);
      WHEN "101100100" => data <= conv_std_logic_vector(712,11);
      WHEN "101100101" => data <= conv_std_logic_vector(710,11);
      WHEN "101100110" => data <= conv_std_logic_vector(708,11);
      WHEN "101100111" => data <= conv_std_logic_vector(707,11);
      WHEN "101101000" => data <= conv_std_logic_vector(705,11);
      WHEN "101101001" => data <= conv_std_logic_vector(704,11);
      WHEN "101101010" => data <= conv_std_logic_vector(702,11);
      WHEN "101101011" => data <= conv_std_logic_vector(700,11);
      WHEN "101101100" => data <= conv_std_logic_vector(699,11);
      WHEN "101101101" => data <= conv_std_logic_vector(697,11);
      WHEN "101101110" => data <= conv_std_logic_vector(696,11);
      WHEN "101101111" => data <= conv_std_logic_vector(694,11);
      WHEN "101110000" => data <= conv_std_logic_vector(692,11);
      WHEN "101110001" => data <= conv_std_logic_vector(691,11);
      WHEN "101110010" => data <= conv_std_logic_vector(689,11);
      WHEN "101110011" => data <= conv_std_logic_vector(688,11);
      WHEN "101110100" => data <= conv_std_logic_vector(686,11);
      WHEN "101110101" => data <= conv_std_logic_vector(685,11);
      WHEN "101110110" => data <= conv_std_logic_vector(683,11);
      WHEN "101110111" => data <= conv_std_logic_vector(682,11);
      WHEN "101111000" => data <= conv_std_logic_vector(680,11);
      WHEN "101111001" => data <= conv_std_logic_vector(679,11);
      WHEN "101111010" => data <= conv_std_logic_vector(677,11);
      WHEN "101111011" => data <= conv_std_logic_vector(676,11);
      WHEN "101111100" => data <= conv_std_logic_vector(674,11);
      WHEN "101111101" => data <= conv_std_logic_vector(672,11);
      WHEN "101111110" => data <= conv_std_logic_vector(671,11);
      WHEN "101111111" => data <= conv_std_logic_vector(669,11);
      WHEN "110000000" => data <= conv_std_logic_vector(668,11);
      WHEN "110000001" => data <= conv_std_logic_vector(667,11);
      WHEN "110000010" => data <= conv_std_logic_vector(665,11);
      WHEN "110000011" => data <= conv_std_logic_vector(664,11);
      WHEN "110000100" => data <= conv_std_logic_vector(662,11);
      WHEN "110000101" => data <= conv_std_logic_vector(661,11);
      WHEN "110000110" => data <= conv_std_logic_vector(659,11);
      WHEN "110000111" => data <= conv_std_logic_vector(658,11);
      WHEN "110001000" => data <= conv_std_logic_vector(656,11);
      WHEN "110001001" => data <= conv_std_logic_vector(655,11);
      WHEN "110001010" => data <= conv_std_logic_vector(653,11);
      WHEN "110001011" => data <= conv_std_logic_vector(652,11);
      WHEN "110001100" => data <= conv_std_logic_vector(650,11);
      WHEN "110001101" => data <= conv_std_logic_vector(649,11);
      WHEN "110001110" => data <= conv_std_logic_vector(648,11);
      WHEN "110001111" => data <= conv_std_logic_vector(646,11);
      WHEN "110010000" => data <= conv_std_logic_vector(645,11);
      WHEN "110010001" => data <= conv_std_logic_vector(643,11);
      WHEN "110010010" => data <= conv_std_logic_vector(642,11);
      WHEN "110010011" => data <= conv_std_logic_vector(641,11);
      WHEN "110010100" => data <= conv_std_logic_vector(639,11);
      WHEN "110010101" => data <= conv_std_logic_vector(638,11);
      WHEN "110010110" => data <= conv_std_logic_vector(636,11);
      WHEN "110010111" => data <= conv_std_logic_vector(635,11);
      WHEN "110011000" => data <= conv_std_logic_vector(634,11);
      WHEN "110011001" => data <= conv_std_logic_vector(632,11);
      WHEN "110011010" => data <= conv_std_logic_vector(631,11);
      WHEN "110011011" => data <= conv_std_logic_vector(630,11);
      WHEN "110011100" => data <= conv_std_logic_vector(628,11);
      WHEN "110011101" => data <= conv_std_logic_vector(627,11);
      WHEN "110011110" => data <= conv_std_logic_vector(625,11);
      WHEN "110011111" => data <= conv_std_logic_vector(624,11);
      WHEN "110100000" => data <= conv_std_logic_vector(623,11);
      WHEN "110100001" => data <= conv_std_logic_vector(621,11);
      WHEN "110100010" => data <= conv_std_logic_vector(620,11);
      WHEN "110100011" => data <= conv_std_logic_vector(619,11);
      WHEN "110100100" => data <= conv_std_logic_vector(617,11);
      WHEN "110100101" => data <= conv_std_logic_vector(616,11);
      WHEN "110100110" => data <= conv_std_logic_vector(615,11);
      WHEN "110100111" => data <= conv_std_logic_vector(613,11);
      WHEN "110101000" => data <= conv_std_logic_vector(612,11);
      WHEN "110101001" => data <= conv_std_logic_vector(611,11);
      WHEN "110101010" => data <= conv_std_logic_vector(610,11);
      WHEN "110101011" => data <= conv_std_logic_vector(608,11);
      WHEN "110101100" => data <= conv_std_logic_vector(607,11);
      WHEN "110101101" => data <= conv_std_logic_vector(606,11);
      WHEN "110101110" => data <= conv_std_logic_vector(604,11);
      WHEN "110101111" => data <= conv_std_logic_vector(603,11);
      WHEN "110110000" => data <= conv_std_logic_vector(602,11);
      WHEN "110110001" => data <= conv_std_logic_vector(601,11);
      WHEN "110110010" => data <= conv_std_logic_vector(599,11);
      WHEN "110110011" => data <= conv_std_logic_vector(598,11);
      WHEN "110110100" => data <= conv_std_logic_vector(597,11);
      WHEN "110110101" => data <= conv_std_logic_vector(595,11);
      WHEN "110110110" => data <= conv_std_logic_vector(594,11);
      WHEN "110110111" => data <= conv_std_logic_vector(593,11);
      WHEN "110111000" => data <= conv_std_logic_vector(592,11);
      WHEN "110111001" => data <= conv_std_logic_vector(591,11);
      WHEN "110111010" => data <= conv_std_logic_vector(589,11);
      WHEN "110111011" => data <= conv_std_logic_vector(588,11);
      WHEN "110111100" => data <= conv_std_logic_vector(587,11);
      WHEN "110111101" => data <= conv_std_logic_vector(586,11);
      WHEN "110111110" => data <= conv_std_logic_vector(584,11);
      WHEN "110111111" => data <= conv_std_logic_vector(583,11);
      WHEN "111000000" => data <= conv_std_logic_vector(582,11);
      WHEN "111000001" => data <= conv_std_logic_vector(581,11);
      WHEN "111000010" => data <= conv_std_logic_vector(580,11);
      WHEN "111000011" => data <= conv_std_logic_vector(578,11);
      WHEN "111000100" => data <= conv_std_logic_vector(577,11);
      WHEN "111000101" => data <= conv_std_logic_vector(576,11);
      WHEN "111000110" => data <= conv_std_logic_vector(575,11);
      WHEN "111000111" => data <= conv_std_logic_vector(574,11);
      WHEN "111001000" => data <= conv_std_logic_vector(572,11);
      WHEN "111001001" => data <= conv_std_logic_vector(571,11);
      WHEN "111001010" => data <= conv_std_logic_vector(570,11);
      WHEN "111001011" => data <= conv_std_logic_vector(569,11);
      WHEN "111001100" => data <= conv_std_logic_vector(568,11);
      WHEN "111001101" => data <= conv_std_logic_vector(566,11);
      WHEN "111001110" => data <= conv_std_logic_vector(565,11);
      WHEN "111001111" => data <= conv_std_logic_vector(564,11);
      WHEN "111010000" => data <= conv_std_logic_vector(563,11);
      WHEN "111010001" => data <= conv_std_logic_vector(562,11);
      WHEN "111010010" => data <= conv_std_logic_vector(561,11);
      WHEN "111010011" => data <= conv_std_logic_vector(560,11);
      WHEN "111010100" => data <= conv_std_logic_vector(558,11);
      WHEN "111010101" => data <= conv_std_logic_vector(557,11);
      WHEN "111010110" => data <= conv_std_logic_vector(556,11);
      WHEN "111010111" => data <= conv_std_logic_vector(555,11);
      WHEN "111011000" => data <= conv_std_logic_vector(554,11);
      WHEN "111011001" => data <= conv_std_logic_vector(553,11);
      WHEN "111011010" => data <= conv_std_logic_vector(552,11);
      WHEN "111011011" => data <= conv_std_logic_vector(551,11);
      WHEN "111011100" => data <= conv_std_logic_vector(549,11);
      WHEN "111011101" => data <= conv_std_logic_vector(548,11);
      WHEN "111011110" => data <= conv_std_logic_vector(547,11);
      WHEN "111011111" => data <= conv_std_logic_vector(546,11);
      WHEN "111100000" => data <= conv_std_logic_vector(545,11);
      WHEN "111100001" => data <= conv_std_logic_vector(544,11);
      WHEN "111100010" => data <= conv_std_logic_vector(543,11);
      WHEN "111100011" => data <= conv_std_logic_vector(542,11);
      WHEN "111100100" => data <= conv_std_logic_vector(541,11);
      WHEN "111100101" => data <= conv_std_logic_vector(540,11);
      WHEN "111100110" => data <= conv_std_logic_vector(538,11);
      WHEN "111100111" => data <= conv_std_logic_vector(537,11);
      WHEN "111101000" => data <= conv_std_logic_vector(536,11);
      WHEN "111101001" => data <= conv_std_logic_vector(535,11);
      WHEN "111101010" => data <= conv_std_logic_vector(534,11);
      WHEN "111101011" => data <= conv_std_logic_vector(533,11);
      WHEN "111101100" => data <= conv_std_logic_vector(532,11);
      WHEN "111101101" => data <= conv_std_logic_vector(531,11);
      WHEN "111101110" => data <= conv_std_logic_vector(530,11);
      WHEN "111101111" => data <= conv_std_logic_vector(529,11);
      WHEN "111110000" => data <= conv_std_logic_vector(528,11);
      WHEN "111110001" => data <= conv_std_logic_vector(527,11);
      WHEN "111110010" => data <= conv_std_logic_vector(526,11);
      WHEN "111110011" => data <= conv_std_logic_vector(525,11);
      WHEN "111110100" => data <= conv_std_logic_vector(524,11);
      WHEN "111110101" => data <= conv_std_logic_vector(523,11);
      WHEN "111110110" => data <= conv_std_logic_vector(522,11);
      WHEN "111110111" => data <= conv_std_logic_vector(521,11);
      WHEN "111111000" => data <= conv_std_logic_vector(520,11);
      WHEN "111111001" => data <= conv_std_logic_vector(519,11);
      WHEN "111111010" => data <= conv_std_logic_vector(518,11);
      WHEN "111111011" => data <= conv_std_logic_vector(517,11);
      WHEN "111111100" => data <= conv_std_logic_vector(516,11);
      WHEN "111111101" => data <= conv_std_logic_vector(515,11);
      WHEN "111111110" => data <= conv_std_logic_vector(514,11);
      WHEN "111111111" => data <= conv_std_logic_vector(513,11);
      WHEN others => data <= conv_std_logic_vector(0,11);
    END CASE;
  END PROCESS;

END rtl;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   SINGLE PRECISION DIVIDER - OUTPUT STAGE   ***
--***                                             ***
--***   FP_DIVRND.VHD                             ***
--***                                             ***
--***   Function: Output Stage, Rounding          ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes: Latency = 2                          ***
--***************************************************

ENTITY fp_divrnd IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentdiv : IN STD_LOGIC_VECTOR (10 DOWNTO 1);
      mantissadiv : IN STD_LOGIC_VECTOR (24 DOWNTO 1); -- includes roundbit
      nanin : IN STD_LOGIC;
      dividebyzeroin : IN STD_LOGIC;

		signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
      --------------------------------------------------
      nanout : OUT STD_LOGIC;
      invalidout : OUT STD_LOGIC;
      dividebyzeroout : OUT STD_LOGIC
		);
END fp_divrnd;

ARCHITECTURE rtl OF fp_divrnd IS
  
  constant expwidth : positive := 8;
  constant manwidth : positive := 23;

  signal zerovec : STD_LOGIC_VECTOR (manwidth-1 DOWNTO 1);
  signal signff : STD_LOGIC_VECTOR (2 DOWNTO 1);
  signal nanff : STD_LOGIC_VECTOR (2 DOWNTO 1);
  signal dividebyzeroff : STD_LOGIC_VECTOR (2 DOWNTO 1);  
  signal roundmantissaff, mantissaff : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal exponentnode : STD_LOGIC_VECTOR (expwidth+2 DOWNTO 1);
  signal exponentoneff : STD_LOGIC_VECTOR (expwidth+2 DOWNTO 1);
  signal exponenttwoff : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal overflowbitff : STD_LOGIC;
  signal manoverflow : STD_LOGIC_VECTOR (manwidth+1 DOWNTO 1);
  
  signal infinitygen : STD_LOGIC_VECTOR (expwidth+1 DOWNTO 1);
  signal zerogen : STD_LOGIC_VECTOR (expwidth+1 DOWNTO 1);  
  signal setmanzero, setmanmax : STD_LOGIC;
  signal setexpzero, setexpmax : STD_LOGIC;
  signal setmanzeroff, setmanmaxff : STD_LOGIC;
  signal setexpzeroff, setexpmaxff : STD_LOGIC;

BEGIN
    
  gzv: FOR k IN 1 TO manwidth-1 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  pra: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN
        
      signff <= "00";
      nanff <= "00";
      dividebyzeroff <= "00";
      FOR k IN 1 TO manwidth LOOP
        roundmantissaff(k) <= '0';
        mantissaff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth+2 LOOP
        exponentoneff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        exponenttwoff(k) <= '0';
      END LOOP;
      overflowbitff <= '0';
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF(enable = '1') THEN 
      
        signff(1) <= signin;
        signff(2) <= signff(1);
        nanff(1) <= nanin;
        nanff(2) <= nanff(1);
        dividebyzeroff(1) <= dividebyzeroin;
        dividebyzeroff(2) <= dividebyzeroff(1);
        
        roundmantissaff <= mantissadiv(manwidth+1 DOWNTO 2) + (zerovec & mantissadiv(1));
        
        overflowbitff <= manoverflow(manwidth+1);
        
        -- nan takes precedence (set max)
        -- nan takes precedence (set max)  
        FOR k IN 1 TO manwidth LOOP
          mantissaff(k) <= (roundmantissaff(k) AND setmanzero) OR setmanmax;
        END LOOP;
        
        exponentoneff(expwidth+2 DOWNTO 1) <= exponentdiv(expwidth+2 DOWNTO 1);                 
        FOR k IN 1 TO expwidth LOOP
          exponenttwoff(k) <= (exponentnode(k) AND setexpzero) OR setexpmax;
        END LOOP;
      
      END IF;
             
    END IF;
      
  END PROCESS;

  exponentnode <= exponentoneff(expwidth+2 DOWNTO 1) + 
                 (zerovec(expwidth+1 DOWNTO 1) & overflowbitff);
                 
--*********************************
--*** PREDICT MANTISSA OVERFLOW ***   
--*********************************
     
  manoverflow(1) <= mantissadiv(1);
  gmoa: FOR k IN 2 TO manwidth+1 GENERATE
    manoverflow(k) <= manoverflow(k-1) AND mantissadiv(k);
  END GENERATE; 
                                                                 
--**********************************
--*** CHECK GENERATED CONDITIONS ***   
--**********************************

  -- infinity if exponent >= 255
  infinitygen(1) <= exponentnode(1);
  gia: FOR k IN 2 TO expwidth GENERATE
    infinitygen(k) <= infinitygen(k-1) AND exponentnode(k);
  END GENERATE;
  infinitygen(expwidth+1) <= infinitygen(expwidth) OR 
                            (exponentnode(expwidth+1) AND 
                             NOT(exponentnode(expwidth+2))); -- ;1' if infinity
                         
  -- zero if exponent <= 0
  zerogen(1) <= exponentnode(1);
  gza: FOR k IN 2 TO expwidth GENERATE
    zerogen(k) <= zerogen(k-1) OR exponentnode(k);
  END GENERATE;
  zerogen(expwidth+1) <= zerogen(expwidth) AND 
                         NOT(exponentnode(expwidth+2)); -- '0' if zero
                    
  -- set mantissa to 0 when infinity or zero condition
  setmanzero <= NOT(infinitygen(expwidth+1)) AND zerogen(expwidth+1) AND NOT(dividebyzeroff(1));
  -- setmantissa to "11..11" when nan
  setmanmax <= nanff(1);
  -- set exponent to 0 when zero condition 
  setexpzero <= zerogen(expwidth+1);
  -- set exponent to "11..11" when nan, infinity, or divide by 0
  setexpmax <= nanff(1) OR infinitygen(expwidth+1) OR dividebyzeroff(1);
                             
--***************
--*** OUTPUTS ***
--***************

  signout <= signff(2);   
  mantissaout <= mantissaff;
  exponentout <= exponenttwoff(expwidth DOWNTO 1); 
  -----------------------------------------------
  nanout <= nanff(2);
  invalidout <= nanff(2);
  dividebyzeroout <= dividebyzeroff(2);

END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   SINGLE PRECISION EXPONENT(e) - TOP LEVEL  ***
--***                                             ***
--***   FP_EXP.VHD                                ***
--***                                             ***
--***   Function: IEEE754 SP EXP()                ***
--***                                             ***
--***   05/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** Latency = 16                                ***
--***************************************************

ENTITY fp_exp IS 
GENERIC (synthesize : integer := 1);
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (23 DOWNTO 1);

		signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
      --------------------------------------------------
      nanout : OUT STD_LOGIC;
      overflowout : OUT STD_LOGIC;
      underflowout : OUT STD_LOGIC
		);
END fp_exp;

ARCHITECTURE rtl OF fp_exp IS
  
  constant expwidth : positive := 8;
  constant manwidth : positive := 23;
  
  constant coredepth : positive := 14;

  signal signinff : STD_LOGIC;
  signal maninff : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal expinff : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal signff : STD_LOGIC_VECTOR (coredepth-1 DOWNTO 1);    
  signal mantissanode : STD_LOGIC_VECTOR (24 DOWNTO 1);
  signal exponentnode : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal rangeerror : STD_LOGIC;
      
  -- conditions
  signal zeroman : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal zeroexp : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal maxexp : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal zeromaninff : STD_LOGIC;
  signal maxexpinff : STD_LOGIC;
  signal naninff : STD_LOGIC;
  signal nanff : STD_LOGIC_VECTOR (coredepth-3 DOWNTO 1);
      
  component fp_exp_core
  GENERIC (synthesize : integer := 1);
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aasgn : IN STD_LOGIC;
        aaman : IN STD_LOGIC_VECTOR (23 DOWNTO 1);
        aaexp : IN STD_LOGIC_VECTOR (8 DOWNTO 1);

        ccman : OUT STD_LOGIC_VECTOR (24 DOWNTO 1);
        ccexp : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
        rangeerror : OUT STD_LOGIC
       );
  end component;
       	
  component fp_exprnd
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        signin : IN STD_LOGIC;
        exponentexp : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
        mantissaexp : IN STD_LOGIC_VECTOR (24 DOWNTO 1);
        nanin : IN STD_LOGIC;
        rangeerror : IN STD_LOGIC;

        exponentout : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
        mantissaout : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
        --------------------------------------------------
        nanout : OUT STD_LOGIC;
        overflowout : OUT STD_LOGIC;
        underflowout : OUT STD_LOGIC
		  );
  end component;
  
BEGIN

  pma: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
  
      signinff <= '0';
      FOR k IN 1 TO manwidth LOOP
        maninff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        expinff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO coredepth-1 LOOP
        signff(k) <= '0';
      END LOOP;
    
    ELSIF (rising_edge(sysclk)) THEN

      IF (enable = '1') THEN
        
        signinff <= signin;
        maninff <= mantissain;
        expinff <= exponentin;

        signff(1) <= signinff;
        FOR k IN 2 TO coredepth-1 LOOP
          signff(k) <= signff(k-1);
        END LOOP;
                                                  
      END IF;
  
    END IF;
  
  END PROCESS;

--********************
--*** CHECK INPUTS ***
--********************

  zeroman(1) <= maninff(1);
  gca: FOR k IN 2 TO manwidth GENERATE
    zeroman(k) <= zeroman(k-1) OR maninff(k);
  END GENERATE; 
  zeroexp(1) <= expinff(1);
  gcb: FOR k IN 2 TO expwidth GENERATE
    zeroexp(k) <= zeroexp(k-1) OR expinff(k);
  END GENERATE;
  maxexp(1) <= expinff(1);
  gcc: FOR k IN 2 TO expwidth GENERATE
    maxexp(k) <= maxexp(k-1) AND expinff(k);
  END GENERATE;

  pcc: PROCESS (sysclk,reset)
  BEGIN
    
    IF (reset = '1') THEN
      
      zeromaninff <= '0';
      maxexpinff <= '0';  
      naninff <= '0';
      FOR k IN 1 TO coredepth-3 LOOP
        nanff(k) <= '0';
      END LOOP;
     
    ELSIF (rising_edge(sysclk)) THEN
            
      IF (enable = '1') THEN
     
        zeromaninff <= zeroman(manwidth);
        maxexpinff <= maxexp(expwidth);
    
        -- zero when man = 0, exp = 0
        -- infinity when man = 0, exp = max
        -- nan when man != 0, exp = max
    
        -- all ffs '1' when condition true
        naninff <= zeromaninff AND maxexpinff;

        -- nan output when nan input
        nanff(1) <= naninff;
        FOR k IN 2 TO coredepth-3 LOOP
          nanff(k) <= nanff(k-1);
        END LOOP;
      
      END IF;
   
    END IF;

  END PROCESS;


--****************
--*** EXP CORE ***
--****************

  expcore: fp_exp_core
  GENERIC MAP (synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aasgn=>signin,aaman=>mantissain,aaexp=>exponentin,
            ccman=>mantissanode,ccexp=>exponentnode,
            rangeerror=>rangeerror);
  
--************************
--*** ROUND AND OUTPUT ***
--************************

  rndout: fp_exprnd
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            signin=>signff(coredepth-1),
            exponentexp=>exponentnode,
            mantissaexp=>mantissanode,
            nanin=>nanff(coredepth-3),
            rangeerror=>rangeerror,

            exponentout=>exponentout,mantissaout=>mantissaout,
            nanout=>nanout,overflowout=>overflowout,underflowout=>underflowout);
              
  signout <= '0';
  
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   SINGLE PRECISION EXPONENT(e) - CORE       ***
--***                                             ***
--***   FP_EXP_CORE.VHD                           ***
--***                                             ***
--***   Function: Single Precision Exponent Core  ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** Latency = 14                                ***
--***************************************************

ENTITY fp_exp_core IS
GENERIC (synthesize : integer := 1);
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      aasgn : IN STD_LOGIC;
      aaman : IN STD_LOGIC_VECTOR (23 DOWNTO 1);
      aaexp : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      
      ccman : OUT STD_LOGIC_VECTOR (24 DOWNTO 1); -- includes round bit
      ccexp : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
      rangeerror : OUT STD_LOGIC
     );
END fp_exp_core;

ARCHITECTURE rtl OF fp_exp_core IS

  -- latency 14
  
  type expcalcfftype IS ARRAY (6 DOWNTO 1) OF STD_LOGIC_VECTOR (8 DOWNTO 1);
  
  signal zerovec : STD_LOGIC_VECTOR (32 DOWNTO 1);
  -- INPUT AND SHIFT STAGE
  signal signff : STD_LOGIC_VECTOR (13 DOWNTO 1);
  signal aamanff, aamandelff : STD_LOGIC_VECTOR (23 DOWNTO 1); 
  signal aaexpff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal selshiftff : STD_LOGIC_VECTOR (2 DOWNTO 1); 
  signal leftshift, rightshift : STD_LOGIC_VECTOR (9 DOWNTO 1);
  signal leftshiftff : STD_LOGIC_VECTOR (7 DOWNTO 1);
  signal rightshiftff : STD_LOGIC_VECTOR (7 DOWNTO 1);
  signal bigexp : STD_LOGIC;
  signal bigexpff : STD_LOGIC_VECTOR(2 DOWNTO 1);
  signal leftff, rightff : STD_LOGIC_VECTOR (32 DOWNTO 1); 
  signal powerff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal fractionalff : STD_LOGIC_VECTOR (25 DOWNTO 1); 
  signal powerbus : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal decimalleft : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal decimalright : STD_LOGIC_VECTOR (7 DOWNTO 1);
  signal fractionalleft, fractionalright : STD_LOGIC_VECTOR (25 DOWNTO 1); 
  signal leftone, rightone : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal lefttwo, righttwo, rightthree : STD_LOGIC_VECTOR (32 DOWNTO 1);
  -- TABLE STAGE
  signal addlutposff, addlutnegff : STD_LOGIC_VECTOR (7 DOWNTO 1);
  signal addlutoneff : STD_LOGIC_VECTOR (7 DOWNTO 1);  
  signal lutposmanff, lutnegmanff : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal lutonemanff : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal lutposexpff, lutnegexpff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal lutoneexpff : STD_LOGIC;
  signal manpos, manneg, manone : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal exppos, expneg : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal expone : STD_LOGIC;
  signal lutmanpowerff, lutmanfractionalff : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal lutexppowerff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal lutexpfractionalff : STD_LOGIC; 
  signal expcalcff : expcalcfftype;
  signal manpowernode, manfractionalnode : STD_LOGIC_VECTOR (32 DOWNTO 1);
  -- MULTIPLY STAGE
  signal manmultone, manmulttwo : STD_LOGIC_VECTOR (32 DOWNTO 1);
  -- RANGE
  signal powercheck : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal rangeff : STD_LOGIC_VECTOR (10 DOWNTO 1);
  -- SERIES STAGE
  signal squareterm : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal scaleterm : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal onesixth : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal cubedterm : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal xtermnode, xterm : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal xxterm, xxxterm : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal seriesoneff, seriesoneterm : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal seriestwoff, seriesterm : STD_LOGIC_VECTOR (32 DOWNTO 1);
  -- NORMALIZE
  signal normshift : STD_LOGIC_VECTOR (2 DOWNTO 1);
  signal mantissaoutff : STD_LOGIC_VECTOR (25 DOWNTO 1);
  signal exponentout, exponentoutff : STD_LOGIC_VECTOR (8 DOWNTO 1);     

  component fp_explutpos 
  PORT (
        address : IN STD_LOGIC_VECTOR (7 DOWNTO 1);
        mantissa : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
        exponent : OUT STD_LOGIC_VECTOR (8 DOWNTO 1)
       );
  end component;
  
  component fp_explutneg 
  PORT (
        address : IN STD_LOGIC_VECTOR (7 DOWNTO 1);
        mantissa : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
        exponent : OUT STD_LOGIC_VECTOR (8 DOWNTO 1)
       );
  end component;
  
  component fp_explut7
  PORT (
        address : IN STD_LOGIC_VECTOR (7 DOWNTO 1);
        mantissa : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
        exponent : OUT STD_LOGIC
       );
  end component;

  component fp_fxmul
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36;
           pipes : positive := 1;
           accuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1); 
      
        result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
       );
  end component;

  component fp_del
  GENERIC (
           width : positive := 64;
           pipes : positive := 2
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
       
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
   end component;  
         
BEGIN
    
  gza: FOR k IN 1 TO 32 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  pin: PROCESS (sysclk,reset)
  BEGIN
  
    IF (reset = '1') THEN
    
      FOR k IN 1 TO 13 LOOP
        signff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 23 LOOP 
        aamanff(k) <= '0';
        aamandelff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 8 LOOP
        aaexpff(k) <= '0';
      END LOOP;
      selshiftff <= "00";
      leftshiftff <= "0000000";
      rightshiftff <= "0000000";
      FOR k IN 1 TO 32 LOOP
        leftff(k) <= '0';
        rightff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 8 LOOP
        powerff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 25 LOOP
        fractionalff(k) <= '0';
      END LOOP;
	  bigexpff <= "00";
     
    ELSIF (rising_edge(sysclk)) THEN
    
      IF (enable = '1') THEN
      
        signff(1) <= aasgn;
        FOR k IN 2 TO 13 LOOP
          signff(k) <= signff(k-1);
        END LOOP;
    
        aamanff <= aaman;  -- level 1
        aamandelff <= aamanff; -- level 2
        
        aaexpff <= aaexp;
    
        selshiftff(1) <= leftshift(9); -- level 2
        selshiftff(2) <= selshiftff(1); -- level 3
            
        leftshiftff <= leftshift(7 DOWNTO 1); -- level 2
        rightshiftff <= rightshift(7 DOWNTO 1); -- level 2
        
        leftff <= lefttwo; -- level 3
        rightff <= rightthree; -- level 3
		-- left barrel shifter overflow is relevent only if using result of left shifted mantissa
		bigexpff(2) <= bigexpff(1) AND NOT (selshiftff(2));
		bigexpff(1) <= bigexp;
        
        -- level 4
        FOR k IN 1 TO 7 LOOP
          powerff(k) <= (decimalleft(k) AND NOT(selshiftff(2))) OR
                        (decimalright(k) AND selshiftff(2));
        END LOOP;
		powerff(8) <= (decimalleft(8) AND NOT(selshiftff(2)));
		-- overflow bit to catch case exp(-127.frac)
        FOR k IN 1 TO 25 LOOP
          fractionalff(k) <= (fractionalleft(k) AND NOT(selshiftff(2))) OR
                             (fractionalright(k) AND selshiftff(2));
        END LOOP;
        
      END IF;
    
    END IF;    
      
  END PROCESS;

  leftshift <= ('0' & aaexpff) - "001111111"; 
  rightshift <= "001111111" - ('0' & aaexpff); 
        
  powerbus <= "0000001" & aamandelff & "00";
  
  decimalleft <= ('0' & leftff(32 DOWNTO 26)) +  ("0000000" & signff(3));
  -- decimalleft may overflow to bit 8 when exp(x), where -128 < x <= -127
  decimalright <= rightff(32 DOWNTO 26) +  ("000000" & signff(3));
  gfa: FOR k IN 1 TO 25 GENERATE
    fractionalleft(k) <= leftff(k) XOR signff(3);
    fractionalright(k) <= rightff(k) XOR signff(3);
  END GENERATE;
  
  --**********************
  --*** BARREL SHIFTER ***
  --**********************
  
  leftone(1) <=  powerbus(1)     AND NOT(leftshiftff(2)) AND NOT(leftshiftff(1));
  leftone(2) <= (powerbus(2)     AND NOT(leftshiftff(2)) AND NOT(leftshiftff(1))) OR
                (powerbus(1)     AND NOT(leftshiftff(2)) AND     leftshiftff(1)); 
  leftone(3) <= (powerbus(3)     AND NOT(leftshiftff(2)) AND NOT(leftshiftff(1))) OR
                (powerbus(2)     AND NOT(leftshiftff(2)) AND     leftshiftff(1)) OR
                (powerbus(1)     AND     leftshiftff(2)  AND NOT(leftshiftff(1))); 
  gla: FOR k IN 4 TO 32 GENERATE
    leftone(k) <= (powerbus(k)   AND NOT(leftshiftff(2)) AND NOT(leftshiftff(1))) OR
                  (powerbus(k-1) AND NOT(leftshiftff(2)) AND     leftshiftff(1)) OR
                  (powerbus(k-2) AND     leftshiftff(2)  AND NOT(leftshiftff(1))) OR
                  (powerbus(k-3) AND     leftshiftff(2)  AND     leftshiftff(1));
  END GENERATE;
             
  glb: FOR k IN 1 TO 4 GENERATE
    lefttwo(k) <=  leftone(k)    AND NOT(leftshiftff(3));
  END GENERATE;
  glc: FOR k IN 5 TO 32 GENERATE
    lefttwo(k) <= (leftone(k)    AND NOT(leftshiftff(3))) OR
                  (leftone(k-4)  AND     leftshiftff(3)); 
  END GENERATE;
  -- has left barrel shifter overflowed? (i.e. leftshiftff >= 7)
  bigexp <= leftshiftff(4) OR leftshiftff(5) OR leftshiftff(6) OR leftshiftff(7) OR
			(leftshiftff(3) AND leftshiftff(2) AND leftshiftff(1));
 
  gra: FOR k IN 1 TO 29 GENERATE
    rightone(k) <= (powerbus(k)   AND NOT(rightshiftff(2)) AND NOT(rightshiftff(1))) OR
                   (powerbus(k+1) AND NOT(rightshiftff(2)) AND     rightshiftff(1)) OR
                   (powerbus(k+2) AND     rightshiftff(2)  AND NOT(rightshiftff(1))) OR
                   (powerbus(k+3) AND     rightshiftff(2)  AND     rightshiftff(1));
  END GENERATE;
  rightone(30) <= (powerbus(30) AND NOT(rightshiftff(2)) AND NOT(rightshiftff(1))) OR
                  (powerbus(31) AND NOT(rightshiftff(2)) AND     rightshiftff(1)) OR
                  (powerbus(32) AND     rightshiftff(2)  AND NOT(rightshiftff(1))); 
  rightone(31) <= (powerbus(31) AND NOT(rightshiftff(2)) AND NOT(rightshiftff(1))) OR
                  (powerbus(32) AND NOT(rightshiftff(2)) AND     rightshiftff(1));
  rightone(32) <=  powerbus(32) AND NOT(rightshiftff(2)) AND NOT(rightshiftff(1));
  
  grb: FOR k IN 1 TO 20 GENERATE
    righttwo(k) <= (rightone(k)    AND NOT(rightshiftff(4)) AND NOT(rightshiftff(3))) OR
                   (rightone(k+4)  AND NOT(rightshiftff(4)) AND     rightshiftff(3)) OR
				   (rightone(k+8)  AND     rightshiftff(4)  AND NOT(rightshiftff(3))) OR
				   (rightone(k+12) AND     rightshiftff(4)  AND     rightshiftff(3));
  END GENERATE;
  grc0: FOR k IN 21 TO 24 GENERATE
    righttwo(k) <= (rightone(k)    AND NOT(rightshiftff(4)) AND NOT(rightshiftff(3))) OR
                   (rightone(k+4)  AND NOT(rightshiftff(4)) AND     rightshiftff(3)) OR
				   (rightone(k+8)  AND     rightshiftff(4)  AND NOT(rightshiftff(3)));
  END GENERATE;
  grc1: FOR k IN 25 TO 28 GENERATE
    righttwo(k) <= (rightone(k)    AND NOT(rightshiftff(4)) AND NOT(rightshiftff(3))) OR
                   (rightone(k+4)  AND NOT(rightshiftff(4)) AND     rightshiftff(3));
  END GENERATE;
  grc2: FOR k IN 29 TO 32 GENERATE
    righttwo(k) <= (rightone(k)    AND NOT(rightshiftff(4)) AND NOT(rightshiftff(3)));
  END GENERATE;

  -- right barrel shifter outputs zero if rightshiftff >= 32
  grd0: FOR k IN 1 TO 16 GENERATE
    rightthree(k) <= ((righttwo(k)    AND NOT(rightshiftff(5))) OR 
                     (righttwo(k+16) AND rightshiftff(5))) AND
					 NOT (rightshiftff(6)) AND NOT(rightshiftff(7));
  END GENERATE;
  grd1: FOR k IN 17 TO 32 GENERATE
    rightthree(k) <= (righttwo(k)    AND NOT(rightshiftff(5))) AND
					   NOT (rightshiftff(6)) AND NOT(rightshiftff(7));
  END GENERATE;
  
  --******************************************
  --*** TABLES - NO RESET, FORCE TO MEMORY ***
  --******************************************
  
  -- level: 4 in, 6 out
  pla: PROCESS (sysclk)
  BEGIN
  
    IF (rising_edge(sysclk)) THEN
        
      IF (enable = '1') THEN
          
        addlutposff <= powerff(7 DOWNTO 1);
        addlutnegff <= powerff(7 DOWNTO 1);
        addlutoneff <= fractionalff(25 DOWNTO 19);
      
        lutposmanff <= manpos;
        lutposexpff <= exppos;
        lutnegmanff <= manneg;
        lutnegexpff <= expneg;
        lutonemanff <= manone;
        lutoneexpff <= expone;
            
      END IF;
      
    END IF;
  
  END PROCESS;
 
  declut: fp_explutpos
  PORT MAP (address=>addlutposff,
            mantissa=>manpos,exponent=>exppos);
            
  neglut: fp_explutneg
  PORT MAP (address=>addlutnegff,
            mantissa=>manneg,exponent=>expneg);
                     
  fraclut: fp_explut7
  PORT MAP (address=>addlutoneff,
            mantissa=>manone,exponent=>expone);
  
  -- level: 6 in, 7 out
  pma: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
    
      FOR k IN 1 TO 23 LOOP
        lutmanpowerff(k) <= '0';
        lutmanfractionalff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 8 LOOP
        lutexppowerff(k) <= '0';
      END LOOP;
      lutexpfractionalff <= '0';
      
      FOR k IN 1 TO 6 LOOP
        expcalcff(k)(8 DOWNTO 1) <= "00000000";
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
        
      IF (enable = '1') THEN
          
        FOR k IN 1 TO 23 LOOP
          lutmanpowerff(k) <= (lutposmanff(k) AND NOT(signff(6))) OR (lutnegmanff(k) AND signff(6));
        END LOOP;
        lutmanfractionalff <= lutonemanff;
        FOR k IN 1 TO 8 LOOP
          lutexppowerff(k) <= (lutposexpff(k) AND NOT(signff(6))) OR (lutnegexpff(k) AND signff(6));
        END LOOP;
        lutexpfractionalff <= lutoneexpff;
        
        -- level: 7 in, 13 out
        expcalcff(1)(8 DOWNTO 1) <= lutexppowerff + ("0000000" & lutexpfractionalff);
        FOR k IN 2 TO 6 LOOP
          expcalcff(k)(8 DOWNTO 1) <= expcalcff(k-1)(8 DOWNTO 1);
        END LOOP;
            
      END IF;
      
    END IF;
          
  END PROCESS;  
  
  manpowernode(32) <= '1';
  manpowernode(31 DOWNTO 9) <= lutmanpowerff;
  manpowernode(8 DOWNTO 1) <= "00000000";
 
  manfractionalnode(32) <= '1';
  manfractionalnode(31 DOWNTO 9) <= lutmanfractionalff;
  manfractionalnode(8 DOWNTO 1) <= "00000000"; 
  
  --*************************************
  --*** MULTIPLY ALL EXP(X) SUBRANGES ***
  --*************************************
  
  -- level 7 in, 10 out
  mulone: fp_fxmul
  GENERIC MAP (widthaa=>32,widthbb=>32,widthcc=>32,
               pipes=>3,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>manpowernode,databb=>manfractionalnode,
            result=>manmultone);

  -- level 10 in, 13 out
  multwo: fp_fxmul
  GENERIC MAP (widthaa=>32,widthbb=>32,widthcc=>32,
               pipes=>3,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>manmultone,databb=>seriesterm,
            result=>manmulttwo);
            
  --**************************************
  --*** PREDICT OVERFLOW AND UNDERFLOW ***
  --**************************************
  
  -- overflow or underflow if power > 88
  -- overflow or underflow if power != 0 and explut = 0
  
  powercheck <= powerff - "01011001";  -- 89
  
  -- level 4 in, level 14 out
  ppca: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
    
      FOR k IN 1 TO 10 LOOP
        rangeff(k) <= '0';
      END LOOP;
    
    ELSIF (rising_edge(sysclk)) THEN
        
      IF (enable = '1') THEN
       
         rangeff(1) <= bigexpff(2) OR NOT(powercheck(8));
		 -- if left barrel shifter has overflowed, or abs(x) >= 89 then exp(x) -> 0 or Inf
         FOR k IN 2 TO 9 LOOP
           rangeff(k) <= rangeff(k-1);
         END LOOP;
		 rangeff(10) <= rangeff(9) AND NOT(signff(13));
		 -- exp(x) can only overflow if x was positive
       
      END IF;
      
    END IF;
          
  END PROCESS;
  
  --***********************
  --*** TAYLOR's SERIES ***
  --***********************
  
  --*** calculate lowest 18 bits ***
  -- sequence is 1 + x + x^2/2 + x^3/6 + x^4/24
  -- x*x/2 term is (7+7+1=15 bits down)
  -- x*x*x/6 is (7+7+7+2=23 bits) down
  
  -- level 4 in, 6 out
  mulsqr: fp_fxmul
  GENERIC MAP (widthaa=>18,widthbb=>18,widthcc=>18,
               pipes=>2,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>fractionalff(18 DOWNTO 1),
            databb=>fractionalff(18 DOWNTO 1),
            result=>squareterm);  
  
  -- level 4 in, 6 out
  mulscl: fp_fxmul
  GENERIC MAP (widthaa=>18,widthbb=>18,widthcc=>18,
               pipes=>2,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>fractionalff(18 DOWNTO 1),
            databb=>onesixth,
            result=>scaleterm); 
                      
  onesixth <= "001010101010101011";
  
  -- level 6 in, 8 out
  mulcub: fp_fxmul
  GENERIC MAP (widthaa=>18,widthbb=>18,widthcc=>18,
               pipes=>2,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>squareterm,
            databb=>scaleterm,
            result=>cubedterm);
       
  xtermnode <= "10000000" & fractionalff(18 DOWNTO 1) & "000000"; -- '1' + x term   
  xxterm <= (zerovec(16 DOWNTO 1) & squareterm(18 DOWNTO 3));
  xxxterm <= (zerovec(22 DOWNTO 1) & cubedterm(18 DOWNTO 9));
  
  -- level 4 in, level 6 out
  delone: fp_del
  GENERIC MAP (width=>32,pipes=>2)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>xtermnode,cc=>xterm);
            
  -- level 7 in, level 8 out
  deltwo: fp_del
  GENERIC MAP (width=>32,pipes=>1)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>seriesoneff,cc=>seriesoneterm);
    
  ptsa: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
    
      FOR k IN 1 TO 32 LOOP
        seriesoneff(k) <= '0';
        seriestwoff(k) <= '0';
      END LOOP;
 
      
    ELSIF (rising_edge(sysclk)) THEN
        
      IF (enable = '1') THEN
          
        seriesoneff <= xterm + xxterm; -- level 7
        seriestwoff <= seriesoneterm + xxxterm; -- level 9
             
      END IF;
      
    END IF;
          
  END PROCESS;            
  
  -- level 9 in, level 10 out
  delthr: fp_del
  GENERIC MAP (width=>32,pipes=>1)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>seriestwoff,cc=>seriesterm);
                      
  --square <= powerfractional(18 DOWNTO 1) * powerfractional(18 DOWNTO 1);
  --scaleterm <= powerfractional(18 DOWNTO 1) * onesixth;
  --onesixth <= "001010101010101011";
  --cubedterm <= square(36 DOWNTO 19) * scaleterm(36 DOWNTO 19);
  --manseries <= ('1' & zerovec(31 DOWNTO 1)) +  -- 1 term
  --             (zerovec(8 DOWNTO 1) & powerfractional(18 DOWNTO 1) & zerovec(6 DOWNTO 1)) + -- x term
  --             (zerovec(16 DOWNTO 1) & square(36 DOWNTO 21)) + 
  --             (zerovec(22 DOWNTO 1) & cubedterm(36 DOWNTO 27));
  --xterm <= (zerovec(7 DOWNTO 1) & powerfractional(18 DOWNTO 1) & zerovec(7 DOWNTO 1));
  --xxterm <= (zerovec(15 DOWNTO 1) & square(36 DOWNTO 20));
  --xxxterm <= (zerovec(21 DOWNTO 1) & cubedterm(36 DOWNTO 26));
  
  --************************
  --*** NORMALIZE OUTPUT ***
  --************************
   
  pns: PROCESS (manmulttwo)
  BEGIN
      
    CASE manmulttwo(32 DOWNTO 30) IS
      WHEN "000" => normshift <= "11";
      WHEN "001" => normshift <= "10";
      WHEN "010" => normshift <= "01";
      WHEN "011" => normshift <= "01";
      WHEN "100" => normshift <= "00";
      WHEN "101" => normshift <= "00";
      WHEN "110" => normshift <= "00";
      WHEN "111" => normshift <= "00"; 
      WHEN others => normshift <= "00";
    END CASE;
        
  END PROCESS;
  
  pna: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
    
      FOR k IN 1 TO 25 LOOP
        mantissaoutff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 8 LOOP
        exponentoutff(k) <= '0';
      END LOOP;
        
 
    ELSIF (rising_edge(sysclk)) THEN
        
      IF (enable = '1') THEN
          
        FOR k IN 1 TO 25 LOOP
          mantissaoutff(k) <= (manmulttwo(k+7) AND NOT(normshift(2)) AND NOT(normshift(1))) OR
                              (manmulttwo(k+6) AND NOT(normshift(2)) AND     normshift(1)) OR
                              (manmulttwo(k+5) AND     normshift(2)  AND NOT(normshift(1))) OR
                              (manmulttwo(k+4) AND     normshift(2)  AND     normshift(1));
        END LOOP;
        -- correction factor of 2 due to two multiplications (double has 3)
        FOR k IN 1 TO 8 LOOP
		  exponentoutff(k) <= exponentout(k) AND NOT(rangeff(9) AND signff(13));
		END LOOP;
		-- set exponent to zero if x = large negative value, exp(x)->0
      END IF;
      
    END IF;
          
  END PROCESS; 
exponentout <= expcalcff(6)(8 DOWNTO 1) - ("000000" & normshift) + "00000010";

  --**************
  --*** OUTPUT ***
  --**************
  
  ccman <= mantissaoutff(24 DOWNTO 1);
  ccexp <= exponentoutff;
  rangeerror <= rangeff(10);
        
END rtl;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_EXPLUT7.VHD                            ***
--***                                             ***
--***   Function: Look Up Table - EXP()           ***
--***                                             ***
--***   Generated by MATLAB Utility               ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_explut7 IS
PORT (
      address : IN STD_LOGIC_VECTOR (7 DOWNTO 1);
      mantissa : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
      exponent : OUT STD_LOGIC
     );
END fp_explut7;

ARCHITECTURE rtl OF fp_explut7 IS

BEGIN

  pca: PROCESS (address)
  BEGIN
    CASE address IS
      WHEN "0000000" =>
            mantissa <= conv_std_logic_vector(0,23);
            exponent <= '0';
      WHEN "0000001" =>
            mantissa <= conv_std_logic_vector(65793,23);
            exponent <= '0';
      WHEN "0000010" =>
            mantissa <= conv_std_logic_vector(132101,23);
            exponent <= '0';
      WHEN "0000011" =>
            mantissa <= conv_std_logic_vector(198930,23);
            exponent <= '0';
      WHEN "0000100" =>
            mantissa <= conv_std_logic_vector(266283,23);
            exponent <= '0';
      WHEN "0000101" =>
            mantissa <= conv_std_logic_vector(334164,23);
            exponent <= '0';
      WHEN "0000110" =>
            mantissa <= conv_std_logic_vector(402578,23);
            exponent <= '0';
      WHEN "0000111" =>
            mantissa <= conv_std_logic_vector(471528,23);
            exponent <= '0';
      WHEN "0001000" =>
            mantissa <= conv_std_logic_vector(541019,23);
            exponent <= '0';
      WHEN "0001001" =>
            mantissa <= conv_std_logic_vector(611055,23);
            exponent <= '0';
      WHEN "0001010" =>
            mantissa <= conv_std_logic_vector(681640,23);
            exponent <= '0';
      WHEN "0001011" =>
            mantissa <= conv_std_logic_vector(752779,23);
            exponent <= '0';
      WHEN "0001100" =>
            mantissa <= conv_std_logic_vector(824476,23);
            exponent <= '0';
      WHEN "0001101" =>
            mantissa <= conv_std_logic_vector(896735,23);
            exponent <= '0';
      WHEN "0001110" =>
            mantissa <= conv_std_logic_vector(969560,23);
            exponent <= '0';
      WHEN "0001111" =>
            mantissa <= conv_std_logic_vector(1042957,23);
            exponent <= '0';
      WHEN "0010000" =>
            mantissa <= conv_std_logic_vector(1116930,23);
            exponent <= '0';
      WHEN "0010001" =>
            mantissa <= conv_std_logic_vector(1191483,23);
            exponent <= '0';
      WHEN "0010010" =>
            mantissa <= conv_std_logic_vector(1266621,23);
            exponent <= '0';
      WHEN "0010011" =>
            mantissa <= conv_std_logic_vector(1342348,23);
            exponent <= '0';
      WHEN "0010100" =>
            mantissa <= conv_std_logic_vector(1418668,23);
            exponent <= '0';
      WHEN "0010101" =>
            mantissa <= conv_std_logic_vector(1495588,23);
            exponent <= '0';
      WHEN "0010110" =>
            mantissa <= conv_std_logic_vector(1573110,23);
            exponent <= '0';
      WHEN "0010111" =>
            mantissa <= conv_std_logic_vector(1651241,23);
            exponent <= '0';
      WHEN "0011000" =>
            mantissa <= conv_std_logic_vector(1729985,23);
            exponent <= '0';
      WHEN "0011001" =>
            mantissa <= conv_std_logic_vector(1809346,23);
            exponent <= '0';
      WHEN "0011010" =>
            mantissa <= conv_std_logic_vector(1889329,23);
            exponent <= '0';
      WHEN "0011011" =>
            mantissa <= conv_std_logic_vector(1969940,23);
            exponent <= '0';
      WHEN "0011100" =>
            mantissa <= conv_std_logic_vector(2051183,23);
            exponent <= '0';
      WHEN "0011101" =>
            mantissa <= conv_std_logic_vector(2133064,23);
            exponent <= '0';
      WHEN "0011110" =>
            mantissa <= conv_std_logic_vector(2215586,23);
            exponent <= '0';
      WHEN "0011111" =>
            mantissa <= conv_std_logic_vector(2298756,23);
            exponent <= '0';
      WHEN "0100000" =>
            mantissa <= conv_std_logic_vector(2382578,23);
            exponent <= '0';
      WHEN "0100001" =>
            mantissa <= conv_std_logic_vector(2467057,23);
            exponent <= '0';
      WHEN "0100010" =>
            mantissa <= conv_std_logic_vector(2552199,23);
            exponent <= '0';
      WHEN "0100011" =>
            mantissa <= conv_std_logic_vector(2638009,23);
            exponent <= '0';
      WHEN "0100100" =>
            mantissa <= conv_std_logic_vector(2724492,23);
            exponent <= '0';
      WHEN "0100101" =>
            mantissa <= conv_std_logic_vector(2811653,23);
            exponent <= '0';
      WHEN "0100110" =>
            mantissa <= conv_std_logic_vector(2899498,23);
            exponent <= '0';
      WHEN "0100111" =>
            mantissa <= conv_std_logic_vector(2988032,23);
            exponent <= '0';
      WHEN "0101000" =>
            mantissa <= conv_std_logic_vector(3077260,23);
            exponent <= '0';
      WHEN "0101001" =>
            mantissa <= conv_std_logic_vector(3167188,23);
            exponent <= '0';
      WHEN "0101010" =>
            mantissa <= conv_std_logic_vector(3257821,23);
            exponent <= '0';
      WHEN "0101011" =>
            mantissa <= conv_std_logic_vector(3349165,23);
            exponent <= '0';
      WHEN "0101100" =>
            mantissa <= conv_std_logic_vector(3441225,23);
            exponent <= '0';
      WHEN "0101101" =>
            mantissa <= conv_std_logic_vector(3534008,23);
            exponent <= '0';
      WHEN "0101110" =>
            mantissa <= conv_std_logic_vector(3627518,23);
            exponent <= '0';
      WHEN "0101111" =>
            mantissa <= conv_std_logic_vector(3721762,23);
            exponent <= '0';
      WHEN "0110000" =>
            mantissa <= conv_std_logic_vector(3816745,23);
            exponent <= '0';
      WHEN "0110001" =>
            mantissa <= conv_std_logic_vector(3912472,23);
            exponent <= '0';
      WHEN "0110010" =>
            mantissa <= conv_std_logic_vector(4008951,23);
            exponent <= '0';
      WHEN "0110011" =>
            mantissa <= conv_std_logic_vector(4106186,23);
            exponent <= '0';
      WHEN "0110100" =>
            mantissa <= conv_std_logic_vector(4204184,23);
            exponent <= '0';
      WHEN "0110101" =>
            mantissa <= conv_std_logic_vector(4302951,23);
            exponent <= '0';
      WHEN "0110110" =>
            mantissa <= conv_std_logic_vector(4402492,23);
            exponent <= '0';
      WHEN "0110111" =>
            mantissa <= conv_std_logic_vector(4502814,23);
            exponent <= '0';
      WHEN "0111000" =>
            mantissa <= conv_std_logic_vector(4603922,23);
            exponent <= '0';
      WHEN "0111001" =>
            mantissa <= conv_std_logic_vector(4705824,23);
            exponent <= '0';
      WHEN "0111010" =>
            mantissa <= conv_std_logic_vector(4808525,23);
            exponent <= '0';
      WHEN "0111011" =>
            mantissa <= conv_std_logic_vector(4912031,23);
            exponent <= '0';
      WHEN "0111100" =>
            mantissa <= conv_std_logic_vector(5016349,23);
            exponent <= '0';
      WHEN "0111101" =>
            mantissa <= conv_std_logic_vector(5121486,23);
            exponent <= '0';
      WHEN "0111110" =>
            mantissa <= conv_std_logic_vector(5227447,23);
            exponent <= '0';
      WHEN "0111111" =>
            mantissa <= conv_std_logic_vector(5334239,23);
            exponent <= '0';
      WHEN "1000000" =>
            mantissa <= conv_std_logic_vector(5441868,23);
            exponent <= '0';
      WHEN "1000001" =>
            mantissa <= conv_std_logic_vector(5550342,23);
            exponent <= '0';
      WHEN "1000010" =>
            mantissa <= conv_std_logic_vector(5659667,23);
            exponent <= '0';
      WHEN "1000011" =>
            mantissa <= conv_std_logic_vector(5769849,23);
            exponent <= '0';
      WHEN "1000100" =>
            mantissa <= conv_std_logic_vector(5880895,23);
            exponent <= '0';
      WHEN "1000101" =>
            mantissa <= conv_std_logic_vector(5992812,23);
            exponent <= '0';
      WHEN "1000110" =>
            mantissa <= conv_std_logic_vector(6105607,23);
            exponent <= '0';
      WHEN "1000111" =>
            mantissa <= conv_std_logic_vector(6219286,23);
            exponent <= '0';
      WHEN "1001000" =>
            mantissa <= conv_std_logic_vector(6333858,23);
            exponent <= '0';
      WHEN "1001001" =>
            mantissa <= conv_std_logic_vector(6449327,23);
            exponent <= '0';
      WHEN "1001010" =>
            mantissa <= conv_std_logic_vector(6565703,23);
            exponent <= '0';
      WHEN "1001011" =>
            mantissa <= conv_std_logic_vector(6682991,23);
            exponent <= '0';
      WHEN "1001100" =>
            mantissa <= conv_std_logic_vector(6801199,23);
            exponent <= '0';
      WHEN "1001101" =>
            mantissa <= conv_std_logic_vector(6920334,23);
            exponent <= '0';
      WHEN "1001110" =>
            mantissa <= conv_std_logic_vector(7040403,23);
            exponent <= '0';
      WHEN "1001111" =>
            mantissa <= conv_std_logic_vector(7161415,23);
            exponent <= '0';
      WHEN "1010000" =>
            mantissa <= conv_std_logic_vector(7283375,23);
            exponent <= '0';
      WHEN "1010001" =>
            mantissa <= conv_std_logic_vector(7406292,23);
            exponent <= '0';
      WHEN "1010010" =>
            mantissa <= conv_std_logic_vector(7530173,23);
            exponent <= '0';
      WHEN "1010011" =>
            mantissa <= conv_std_logic_vector(7655025,23);
            exponent <= '0';
      WHEN "1010100" =>
            mantissa <= conv_std_logic_vector(7780857,23);
            exponent <= '0';
      WHEN "1010101" =>
            mantissa <= conv_std_logic_vector(7907676,23);
            exponent <= '0';
      WHEN "1010110" =>
            mantissa <= conv_std_logic_vector(8035489,23);
            exponent <= '0';
      WHEN "1010111" =>
            mantissa <= conv_std_logic_vector(8164305,23);
            exponent <= '0';
      WHEN "1011000" =>
            mantissa <= conv_std_logic_vector(8294131,23);
            exponent <= '0';
      WHEN "1011001" =>
            mantissa <= conv_std_logic_vector(18184,23);
            exponent <= '1';
      WHEN "1011010" =>
            mantissa <= conv_std_logic_vector(84119,23);
            exponent <= '1';
      WHEN "1011011" =>
            mantissa <= conv_std_logic_vector(150571,23);
            exponent <= '1';
      WHEN "1011100" =>
            mantissa <= conv_std_logic_vector(217545,23);
            exponent <= '1';
      WHEN "1011101" =>
            mantissa <= conv_std_logic_vector(285044,23);
            exponent <= '1';
      WHEN "1011110" =>
            mantissa <= conv_std_logic_vector(353072,23);
            exponent <= '1';
      WHEN "1011111" =>
            mantissa <= conv_std_logic_vector(421634,23);
            exponent <= '1';
      WHEN "1100000" =>
            mantissa <= conv_std_logic_vector(490734,23);
            exponent <= '1';
      WHEN "1100001" =>
            mantissa <= conv_std_logic_vector(560375,23);
            exponent <= '1';
      WHEN "1100010" =>
            mantissa <= conv_std_logic_vector(630563,23);
            exponent <= '1';
      WHEN "1100011" =>
            mantissa <= conv_std_logic_vector(701301,23);
            exponent <= '1';
      WHEN "1100100" =>
            mantissa <= conv_std_logic_vector(772594,23);
            exponent <= '1';
      WHEN "1100101" =>
            mantissa <= conv_std_logic_vector(844446,23);
            exponent <= '1';
      WHEN "1100110" =>
            mantissa <= conv_std_logic_vector(916862,23);
            exponent <= '1';
      WHEN "1100111" =>
            mantissa <= conv_std_logic_vector(989846,23);
            exponent <= '1';
      WHEN "1101000" =>
            mantissa <= conv_std_logic_vector(1063402,23);
            exponent <= '1';
      WHEN "1101001" =>
            mantissa <= conv_std_logic_vector(1137535,23);
            exponent <= '1';
      WHEN "1101010" =>
            mantissa <= conv_std_logic_vector(1212249,23);
            exponent <= '1';
      WHEN "1101011" =>
            mantissa <= conv_std_logic_vector(1287550,23);
            exponent <= '1';
      WHEN "1101100" =>
            mantissa <= conv_std_logic_vector(1363441,23);
            exponent <= '1';
      WHEN "1101101" =>
            mantissa <= conv_std_logic_vector(1439927,23);
            exponent <= '1';
      WHEN "1101110" =>
            mantissa <= conv_std_logic_vector(1517013,23);
            exponent <= '1';
      WHEN "1101111" =>
            mantissa <= conv_std_logic_vector(1594704,23);
            exponent <= '1';
      WHEN "1110000" =>
            mantissa <= conv_std_logic_vector(1673004,23);
            exponent <= '1';
      WHEN "1110001" =>
            mantissa <= conv_std_logic_vector(1751918,23);
            exponent <= '1';
      WHEN "1110010" =>
            mantissa <= conv_std_logic_vector(1831452,23);
            exponent <= '1';
      WHEN "1110011" =>
            mantissa <= conv_std_logic_vector(1911608,23);
            exponent <= '1';
      WHEN "1110100" =>
            mantissa <= conv_std_logic_vector(1992394,23);
            exponent <= '1';
      WHEN "1110101" =>
            mantissa <= conv_std_logic_vector(2073813,23);
            exponent <= '1';
      WHEN "1110110" =>
            mantissa <= conv_std_logic_vector(2155871,23);
            exponent <= '1';
      WHEN "1110111" =>
            mantissa <= conv_std_logic_vector(2238572,23);
            exponent <= '1';
      WHEN "1111000" =>
            mantissa <= conv_std_logic_vector(2321922,23);
            exponent <= '1';
      WHEN "1111001" =>
            mantissa <= conv_std_logic_vector(2405926,23);
            exponent <= '1';
      WHEN "1111010" =>
            mantissa <= conv_std_logic_vector(2490589,23);
            exponent <= '1';
      WHEN "1111011" =>
            mantissa <= conv_std_logic_vector(2575915,23);
            exponent <= '1';
      WHEN "1111100" =>
            mantissa <= conv_std_logic_vector(2661911,23);
            exponent <= '1';
      WHEN "1111101" =>
            mantissa <= conv_std_logic_vector(2748582,23);
            exponent <= '1';
      WHEN "1111110" =>
            mantissa <= conv_std_logic_vector(2835932,23);
            exponent <= '1';
      WHEN "1111111" =>
            mantissa <= conv_std_logic_vector(2923967,23);
            exponent <= '1';
      WHEN others =>
           mantissa <= conv_std_logic_vector(0,23);
           exponent <= '0';
    END CASE;
  END PROCESS;

END rtl;
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_EXPLUT8.VHD                            ***
--***                                             ***
--***   Function: Look Up Table - EXP()           ***
--***                                             ***
--***   Generated by MATLAB Utility               ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_explut8 IS
PORT (
      address : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissa : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
      exponent : OUT STD_LOGIC_VECTOR (8 DOWNTO 1)
     );
END fp_explut8;

ARCHITECTURE rtl OF fp_explut8 IS

BEGIN

  pca: PROCESS (address)
  BEGIN
    CASE address IS
      WHEN "00000000" =>
            mantissa <= conv_std_logic_vector(0,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00000001" =>
            mantissa <= conv_std_logic_vector(32832,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00000010" =>
            mantissa <= conv_std_logic_vector(65793,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00000011" =>
            mantissa <= conv_std_logic_vector(98882,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00000100" =>
            mantissa <= conv_std_logic_vector(132101,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00000101" =>
            mantissa <= conv_std_logic_vector(165450,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00000110" =>
            mantissa <= conv_std_logic_vector(198930,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00000111" =>
            mantissa <= conv_std_logic_vector(232541,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00001000" =>
            mantissa <= conv_std_logic_vector(266283,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00001001" =>
            mantissa <= conv_std_logic_vector(300157,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00001010" =>
            mantissa <= conv_std_logic_vector(334164,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00001011" =>
            mantissa <= conv_std_logic_vector(368304,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00001100" =>
            mantissa <= conv_std_logic_vector(402578,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00001101" =>
            mantissa <= conv_std_logic_vector(436985,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00001110" =>
            mantissa <= conv_std_logic_vector(471528,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00001111" =>
            mantissa <= conv_std_logic_vector(506205,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00010000" =>
            mantissa <= conv_std_logic_vector(541019,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00010001" =>
            mantissa <= conv_std_logic_vector(575968,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00010010" =>
            mantissa <= conv_std_logic_vector(611055,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00010011" =>
            mantissa <= conv_std_logic_vector(646278,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00010100" =>
            mantissa <= conv_std_logic_vector(681640,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00010101" =>
            mantissa <= conv_std_logic_vector(717140,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00010110" =>
            mantissa <= conv_std_logic_vector(752779,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00010111" =>
            mantissa <= conv_std_logic_vector(788557,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00011000" =>
            mantissa <= conv_std_logic_vector(824476,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00011001" =>
            mantissa <= conv_std_logic_vector(860535,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00011010" =>
            mantissa <= conv_std_logic_vector(896735,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00011011" =>
            mantissa <= conv_std_logic_vector(933076,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00011100" =>
            mantissa <= conv_std_logic_vector(969560,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00011101" =>
            mantissa <= conv_std_logic_vector(1006187,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00011110" =>
            mantissa <= conv_std_logic_vector(1042957,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00011111" =>
            mantissa <= conv_std_logic_vector(1079872,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00100000" =>
            mantissa <= conv_std_logic_vector(1116930,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00100001" =>
            mantissa <= conv_std_logic_vector(1154134,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00100010" =>
            mantissa <= conv_std_logic_vector(1191483,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00100011" =>
            mantissa <= conv_std_logic_vector(1228978,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00100100" =>
            mantissa <= conv_std_logic_vector(1266621,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00100101" =>
            mantissa <= conv_std_logic_vector(1304410,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00100110" =>
            mantissa <= conv_std_logic_vector(1342348,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00100111" =>
            mantissa <= conv_std_logic_vector(1380433,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00101000" =>
            mantissa <= conv_std_logic_vector(1418668,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00101001" =>
            mantissa <= conv_std_logic_vector(1457053,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00101010" =>
            mantissa <= conv_std_logic_vector(1495588,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00101011" =>
            mantissa <= conv_std_logic_vector(1534273,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00101100" =>
            mantissa <= conv_std_logic_vector(1573110,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00101101" =>
            mantissa <= conv_std_logic_vector(1612100,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00101110" =>
            mantissa <= conv_std_logic_vector(1651241,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00101111" =>
            mantissa <= conv_std_logic_vector(1690536,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00110000" =>
            mantissa <= conv_std_logic_vector(1729985,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00110001" =>
            mantissa <= conv_std_logic_vector(1769588,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00110010" =>
            mantissa <= conv_std_logic_vector(1809346,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00110011" =>
            mantissa <= conv_std_logic_vector(1849259,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00110100" =>
            mantissa <= conv_std_logic_vector(1889329,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00110101" =>
            mantissa <= conv_std_logic_vector(1929556,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00110110" =>
            mantissa <= conv_std_logic_vector(1969940,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00110111" =>
            mantissa <= conv_std_logic_vector(2010482,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00111000" =>
            mantissa <= conv_std_logic_vector(2051183,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00111001" =>
            mantissa <= conv_std_logic_vector(2092044,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00111010" =>
            mantissa <= conv_std_logic_vector(2133064,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00111011" =>
            mantissa <= conv_std_logic_vector(2174244,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00111100" =>
            mantissa <= conv_std_logic_vector(2215586,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00111101" =>
            mantissa <= conv_std_logic_vector(2257090,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00111110" =>
            mantissa <= conv_std_logic_vector(2298756,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "00111111" =>
            mantissa <= conv_std_logic_vector(2340585,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01000000" =>
            mantissa <= conv_std_logic_vector(2382578,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01000001" =>
            mantissa <= conv_std_logic_vector(2424735,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01000010" =>
            mantissa <= conv_std_logic_vector(2467057,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01000011" =>
            mantissa <= conv_std_logic_vector(2509545,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01000100" =>
            mantissa <= conv_std_logic_vector(2552199,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01000101" =>
            mantissa <= conv_std_logic_vector(2595020,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01000110" =>
            mantissa <= conv_std_logic_vector(2638009,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01000111" =>
            mantissa <= conv_std_logic_vector(2681166,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01001000" =>
            mantissa <= conv_std_logic_vector(2724492,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01001001" =>
            mantissa <= conv_std_logic_vector(2767987,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01001010" =>
            mantissa <= conv_std_logic_vector(2811653,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01001011" =>
            mantissa <= conv_std_logic_vector(2855490,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01001100" =>
            mantissa <= conv_std_logic_vector(2899498,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01001101" =>
            mantissa <= conv_std_logic_vector(2943678,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01001110" =>
            mantissa <= conv_std_logic_vector(2988032,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01001111" =>
            mantissa <= conv_std_logic_vector(3032559,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01010000" =>
            mantissa <= conv_std_logic_vector(3077260,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01010001" =>
            mantissa <= conv_std_logic_vector(3122136,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01010010" =>
            mantissa <= conv_std_logic_vector(3167188,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01010011" =>
            mantissa <= conv_std_logic_vector(3212416,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01010100" =>
            mantissa <= conv_std_logic_vector(3257821,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01010101" =>
            mantissa <= conv_std_logic_vector(3303404,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01010110" =>
            mantissa <= conv_std_logic_vector(3349165,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01010111" =>
            mantissa <= conv_std_logic_vector(3395105,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01011000" =>
            mantissa <= conv_std_logic_vector(3441225,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01011001" =>
            mantissa <= conv_std_logic_vector(3487526,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01011010" =>
            mantissa <= conv_std_logic_vector(3534008,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01011011" =>
            mantissa <= conv_std_logic_vector(3580672,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01011100" =>
            mantissa <= conv_std_logic_vector(3627518,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01011101" =>
            mantissa <= conv_std_logic_vector(3674548,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01011110" =>
            mantissa <= conv_std_logic_vector(3721762,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01011111" =>
            mantissa <= conv_std_logic_vector(3769160,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01100000" =>
            mantissa <= conv_std_logic_vector(3816745,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01100001" =>
            mantissa <= conv_std_logic_vector(3864515,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01100010" =>
            mantissa <= conv_std_logic_vector(3912472,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01100011" =>
            mantissa <= conv_std_logic_vector(3960617,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01100100" =>
            mantissa <= conv_std_logic_vector(4008951,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01100101" =>
            mantissa <= conv_std_logic_vector(4057474,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01100110" =>
            mantissa <= conv_std_logic_vector(4106186,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01100111" =>
            mantissa <= conv_std_logic_vector(4155089,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01101000" =>
            mantissa <= conv_std_logic_vector(4204184,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01101001" =>
            mantissa <= conv_std_logic_vector(4253471,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01101010" =>
            mantissa <= conv_std_logic_vector(4302951,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01101011" =>
            mantissa <= conv_std_logic_vector(4352624,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01101100" =>
            mantissa <= conv_std_logic_vector(4402492,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01101101" =>
            mantissa <= conv_std_logic_vector(4452555,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01101110" =>
            mantissa <= conv_std_logic_vector(4502814,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01101111" =>
            mantissa <= conv_std_logic_vector(4553269,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01110000" =>
            mantissa <= conv_std_logic_vector(4603922,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01110001" =>
            mantissa <= conv_std_logic_vector(4654774,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01110010" =>
            mantissa <= conv_std_logic_vector(4705824,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01110011" =>
            mantissa <= conv_std_logic_vector(4757074,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01110100" =>
            mantissa <= conv_std_logic_vector(4808525,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01110101" =>
            mantissa <= conv_std_logic_vector(4860177,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01110110" =>
            mantissa <= conv_std_logic_vector(4912031,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01110111" =>
            mantissa <= conv_std_logic_vector(4964088,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01111000" =>
            mantissa <= conv_std_logic_vector(5016349,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01111001" =>
            mantissa <= conv_std_logic_vector(5068815,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01111010" =>
            mantissa <= conv_std_logic_vector(5121486,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01111011" =>
            mantissa <= conv_std_logic_vector(5174363,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01111100" =>
            mantissa <= conv_std_logic_vector(5227447,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01111101" =>
            mantissa <= conv_std_logic_vector(5280739,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01111110" =>
            mantissa <= conv_std_logic_vector(5334239,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "01111111" =>
            mantissa <= conv_std_logic_vector(5387949,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10000000" =>
            mantissa <= conv_std_logic_vector(5441868,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10000001" =>
            mantissa <= conv_std_logic_vector(5495999,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10000010" =>
            mantissa <= conv_std_logic_vector(5550342,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10000011" =>
            mantissa <= conv_std_logic_vector(5604898,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10000100" =>
            mantissa <= conv_std_logic_vector(5659667,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10000101" =>
            mantissa <= conv_std_logic_vector(5714650,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10000110" =>
            mantissa <= conv_std_logic_vector(5769849,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10000111" =>
            mantissa <= conv_std_logic_vector(5825263,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10001000" =>
            mantissa <= conv_std_logic_vector(5880895,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10001001" =>
            mantissa <= conv_std_logic_vector(5936744,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10001010" =>
            mantissa <= conv_std_logic_vector(5992812,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10001011" =>
            mantissa <= conv_std_logic_vector(6049099,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10001100" =>
            mantissa <= conv_std_logic_vector(6105607,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10001101" =>
            mantissa <= conv_std_logic_vector(6162336,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10001110" =>
            mantissa <= conv_std_logic_vector(6219286,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10001111" =>
            mantissa <= conv_std_logic_vector(6276460,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10010000" =>
            mantissa <= conv_std_logic_vector(6333858,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10010001" =>
            mantissa <= conv_std_logic_vector(6391480,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10010010" =>
            mantissa <= conv_std_logic_vector(6449327,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10010011" =>
            mantissa <= conv_std_logic_vector(6507401,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10010100" =>
            mantissa <= conv_std_logic_vector(6565703,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10010101" =>
            mantissa <= conv_std_logic_vector(6624232,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10010110" =>
            mantissa <= conv_std_logic_vector(6682991,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10010111" =>
            mantissa <= conv_std_logic_vector(6741979,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10011000" =>
            mantissa <= conv_std_logic_vector(6801199,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10011001" =>
            mantissa <= conv_std_logic_vector(6860650,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10011010" =>
            mantissa <= conv_std_logic_vector(6920334,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10011011" =>
            mantissa <= conv_std_logic_vector(6980251,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10011100" =>
            mantissa <= conv_std_logic_vector(7040403,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10011101" =>
            mantissa <= conv_std_logic_vector(7100791,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10011110" =>
            mantissa <= conv_std_logic_vector(7161415,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10011111" =>
            mantissa <= conv_std_logic_vector(7222276,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10100000" =>
            mantissa <= conv_std_logic_vector(7283375,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10100001" =>
            mantissa <= conv_std_logic_vector(7344713,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10100010" =>
            mantissa <= conv_std_logic_vector(7406292,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10100011" =>
            mantissa <= conv_std_logic_vector(7468111,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10100100" =>
            mantissa <= conv_std_logic_vector(7530173,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10100101" =>
            mantissa <= conv_std_logic_vector(7592477,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10100110" =>
            mantissa <= conv_std_logic_vector(7655025,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10100111" =>
            mantissa <= conv_std_logic_vector(7717818,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10101000" =>
            mantissa <= conv_std_logic_vector(7780857,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10101001" =>
            mantissa <= conv_std_logic_vector(7844143,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10101010" =>
            mantissa <= conv_std_logic_vector(7907676,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10101011" =>
            mantissa <= conv_std_logic_vector(7971458,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10101100" =>
            mantissa <= conv_std_logic_vector(8035489,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10101101" =>
            mantissa <= conv_std_logic_vector(8099771,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10101110" =>
            mantissa <= conv_std_logic_vector(8164305,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10101111" =>
            mantissa <= conv_std_logic_vector(8229091,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10110000" =>
            mantissa <= conv_std_logic_vector(8294131,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10110001" =>
            mantissa <= conv_std_logic_vector(8359425,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "10110010" =>
            mantissa <= conv_std_logic_vector(18184,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "10110011" =>
            mantissa <= conv_std_logic_vector(51087,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "10110100" =>
            mantissa <= conv_std_logic_vector(84119,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "10110101" =>
            mantissa <= conv_std_logic_vector(117280,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "10110110" =>
            mantissa <= conv_std_logic_vector(150571,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "10110111" =>
            mantissa <= conv_std_logic_vector(183993,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "10111000" =>
            mantissa <= conv_std_logic_vector(217545,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "10111001" =>
            mantissa <= conv_std_logic_vector(251229,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "10111010" =>
            mantissa <= conv_std_logic_vector(285044,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "10111011" =>
            mantissa <= conv_std_logic_vector(318992,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "10111100" =>
            mantissa <= conv_std_logic_vector(353072,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "10111101" =>
            mantissa <= conv_std_logic_vector(387286,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "10111110" =>
            mantissa <= conv_std_logic_vector(421634,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "10111111" =>
            mantissa <= conv_std_logic_vector(456116,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11000000" =>
            mantissa <= conv_std_logic_vector(490734,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11000001" =>
            mantissa <= conv_std_logic_vector(525486,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11000010" =>
            mantissa <= conv_std_logic_vector(560375,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11000011" =>
            mantissa <= conv_std_logic_vector(595401,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11000100" =>
            mantissa <= conv_std_logic_vector(630563,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11000101" =>
            mantissa <= conv_std_logic_vector(665863,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11000110" =>
            mantissa <= conv_std_logic_vector(701301,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11000111" =>
            mantissa <= conv_std_logic_vector(736878,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11001000" =>
            mantissa <= conv_std_logic_vector(772594,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11001001" =>
            mantissa <= conv_std_logic_vector(808450,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11001010" =>
            mantissa <= conv_std_logic_vector(844446,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11001011" =>
            mantissa <= conv_std_logic_vector(880584,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11001100" =>
            mantissa <= conv_std_logic_vector(916862,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11001101" =>
            mantissa <= conv_std_logic_vector(953283,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11001110" =>
            mantissa <= conv_std_logic_vector(989846,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11001111" =>
            mantissa <= conv_std_logic_vector(1026552,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11010000" =>
            mantissa <= conv_std_logic_vector(1063402,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11010001" =>
            mantissa <= conv_std_logic_vector(1100396,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11010010" =>
            mantissa <= conv_std_logic_vector(1137535,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11010011" =>
            mantissa <= conv_std_logic_vector(1174819,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11010100" =>
            mantissa <= conv_std_logic_vector(1212249,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11010101" =>
            mantissa <= conv_std_logic_vector(1249826,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11010110" =>
            mantissa <= conv_std_logic_vector(1287550,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11010111" =>
            mantissa <= conv_std_logic_vector(1325421,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11011000" =>
            mantissa <= conv_std_logic_vector(1363441,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11011001" =>
            mantissa <= conv_std_logic_vector(1401609,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11011010" =>
            mantissa <= conv_std_logic_vector(1439927,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11011011" =>
            mantissa <= conv_std_logic_vector(1478395,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11011100" =>
            mantissa <= conv_std_logic_vector(1517013,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11011101" =>
            mantissa <= conv_std_logic_vector(1555783,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11011110" =>
            mantissa <= conv_std_logic_vector(1594704,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11011111" =>
            mantissa <= conv_std_logic_vector(1633778,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11100000" =>
            mantissa <= conv_std_logic_vector(1673004,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11100001" =>
            mantissa <= conv_std_logic_vector(1712384,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11100010" =>
            mantissa <= conv_std_logic_vector(1751918,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11100011" =>
            mantissa <= conv_std_logic_vector(1791607,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11100100" =>
            mantissa <= conv_std_logic_vector(1831452,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11100101" =>
            mantissa <= conv_std_logic_vector(1871452,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11100110" =>
            mantissa <= conv_std_logic_vector(1911608,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11100111" =>
            mantissa <= conv_std_logic_vector(1951922,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11101000" =>
            mantissa <= conv_std_logic_vector(1992394,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11101001" =>
            mantissa <= conv_std_logic_vector(2033024,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11101010" =>
            mantissa <= conv_std_logic_vector(2073813,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11101011" =>
            mantissa <= conv_std_logic_vector(2114762,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11101100" =>
            mantissa <= conv_std_logic_vector(2155871,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11101101" =>
            mantissa <= conv_std_logic_vector(2197141,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11101110" =>
            mantissa <= conv_std_logic_vector(2238572,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11101111" =>
            mantissa <= conv_std_logic_vector(2280166,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11110000" =>
            mantissa <= conv_std_logic_vector(2321922,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11110001" =>
            mantissa <= conv_std_logic_vector(2363842,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11110010" =>
            mantissa <= conv_std_logic_vector(2405926,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11110011" =>
            mantissa <= conv_std_logic_vector(2448175,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11110100" =>
            mantissa <= conv_std_logic_vector(2490589,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11110101" =>
            mantissa <= conv_std_logic_vector(2533169,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11110110" =>
            mantissa <= conv_std_logic_vector(2575915,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11110111" =>
            mantissa <= conv_std_logic_vector(2618829,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11111000" =>
            mantissa <= conv_std_logic_vector(2661911,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11111001" =>
            mantissa <= conv_std_logic_vector(2705162,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11111010" =>
            mantissa <= conv_std_logic_vector(2748582,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11111011" =>
            mantissa <= conv_std_logic_vector(2792171,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11111100" =>
            mantissa <= conv_std_logic_vector(2835932,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11111101" =>
            mantissa <= conv_std_logic_vector(2879863,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11111110" =>
            mantissa <= conv_std_logic_vector(2923967,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "11111111" =>
            mantissa <= conv_std_logic_vector(2968243,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN others =>
           mantissa <= conv_std_logic_vector(0,23);
           exponent <= conv_std_logic_vector(0,8);
    END CASE;
  END PROCESS;

END rtl;
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_EXPLUTNEG.VHD                          ***
--***                                             ***
--***   Function: Look Up Table - EXP()           ***
--***                                             ***
--***   Generated by MATLAB Utility               ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_explutneg IS
PORT (
      address : IN STD_LOGIC_VECTOR (7 DOWNTO 1);
      mantissa : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
      exponent : OUT STD_LOGIC_VECTOR (8 DOWNTO 1)
     );
END fp_explutneg;

ARCHITECTURE rtl OF fp_explutneg IS

BEGIN

  pca: PROCESS (address)
  BEGIN
    CASE address IS
      WHEN "0000000" =>
            mantissa <= conv_std_logic_vector(0,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "0000001" =>
            mantissa <= conv_std_logic_vector(3955378,23);
            exponent <= conv_std_logic_vector(125,8);
      WHEN "0000010" =>
            mantissa <= conv_std_logic_vector(693589,23);
            exponent <= conv_std_logic_vector(124,8);
      WHEN "0000011" =>
            mantissa <= conv_std_logic_vector(4976006,23);
            exponent <= conv_std_logic_vector(122,8);
      WHEN "0000100" =>
            mantissa <= conv_std_logic_vector(1444526,23);
            exponent <= conv_std_logic_vector(121,8);
      WHEN "0000101" =>
            mantissa <= conv_std_logic_vector(6081023,23);
            exponent <= conv_std_logic_vector(119,8);
      WHEN "0000110" =>
            mantissa <= conv_std_logic_vector(2257552,23);
            exponent <= conv_std_logic_vector(118,8);
      WHEN "0000111" =>
            mantissa <= conv_std_logic_vector(7277405,23);
            exponent <= conv_std_logic_vector(116,8);
      WHEN "0001000" =>
            mantissa <= conv_std_logic_vector(3137800,23);
            exponent <= conv_std_logic_vector(115,8);
      WHEN "0001001" =>
            mantissa <= conv_std_logic_vector(92049,23);
            exponent <= conv_std_logic_vector(114,8);
      WHEN "0001010" =>
            mantissa <= conv_std_logic_vector(4090830,23);
            exponent <= conv_std_logic_vector(112,8);
      WHEN "0001011" =>
            mantissa <= conv_std_logic_vector(793249,23);
            exponent <= conv_std_logic_vector(111,8);
      WHEN "0001100" =>
            mantissa <= conv_std_logic_vector(5122658,23);
            exponent <= conv_std_logic_vector(109,8);
      WHEN "0001101" =>
            mantissa <= conv_std_logic_vector(1552426,23);
            exponent <= conv_std_logic_vector(108,8);
      WHEN "0001110" =>
            mantissa <= conv_std_logic_vector(6239800,23);
            exponent <= conv_std_logic_vector(106,8);
      WHEN "0001111" =>
            mantissa <= conv_std_logic_vector(2374373,23);
            exponent <= conv_std_logic_vector(105,8);
      WHEN "0010000" =>
            mantissa <= conv_std_logic_vector(7449310,23);
            exponent <= conv_std_logic_vector(103,8);
      WHEN "0010001" =>
            mantissa <= conv_std_logic_vector(3264281,23);
            exponent <= conv_std_logic_vector(102,8);
      WHEN "0010010" =>
            mantissa <= conv_std_logic_vector(185108,23);
            exponent <= conv_std_logic_vector(101,8);
      WHEN "0010011" =>
            mantissa <= conv_std_logic_vector(4227768,23);
            exponent <= conv_std_logic_vector(99,8);
      WHEN "0010100" =>
            mantissa <= conv_std_logic_vector(894003,23);
            exponent <= conv_std_logic_vector(98,8);
      WHEN "0010101" =>
            mantissa <= conv_std_logic_vector(5270919,23);
            exponent <= conv_std_logic_vector(96,8);
      WHEN "0010110" =>
            mantissa <= conv_std_logic_vector(1661510,23);
            exponent <= conv_std_logic_vector(95,8);
      WHEN "0010111" =>
            mantissa <= conv_std_logic_vector(6400319,23);
            exponent <= conv_std_logic_vector(93,8);
      WHEN "0011000" =>
            mantissa <= conv_std_logic_vector(2492476,23);
            exponent <= conv_std_logic_vector(92,8);
      WHEN "0011001" =>
            mantissa <= conv_std_logic_vector(7623101,23);
            exponent <= conv_std_logic_vector(90,8);
      WHEN "0011010" =>
            mantissa <= conv_std_logic_vector(3392149,23);
            exponent <= conv_std_logic_vector(89,8);
      WHEN "0011011" =>
            mantissa <= conv_std_logic_vector(279189,23);
            exponent <= conv_std_logic_vector(88,8);
      WHEN "0011100" =>
            mantissa <= conv_std_logic_vector(4366209,23);
            exponent <= conv_std_logic_vector(86,8);
      WHEN "0011101" =>
            mantissa <= conv_std_logic_vector(995862,23);
            exponent <= conv_std_logic_vector(85,8);
      WHEN "0011110" =>
            mantissa <= conv_std_logic_vector(5420806,23);
            exponent <= conv_std_logic_vector(83,8);
      WHEN "0011111" =>
            mantissa <= conv_std_logic_vector(1771791,23);
            exponent <= conv_std_logic_vector(82,8);
      WHEN "0100000" =>
            mantissa <= conv_std_logic_vector(6562600,23);
            exponent <= conv_std_logic_vector(80,8);
      WHEN "0100001" =>
            mantissa <= conv_std_logic_vector(2611876,23);
            exponent <= conv_std_logic_vector(79,8);
      WHEN "0100010" =>
            mantissa <= conv_std_logic_vector(7798799,23);
            exponent <= conv_std_logic_vector(77,8);
      WHEN "0100011" =>
            mantissa <= conv_std_logic_vector(3521421,23);
            exponent <= conv_std_logic_vector(76,8);
      WHEN "0100100" =>
            mantissa <= conv_std_logic_vector(374301,23);
            exponent <= conv_std_logic_vector(75,8);
      WHEN "0100101" =>
            mantissa <= conv_std_logic_vector(4506169,23);
            exponent <= conv_std_logic_vector(73,8);
      WHEN "0100110" =>
            mantissa <= conv_std_logic_vector(1098839,23);
            exponent <= conv_std_logic_vector(72,8);
      WHEN "0100111" =>
            mantissa <= conv_std_logic_vector(5572338,23);
            exponent <= conv_std_logic_vector(70,8);
      WHEN "0101000" =>
            mantissa <= conv_std_logic_vector(1883282,23);
            exponent <= conv_std_logic_vector(69,8);
      WHEN "0101001" =>
            mantissa <= conv_std_logic_vector(6726661,23);
            exponent <= conv_std_logic_vector(67,8);
      WHEN "0101010" =>
            mantissa <= conv_std_logic_vector(2732585,23);
            exponent <= conv_std_logic_vector(66,8);
      WHEN "0101011" =>
            mantissa <= conv_std_logic_vector(7976426,23);
            exponent <= conv_std_logic_vector(64,8);
      WHEN "0101100" =>
            mantissa <= conv_std_logic_vector(3652111,23);
            exponent <= conv_std_logic_vector(63,8);
      WHEN "0101101" =>
            mantissa <= conv_std_logic_vector(470458,23);
            exponent <= conv_std_logic_vector(62,8);
      WHEN "0101110" =>
            mantissa <= conv_std_logic_vector(4647665,23);
            exponent <= conv_std_logic_vector(60,8);
      WHEN "0101111" =>
            mantissa <= conv_std_logic_vector(1202946,23);
            exponent <= conv_std_logic_vector(59,8);
      WHEN "0110000" =>
            mantissa <= conv_std_logic_vector(5725533,23);
            exponent <= conv_std_logic_vector(57,8);
      WHEN "0110001" =>
            mantissa <= conv_std_logic_vector(1995997,23);
            exponent <= conv_std_logic_vector(56,8);
      WHEN "0110010" =>
            mantissa <= conv_std_logic_vector(6892523,23);
            exponent <= conv_std_logic_vector(54,8);
      WHEN "0110011" =>
            mantissa <= conv_std_logic_vector(2854620,23);
            exponent <= conv_std_logic_vector(53,8);
      WHEN "0110100" =>
            mantissa <= conv_std_logic_vector(8156001,23);
            exponent <= conv_std_logic_vector(51,8);
      WHEN "0110101" =>
            mantissa <= conv_std_logic_vector(3784235,23);
            exponent <= conv_std_logic_vector(50,8);
      WHEN "0110110" =>
            mantissa <= conv_std_logic_vector(567669,23);
            exponent <= conv_std_logic_vector(49,8);
      WHEN "0110111" =>
            mantissa <= conv_std_logic_vector(4790713,23);
            exponent <= conv_std_logic_vector(47,8);
      WHEN "0111000" =>
            mantissa <= conv_std_logic_vector(1308195,23);
            exponent <= conv_std_logic_vector(46,8);
      WHEN "0111001" =>
            mantissa <= conv_std_logic_vector(5880410,23);
            exponent <= conv_std_logic_vector(44,8);
      WHEN "0111010" =>
            mantissa <= conv_std_logic_vector(2109948,23);
            exponent <= conv_std_logic_vector(43,8);
      WHEN "0111011" =>
            mantissa <= conv_std_logic_vector(7060204,23);
            exponent <= conv_std_logic_vector(41,8);
      WHEN "0111100" =>
            mantissa <= conv_std_logic_vector(2977993,23);
            exponent <= conv_std_logic_vector(40,8);
      WHEN "0111101" =>
            mantissa <= conv_std_logic_vector(8337547,23);
            exponent <= conv_std_logic_vector(38,8);
      WHEN "0111110" =>
            mantissa <= conv_std_logic_vector(3917809,23);
            exponent <= conv_std_logic_vector(37,8);
      WHEN "0111111" =>
            mantissa <= conv_std_logic_vector(665948,23);
            exponent <= conv_std_logic_vector(36,8);
      WHEN "1000000" =>
            mantissa <= conv_std_logic_vector(4935332,23);
            exponent <= conv_std_logic_vector(34,8);
      WHEN "1000001" =>
            mantissa <= conv_std_logic_vector(1414599,23);
            exponent <= conv_std_logic_vector(33,8);
      WHEN "1000010" =>
            mantissa <= conv_std_logic_vector(6036985,23);
            exponent <= conv_std_logic_vector(31,8);
      WHEN "1000011" =>
            mantissa <= conv_std_logic_vector(2225150,23);
            exponent <= conv_std_logic_vector(30,8);
      WHEN "1000100" =>
            mantissa <= conv_std_logic_vector(7229726,23);
            exponent <= conv_std_logic_vector(28,8);
      WHEN "1000101" =>
            mantissa <= conv_std_logic_vector(3102720,23);
            exponent <= conv_std_logic_vector(27,8);
      WHEN "1000110" =>
            mantissa <= conv_std_logic_vector(66239,23);
            exponent <= conv_std_logic_vector(26,8);
      WHEN "1000111" =>
            mantissa <= conv_std_logic_vector(4052849,23);
            exponent <= conv_std_logic_vector(24,8);
      WHEN "1001000" =>
            mantissa <= conv_std_logic_vector(765304,23);
            exponent <= conv_std_logic_vector(23,8);
      WHEN "1001001" =>
            mantissa <= conv_std_logic_vector(5081537,23);
            exponent <= conv_std_logic_vector(21,8);
      WHEN "1001010" =>
            mantissa <= conv_std_logic_vector(1522171,23);
            exponent <= conv_std_logic_vector(20,8);
      WHEN "1001011" =>
            mantissa <= conv_std_logic_vector(6195279,23);
            exponent <= conv_std_logic_vector(18,8);
      WHEN "1001100" =>
            mantissa <= conv_std_logic_vector(2341616,23);
            exponent <= conv_std_logic_vector(17,8);
      WHEN "1001101" =>
            mantissa <= conv_std_logic_vector(7401108,23);
            exponent <= conv_std_logic_vector(15,8);
      WHEN "1001110" =>
            mantissa <= conv_std_logic_vector(3228816,23);
            exponent <= conv_std_logic_vector(14,8);
      WHEN "1001111" =>
            mantissa <= conv_std_logic_vector(159015,23);
            exponent <= conv_std_logic_vector(13,8);
      WHEN "1010000" =>
            mantissa <= conv_std_logic_vector(4189370,23);
            exponent <= conv_std_logic_vector(11,8);
      WHEN "1010001" =>
            mantissa <= conv_std_logic_vector(865751,23);
            exponent <= conv_std_logic_vector(10,8);
      WHEN "1010010" =>
            mantissa <= conv_std_logic_vector(5229346,23);
            exponent <= conv_std_logic_vector(8,8);
      WHEN "1010011" =>
            mantissa <= conv_std_logic_vector(1630923,23);
            exponent <= conv_std_logic_vector(7,8);
      WHEN "1010100" =>
            mantissa <= conv_std_logic_vector(6355309,23);
            exponent <= conv_std_logic_vector(5,8);
      WHEN "1010101" =>
            mantissa <= conv_std_logic_vector(2459360,23);
            exponent <= conv_std_logic_vector(4,8);
      WHEN "1010110" =>
            mantissa <= conv_std_logic_vector(7574370,23);
            exponent <= conv_std_logic_vector(2,8);
      WHEN "1010111" =>
            mantissa <= conv_std_logic_vector(3356295,23);
            exponent <= conv_std_logic_vector(1,8);
      WHEN "1011000" =>
            mantissa <= conv_std_logic_vector(252809,23);
            exponent <= conv_std_logic_vector(0,8);
      WHEN "1011001" =>
            mantissa <= conv_std_logic_vector(4327390,23);
            exponent <= conv_std_logic_vector(-2,8);
      WHEN others =>
           mantissa <= conv_std_logic_vector(0,23);
           exponent <= conv_std_logic_vector(0,8);
    END CASE;
  END PROCESS;

END rtl;
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_EXPLUTPOS.VHD                          ***
--***                                             ***
--***   Function: Look Up Table - EXP()           ***
--***                                             ***
--***   Generated by MATLAB Utility               ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_explutpos IS
PORT (
      address : IN STD_LOGIC_VECTOR (7 DOWNTO 1);
      mantissa : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
      exponent : OUT STD_LOGIC_VECTOR (8 DOWNTO 1)
     );
END fp_explutpos;

ARCHITECTURE rtl OF fp_explutpos IS

BEGIN

  pca: PROCESS (address)
  BEGIN
    CASE address IS
      WHEN "0000000" =>
            mantissa <= conv_std_logic_vector(0,23);
            exponent <= conv_std_logic_vector(127,8);
      WHEN "0000001" =>
            mantissa <= conv_std_logic_vector(3012692,23);
            exponent <= conv_std_logic_vector(128,8);
      WHEN "0000010" =>
            mantissa <= conv_std_logic_vector(7107366,23);
            exponent <= conv_std_logic_vector(129,8);
      WHEN "0000011" =>
            mantissa <= conv_std_logic_vector(2141998,23);
            exponent <= conv_std_logic_vector(131,8);
      WHEN "0000100" =>
            mantissa <= conv_std_logic_vector(5923969,23);
            exponent <= conv_std_logic_vector(132,8);
      WHEN "0000101" =>
            mantissa <= conv_std_logic_vector(1337797,23);
            exponent <= conv_std_logic_vector(134,8);
      WHEN "0000110" =>
            mantissa <= conv_std_logic_vector(4830947,23);
            exponent <= conv_std_logic_vector(135,8);
      WHEN "0000111" =>
            mantissa <= conv_std_logic_vector(595011,23);
            exponent <= conv_std_logic_vector(137,8);
      WHEN "0001000" =>
            mantissa <= conv_std_logic_vector(3821396,23);
            exponent <= conv_std_logic_vector(138,8);
      WHEN "0001001" =>
            mantissa <= conv_std_logic_vector(8206508,23);
            exponent <= conv_std_logic_vector(139,8);
      WHEN "0001010" =>
            mantissa <= conv_std_logic_vector(2888942,23);
            exponent <= conv_std_logic_vector(141,8);
      WHEN "0001011" =>
            mantissa <= conv_std_logic_vector(6939172,23);
            exponent <= conv_std_logic_vector(142,8);
      WHEN "0001100" =>
            mantissa <= conv_std_logic_vector(2027699,23);
            exponent <= conv_std_logic_vector(144,8);
      WHEN "0001101" =>
            mantissa <= conv_std_logic_vector(5768621,23);
            exponent <= conv_std_logic_vector(145,8);
      WHEN "0001110" =>
            mantissa <= conv_std_logic_vector(1232226,23);
            exponent <= conv_std_logic_vector(147,8);
      WHEN "0001111" =>
            mantissa <= conv_std_logic_vector(4687461,23);
            exponent <= conv_std_logic_vector(148,8);
      WHEN "0010000" =>
            mantissa <= conv_std_logic_vector(497503,23);
            exponent <= conv_std_logic_vector(150,8);
      WHEN "0010001" =>
            mantissa <= conv_std_logic_vector(3688868,23);
            exponent <= conv_std_logic_vector(151,8);
      WHEN "0010010" =>
            mantissa <= conv_std_logic_vector(8026384,23);
            exponent <= conv_std_logic_vector(152,8);
      WHEN "0010011" =>
            mantissa <= conv_std_logic_vector(2766536,23);
            exponent <= conv_std_logic_vector(154,8);
      WHEN "0010100" =>
            mantissa <= conv_std_logic_vector(6772804,23);
            exponent <= conv_std_logic_vector(155,8);
      WHEN "0010101" =>
            mantissa <= conv_std_logic_vector(1914640,23);
            exponent <= conv_std_logic_vector(157,8);
      WHEN "0010110" =>
            mantissa <= conv_std_logic_vector(5614958,23);
            exponent <= conv_std_logic_vector(158,8);
      WHEN "0010111" =>
            mantissa <= conv_std_logic_vector(1127802,23);
            exponent <= conv_std_logic_vector(160,8);
      WHEN "0011000" =>
            mantissa <= conv_std_logic_vector(4545534,23);
            exponent <= conv_std_logic_vector(161,8);
      WHEN "0011001" =>
            mantissa <= conv_std_logic_vector(401053,23);
            exponent <= conv_std_logic_vector(163,8);
      WHEN "0011010" =>
            mantissa <= conv_std_logic_vector(3557779,23);
            exponent <= conv_std_logic_vector(164,8);
      WHEN "0011011" =>
            mantissa <= conv_std_logic_vector(7848216,23);
            exponent <= conv_std_logic_vector(165,8);
      WHEN "0011100" =>
            mantissa <= conv_std_logic_vector(2645458,23);
            exponent <= conv_std_logic_vector(167,8);
      WHEN "0011101" =>
            mantissa <= conv_std_logic_vector(6608242,23);
            exponent <= conv_std_logic_vector(168,8);
      WHEN "0011110" =>
            mantissa <= conv_std_logic_vector(1802808,23);
            exponent <= conv_std_logic_vector(170,8);
      WHEN "0011111" =>
            mantissa <= conv_std_logic_vector(5462963,23);
            exponent <= conv_std_logic_vector(171,8);
      WHEN "0100000" =>
            mantissa <= conv_std_logic_vector(1024510,23);
            exponent <= conv_std_logic_vector(173,8);
      WHEN "0100001" =>
            mantissa <= conv_std_logic_vector(4405146,23);
            exponent <= conv_std_logic_vector(174,8);
      WHEN "0100010" =>
            mantissa <= conv_std_logic_vector(305649,23);
            exponent <= conv_std_logic_vector(176,8);
      WHEN "0100011" =>
            mantissa <= conv_std_logic_vector(3428113,23);
            exponent <= conv_std_logic_vector(177,8);
      WHEN "0100100" =>
            mantissa <= conv_std_logic_vector(7671981,23);
            exponent <= conv_std_logic_vector(178,8);
      WHEN "0100101" =>
            mantissa <= conv_std_logic_vector(2525694,23);
            exponent <= conv_std_logic_vector(180,8);
      WHEN "0100110" =>
            mantissa <= conv_std_logic_vector(6445466,23);
            exponent <= conv_std_logic_vector(181,8);
      WHEN "0100111" =>
            mantissa <= conv_std_logic_vector(1692191,23);
            exponent <= conv_std_logic_vector(183,8);
      WHEN "0101000" =>
            mantissa <= conv_std_logic_vector(5312618,23);
            exponent <= conv_std_logic_vector(184,8);
      WHEN "0101001" =>
            mantissa <= conv_std_logic_vector(922340,23);
            exponent <= conv_std_logic_vector(186,8);
      WHEN "0101010" =>
            mantissa <= conv_std_logic_vector(4266283,23);
            exponent <= conv_std_logic_vector(187,8);
      WHEN "0101011" =>
            mantissa <= conv_std_logic_vector(211282,23);
            exponent <= conv_std_logic_vector(189,8);
      WHEN "0101100" =>
            mantissa <= conv_std_logic_vector(3299854,23);
            exponent <= conv_std_logic_vector(190,8);
      WHEN "0101101" =>
            mantissa <= conv_std_logic_vector(7497659,23);
            exponent <= conv_std_logic_vector(191,8);
      WHEN "0101110" =>
            mantissa <= conv_std_logic_vector(2407230,23);
            exponent <= conv_std_logic_vector(193,8);
      WHEN "0101111" =>
            mantissa <= conv_std_logic_vector(6284457,23);
            exponent <= conv_std_logic_vector(194,8);
      WHEN "0110000" =>
            mantissa <= conv_std_logic_vector(1582773,23);
            exponent <= conv_std_logic_vector(196,8);
      WHEN "0110001" =>
            mantissa <= conv_std_logic_vector(5163905,23);
            exponent <= conv_std_logic_vector(197,8);
      WHEN "0110010" =>
            mantissa <= conv_std_logic_vector(821279,23);
            exponent <= conv_std_logic_vector(199,8);
      WHEN "0110011" =>
            mantissa <= conv_std_logic_vector(4128926,23);
            exponent <= conv_std_logic_vector(200,8);
      WHEN "0110100" =>
            mantissa <= conv_std_logic_vector(117939,23);
            exponent <= conv_std_logic_vector(202,8);
      WHEN "0110101" =>
            mantissa <= conv_std_logic_vector(3172987,23);
            exponent <= conv_std_logic_vector(203,8);
      WHEN "0110110" =>
            mantissa <= conv_std_logic_vector(7325229,23);
            exponent <= conv_std_logic_vector(204,8);
      WHEN "0110111" =>
            mantissa <= conv_std_logic_vector(2290052,23);
            exponent <= conv_std_logic_vector(206,8);
      WHEN "0111000" =>
            mantissa <= conv_std_logic_vector(6125195,23);
            exponent <= conv_std_logic_vector(207,8);
      WHEN "0111001" =>
            mantissa <= conv_std_logic_vector(1474544,23);
            exponent <= conv_std_logic_vector(209,8);
      WHEN "0111010" =>
            mantissa <= conv_std_logic_vector(5016805,23);
            exponent <= conv_std_logic_vector(210,8);
      WHEN "0111011" =>
            mantissa <= conv_std_logic_vector(721315,23);
            exponent <= conv_std_logic_vector(212,8);
      WHEN "0111100" =>
            mantissa <= conv_std_logic_vector(3993061,23);
            exponent <= conv_std_logic_vector(213,8);
      WHEN "0111101" =>
            mantissa <= conv_std_logic_vector(25608,23);
            exponent <= conv_std_logic_vector(215,8);
      WHEN "0111110" =>
            mantissa <= conv_std_logic_vector(3047498,23);
            exponent <= conv_std_logic_vector(216,8);
      WHEN "0111111" =>
            mantissa <= conv_std_logic_vector(7154671,23);
            exponent <= conv_std_logic_vector(217,8);
      WHEN "1000000" =>
            mantissa <= conv_std_logic_vector(2174145,23);
            exponent <= conv_std_logic_vector(219,8);
      WHEN "1000001" =>
            mantissa <= conv_std_logic_vector(5967662,23);
            exponent <= conv_std_logic_vector(220,8);
      WHEN "1000010" =>
            mantissa <= conv_std_logic_vector(1367489,23);
            exponent <= conv_std_logic_vector(222,8);
      WHEN "1000011" =>
            mantissa <= conv_std_logic_vector(4871303,23);
            exponent <= conv_std_logic_vector(223,8);
      WHEN "1000100" =>
            mantissa <= conv_std_logic_vector(622436,23);
            exponent <= conv_std_logic_vector(225,8);
      WHEN "1000101" =>
            mantissa <= conv_std_logic_vector(3858670,23);
            exponent <= conv_std_logic_vector(226,8);
      WHEN "1000110" =>
            mantissa <= conv_std_logic_vector(8257169,23);
            exponent <= conv_std_logic_vector(227,8);
      WHEN "1000111" =>
            mantissa <= conv_std_logic_vector(2923370,23);
            exponent <= conv_std_logic_vector(229,8);
      WHEN "1001000" =>
            mantissa <= conv_std_logic_vector(6985964,23);
            exponent <= conv_std_logic_vector(230,8);
      WHEN "1001001" =>
            mantissa <= conv_std_logic_vector(2059497,23);
            exponent <= conv_std_logic_vector(232,8);
      WHEN "1001010" =>
            mantissa <= conv_std_logic_vector(5811839,23);
            exponent <= conv_std_logic_vector(233,8);
      WHEN "1001011" =>
            mantissa <= conv_std_logic_vector(1261596,23);
            exponent <= conv_std_logic_vector(235,8);
      WHEN "1001100" =>
            mantissa <= conv_std_logic_vector(4727380,23);
            exponent <= conv_std_logic_vector(236,8);
      WHEN "1001101" =>
            mantissa <= conv_std_logic_vector(524630,23);
            exponent <= conv_std_logic_vector(238,8);
      WHEN "1001110" =>
            mantissa <= conv_std_logic_vector(3725738,23);
            exponent <= conv_std_logic_vector(239,8);
      WHEN "1001111" =>
            mantissa <= conv_std_logic_vector(8076495,23);
            exponent <= conv_std_logic_vector(240,8);
      WHEN "1010000" =>
            mantissa <= conv_std_logic_vector(2800590,23);
            exponent <= conv_std_logic_vector(242,8);
      WHEN "1010001" =>
            mantissa <= conv_std_logic_vector(6819089,23);
            exponent <= conv_std_logic_vector(243,8);
      WHEN "1010010" =>
            mantissa <= conv_std_logic_vector(1946093,23);
            exponent <= conv_std_logic_vector(245,8);
      WHEN "1010011" =>
            mantissa <= conv_std_logic_vector(5657707,23);
            exponent <= conv_std_logic_vector(246,8);
      WHEN "1010100" =>
            mantissa <= conv_std_logic_vector(1156853,23);
            exponent <= conv_std_logic_vector(248,8);
      WHEN "1010101" =>
            mantissa <= conv_std_logic_vector(4585019,23);
            exponent <= conv_std_logic_vector(249,8);
      WHEN "1010110" =>
            mantissa <= conv_std_logic_vector(427885,23);
            exponent <= conv_std_logic_vector(251,8);
      WHEN "1010111" =>
            mantissa <= conv_std_logic_vector(3594249,23);
            exponent <= conv_std_logic_vector(252,8);
      WHEN "1011000" =>
            mantissa <= conv_std_logic_vector(7897783,23);
            exponent <= conv_std_logic_vector(253,8);
      WHEN "1011001" =>
            mantissa <= conv_std_logic_vector(2679142,23);
            exponent <= conv_std_logic_vector(255,8);
      WHEN others =>
           mantissa <= conv_std_logic_vector(0,23);
           exponent <= conv_std_logic_vector(0,8);
    END CASE;
  END PROCESS;

END rtl;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_EXPRND.VHD                             ***
--***                                             ***
--***   Function: FP Exponent Output Block -      ***
--***   Rounded                                   ***
--***                                             ***
--***   Generated by MATLAB Utility               ***
--***                                             ***
--***   18/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_exprnd IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentexp : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissaexp : IN STD_LOGIC_VECTOR (24 DOWNTO 1); -- includes roundbit
      nanin : IN STD_LOGIC;
      rangeerror : IN STD_LOGIC;

		  signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
      --------------------------------------------------
      nanout : OUT STD_LOGIC;
      overflowout : OUT STD_LOGIC;
      underflowout : OUT STD_LOGIC
		);
END fp_exprnd;

ARCHITECTURE rtl OF fp_exprnd IS

  constant expwidth : positive := 8;
  constant manwidth : positive := 23;
  
  type exponentfftype IS ARRAY (2 DOWNTO 1) OF STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  
  signal zerovec : STD_LOGIC_VECTOR (manwidth-1 DOWNTO 1);
  signal nanff : STD_LOGIC_VECTOR (2 DOWNTO 1);
  signal rangeerrorff : STD_LOGIC;
  signal overflownode, underflownode : STD_LOGIC;
  signal overflowff, underflowff : STD_LOGIC_VECTOR (2 DOWNTO 1);
  signal manoverflowbitff : STD_LOGIC; 
  signal roundmantissaff, mantissaff : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal exponentnode : STD_LOGIC_VECTOR (expwidth+2 DOWNTO 1);
  signal exponentoneff : STD_LOGIC_VECTOR (expwidth+2 DOWNTO 1);
  signal exponenttwoff : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
    
  signal manoverflow : STD_LOGIC_VECTOR (manwidth+1 DOWNTO 1);
  signal infinitygen : STD_LOGIC_VECTOR (expwidth+1 DOWNTO 1);
  signal zerogen : STD_LOGIC_VECTOR (expwidth+1 DOWNTO 1);  
  signal setmanzero, setmanmax : STD_LOGIC;
  signal setexpzero, setexpmax : STD_LOGIC;

BEGIN
    
  gzv: FOR k IN 1 TO manwidth-1 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  pra: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN
        
      nanff <= "00";
      rangeerrorff <= '0';
      overflowff <= "00";
      underflowff <= "00";
      manoverflowbitff <= '0';
      FOR k IN 1 TO manwidth LOOP
        roundmantissaff(k) <= '0';
        mantissaff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth+2 LOOP
        exponentoneff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        exponenttwoff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF(enable = '1') THEN 
      
        nanff(1) <= nanin;
        nanff(2) <= nanff(1);
        rangeerrorff <= rangeerror;
        overflowff(1) <= overflownode;
        overflowff(2) <= overflowff(1);
        underflowff(1) <= underflownode;
        underflowff(2) <= underflowff(1);
        
        manoverflowbitff <= manoverflow(manwidth+1);
        
        roundmantissaff <= mantissaexp(manwidth+1 DOWNTO 2) + (zerovec & mantissaexp(1));
        
        -- nan takes precedence (set max)
        -- nan takes precedence (set max)  
        FOR k IN 1 TO manwidth LOOP
          mantissaff(k) <= (roundmantissaff(k) AND setmanzero) OR setmanmax;
        END LOOP;
        
        exponentoneff(expwidth+2 DOWNTO 1) <= "00" & exponentexp;                 
        FOR k IN 1 TO expwidth LOOP
          exponenttwoff(k) <= (exponentnode(k) AND setexpzero) OR setexpmax;
        END LOOP;
      
      END IF;
             
    END IF;
      
  END PROCESS;
  
  exponentnode <= exponentoneff(expwidth+2 DOWNTO 1) + 
                 (zerovec(expwidth+1 DOWNTO 1) & manoverflowbitff);

--*********************************
--*** PREDICT MANTISSA OVERFLOW ***   
--*********************************
     
  manoverflow(1) <= mantissaexp(1);
  gmoa: FOR k IN 2 TO manwidth+1 GENERATE
    manoverflow(k) <= manoverflow(k-1) AND mantissaexp(k);
  END GENERATE; 
                                                                 
--**********************************
--*** CHECK GENERATED CONDITIONS ***   
--**********************************

  -- infinity if exponent == 255
  infinitygen(1) <= exponentnode(1);
  gia: FOR k IN 2 TO expwidth GENERATE
    infinitygen(k) <= infinitygen(k-1) AND exponentnode(k);
  END GENERATE;
  infinitygen(expwidth+1) <= infinitygen(expwidth) OR 
                            (exponentnode(expwidth+1) AND 
                             NOT(exponentnode(expwidth+2))); -- '1' if infinity
                                                    
  -- zero if exponent == 0
  zerogen(1) <= exponentnode(1);
  gza: FOR k IN 2 TO expwidth GENERATE
    zerogen(k) <= zerogen(k-1) OR exponentnode(k);
  END GENERATE;
  zerogen(expwidth+1) <= zerogen(expwidth) AND 
                         NOT(exponentnode(expwidth+2)); -- '0' if zero
                                           
  -- trap any other overflow errors
  -- when sign = 0 and rangeerror = 1, overflow
  -- when sign = 1 and rangeerror = 1, underflow
  overflownode <= NOT(signin) AND rangeerror;
  underflownode <= signin AND rangeerror;
  
  -- set mantissa to 0 when infinity or zero condition
  setmanzero <= NOT(infinitygen(expwidth+1)) AND zerogen(expwidth+1) AND NOT(rangeerrorff);
  -- setmantissa to "11..11" when nan
  setmanmax <= nanin;
  -- set exponent to 0 when zero condition 
  setexpzero <= zerogen(expwidth+1);
  -- set exponent to "11..11" when nan, infinity, or divide by 0
  setexpmax <= nanin OR infinitygen(expwidth+1) OR rangeerrorff;
                             
--***************
--*** OUTPUTS ***
--***************
  
  signout <= '0';   
  mantissaout <= mantissaff;
  exponentout <= exponenttwoff; 
  -----------------------------------------------
  nanout <= nanff(2);
  overflowout <= overflowff(2);
  underflowout <= underflowff(2);

END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   ALTERA FLOATING POINT DATAPATH COMPILER   ***
--***                                             ***
--***   FP_FABS.VHD                               ***
--***                                             ***
--***   Function: Single Precision Absolute Value ***
--***                                             ***
--***   abs(x)                                    ***
--***                                             ***
--***   Created 11/09/09                          ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_fabs IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (23 DOWNTO 1);

		  signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
		  satout, zeroout, nanout : OUT STD_LOGIC
		);
END fp_fabs;

ARCHITECTURE rtl OF fp_fabs IS
 
  signal signff : STD_LOGIC;
  signal exponentff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal mantissaff : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal expnode : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal expzerochk, expmaxchk : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal expzero, expmax : STD_LOGIC;
  signal manzerochk : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal manzero, mannonzero : STD_LOGIC; 

BEGIN
    
  pin: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
    
      signff <= '0';
      FOR k IN 1 TO 8 LOOP
        exponentff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 23 LOOP
        mantissaff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF (enable = '1') THEN
          
        signff <= '0';
        exponentff <= exponentin;
        mantissaff <= mantissain;
        
      END IF;
    
    END IF;  
      
  END PROCESS;

  expzerochk(1) <= exponentff(1);
  expmaxchk(1) <= exponentff(1);
  gxa: FOR k IN 2 TO 8 GENERATE
    expzerochk(k) <= expzerochk(k-1) OR exponentff(k);
    expmaxchk(k) <= expmaxchk(k-1) AND exponentff(k);
  END GENERATE;
  expzero <= NOT(expzerochk(8));
  expmax <= expmaxchk(8);
  
  manzerochk(1) <= mantissaff(1);
  gma: FOR k IN 2 TO 23 GENERATE
    manzerochk(k) <= manzerochk(k-1) OR mantissaff(k);
  END GENERATE;
  manzero <= NOT(manzerochk(23));
  mannonzero <= manzerochk(23);
  
  signout <= signff;
  exponentout <= exponentff;
  mantissaout <= mantissaff;
  satout <= expmax AND manzero;
  zeroout <= expzero;
  nanout <= expmax AND mannonzero;

END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_FXMUL.VHD                              ***
--***                                             ***
--***   Function: Parameterized Fixed Point       ***
--***   Multiplier                                ***
--***   (behavioral and synthesizable support)    ***
--***                                             ***
--***   09/12/07 ML                               ***
--***                                             ***
--***   (c) 2007 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***   15/01/08 - change 54x18 to >54 outputs    ***
--***   23/04/09 - change 54x54 to SII & SIII     ***
--***   versions with both 8&9(10) multipliers    ***
--***                                             ***
--***************************************************

--***************************************************
--*** valid supported cores                       ***
--***                                             ***
--*** 1: SII/SIII, 18-36 bit inputs,              ***
--***    any output width, 2 pipes                ***
--*** 2: SII/SIII, 18-36 bit inputs,              ***
--***    any output width, 3 pipes                ***
--*** 3: SII/SIII 54x18 inputs,                   ***
--***    up to 72 bit output, 3 or 4 pipes        ***
--*** 4: SII 54x54 inputs, 72 bit outputs,        ***
--***    8 or 9 multiplier core 5 or 6 pipes      ***
--*** 5: SIII/IV 54x54 inputs, 72 bit outputs,    ***
--***    8 or 9 (10) multiplier core 4 pipes      ***
--***                                             ***
--***************************************************

ENTITY fp_fxmul IS 
GENERIC (
         widthaa : positive := 18;
         widthbb : positive := 18;
         widthcc : positive := 36;
         pipes : positive := 1;
         accuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
         device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
         synthesize : integer := 0
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
      databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1); 
      
      result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
     );
END fp_fxmul;

ARCHITECTURE rtl OF fp_fxmul IS

  component fp_mul2s
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36
          );
  PORT
	   (
       sysclk : IN STD_LOGIC;
       reset : IN STD_LOGIC;
       enable : IN STD_LOGIC;
       dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
       databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1);

	    result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
	  );
  end component;
  
  component fp_mul3s
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36
          );
  PORT
	   (
       sysclk : IN STD_LOGIC;
       reset : IN STD_LOGIC;
       enable : IN STD_LOGIC;
       dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
       databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1);

	    result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
	  );
  end component;
  
  component fp_mul5418s 
  GENERIC (
           widthcc : positive := 36;
           pipes : positive := 3  --3/4
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (54 DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (18 DOWNTO 1);
      
		  result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
		  );
  end component;
  
  component fp_mul54us_3xs
  PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      mulaa, mulbb : IN STD_LOGIC_VECTOR (54 DOWNTO 1);      

      mulcc : OUT STD_LOGIC_VECTOR (72 DOWNTO 1)  
     );
  end component;
  
  component fp_mul54us_28s 
  GENERIC (latency : positive := 5);
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        mulaa, mulbb : IN STD_LOGIC_VECTOR (54 DOWNTO 1);      

        mulcc : OUT STD_LOGIC_VECTOR (72 DOWNTO 1)  
       );
  end component;
  
  component fp_mul54us_29s 
  GENERIC (latency : positive := 5);
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        mulaa, mulbb : IN STD_LOGIC_VECTOR (54 DOWNTO 1);      

        mulcc : OUT STD_LOGIC_VECTOR (72 DOWNTO 1)  
       );
  end component;
  
  component fp_mul54us_38s
  PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      mulaa, mulbb : IN STD_LOGIC_VECTOR (54 DOWNTO 1);      

      mulcc : OUT STD_LOGIC_VECTOR (72 DOWNTO 1)  
     );
  end component;
  
  component fp_mul54usb 
  GENERIC (
           latency : positive := 5; -- 4/5/6
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           prune : integer := 0 -- 0 = pruned multiplier, 1 = normal multiplier
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa, bb : IN STD_LOGIC_VECTOR (54 DOWNTO 1);
      
		  cc : OUT STD_LOGIC_VECTOR (72 DOWNTO 1)
		  );
  end component;		
  
  component fp_mul7218s 
  GENERIC (
           widthcc : positive := 36;
           pipes : positive := 3  --3/4
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (72 DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (18 DOWNTO 1);
      
		  result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
		  );
  end component;
    		 
BEGIN
  
  gone: IF ((widthaa < 37) AND 
            (widthbb < 37) AND 
            (widthcc <= (widthaa + widthbb)) AND
            (pipes = 2)) GENERATE
            
    mulone: fp_mul2s
    GENERIC MAP (widthaa=>widthaa,widthbb=>widthbb,widthcc=>widthcc)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              dataaa=>dataaa,databb=>databb,
              result=>result);
          
  END GENERATE;

  gtwo: IF ((widthaa < 37) AND 
            (widthbb < 37) AND 
            (widthcc <= (widthaa + widthbb)) AND
            (pipes = 3)) GENERATE
            
    multwo: fp_mul3s
    GENERIC MAP (widthaa=>widthaa,widthbb=>widthbb,widthcc=>widthcc)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              dataaa=>dataaa,databb=>databb,
              result=>result);
          
  END GENERATE;

  gthr: IF ((widthaa = 54) AND 
            (widthbb = 18) AND 
            (widthcc < 73) AND
            ((pipes = 3) OR (pipes = 4))) GENERATE
            
    multhr: fp_mul5418s
    GENERIC MAP (widthcc=>widthcc,pipes=>pipes)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              dataaa=>dataaa,databb=>databb,
              result=>result);
              
  END GENERATE;
  
  gforone: IF ((widthaa = 54) AND 
               (widthbb = 54) AND 
               (widthcc = 72) AND
               (accuracy = 1) AND
               (device = 1) AND
               (synthesize = 1)) GENERATE
            
    mulforone: fp_mul54us_3xs
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              mulaa=>dataaa,mulbb=>databb,
              mulcc=>result);
          
  END GENERATE;
  
  gfortwo: IF ((widthaa = 54) AND 
               (widthbb = 54) AND 
               (widthcc = 72) AND
               (accuracy = 0) AND
               (device = 1) AND
               (synthesize = 1)) GENERATE
            
    mulfortwo: fp_mul54us_38s
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              mulaa=>dataaa,mulbb=>databb,
              mulcc=>result);
          
  END GENERATE;
  
  gforthr: IF ((widthaa = 54) AND 
               (widthbb = 54) AND 
               (widthcc = 72) AND
               (accuracy = 0) AND
               (device = 0) AND
               (synthesize = 1) AND
               ((pipes = 5) OR (pipes = 6))) GENERATE
            
    mulforthr: fp_mul54us_28s
    GENERIC MAP (latency=>pipes)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              mulaa=>dataaa,mulbb=>databb,
              mulcc=>result);
          
  END GENERATE;
  
  gforfor: IF ((widthaa = 54) AND 
               (widthbb = 54) AND 
               (widthcc = 72) AND
               (accuracy = 1) AND
               (device = 0) AND
               (synthesize = 1) AND
               ((pipes = 5) OR (pipes = 6))) GENERATE
            
    mulforfor: fp_mul54us_29s
    GENERIC MAP (latency=>pipes)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              mulaa=>dataaa,mulbb=>databb,
              mulcc=>result);
          
  END GENERATE;

  gforfiv: IF ((widthaa = 54) AND 
               (widthbb = 54) AND 
               (widthcc = 72) AND
               (synthesize = 0)) GENERATE
            
    mulforfiv: fp_mul54usb
    GENERIC MAP (latency=>pipes,device=>device,prune=>accuracy)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>dataaa,bb=>databb,
              cc=>result);
          
  END GENERATE;
		  
  gfiv: IF ((widthaa = 72) AND 
            (widthbb = 18) AND 
            (widthcc < 90) AND
            ((pipes = 3) OR (pipes = 4))) GENERATE
            
    multhr: fp_mul7218s
    GENERIC MAP (widthcc=>widthcc,pipes=>pipes)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              dataaa=>dataaa,databb=>databb,
              result=>result);
              
  END GENERATE;
  		          
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   SINGLE PRECISION INVERSE - TOP LEVEL      ***
--***                                             ***
--***   FP_INV.VHD                                ***
--***                                             ***
--***   Function: IEEE754 SP Inverse              ***
--***   (multiplicative iterative algorithm)      ***
--***                                             ***
--***   09/12/07 ML                               ***
--***                                             ***
--***   (c) 2007 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes: Latency = 14                         ***
--***************************************************

ENTITY fp_inv IS 
GENERIC (synthesize : integer := 1);
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (23 DOWNTO 1);

		signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
      --------------------------------------------------
      nanout : OUT STD_LOGIC;
      invalidout : OUT STD_LOGIC;
      dividebyzeroout : OUT STD_LOGIC
		);
END fp_inv;

ARCHITECTURE div OF fp_inv IS
  
  constant expwidth : positive := 8;
  constant manwidth : positive := 23;
  
  constant coredepth : positive := 12;
  
  type expfftype IS ARRAY (coredepth-1 DOWNTO 1) OF STD_LOGIC_VECTOR (expwidth+2 DOWNTO 1);
  
  signal zerovec : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
    
  signal signinff : STD_LOGIC;
  signal manff : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal expinff : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal expoffset : STD_LOGIC_VECTOR (expwidth+2 DOWNTO 1);
  signal invertnum : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal quotient : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal signff : STD_LOGIC_VECTOR (coredepth-1 DOWNTO 1);  
  signal expff : expfftype; 

  -- conditions
  signal zeroman : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal zeroexp : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal maxexp : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal zeromaninff : STD_LOGIC;
  signal zeroexpinff : STD_LOGIC;
  signal maxexpinff : STD_LOGIC;
  signal zeroinff : STD_LOGIC;
  signal infinityinff : STD_LOGIC;
  signal naninff : STD_LOGIC;
  signal dividebyzeroff, nanff : STD_LOGIC_VECTOR (coredepth-3 DOWNTO 1);

  component fp_inv_core IS 
  GENERIC (synthesize : integer := 1); 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        divisor : IN STD_LOGIC_VECTOR (36 DOWNTO 1);

		  quotient : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
		  );
  end component;
  
  component fp_divrnd 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        signin : IN STD_LOGIC;
        exponentdiv : IN STD_LOGIC_VECTOR (expwidth+2 DOWNTO 1);
        mantissadiv : IN STD_LOGIC_VECTOR (manwidth+1 DOWNTO 1);
        nanin : IN STD_LOGIC;
        dividebyzeroin : IN STD_LOGIC;

		  signout : OUT STD_LOGIC;
        exponentout : OUT STD_LOGIC_VECTOR (expwidth DOWNTO 1);
        mantissaout : OUT STD_LOGIC_VECTOR (manwidth DOWNTO 1);
        --------------------------------------------------
        nanout : OUT STD_LOGIC;
        invalidout : OUT STD_LOGIC;
        dividebyzeroout : OUT STD_LOGIC
		  );
  end component;
  
BEGIN
    
  gzva: FOR k IN 1 TO manwidth GENERATE
    zerovec(k) <= '0';
  END GENERATE;

  gxa: FOR k IN 1 TO expwidth-1 GENERATE
    expoffset(k) <= '1';
  END GENERATE;
  expoffset(expwidth+2 DOWNTO expwidth) <= "000";

  pma: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
  
      FOR k IN 1 TO manwidth LOOP
        manff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        expinff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO coredepth-1 LOOP
        signff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO coredepth-1 LOOP
        FOR j IN 1 TO expwidth+2 LOOP
          expff(k)(j) <= '0';
        END LOOP;
      END LOOP;
    
    ELSIF (rising_edge(sysclk)) THEN

      IF (enable = '1') THEN
        
        signinff <= signin;
        manff <= mantissain;
        expinff <= exponentin;

        signff(1) <= signinff;
        FOR k IN 2 TO coredepth-1 LOOP
          signff(k) <= signff(k-1);
        END LOOP;
    
        expff(1)(expwidth+2 DOWNTO 1) <= expoffset - ("00" & expinff);
        expff(2)(expwidth+2 DOWNTO 1) <= expff(1)(expwidth+2 DOWNTO 1) + expoffset;
        FOR k IN 3 TO coredepth-2 LOOP
          expff(k)(expwidth+2 DOWNTO 1) <= expff(k-1)(expwidth+2 DOWNTO 1);
        END LOOP;
        -- inverse always less than 1, decrement exponent
        expff(coredepth-1)(expwidth+2 DOWNTO 1) <= expff(coredepth-2)(expwidth+2 DOWNTO 1) - 
                                                  (zerovec(expwidth+1 DOWNTO 1) & '1');   
    
      END IF;
  
    END IF;
  
  END PROCESS;

--********************
--*** CHECK INPUTS ***
--********************

  zeroman(1) <= manff(1);
  gca: FOR k IN 2 TO manwidth GENERATE
    zeroman(k) <= zeroman(k-1) OR manff(k);
  END GENERATE; 
  zeroexp(1) <= expinff(1);
  gcb: FOR k IN 2 TO expwidth GENERATE
    zeroexp(k) <= zeroexp(k-1) OR expinff(k);
  END GENERATE;
  maxexp(1) <= expinff(1);
  gcc: FOR k IN 2 TO expwidth GENERATE
    maxexp(k) <= maxexp(k-1) AND expinff(k);
  END GENERATE;

  pcc: PROCESS (sysclk,reset)
  BEGIN
    
    IF (reset = '1') THEN
      
      zeromaninff <= '0';  
      zeroexpinff <= '0'; 
      maxexpinff <= '0';  
      zeroinff <= '0';
      infinityinff <= '0';
      naninff <= '0';
      FOR k IN 1 TO coredepth-3 LOOP
        dividebyzeroff(k) <= '0';
        nanff(k) <= '0';
      END LOOP;
     
    ELSIF (rising_edge(sysclk)) THEN
            
      IF (enable = '1') THEN
     
        zeromaninff <= zeroman(manwidth);
        zeroexpinff <= zeroexp(expwidth);
        maxexpinff <= maxexp(expwidth);
    
        -- zero when man = 0, exp = 0
        -- infinity when man = 0, exp = max
        -- nan when man != 0, exp = max
    
        -- all ffs '1' when condition true
        zeroinff <= NOT(zeromaninff OR zeroexpinff); 
        infinityinff <= NOT(zeromaninff) AND maxexpinff;
        naninff <= zeromaninff AND maxexpinff;

        -- nan output when nan input
        nanff(1) <= naninff;
        FOR k IN 2 TO coredepth-3 LOOP
          nanff(k) <= nanff(k-1);
        END LOOP;
        
        dividebyzeroff(1) <= zeroinff;
        FOR k IN 2 TO coredepth-3 LOOP
          dividebyzeroff(k) <= dividebyzeroff(k-1);
        END LOOP;
      
      END IF;
   
    END IF;

  END PROCESS;


--*******************
--*** DIVIDE CORE ***
--*******************

  invertnum <= '1' & mantissain & "000000000000";

  -- will give output between 0.5 and 0.99999...
  -- will always need to be normalized
  invcore: fp_inv_core
  GENERIC MAP (synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            divisor=>invertnum,
            quotient=>quotient);

--************************
--*** ROUND AND OUTPUT ***
--************************

  rndout: fp_divrnd
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            signin=>signff(coredepth-1),
            exponentdiv=>expff(coredepth-1)(expwidth+2 DOWNTO 1),
            mantissadiv=>quotient(34 DOWNTO 11),
            nanin=>nanff(coredepth-3),dividebyzeroin=>dividebyzeroff(coredepth-3),

            signout=>signout,exponentout=>exponentout,mantissaout=>mantissaout,
            nanout=>nanout,invalidout=>invalidout,dividebyzeroout=>dividebyzeroout);
  
END div;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   SINGLE PRECISION INVERSE - CORE           ***
--***                                             ***
--***   FP_INV_CORE.VHD                           ***
--***                                             ***
--***   Function: 36 bit Inverse                  ***
--***   (multiplicative iterative algorithm)      ***
--***                                             ***
--***   09/12/07 ML                               ***
--***                                             ***
--***   (c) 2007 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes: Latency = 12                         ***
--***************************************************

ENTITY fp_inv_core IS 
GENERIC (synthesize : integer := 1); 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      divisor : IN STD_LOGIC_VECTOR (36 DOWNTO 1);

		quotient : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
		);
END fp_inv_core;

ARCHITECTURE rtl OF fp_inv_core IS

  signal zerovec : STD_LOGIC_VECTOR (36 DOWNTO 1);
  
  signal divisordel : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal invdivisor : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal delinvdivisor : STD_LOGIC_VECTOR (18 DOWNTO 1);
  
  signal scaleden : STD_LOGIC_VECTOR (36 DOWNTO 1);
  
  signal twonode : STD_LOGIC_VECTOR (37 DOWNTO 1);
  signal nextguessff : STD_LOGIC_VECTOR (37 DOWNTO 1);
          
  signal quotientnode : STD_LOGIC_VECTOR (36 DOWNTO 1);
  
  component fp_div_est IS 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        divisor : IN STD_LOGIC_VECTOR (19 DOWNTO 1);

		  invdivisor : OUT STD_LOGIC_VECTOR (18 DOWNTO 1)
		  );
  end component;
  
  component fp_fxmul IS 
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36;
           pipes : positive := 1;
           accuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1); 
      
        result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
       );
  end component;

  component fp_del
  GENERIC (
           width : positive := 64;
           pipes : positive := 2
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
       
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
   end component;  
       
BEGIN
  
  gza: FOR k IN 1 TO 36 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  invcore: fp_div_est
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            divisor=>divisor(36 DOWNTO 18),invdivisor=>invdivisor);
  
  delinone: fp_del
  GENERIC MAP (width=>36,pipes=>5)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>divisor,cc=>divisordel);

  --**********************************
  --*** ITERATION 0 - SCALE INPUTS ***
  --**********************************
  
  -- in level 5, out level 8
  mulscaleone: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>18,widthcc=>36,
               pipes=>3,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>divisordel,databb=>invdivisor,
            result=>scaleden);
              
  --********************
  --*** ITERATION 1  ***
  --********************

  twonode <= '1' & zerovec(36 DOWNTO 1);
  
  pita: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN

      FOR k IN 1 TO 37 LOOP
        nextguessff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN
        nextguessff <= twonode - ('0' & scaleden); -- level 9
      END IF;
    
    END IF;
    
  END PROCESS;
  
  deloneone: fp_del
  GENERIC MAP (width=>18,pipes=>4)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>invdivisor,
            cc=>delinvdivisor);
 
  -- in level 9, out level 12
  muloneone: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>18,widthcc=>36,
               pipes=>3,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>nextguessff(36 DOWNTO 1),databb=>delinvdivisor,
            result=>quotientnode);
 
  quotient <= quotientnode(36 DOWNTO 1);
                  
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   SINGLE PRECISION INVERSE SQUARE ROOT      ***
--***               TOP LEVEL                     ***
--***                                             ***
--***   FP_INV.VHD                                ***
--***                                             ***
--***   Function: IEEE754 SP Inverse Square Root  ***
--***   (multiplicative iterative algorithm)      ***
--***                                             ***
--***   09/12/07 ML                               ***
--***                                             ***
--***   (c) 2007 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes: Latency = 19                         ***
--***************************************************

ENTITY fp_invsqr IS 
GENERIC (synthesize : integer := 1); 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin: IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (23 DOWNTO 1);

		signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
      --------------------------------------------------
      nanout : OUT STD_LOGIC;
      invalidout : OUT STD_LOGIC
		);
END fp_invsqr;

ARCHITECTURE rtl OF fp_invsqr IS
  
  constant manwidth : positive := 23;
  constant expwidth : positive := 8;
  
  constant coredepth : positive := 17;
  
  type expfftype IS ARRAY (coredepth+2 DOWNTO 1) OF STD_LOGIC_VECTOR (expwidth DOWNTO 1);

  signal maninff : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal expinff : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal signff : STD_LOGIC_VECTOR (coredepth+2 DOWNTO 1);
  signal correctff : STD_LOGIC_VECTOR (3 DOWNTO 1);  -- 09/03/11 ML
  signal expff : expfftype;
  signal radicand : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal oddexponent : STD_LOGIC;
  signal invroot : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal roundff : STD_LOGIC_VECTOR (manwidth DOWNTO 1); 
  signal manff : STD_LOGIC_VECTOR (manwidth DOWNTO 1); 
  signal zerovec : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal offset : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
    
  -- conditions
  signal nanmanff, nanexpff : STD_LOGIC_VECTOR (coredepth DOWNTO 1);
  signal zeroexpff, zeromanff : STD_LOGIC_VECTOR (coredepth-1 DOWNTO 1); 
  signal expinzero, expinmax : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal maninzero : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal expzero, expmax, manzero : STD_LOGIC;
  signal infinityconditionff, nanconditionff, expzeroff : STD_LOGIC;
  signal correct_powers_of_two : STD_LOGIC;  -- 09/03/11 ML
    
  component fp_invsqr_core IS 
  GENERIC (synthesize : integer := 1); -- 0/1 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        radicand : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
        odd : IN STD_LOGIC;

		  invroot : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
		  );
  end component;
	
BEGIN
    
  gzva: FOR k IN 1 TO manwidth GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  gxoa: FOR k IN 1 TO expwidth-1 GENERATE
    offset(k) <= '1';
  END GENERATE;
  offset(expwidth) <= '0';

  pma: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN

      FOR k IN 1 TO manwidth LOOP
        maninff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        expinff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO coredepth+2 LOOP
        signff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO coredepth+2 LOOP
        FOR j IN 1 TO expwidth LOOP
          expff(k)(j) <= '0';
        END LOOP;
      END LOOP;
      FOR k IN 1 TO manwidth LOOP
        roundff(k) <= '0';
        manff(k) <= '0';
      END LOOP;
      correctff <= "000";  -- 09/03/11 ML
  
    ELSIF (rising_edge(sysclk)) THEN

      maninff <= mantissain;
      expinff <= exponentin;
    
      signff(1) <= signin;
      FOR k IN 2 TO coredepth+2 LOOP
        signff(k) <= signff(k-1);
      END LOOP;
  
      expff(1)(expwidth DOWNTO 1) <= exponentin;
      expff(2)(expwidth DOWNTO 1) <= expff(1)(expwidth DOWNTO 1) - offset;
      expff(3)(expwidth DOWNTO 1) <= expff(2)(expwidth) & expff(2)(expwidth DOWNTO 2);
      expff(4)(expwidth DOWNTO 1) <= offset - expff(3)(expwidth DOWNTO 1);
      expff(5)(expwidth DOWNTO 1) <= expff(4)(expwidth DOWNTO 1) - 1 + correctff(3);  -- 09/03/11 ML
      FOR k IN 6 TO coredepth+1 LOOP
        expff(k)(expwidth DOWNTO 1) <= expff(k-1)(expwidth DOWNTO 1);
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        expff(coredepth+2)(k) <= (expff(coredepth+1)(k) AND zeroexpff(coredepth-1)) OR nanexpff(coredepth-1);
      END LOOP;
      
      -- 09/03/11 ML
      correctff(1) <= correct_powers_of_two;
      correctff(2) <= correctff(1);
      correctff(3) <= correctff(2);
    
      roundff <= invroot(35 DOWNTO 13) + (zerovec(22 DOWNTO 1) & invroot(12));
    
      -- invroot 36, so mantissa is at 35:13
      FOR k IN 1 TO manwidth LOOP
        manff(k) <= (roundff(k) AND zeromanff(coredepth-1)) OR nanmanff(coredepth-1);
      END LOOP;
  
    END IF;
  
  END PROCESS;

--*******************
--*** CONDITIONS ***
--*******************

  pcc: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
      
      FOR k IN 1 TO coredepth LOOP
        nanmanff(k) <= '0';
        nanexpff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO coredepth-1 LOOP
        zeroexpff(k) <= '0';
        zeromanff(k) <= '0';
      END LOOP;
      infinityconditionff <= '0'; 
      nanconditionff <= '0';
      expzeroff <= '0';

    ELSIF (rising_edge(sysclk)) THEN
     
      infinityconditionff <= manzero AND expmax;
      nanconditionff <= signff(1) OR expzero OR (expmax AND manzero);
      expzeroff <= expzero;
 
      nanmanff(1) <= nanconditionff; -- level 3
      nanexpff(1) <= nanconditionff OR infinityconditionff; -- also max exp when infinity
      FOR k IN 2 TO coredepth LOOP
        nanmanff(k) <= nanmanff(k-1);
        nanexpff(k) <= nanexpff(k-1);
      END LOOP;

      zeromanff(1) <= NOT(expzeroff) AND NOT(infinityconditionff); -- level 3
      zeroexpff(1) <= NOT(expzeroff); -- level 3
      FOR k IN 2 TO coredepth-1 LOOP
        zeromanff(k) <= zeromanff(k-1);
        zeroexpff(k) <= zeroexpff(k-1);
      END LOOP;
    
    END IF;
  
  END PROCESS;

--*******************
--*** SQUARE ROOT ***
--*******************

  radicand <= '1' & mantissain & "000000000000";
  -- sub 127, so 127 (odd) = 2^0 => even
  oddexponent <= NOT(exponentin(1));

  -- does not require rounding, output of core rounded already, LSB always 0
  isqr: fp_invsqr_core
  GENERIC MAP (synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            radicand=>radicand,odd=>oddexponent,
            invroot=>invroot);
		
--*********************
--*** SPECIAL CASES ***
--*********************
-- 1. if negative input, invalid operation, NAN 
-- 2. 0 in, invalid operation, NAN
-- 3. infinity in, invalid operation, infinity out
-- 4. NAN in, invalid operation, NAN

  -- '1' if 0 
  expinzero(1) <= expinff(1);
  gxza: FOR k IN 2 TO expwidth GENERATE
    expinzero(k) <= expinzero(k-1) OR expinff(k);
  END GENERATE;
  expzero <= NOT(expinzero(expwidth)); -- '0' when zero
                 
  -- '1' if nan or infinity
  expinmax(1) <= expinff(1);
  gxia: FOR k IN 2 TO expwidth GENERATE
    expinmax(k) <= expinmax(k-1) AND expinff(k);
  END GENERATE;
  expmax <= expinmax(expwidth); -- '1' when true
          
  -- '1' if zero or infinity
  maninzero(1) <= maninff(1);
  gmza: FOR k IN 2 TO manwidth GENERATE
    maninzero(k) <= maninzero(k-1) OR maninff(k);
  END GENERATE;
  manzero <= NOT(maninzero(manwidth)); 
  
  -- 09/03/11 ML
  -- if mantissa is 0 and exponent is odd (...123,125,127,129,131...) then dont subtract 1 from offset corrected exponent
  -- '1' is subtracted as any value, no matter how small, in the mantissa will reduce the inverse below the mirrored exponent (around 127)
  -- if the exponent is odd (with mantissa 0) the value is a power of 2 (...0.25,0.5,1,2,4...) and the mirrored exponent is correct
  -- if the exponent is even (with mantissa 0), the inverse square root will have a non zero mantissa and can be handled normally
  correct_powers_of_two <= manzero AND expinff(1);
       
--***************
--*** OUTPUTS ***
--***************

  signout <= signff(coredepth+2);
  exponentout <= expff(coredepth+2)(expwidth DOWNTO 1);   
  mantissaout <= manff;  
  -----------------------------------------------
  nanout <= nanmanff(coredepth);
  invalidout <= nanmanff(coredepth);

END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   SINGLE PRECISION INVERSE SQUARE ROOT      ***
--***                 CORE                        ***
--***                                             ***
--***   FP_INVSQR_CORE.VHD                        ***
--***                                             ***
--***   Function: 36 bit Inverse Square Root      ***
--***   (multiplicative iterative algorithm)      ***
--***                                             ***
--***   09/12/07 ML                               ***
--***                                             ***
--***   (c) 2007 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes: Latency = 17                         ***
--***************************************************

ENTITY fp_invsqr_core IS 
GENERIC (
         synthesize : integer := 1      -- 0/1      
        ); 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      radicand : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
      odd : IN STD_LOGIC;

		invroot : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
		);
END fp_invsqr_core;

ARCHITECTURE rtl OF fp_invsqr_core IS
  
  signal zerovec : STD_LOGIC_VECTOR (36 DOWNTO 1);
  
  signal evennum : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal oddnum : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal guessvec : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal oddff : STD_LOGIC_VECTOR (12 DOWNTO 1);
  signal scalenumff : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal guess : STD_LOGIC_VECTOR (18 DOWNTO 1);

  -- 1st iteration
  signal radicanddelone : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal guessdel : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal multoneone : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal multonetwo : STD_LOGIC_VECTOR (37 DOWNTO 1);
  signal multonetwoff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal suboneff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal multonethr : STD_LOGIC_VECTOR (37 DOWNTO 1);

  component fp_invsqr_est IS 
  GENERIC (synthesize : integer := 0); -- 0 = behavioral, 1 = syntheziable
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        radicand : IN STD_LOGIC_VECTOR (19 DOWNTO 1);

		  invroot : OUT STD_LOGIC_VECTOR (18 DOWNTO 1)
		  );
  end component;
  
  component fp_fxmul IS 
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36;
           pipes : positive := 1;
           accuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1); 
      
        result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
       ); 
  end component;
 
  component fp_del
  GENERIC (
           width : positive := 64;
           pipes : positive := 2
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
       
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
   end component;
   		 
BEGIN
    
  oddnum <= conv_std_logic_vector(185363,18); -- mult by 2^-.5 (odd exp)
  evennum <= conv_std_logic_vector(262143,18); -- mult by 1 (even exp)
  
  gza: FOR k IN 1 TO 36 GENERATE
    zerovec(k) <= '0';
  END GENERATE;

  -- in level 0, out level 5
  look: fp_invsqr_est
  GENERIC MAP (synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            radicand=>radicand(36 DOWNTO 18),invroot=>guessvec);
              
  pta: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN
    
      FOR k IN 1 TO 12 LOOP
        oddff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 18 LOOP
        scalenumff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF (enable = '1') THEN
        
        oddff(1) <= odd;
        FOR k IN 2 TO 12 LOOP
          oddff(k) <= oddff(k-1);
        END LOOP; 
        
        FOR k IN 1 TO 18 LOOP
          scalenumff(k) <= (oddnum(k) AND oddff(4)) OR (evennum(k) AND NOT(oddff(4)));
        END LOOP;
          
      END IF;
    
    END IF;    
      
  END PROCESS;

  -- in level 5, out level 7
  mulscale: fp_fxmul
  GENERIC MAP (widthaa=>18,widthbb=>18,widthcc=>18,pipes=>2,
               synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>guessvec,databb=>scalenumff,
            result=>guess);

  --*********************
  --*** ITERATION ONE ***
  --*********************
  --X' = X/2(3-YXX)
  
  deloneone: fp_del
  GENERIC MAP(width=>36,pipes=>9)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>radicand,cc=>radicanddelone);
            
  delonetwo: fp_del
  GENERIC MAP(width=>18,pipes=>7)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>guess,cc=>guessdel);
            
  -- in level 7, out level 9 (18x18=36)
  oneone: fp_fxmul
  GENERIC MAP (widthaa=>18,widthbb=>18,widthcc=>36,pipes=>2,
               synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>guess,databb=>guess,
            result=>multoneone);
                   
  -- in level 9, out level 12 (36x36=37)
  onetwo: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>36,widthcc=>37,pipes=>3,
               synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>radicanddelone,databb=>multoneone,
            result=>multonetwo);
                   
  -- multonetwo is about 1 - either 1.000000XXX or 0.9999999
  -- mult by 2 if odd exponent (37 DOWNTO 2), otherwise (38 DOWNTO 3)
  -- round bit in position 1 or 2
  pone: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN

      FOR k IN 1 TO 36 LOOP
        multonetwoff(k) <= '0';
        suboneff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF (enable = '1') THEN
        
        --invert here so that borrow can be added in simple expression
        -- level 13
        FOR k IN 1 TO 36 LOOP
          multonetwoff(k) <= NOT((multonetwo(k) AND oddff(12)) OR (multonetwo(k+1) AND NOT(oddff(12))));
        END LOOP;
        -- level 14
        suboneff <= ("11" & zerovec(34 DOWNTO 1)) + 
                    ('1' & multonetwoff(36 DOWNTO 2)) +
                    (zerovec(35 DOWNTO 1) & multonetwoff(1));
          
      END IF;
    
    END IF;    
      
  END PROCESS;    

  -- in level 14, out level 17 (36x18=37)
  onethr: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>18,widthcc=>37,pipes=>3,
               synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>suboneff,databb=>guessdel,
            result=>multonethr); 

  invroot <= multonethr(36 DOWNTO 1);
   
END rtl;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_INVSQR_EST.VHD                         ***
--***                                             ***
--***   Function: Estimates 18 Bit Inverse Root   ***
--***                                             ***
--***   Used by both single and double inverse    ***
--***   square root cores                         ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** 1. Inverse square root of 18 bit header     ***
--*** (not including leading '1')                 ***
--*** 2. Uses 20 bit precision tables - 18 bits   ***
--*** drops a bit occasionally                    ***
--***************************************************

ENTITY fp_invsqr_est IS 
GENERIC (synthesize : integer := 0); -- 0 = behavioral, 1 = syntheziable
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      radicand : IN STD_LOGIC_VECTOR (19 DOWNTO 1);

		invroot : OUT STD_LOGIC_VECTOR (18 DOWNTO 1)
		);
END fp_invsqr_est;

ARCHITECTURE rtl OF fp_invsqr_est IS

  type smalldelfftype IS ARRAY (2 DOWNTO 1) OF STD_LOGIC_VECTOR (9 DOWNTO 1);
  type largedelfftype IS ARRAY (2 DOWNTO 1) OF STD_LOGIC_VECTOR (20 DOWNTO 1);
  
  signal zerovec : STD_LOGIC_VECTOR (9 DOWNTO 1);
  signal one, two : STD_LOGIC_VECTOR (9 DOWNTO 1);
  signal oneaddff, zipaddff : STD_LOGIC_VECTOR (9 DOWNTO 1);
  signal twodelff : smalldelfftype;
  signal onelut, onelutff : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal ziplut, ziplutff : STD_LOGIC_VECTOR (20 DOWNTO 1);
  signal ziplutdelff : largedelfftype;
  signal onetwo : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal invrootff : STD_LOGIC_VECTOR (20 DOWNTO 1);

  component fp_invsqr_lut1 IS
  PORT (
        add : IN STD_LOGIC_VECTOR (9 DOWNTO 1);
		  data : OUT STD_LOGIC_VECTOR (11 DOWNTO 1)
       );
  end component;
    
  component fp_invsqr_lut0 IS
  PORT (
        add : IN STD_LOGIC_VECTOR (9 DOWNTO 1);
		  data : OUT STD_LOGIC_VECTOR (20 DOWNTO 1)
       );
  end component;
  
  component fp_fxmul IS 
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36;
           pipes : positive := 1;
           accuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1); 
      
        result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
       ); 
  end component;
		    
BEGIN
  
  gza: FOR k IN 1 TO 9 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  one <= radicand(18 DOWNTO 10);
  two <= radicand(9 DOWNTO 1);
  
  ppa: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN
    
      FOR k IN 1 TO 9 LOOP
        oneaddff(k) <= '0';
        zipaddff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 2 LOOP
        FOR j IN 1 TO 9 LOOP
          twodelff(k)(j) <= '0';
        END LOOP;
      END LOOP;
      FOR k IN 1 TO 11 LOOP
        onelutff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 20 LOOP
        ziplutff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 2 LOOP
        FOR j IN 1 TO 20 LOOP
          ziplutdelff(k)(j) <= '0';
        END LOOP;
      END LOOP;
      FOR k IN 1 TO 18 LOOP
        invrootff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF (enable = '1') THEN
      
        oneaddff <= one;
        zipaddff <= one;
      
        twodelff(1)(9 DOWNTO 1) <= two;
        twodelff(2)(9 DOWNTO 1) <= twodelff(1)(9 DOWNTO 1);
      
        onelutff <= onelut;
        ziplutff <= ziplut;
        
        ziplutdelff(1)(20 DOWNTO 1) <= ziplutff;
        ziplutdelff(2)(20 DOWNTO 1) <= ziplutdelff(1)(20 DOWNTO 1);
        
        invrootff <= ziplutdelff(2)(20 DOWNTO 1) - (zerovec(9 DOWNTO 1) & onetwo);
        
      END IF;
      
    END IF;
    
      
  END PROCESS;
     
  upper: fp_invsqr_lut1 PORT MAP (add=>oneaddff,data=>onelut);
  
  lower: fp_invsqr_lut0 PORT MAP (add=>zipaddff,data=>ziplut);
  
  mulcore: fp_fxmul
  GENERIC MAP (widthaa=>11,widthbb=>9,widthcc=>11,pipes=>2)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>onelutff,databb=>twodelff(2)(9 DOWNTO 1),
            result=>onetwo);
  
  --**************
  --*** OUTPUT ***
  --**************
  
  invroot <= invrootff(20 DOWNTO 3);  
    
END rtl;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_INVSQR_LUT0.VHD                        ***
--***                                             ***
--***   Function: Look Up Table - Inverse Root    ***
--***                                             ***
--***   Generated by MATLAB Utility               ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_invsqr_lut0 IS
PORT (
      add : IN STD_LOGIC_VECTOR (9 DOWNTO 1);
		data : OUT STD_LOGIC_VECTOR (20 DOWNTO 1)
);
END fp_invsqr_lut0;

ARCHITECTURE rtl OF fp_invsqr_lut0 IS

BEGIN

  pca: PROCESS (add)
  BEGIN
    CASE add IS
      WHEN "000000000" => data <= conv_std_logic_vector(1048575,20);
      WHEN "000000001" => data <= conv_std_logic_vector(1047553,20);
      WHEN "000000010" => data <= conv_std_logic_vector(1046534,20);
      WHEN "000000011" => data <= conv_std_logic_vector(1045517,20);
      WHEN "000000100" => data <= conv_std_logic_vector(1044503,20);
      WHEN "000000101" => data <= conv_std_logic_vector(1043493,20);
      WHEN "000000110" => data <= conv_std_logic_vector(1042485,20);
      WHEN "000000111" => data <= conv_std_logic_vector(1041480,20);
      WHEN "000001000" => data <= conv_std_logic_vector(1040478,20);
      WHEN "000001001" => data <= conv_std_logic_vector(1039479,20);
      WHEN "000001010" => data <= conv_std_logic_vector(1038483,20);
      WHEN "000001011" => data <= conv_std_logic_vector(1037490,20);
      WHEN "000001100" => data <= conv_std_logic_vector(1036500,20);
      WHEN "000001101" => data <= conv_std_logic_vector(1035512,20);
      WHEN "000001110" => data <= conv_std_logic_vector(1034527,20);
      WHEN "000001111" => data <= conv_std_logic_vector(1033545,20);
      WHEN "000010000" => data <= conv_std_logic_vector(1032566,20);
      WHEN "000010001" => data <= conv_std_logic_vector(1031589,20);
      WHEN "000010010" => data <= conv_std_logic_vector(1030616,20);
      WHEN "000010011" => data <= conv_std_logic_vector(1029645,20);
      WHEN "000010100" => data <= conv_std_logic_vector(1028677,20);
      WHEN "000010101" => data <= conv_std_logic_vector(1027711,20);
      WHEN "000010110" => data <= conv_std_logic_vector(1026749,20);
      WHEN "000010111" => data <= conv_std_logic_vector(1025789,20);
      WHEN "000011000" => data <= conv_std_logic_vector(1024831,20);
      WHEN "000011001" => data <= conv_std_logic_vector(1023877,20);
      WHEN "000011010" => data <= conv_std_logic_vector(1022925,20);
      WHEN "000011011" => data <= conv_std_logic_vector(1021975,20);
      WHEN "000011100" => data <= conv_std_logic_vector(1021029,20);
      WHEN "000011101" => data <= conv_std_logic_vector(1020084,20);
      WHEN "000011110" => data <= conv_std_logic_vector(1019143,20);
      WHEN "000011111" => data <= conv_std_logic_vector(1018204,20);
      WHEN "000100000" => data <= conv_std_logic_vector(1017268,20);
      WHEN "000100001" => data <= conv_std_logic_vector(1016334,20);
      WHEN "000100010" => data <= conv_std_logic_vector(1015403,20);
      WHEN "000100011" => data <= conv_std_logic_vector(1014474,20);
      WHEN "000100100" => data <= conv_std_logic_vector(1013548,20);
      WHEN "000100101" => data <= conv_std_logic_vector(1012625,20);
      WHEN "000100110" => data <= conv_std_logic_vector(1011704,20);
      WHEN "000100111" => data <= conv_std_logic_vector(1010785,20);
      WHEN "000101000" => data <= conv_std_logic_vector(1009869,20);
      WHEN "000101001" => data <= conv_std_logic_vector(1008956,20);
      WHEN "000101010" => data <= conv_std_logic_vector(1008045,20);
      WHEN "000101011" => data <= conv_std_logic_vector(1007136,20);
      WHEN "000101100" => data <= conv_std_logic_vector(1006230,20);
      WHEN "000101101" => data <= conv_std_logic_vector(1005327,20);
      WHEN "000101110" => data <= conv_std_logic_vector(1004425,20);
      WHEN "000101111" => data <= conv_std_logic_vector(1003527,20);
      WHEN "000110000" => data <= conv_std_logic_vector(1002630,20);
      WHEN "000110001" => data <= conv_std_logic_vector(1001736,20);
      WHEN "000110010" => data <= conv_std_logic_vector(1000845,20);
      WHEN "000110011" => data <= conv_std_logic_vector(999955,20);
      WHEN "000110100" => data <= conv_std_logic_vector(999068,20);
      WHEN "000110101" => data <= conv_std_logic_vector(998184,20);
      WHEN "000110110" => data <= conv_std_logic_vector(997302,20);
      WHEN "000110111" => data <= conv_std_logic_vector(996422,20);
      WHEN "000111000" => data <= conv_std_logic_vector(995544,20);
      WHEN "000111001" => data <= conv_std_logic_vector(994669,20);
      WHEN "000111010" => data <= conv_std_logic_vector(993796,20);
      WHEN "000111011" => data <= conv_std_logic_vector(992926,20);
      WHEN "000111100" => data <= conv_std_logic_vector(992057,20);
      WHEN "000111101" => data <= conv_std_logic_vector(991191,20);
      WHEN "000111110" => data <= conv_std_logic_vector(990327,20);
      WHEN "000111111" => data <= conv_std_logic_vector(989466,20);
      WHEN "001000000" => data <= conv_std_logic_vector(988607,20);
      WHEN "001000001" => data <= conv_std_logic_vector(987750,20);
      WHEN "001000010" => data <= conv_std_logic_vector(986895,20);
      WHEN "001000011" => data <= conv_std_logic_vector(986042,20);
      WHEN "001000100" => data <= conv_std_logic_vector(985192,20);
      WHEN "001000101" => data <= conv_std_logic_vector(984344,20);
      WHEN "001000110" => data <= conv_std_logic_vector(983498,20);
      WHEN "001000111" => data <= conv_std_logic_vector(982654,20);
      WHEN "001001000" => data <= conv_std_logic_vector(981812,20);
      WHEN "001001001" => data <= conv_std_logic_vector(980973,20);
      WHEN "001001010" => data <= conv_std_logic_vector(980135,20);
      WHEN "001001011" => data <= conv_std_logic_vector(979300,20);
      WHEN "001001100" => data <= conv_std_logic_vector(978467,20);
      WHEN "001001101" => data <= conv_std_logic_vector(977636,20);
      WHEN "001001110" => data <= conv_std_logic_vector(976807,20);
      WHEN "001001111" => data <= conv_std_logic_vector(975980,20);
      WHEN "001010000" => data <= conv_std_logic_vector(975156,20);
      WHEN "001010001" => data <= conv_std_logic_vector(974333,20);
      WHEN "001010010" => data <= conv_std_logic_vector(973513,20);
      WHEN "001010011" => data <= conv_std_logic_vector(972694,20);
      WHEN "001010100" => data <= conv_std_logic_vector(971878,20);
      WHEN "001010101" => data <= conv_std_logic_vector(971063,20);
      WHEN "001010110" => data <= conv_std_logic_vector(970251,20);
      WHEN "001010111" => data <= conv_std_logic_vector(969441,20);
      WHEN "001011000" => data <= conv_std_logic_vector(968633,20);
      WHEN "001011001" => data <= conv_std_logic_vector(967827,20);
      WHEN "001011010" => data <= conv_std_logic_vector(967022,20);
      WHEN "001011011" => data <= conv_std_logic_vector(966220,20);
      WHEN "001011100" => data <= conv_std_logic_vector(965420,20);
      WHEN "001011101" => data <= conv_std_logic_vector(964622,20);
      WHEN "001011110" => data <= conv_std_logic_vector(963826,20);
      WHEN "001011111" => data <= conv_std_logic_vector(963031,20);
      WHEN "001100000" => data <= conv_std_logic_vector(962239,20);
      WHEN "001100001" => data <= conv_std_logic_vector(961449,20);
      WHEN "001100010" => data <= conv_std_logic_vector(960660,20);
      WHEN "001100011" => data <= conv_std_logic_vector(959874,20);
      WHEN "001100100" => data <= conv_std_logic_vector(959089,20);
      WHEN "001100101" => data <= conv_std_logic_vector(958307,20);
      WHEN "001100110" => data <= conv_std_logic_vector(957526,20);
      WHEN "001100111" => data <= conv_std_logic_vector(956747,20);
      WHEN "001101000" => data <= conv_std_logic_vector(955970,20);
      WHEN "001101001" => data <= conv_std_logic_vector(955195,20);
      WHEN "001101010" => data <= conv_std_logic_vector(954422,20);
      WHEN "001101011" => data <= conv_std_logic_vector(953651,20);
      WHEN "001101100" => data <= conv_std_logic_vector(952882,20);
      WHEN "001101101" => data <= conv_std_logic_vector(952114,20);
      WHEN "001101110" => data <= conv_std_logic_vector(951348,20);
      WHEN "001101111" => data <= conv_std_logic_vector(950585,20);
      WHEN "001110000" => data <= conv_std_logic_vector(949823,20);
      WHEN "001110001" => data <= conv_std_logic_vector(949062,20);
      WHEN "001110010" => data <= conv_std_logic_vector(948304,20);
      WHEN "001110011" => data <= conv_std_logic_vector(947548,20);
      WHEN "001110100" => data <= conv_std_logic_vector(946793,20);
      WHEN "001110101" => data <= conv_std_logic_vector(946040,20);
      WHEN "001110110" => data <= conv_std_logic_vector(945289,20);
      WHEN "001110111" => data <= conv_std_logic_vector(944539,20);
      WHEN "001111000" => data <= conv_std_logic_vector(943792,20);
      WHEN "001111001" => data <= conv_std_logic_vector(943046,20);
      WHEN "001111010" => data <= conv_std_logic_vector(942302,20);
      WHEN "001111011" => data <= conv_std_logic_vector(941560,20);
      WHEN "001111100" => data <= conv_std_logic_vector(940819,20);
      WHEN "001111101" => data <= conv_std_logic_vector(940081,20);
      WHEN "001111110" => data <= conv_std_logic_vector(939344,20);
      WHEN "001111111" => data <= conv_std_logic_vector(938608,20);
      WHEN "010000000" => data <= conv_std_logic_vector(937875,20);
      WHEN "010000001" => data <= conv_std_logic_vector(937143,20);
      WHEN "010000010" => data <= conv_std_logic_vector(936413,20);
      WHEN "010000011" => data <= conv_std_logic_vector(935684,20);
      WHEN "010000100" => data <= conv_std_logic_vector(934957,20);
      WHEN "010000101" => data <= conv_std_logic_vector(934232,20);
      WHEN "010000110" => data <= conv_std_logic_vector(933509,20);
      WHEN "010000111" => data <= conv_std_logic_vector(932787,20);
      WHEN "010001000" => data <= conv_std_logic_vector(932067,20);
      WHEN "010001001" => data <= conv_std_logic_vector(931349,20);
      WHEN "010001010" => data <= conv_std_logic_vector(930632,20);
      WHEN "010001011" => data <= conv_std_logic_vector(929917,20);
      WHEN "010001100" => data <= conv_std_logic_vector(929204,20);
      WHEN "010001101" => data <= conv_std_logic_vector(928492,20);
      WHEN "010001110" => data <= conv_std_logic_vector(927782,20);
      WHEN "010001111" => data <= conv_std_logic_vector(927073,20);
      WHEN "010010000" => data <= conv_std_logic_vector(926367,20);
      WHEN "010010001" => data <= conv_std_logic_vector(925661,20);
      WHEN "010010010" => data <= conv_std_logic_vector(924958,20);
      WHEN "010010011" => data <= conv_std_logic_vector(924256,20);
      WHEN "010010100" => data <= conv_std_logic_vector(923555,20);
      WHEN "010010101" => data <= conv_std_logic_vector(922856,20);
      WHEN "010010110" => data <= conv_std_logic_vector(922159,20);
      WHEN "010010111" => data <= conv_std_logic_vector(921463,20);
      WHEN "010011000" => data <= conv_std_logic_vector(920769,20);
      WHEN "010011001" => data <= conv_std_logic_vector(920077,20);
      WHEN "010011010" => data <= conv_std_logic_vector(919386,20);
      WHEN "010011011" => data <= conv_std_logic_vector(918696,20);
      WHEN "010011100" => data <= conv_std_logic_vector(918008,20);
      WHEN "010011101" => data <= conv_std_logic_vector(917322,20);
      WHEN "010011110" => data <= conv_std_logic_vector(916637,20);
      WHEN "010011111" => data <= conv_std_logic_vector(915954,20);
      WHEN "010100000" => data <= conv_std_logic_vector(915272,20);
      WHEN "010100001" => data <= conv_std_logic_vector(914592,20);
      WHEN "010100010" => data <= conv_std_logic_vector(913913,20);
      WHEN "010100011" => data <= conv_std_logic_vector(913236,20);
      WHEN "010100100" => data <= conv_std_logic_vector(912560,20);
      WHEN "010100101" => data <= conv_std_logic_vector(911886,20);
      WHEN "010100110" => data <= conv_std_logic_vector(911213,20);
      WHEN "010100111" => data <= conv_std_logic_vector(910542,20);
      WHEN "010101000" => data <= conv_std_logic_vector(909872,20);
      WHEN "010101001" => data <= conv_std_logic_vector(909204,20);
      WHEN "010101010" => data <= conv_std_logic_vector(908537,20);
      WHEN "010101011" => data <= conv_std_logic_vector(907872,20);
      WHEN "010101100" => data <= conv_std_logic_vector(907208,20);
      WHEN "010101101" => data <= conv_std_logic_vector(906545,20);
      WHEN "010101110" => data <= conv_std_logic_vector(905884,20);
      WHEN "010101111" => data <= conv_std_logic_vector(905225,20);
      WHEN "010110000" => data <= conv_std_logic_vector(904567,20);
      WHEN "010110001" => data <= conv_std_logic_vector(903910,20);
      WHEN "010110010" => data <= conv_std_logic_vector(903255,20);
      WHEN "010110011" => data <= conv_std_logic_vector(902601,20);
      WHEN "010110100" => data <= conv_std_logic_vector(901949,20);
      WHEN "010110101" => data <= conv_std_logic_vector(901298,20);
      WHEN "010110110" => data <= conv_std_logic_vector(900648,20);
      WHEN "010110111" => data <= conv_std_logic_vector(900000,20);
      WHEN "010111000" => data <= conv_std_logic_vector(899353,20);
      WHEN "010111001" => data <= conv_std_logic_vector(898708,20);
      WHEN "010111010" => data <= conv_std_logic_vector(898064,20);
      WHEN "010111011" => data <= conv_std_logic_vector(897421,20);
      WHEN "010111100" => data <= conv_std_logic_vector(896780,20);
      WHEN "010111101" => data <= conv_std_logic_vector(896140,20);
      WHEN "010111110" => data <= conv_std_logic_vector(895501,20);
      WHEN "010111111" => data <= conv_std_logic_vector(894864,20);
      WHEN "011000000" => data <= conv_std_logic_vector(894228,20);
      WHEN "011000001" => data <= conv_std_logic_vector(893594,20);
      WHEN "011000010" => data <= conv_std_logic_vector(892961,20);
      WHEN "011000011" => data <= conv_std_logic_vector(892329,20);
      WHEN "011000100" => data <= conv_std_logic_vector(891699,20);
      WHEN "011000101" => data <= conv_std_logic_vector(891070,20);
      WHEN "011000110" => data <= conv_std_logic_vector(890442,20);
      WHEN "011000111" => data <= conv_std_logic_vector(889816,20);
      WHEN "011001000" => data <= conv_std_logic_vector(889191,20);
      WHEN "011001001" => data <= conv_std_logic_vector(888567,20);
      WHEN "011001010" => data <= conv_std_logic_vector(887944,20);
      WHEN "011001011" => data <= conv_std_logic_vector(887323,20);
      WHEN "011001100" => data <= conv_std_logic_vector(886703,20);
      WHEN "011001101" => data <= conv_std_logic_vector(886085,20);
      WHEN "011001110" => data <= conv_std_logic_vector(885467,20);
      WHEN "011001111" => data <= conv_std_logic_vector(884851,20);
      WHEN "011010000" => data <= conv_std_logic_vector(884237,20);
      WHEN "011010001" => data <= conv_std_logic_vector(883623,20);
      WHEN "011010010" => data <= conv_std_logic_vector(883011,20);
      WHEN "011010011" => data <= conv_std_logic_vector(882400,20);
      WHEN "011010100" => data <= conv_std_logic_vector(881791,20);
      WHEN "011010101" => data <= conv_std_logic_vector(881182,20);
      WHEN "011010110" => data <= conv_std_logic_vector(880575,20);
      WHEN "011010111" => data <= conv_std_logic_vector(879969,20);
      WHEN "011011000" => data <= conv_std_logic_vector(879365,20);
      WHEN "011011001" => data <= conv_std_logic_vector(878762,20);
      WHEN "011011010" => data <= conv_std_logic_vector(878159,20);
      WHEN "011011011" => data <= conv_std_logic_vector(877559,20);
      WHEN "011011100" => data <= conv_std_logic_vector(876959,20);
      WHEN "011011101" => data <= conv_std_logic_vector(876361,20);
      WHEN "011011110" => data <= conv_std_logic_vector(875763,20);
      WHEN "011011111" => data <= conv_std_logic_vector(875167,20);
      WHEN "011100000" => data <= conv_std_logic_vector(874573,20);
      WHEN "011100001" => data <= conv_std_logic_vector(873979,20);
      WHEN "011100010" => data <= conv_std_logic_vector(873387,20);
      WHEN "011100011" => data <= conv_std_logic_vector(872796,20);
      WHEN "011100100" => data <= conv_std_logic_vector(872206,20);
      WHEN "011100101" => data <= conv_std_logic_vector(871617,20);
      WHEN "011100110" => data <= conv_std_logic_vector(871030,20);
      WHEN "011100111" => data <= conv_std_logic_vector(870443,20);
      WHEN "011101000" => data <= conv_std_logic_vector(869858,20);
      WHEN "011101001" => data <= conv_std_logic_vector(869274,20);
      WHEN "011101010" => data <= conv_std_logic_vector(868691,20);
      WHEN "011101011" => data <= conv_std_logic_vector(868110,20);
      WHEN "011101100" => data <= conv_std_logic_vector(867529,20);
      WHEN "011101101" => data <= conv_std_logic_vector(866950,20);
      WHEN "011101110" => data <= conv_std_logic_vector(866372,20);
      WHEN "011101111" => data <= conv_std_logic_vector(865795,20);
      WHEN "011110000" => data <= conv_std_logic_vector(865219,20);
      WHEN "011110001" => data <= conv_std_logic_vector(864644,20);
      WHEN "011110010" => data <= conv_std_logic_vector(864070,20);
      WHEN "011110011" => data <= conv_std_logic_vector(863498,20);
      WHEN "011110100" => data <= conv_std_logic_vector(862927,20);
      WHEN "011110101" => data <= conv_std_logic_vector(862357,20);
      WHEN "011110110" => data <= conv_std_logic_vector(861788,20);
      WHEN "011110111" => data <= conv_std_logic_vector(861220,20);
      WHEN "011111000" => data <= conv_std_logic_vector(860653,20);
      WHEN "011111001" => data <= conv_std_logic_vector(860087,20);
      WHEN "011111010" => data <= conv_std_logic_vector(859523,20);
      WHEN "011111011" => data <= conv_std_logic_vector(858959,20);
      WHEN "011111100" => data <= conv_std_logic_vector(858397,20);
      WHEN "011111101" => data <= conv_std_logic_vector(857836,20);
      WHEN "011111110" => data <= conv_std_logic_vector(857276,20);
      WHEN "011111111" => data <= conv_std_logic_vector(856717,20);
      WHEN "100000000" => data <= conv_std_logic_vector(856159,20);
      WHEN "100000001" => data <= conv_std_logic_vector(855602,20);
      WHEN "100000010" => data <= conv_std_logic_vector(855046,20);
      WHEN "100000011" => data <= conv_std_logic_vector(854491,20);
      WHEN "100000100" => data <= conv_std_logic_vector(853938,20);
      WHEN "100000101" => data <= conv_std_logic_vector(853385,20);
      WHEN "100000110" => data <= conv_std_logic_vector(852834,20);
      WHEN "100000111" => data <= conv_std_logic_vector(852283,20);
      WHEN "100001000" => data <= conv_std_logic_vector(851734,20);
      WHEN "100001001" => data <= conv_std_logic_vector(851186,20);
      WHEN "100001010" => data <= conv_std_logic_vector(850638,20);
      WHEN "100001011" => data <= conv_std_logic_vector(850092,20);
      WHEN "100001100" => data <= conv_std_logic_vector(849547,20);
      WHEN "100001101" => data <= conv_std_logic_vector(849003,20);
      WHEN "100001110" => data <= conv_std_logic_vector(848460,20);
      WHEN "100001111" => data <= conv_std_logic_vector(847918,20);
      WHEN "100010000" => data <= conv_std_logic_vector(847377,20);
      WHEN "100010001" => data <= conv_std_logic_vector(846837,20);
      WHEN "100010010" => data <= conv_std_logic_vector(846298,20);
      WHEN "100010011" => data <= conv_std_logic_vector(845761,20);
      WHEN "100010100" => data <= conv_std_logic_vector(845224,20);
      WHEN "100010101" => data <= conv_std_logic_vector(844688,20);
      WHEN "100010110" => data <= conv_std_logic_vector(844153,20);
      WHEN "100010111" => data <= conv_std_logic_vector(843619,20);
      WHEN "100011000" => data <= conv_std_logic_vector(843087,20);
      WHEN "100011001" => data <= conv_std_logic_vector(842555,20);
      WHEN "100011010" => data <= conv_std_logic_vector(842024,20);
      WHEN "100011011" => data <= conv_std_logic_vector(841494,20);
      WHEN "100011100" => data <= conv_std_logic_vector(840966,20);
      WHEN "100011101" => data <= conv_std_logic_vector(840438,20);
      WHEN "100011110" => data <= conv_std_logic_vector(839911,20);
      WHEN "100011111" => data <= conv_std_logic_vector(839385,20);
      WHEN "100100000" => data <= conv_std_logic_vector(838861,20);
      WHEN "100100001" => data <= conv_std_logic_vector(838337,20);
      WHEN "100100010" => data <= conv_std_logic_vector(837814,20);
      WHEN "100100011" => data <= conv_std_logic_vector(837292,20);
      WHEN "100100100" => data <= conv_std_logic_vector(836771,20);
      WHEN "100100101" => data <= conv_std_logic_vector(836251,20);
      WHEN "100100110" => data <= conv_std_logic_vector(835733,20);
      WHEN "100100111" => data <= conv_std_logic_vector(835215,20);
      WHEN "100101000" => data <= conv_std_logic_vector(834698,20);
      WHEN "100101001" => data <= conv_std_logic_vector(834182,20);
      WHEN "100101010" => data <= conv_std_logic_vector(833666,20);
      WHEN "100101011" => data <= conv_std_logic_vector(833152,20);
      WHEN "100101100" => data <= conv_std_logic_vector(832639,20);
      WHEN "100101101" => data <= conv_std_logic_vector(832127,20);
      WHEN "100101110" => data <= conv_std_logic_vector(831616,20);
      WHEN "100101111" => data <= conv_std_logic_vector(831105,20);
      WHEN "100110000" => data <= conv_std_logic_vector(830596,20);
      WHEN "100110001" => data <= conv_std_logic_vector(830087,20);
      WHEN "100110010" => data <= conv_std_logic_vector(829580,20);
      WHEN "100110011" => data <= conv_std_logic_vector(829073,20);
      WHEN "100110100" => data <= conv_std_logic_vector(828568,20);
      WHEN "100110101" => data <= conv_std_logic_vector(828063,20);
      WHEN "100110110" => data <= conv_std_logic_vector(827559,20);
      WHEN "100110111" => data <= conv_std_logic_vector(827056,20);
      WHEN "100111000" => data <= conv_std_logic_vector(826554,20);
      WHEN "100111001" => data <= conv_std_logic_vector(826053,20);
      WHEN "100111010" => data <= conv_std_logic_vector(825553,20);
      WHEN "100111011" => data <= conv_std_logic_vector(825053,20);
      WHEN "100111100" => data <= conv_std_logic_vector(824555,20);
      WHEN "100111101" => data <= conv_std_logic_vector(824058,20);
      WHEN "100111110" => data <= conv_std_logic_vector(823561,20);
      WHEN "100111111" => data <= conv_std_logic_vector(823065,20);
      WHEN "101000000" => data <= conv_std_logic_vector(822571,20);
      WHEN "101000001" => data <= conv_std_logic_vector(822077,20);
      WHEN "101000010" => data <= conv_std_logic_vector(821584,20);
      WHEN "101000011" => data <= conv_std_logic_vector(821092,20);
      WHEN "101000100" => data <= conv_std_logic_vector(820600,20);
      WHEN "101000101" => data <= conv_std_logic_vector(820110,20);
      WHEN "101000110" => data <= conv_std_logic_vector(819621,20);
      WHEN "101000111" => data <= conv_std_logic_vector(819132,20);
      WHEN "101001000" => data <= conv_std_logic_vector(818644,20);
      WHEN "101001001" => data <= conv_std_logic_vector(818157,20);
      WHEN "101001010" => data <= conv_std_logic_vector(817671,20);
      WHEN "101001011" => data <= conv_std_logic_vector(817186,20);
      WHEN "101001100" => data <= conv_std_logic_vector(816702,20);
      WHEN "101001101" => data <= conv_std_logic_vector(816219,20);
      WHEN "101001110" => data <= conv_std_logic_vector(815736,20);
      WHEN "101001111" => data <= conv_std_logic_vector(815254,20);
      WHEN "101010000" => data <= conv_std_logic_vector(814774,20);
      WHEN "101010001" => data <= conv_std_logic_vector(814294,20);
      WHEN "101010010" => data <= conv_std_logic_vector(813814,20);
      WHEN "101010011" => data <= conv_std_logic_vector(813336,20);
      WHEN "101010100" => data <= conv_std_logic_vector(812859,20);
      WHEN "101010101" => data <= conv_std_logic_vector(812382,20);
      WHEN "101010110" => data <= conv_std_logic_vector(811906,20);
      WHEN "101010111" => data <= conv_std_logic_vector(811431,20);
      WHEN "101011000" => data <= conv_std_logic_vector(810957,20);
      WHEN "101011001" => data <= conv_std_logic_vector(810484,20);
      WHEN "101011010" => data <= conv_std_logic_vector(810012,20);
      WHEN "101011011" => data <= conv_std_logic_vector(809540,20);
      WHEN "101011100" => data <= conv_std_logic_vector(809069,20);
      WHEN "101011101" => data <= conv_std_logic_vector(808599,20);
      WHEN "101011110" => data <= conv_std_logic_vector(808130,20);
      WHEN "101011111" => data <= conv_std_logic_vector(807662,20);
      WHEN "101100000" => data <= conv_std_logic_vector(807194,20);
      WHEN "101100001" => data <= conv_std_logic_vector(806727,20);
      WHEN "101100010" => data <= conv_std_logic_vector(806261,20);
      WHEN "101100011" => data <= conv_std_logic_vector(805796,20);
      WHEN "101100100" => data <= conv_std_logic_vector(805332,20);
      WHEN "101100101" => data <= conv_std_logic_vector(804869,20);
      WHEN "101100110" => data <= conv_std_logic_vector(804406,20);
      WHEN "101100111" => data <= conv_std_logic_vector(803944,20);
      WHEN "101101000" => data <= conv_std_logic_vector(803483,20);
      WHEN "101101001" => data <= conv_std_logic_vector(803023,20);
      WHEN "101101010" => data <= conv_std_logic_vector(802563,20);
      WHEN "101101011" => data <= conv_std_logic_vector(802104,20);
      WHEN "101101100" => data <= conv_std_logic_vector(801646,20);
      WHEN "101101101" => data <= conv_std_logic_vector(801189,20);
      WHEN "101101110" => data <= conv_std_logic_vector(800733,20);
      WHEN "101101111" => data <= conv_std_logic_vector(800277,20);
      WHEN "101110000" => data <= conv_std_logic_vector(799822,20);
      WHEN "101110001" => data <= conv_std_logic_vector(799368,20);
      WHEN "101110010" => data <= conv_std_logic_vector(798915,20);
      WHEN "101110011" => data <= conv_std_logic_vector(798462,20);
      WHEN "101110100" => data <= conv_std_logic_vector(798011,20);
      WHEN "101110101" => data <= conv_std_logic_vector(797560,20);
      WHEN "101110110" => data <= conv_std_logic_vector(797109,20);
      WHEN "101110111" => data <= conv_std_logic_vector(796660,20);
      WHEN "101111000" => data <= conv_std_logic_vector(796211,20);
      WHEN "101111001" => data <= conv_std_logic_vector(795763,20);
      WHEN "101111010" => data <= conv_std_logic_vector(795316,20);
      WHEN "101111011" => data <= conv_std_logic_vector(794870,20);
      WHEN "101111100" => data <= conv_std_logic_vector(794424,20);
      WHEN "101111101" => data <= conv_std_logic_vector(793979,20);
      WHEN "101111110" => data <= conv_std_logic_vector(793535,20);
      WHEN "101111111" => data <= conv_std_logic_vector(793092,20);
      WHEN "110000000" => data <= conv_std_logic_vector(792649,20);
      WHEN "110000001" => data <= conv_std_logic_vector(792207,20);
      WHEN "110000010" => data <= conv_std_logic_vector(791766,20);
      WHEN "110000011" => data <= conv_std_logic_vector(791325,20);
      WHEN "110000100" => data <= conv_std_logic_vector(790885,20);
      WHEN "110000101" => data <= conv_std_logic_vector(790446,20);
      WHEN "110000110" => data <= conv_std_logic_vector(790008,20);
      WHEN "110000111" => data <= conv_std_logic_vector(789571,20);
      WHEN "110001000" => data <= conv_std_logic_vector(789134,20);
      WHEN "110001001" => data <= conv_std_logic_vector(788698,20);
      WHEN "110001010" => data <= conv_std_logic_vector(788262,20);
      WHEN "110001011" => data <= conv_std_logic_vector(787828,20);
      WHEN "110001100" => data <= conv_std_logic_vector(787394,20);
      WHEN "110001101" => data <= conv_std_logic_vector(786960,20);
      WHEN "110001110" => data <= conv_std_logic_vector(786528,20);
      WHEN "110001111" => data <= conv_std_logic_vector(786096,20);
      WHEN "110010000" => data <= conv_std_logic_vector(785665,20);
      WHEN "110010001" => data <= conv_std_logic_vector(785235,20);
      WHEN "110010010" => data <= conv_std_logic_vector(784805,20);
      WHEN "110010011" => data <= conv_std_logic_vector(784376,20);
      WHEN "110010100" => data <= conv_std_logic_vector(783948,20);
      WHEN "110010101" => data <= conv_std_logic_vector(783520,20);
      WHEN "110010110" => data <= conv_std_logic_vector(783093,20);
      WHEN "110010111" => data <= conv_std_logic_vector(782667,20);
      WHEN "110011000" => data <= conv_std_logic_vector(782242,20);
      WHEN "110011001" => data <= conv_std_logic_vector(781817,20);
      WHEN "110011010" => data <= conv_std_logic_vector(781393,20);
      WHEN "110011011" => data <= conv_std_logic_vector(780969,20);
      WHEN "110011100" => data <= conv_std_logic_vector(780547,20);
      WHEN "110011101" => data <= conv_std_logic_vector(780125,20);
      WHEN "110011110" => data <= conv_std_logic_vector(779703,20);
      WHEN "110011111" => data <= conv_std_logic_vector(779283,20);
      WHEN "110100000" => data <= conv_std_logic_vector(778863,20);
      WHEN "110100001" => data <= conv_std_logic_vector(778443,20);
      WHEN "110100010" => data <= conv_std_logic_vector(778025,20);
      WHEN "110100011" => data <= conv_std_logic_vector(777607,20);
      WHEN "110100100" => data <= conv_std_logic_vector(777189,20);
      WHEN "110100101" => data <= conv_std_logic_vector(776773,20);
      WHEN "110100110" => data <= conv_std_logic_vector(776357,20);
      WHEN "110100111" => data <= conv_std_logic_vector(775942,20);
      WHEN "110101000" => data <= conv_std_logic_vector(775527,20);
      WHEN "110101001" => data <= conv_std_logic_vector(775113,20);
      WHEN "110101010" => data <= conv_std_logic_vector(774700,20);
      WHEN "110101011" => data <= conv_std_logic_vector(774287,20);
      WHEN "110101100" => data <= conv_std_logic_vector(773875,20);
      WHEN "110101101" => data <= conv_std_logic_vector(773464,20);
      WHEN "110101110" => data <= conv_std_logic_vector(773053,20);
      WHEN "110101111" => data <= conv_std_logic_vector(772643,20);
      WHEN "110110000" => data <= conv_std_logic_vector(772234,20);
      WHEN "110110001" => data <= conv_std_logic_vector(771825,20);
      WHEN "110110010" => data <= conv_std_logic_vector(771417,20);
      WHEN "110110011" => data <= conv_std_logic_vector(771010,20);
      WHEN "110110100" => data <= conv_std_logic_vector(770603,20);
      WHEN "110110101" => data <= conv_std_logic_vector(770197,20);
      WHEN "110110110" => data <= conv_std_logic_vector(769791,20);
      WHEN "110110111" => data <= conv_std_logic_vector(769387,20);
      WHEN "110111000" => data <= conv_std_logic_vector(768982,20);
      WHEN "110111001" => data <= conv_std_logic_vector(768579,20);
      WHEN "110111010" => data <= conv_std_logic_vector(768176,20);
      WHEN "110111011" => data <= conv_std_logic_vector(767774,20);
      WHEN "110111100" => data <= conv_std_logic_vector(767372,20);
      WHEN "110111101" => data <= conv_std_logic_vector(766971,20);
      WHEN "110111110" => data <= conv_std_logic_vector(766570,20);
      WHEN "110111111" => data <= conv_std_logic_vector(766171,20);
      WHEN "111000000" => data <= conv_std_logic_vector(765772,20);
      WHEN "111000001" => data <= conv_std_logic_vector(765373,20);
      WHEN "111000010" => data <= conv_std_logic_vector(764975,20);
      WHEN "111000011" => data <= conv_std_logic_vector(764578,20);
      WHEN "111000100" => data <= conv_std_logic_vector(764181,20);
      WHEN "111000101" => data <= conv_std_logic_vector(763785,20);
      WHEN "111000110" => data <= conv_std_logic_vector(763390,20);
      WHEN "111000111" => data <= conv_std_logic_vector(762995,20);
      WHEN "111001000" => data <= conv_std_logic_vector(762601,20);
      WHEN "111001001" => data <= conv_std_logic_vector(762207,20);
      WHEN "111001010" => data <= conv_std_logic_vector(761814,20);
      WHEN "111001011" => data <= conv_std_logic_vector(761422,20);
      WHEN "111001100" => data <= conv_std_logic_vector(761030,20);
      WHEN "111001101" => data <= conv_std_logic_vector(760639,20);
      WHEN "111001110" => data <= conv_std_logic_vector(760248,20);
      WHEN "111001111" => data <= conv_std_logic_vector(759858,20);
      WHEN "111010000" => data <= conv_std_logic_vector(759469,20);
      WHEN "111010001" => data <= conv_std_logic_vector(759080,20);
      WHEN "111010010" => data <= conv_std_logic_vector(758692,20);
      WHEN "111010011" => data <= conv_std_logic_vector(758304,20);
      WHEN "111010100" => data <= conv_std_logic_vector(757917,20);
      WHEN "111010101" => data <= conv_std_logic_vector(757531,20);
      WHEN "111010110" => data <= conv_std_logic_vector(757145,20);
      WHEN "111010111" => data <= conv_std_logic_vector(756760,20);
      WHEN "111011000" => data <= conv_std_logic_vector(756375,20);
      WHEN "111011001" => data <= conv_std_logic_vector(755991,20);
      WHEN "111011010" => data <= conv_std_logic_vector(755608,20);
      WHEN "111011011" => data <= conv_std_logic_vector(755225,20);
      WHEN "111011100" => data <= conv_std_logic_vector(754843,20);
      WHEN "111011101" => data <= conv_std_logic_vector(754461,20);
      WHEN "111011110" => data <= conv_std_logic_vector(754080,20);
      WHEN "111011111" => data <= conv_std_logic_vector(753699,20);
      WHEN "111100000" => data <= conv_std_logic_vector(753319,20);
      WHEN "111100001" => data <= conv_std_logic_vector(752940,20);
      WHEN "111100010" => data <= conv_std_logic_vector(752561,20);
      WHEN "111100011" => data <= conv_std_logic_vector(752183,20);
      WHEN "111100100" => data <= conv_std_logic_vector(751805,20);
      WHEN "111100101" => data <= conv_std_logic_vector(751428,20);
      WHEN "111100110" => data <= conv_std_logic_vector(751051,20);
      WHEN "111100111" => data <= conv_std_logic_vector(750675,20);
      WHEN "111101000" => data <= conv_std_logic_vector(750300,20);
      WHEN "111101001" => data <= conv_std_logic_vector(749925,20);
      WHEN "111101010" => data <= conv_std_logic_vector(749551,20);
      WHEN "111101011" => data <= conv_std_logic_vector(749177,20);
      WHEN "111101100" => data <= conv_std_logic_vector(748804,20);
      WHEN "111101101" => data <= conv_std_logic_vector(748431,20);
      WHEN "111101110" => data <= conv_std_logic_vector(748059,20);
      WHEN "111101111" => data <= conv_std_logic_vector(747687,20);
      WHEN "111110000" => data <= conv_std_logic_vector(747317,20);
      WHEN "111110001" => data <= conv_std_logic_vector(746946,20);
      WHEN "111110010" => data <= conv_std_logic_vector(746576,20);
      WHEN "111110011" => data <= conv_std_logic_vector(746207,20);
      WHEN "111110100" => data <= conv_std_logic_vector(745838,20);
      WHEN "111110101" => data <= conv_std_logic_vector(745470,20);
      WHEN "111110110" => data <= conv_std_logic_vector(745102,20);
      WHEN "111110111" => data <= conv_std_logic_vector(744735,20);
      WHEN "111111000" => data <= conv_std_logic_vector(744369,20);
      WHEN "111111001" => data <= conv_std_logic_vector(744002,20);
      WHEN "111111010" => data <= conv_std_logic_vector(743637,20);
      WHEN "111111011" => data <= conv_std_logic_vector(743272,20);
      WHEN "111111100" => data <= conv_std_logic_vector(742908,20);
      WHEN "111111101" => data <= conv_std_logic_vector(742544,20);
      WHEN "111111110" => data <= conv_std_logic_vector(742180,20);
      WHEN "111111111" => data <= conv_std_logic_vector(741817,20);
      WHEN others => data <= conv_std_logic_vector(0,20);
    END CASE;
  END PROCESS;

END rtl;
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_INVSQR_LUT1.VHD                        ***
--***                                             ***
--***   Function: Look Up Table - Inverse Root    ***
--***                                             ***
--***   Generated by MATLAB Utility               ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_invsqr_lut1 IS
PORT (
      add : IN STD_LOGIC_VECTOR (9 DOWNTO 1);
		data : OUT STD_LOGIC_VECTOR (11 DOWNTO 1)
);
END fp_invsqr_lut1;

ARCHITECTURE rtl OF fp_invsqr_lut1 IS

BEGIN

  pca: PROCESS (add)
  BEGIN
    CASE add IS
      WHEN "000000000" => data <= conv_std_logic_vector(1023,11);
      WHEN "000000001" => data <= conv_std_logic_vector(1020,11);
      WHEN "000000010" => data <= conv_std_logic_vector(1017,11);
      WHEN "000000011" => data <= conv_std_logic_vector(1014,11);
      WHEN "000000100" => data <= conv_std_logic_vector(1011,11);
      WHEN "000000101" => data <= conv_std_logic_vector(1008,11);
      WHEN "000000110" => data <= conv_std_logic_vector(1005,11);
      WHEN "000000111" => data <= conv_std_logic_vector(1002,11);
      WHEN "000001000" => data <= conv_std_logic_vector(999,11);
      WHEN "000001001" => data <= conv_std_logic_vector(996,11);
      WHEN "000001010" => data <= conv_std_logic_vector(993,11);
      WHEN "000001011" => data <= conv_std_logic_vector(990,11);
      WHEN "000001100" => data <= conv_std_logic_vector(988,11);
      WHEN "000001101" => data <= conv_std_logic_vector(985,11);
      WHEN "000001110" => data <= conv_std_logic_vector(982,11);
      WHEN "000001111" => data <= conv_std_logic_vector(979,11);
      WHEN "000010000" => data <= conv_std_logic_vector(976,11);
      WHEN "000010001" => data <= conv_std_logic_vector(974,11);
      WHEN "000010010" => data <= conv_std_logic_vector(971,11);
      WHEN "000010011" => data <= conv_std_logic_vector(968,11);
      WHEN "000010100" => data <= conv_std_logic_vector(965,11);
      WHEN "000010101" => data <= conv_std_logic_vector(963,11);
      WHEN "000010110" => data <= conv_std_logic_vector(960,11);
      WHEN "000010111" => data <= conv_std_logic_vector(957,11);
      WHEN "000011000" => data <= conv_std_logic_vector(955,11);
      WHEN "000011001" => data <= conv_std_logic_vector(952,11);
      WHEN "000011010" => data <= conv_std_logic_vector(949,11);
      WHEN "000011011" => data <= conv_std_logic_vector(947,11);
      WHEN "000011100" => data <= conv_std_logic_vector(944,11);
      WHEN "000011101" => data <= conv_std_logic_vector(941,11);
      WHEN "000011110" => data <= conv_std_logic_vector(939,11);
      WHEN "000011111" => data <= conv_std_logic_vector(936,11);
      WHEN "000100000" => data <= conv_std_logic_vector(934,11);
      WHEN "000100001" => data <= conv_std_logic_vector(931,11);
      WHEN "000100010" => data <= conv_std_logic_vector(929,11);
      WHEN "000100011" => data <= conv_std_logic_vector(926,11);
      WHEN "000100100" => data <= conv_std_logic_vector(924,11);
      WHEN "000100101" => data <= conv_std_logic_vector(921,11);
      WHEN "000100110" => data <= conv_std_logic_vector(918,11);
      WHEN "000100111" => data <= conv_std_logic_vector(916,11);
      WHEN "000101000" => data <= conv_std_logic_vector(913,11);
      WHEN "000101001" => data <= conv_std_logic_vector(911,11);
      WHEN "000101010" => data <= conv_std_logic_vector(909,11);
      WHEN "000101011" => data <= conv_std_logic_vector(906,11);
      WHEN "000101100" => data <= conv_std_logic_vector(904,11);
      WHEN "000101101" => data <= conv_std_logic_vector(901,11);
      WHEN "000101110" => data <= conv_std_logic_vector(899,11);
      WHEN "000101111" => data <= conv_std_logic_vector(896,11);
      WHEN "000110000" => data <= conv_std_logic_vector(894,11);
      WHEN "000110001" => data <= conv_std_logic_vector(892,11);
      WHEN "000110010" => data <= conv_std_logic_vector(889,11);
      WHEN "000110011" => data <= conv_std_logic_vector(887,11);
      WHEN "000110100" => data <= conv_std_logic_vector(885,11);
      WHEN "000110101" => data <= conv_std_logic_vector(882,11);
      WHEN "000110110" => data <= conv_std_logic_vector(880,11);
      WHEN "000110111" => data <= conv_std_logic_vector(878,11);
      WHEN "000111000" => data <= conv_std_logic_vector(875,11);
      WHEN "000111001" => data <= conv_std_logic_vector(873,11);
      WHEN "000111010" => data <= conv_std_logic_vector(871,11);
      WHEN "000111011" => data <= conv_std_logic_vector(868,11);
      WHEN "000111100" => data <= conv_std_logic_vector(866,11);
      WHEN "000111101" => data <= conv_std_logic_vector(864,11);
      WHEN "000111110" => data <= conv_std_logic_vector(862,11);
      WHEN "000111111" => data <= conv_std_logic_vector(859,11);
      WHEN "001000000" => data <= conv_std_logic_vector(857,11);
      WHEN "001000001" => data <= conv_std_logic_vector(855,11);
      WHEN "001000010" => data <= conv_std_logic_vector(853,11);
      WHEN "001000011" => data <= conv_std_logic_vector(850,11);
      WHEN "001000100" => data <= conv_std_logic_vector(848,11);
      WHEN "001000101" => data <= conv_std_logic_vector(846,11);
      WHEN "001000110" => data <= conv_std_logic_vector(844,11);
      WHEN "001000111" => data <= conv_std_logic_vector(842,11);
      WHEN "001001000" => data <= conv_std_logic_vector(840,11);
      WHEN "001001001" => data <= conv_std_logic_vector(837,11);
      WHEN "001001010" => data <= conv_std_logic_vector(835,11);
      WHEN "001001011" => data <= conv_std_logic_vector(833,11);
      WHEN "001001100" => data <= conv_std_logic_vector(831,11);
      WHEN "001001101" => data <= conv_std_logic_vector(829,11);
      WHEN "001001110" => data <= conv_std_logic_vector(827,11);
      WHEN "001001111" => data <= conv_std_logic_vector(825,11);
      WHEN "001010000" => data <= conv_std_logic_vector(823,11);
      WHEN "001010001" => data <= conv_std_logic_vector(820,11);
      WHEN "001010010" => data <= conv_std_logic_vector(818,11);
      WHEN "001010011" => data <= conv_std_logic_vector(816,11);
      WHEN "001010100" => data <= conv_std_logic_vector(814,11);
      WHEN "001010101" => data <= conv_std_logic_vector(812,11);
      WHEN "001010110" => data <= conv_std_logic_vector(810,11);
      WHEN "001010111" => data <= conv_std_logic_vector(808,11);
      WHEN "001011000" => data <= conv_std_logic_vector(806,11);
      WHEN "001011001" => data <= conv_std_logic_vector(804,11);
      WHEN "001011010" => data <= conv_std_logic_vector(802,11);
      WHEN "001011011" => data <= conv_std_logic_vector(800,11);
      WHEN "001011100" => data <= conv_std_logic_vector(798,11);
      WHEN "001011101" => data <= conv_std_logic_vector(796,11);
      WHEN "001011110" => data <= conv_std_logic_vector(794,11);
      WHEN "001011111" => data <= conv_std_logic_vector(792,11);
      WHEN "001100000" => data <= conv_std_logic_vector(790,11);
      WHEN "001100001" => data <= conv_std_logic_vector(788,11);
      WHEN "001100010" => data <= conv_std_logic_vector(786,11);
      WHEN "001100011" => data <= conv_std_logic_vector(785,11);
      WHEN "001100100" => data <= conv_std_logic_vector(783,11);
      WHEN "001100101" => data <= conv_std_logic_vector(781,11);
      WHEN "001100110" => data <= conv_std_logic_vector(779,11);
      WHEN "001100111" => data <= conv_std_logic_vector(777,11);
      WHEN "001101000" => data <= conv_std_logic_vector(775,11);
      WHEN "001101001" => data <= conv_std_logic_vector(773,11);
      WHEN "001101010" => data <= conv_std_logic_vector(771,11);
      WHEN "001101011" => data <= conv_std_logic_vector(769,11);
      WHEN "001101100" => data <= conv_std_logic_vector(768,11);
      WHEN "001101101" => data <= conv_std_logic_vector(766,11);
      WHEN "001101110" => data <= conv_std_logic_vector(764,11);
      WHEN "001101111" => data <= conv_std_logic_vector(762,11);
      WHEN "001110000" => data <= conv_std_logic_vector(760,11);
      WHEN "001110001" => data <= conv_std_logic_vector(758,11);
      WHEN "001110010" => data <= conv_std_logic_vector(757,11);
      WHEN "001110011" => data <= conv_std_logic_vector(755,11);
      WHEN "001110100" => data <= conv_std_logic_vector(753,11);
      WHEN "001110101" => data <= conv_std_logic_vector(751,11);
      WHEN "001110110" => data <= conv_std_logic_vector(749,11);
      WHEN "001110111" => data <= conv_std_logic_vector(748,11);
      WHEN "001111000" => data <= conv_std_logic_vector(746,11);
      WHEN "001111001" => data <= conv_std_logic_vector(744,11);
      WHEN "001111010" => data <= conv_std_logic_vector(742,11);
      WHEN "001111011" => data <= conv_std_logic_vector(741,11);
      WHEN "001111100" => data <= conv_std_logic_vector(739,11);
      WHEN "001111101" => data <= conv_std_logic_vector(737,11);
      WHEN "001111110" => data <= conv_std_logic_vector(735,11);
      WHEN "001111111" => data <= conv_std_logic_vector(734,11);
      WHEN "010000000" => data <= conv_std_logic_vector(732,11);
      WHEN "010000001" => data <= conv_std_logic_vector(730,11);
      WHEN "010000010" => data <= conv_std_logic_vector(728,11);
      WHEN "010000011" => data <= conv_std_logic_vector(727,11);
      WHEN "010000100" => data <= conv_std_logic_vector(725,11);
      WHEN "010000101" => data <= conv_std_logic_vector(723,11);
      WHEN "010000110" => data <= conv_std_logic_vector(722,11);
      WHEN "010000111" => data <= conv_std_logic_vector(720,11);
      WHEN "010001000" => data <= conv_std_logic_vector(718,11);
      WHEN "010001001" => data <= conv_std_logic_vector(717,11);
      WHEN "010001010" => data <= conv_std_logic_vector(715,11);
      WHEN "010001011" => data <= conv_std_logic_vector(713,11);
      WHEN "010001100" => data <= conv_std_logic_vector(712,11);
      WHEN "010001101" => data <= conv_std_logic_vector(710,11);
      WHEN "010001110" => data <= conv_std_logic_vector(709,11);
      WHEN "010001111" => data <= conv_std_logic_vector(707,11);
      WHEN "010010000" => data <= conv_std_logic_vector(705,11);
      WHEN "010010001" => data <= conv_std_logic_vector(704,11);
      WHEN "010010010" => data <= conv_std_logic_vector(702,11);
      WHEN "010010011" => data <= conv_std_logic_vector(700,11);
      WHEN "010010100" => data <= conv_std_logic_vector(699,11);
      WHEN "010010101" => data <= conv_std_logic_vector(697,11);
      WHEN "010010110" => data <= conv_std_logic_vector(696,11);
      WHEN "010010111" => data <= conv_std_logic_vector(694,11);
      WHEN "010011000" => data <= conv_std_logic_vector(693,11);
      WHEN "010011001" => data <= conv_std_logic_vector(691,11);
      WHEN "010011010" => data <= conv_std_logic_vector(689,11);
      WHEN "010011011" => data <= conv_std_logic_vector(688,11);
      WHEN "010011100" => data <= conv_std_logic_vector(686,11);
      WHEN "010011101" => data <= conv_std_logic_vector(685,11);
      WHEN "010011110" => data <= conv_std_logic_vector(683,11);
      WHEN "010011111" => data <= conv_std_logic_vector(682,11);
      WHEN "010100000" => data <= conv_std_logic_vector(680,11);
      WHEN "010100001" => data <= conv_std_logic_vector(679,11);
      WHEN "010100010" => data <= conv_std_logic_vector(677,11);
      WHEN "010100011" => data <= conv_std_logic_vector(676,11);
      WHEN "010100100" => data <= conv_std_logic_vector(674,11);
      WHEN "010100101" => data <= conv_std_logic_vector(673,11);
      WHEN "010100110" => data <= conv_std_logic_vector(671,11);
      WHEN "010100111" => data <= conv_std_logic_vector(670,11);
      WHEN "010101000" => data <= conv_std_logic_vector(668,11);
      WHEN "010101001" => data <= conv_std_logic_vector(667,11);
      WHEN "010101010" => data <= conv_std_logic_vector(665,11);
      WHEN "010101011" => data <= conv_std_logic_vector(664,11);
      WHEN "010101100" => data <= conv_std_logic_vector(662,11);
      WHEN "010101101" => data <= conv_std_logic_vector(661,11);
      WHEN "010101110" => data <= conv_std_logic_vector(660,11);
      WHEN "010101111" => data <= conv_std_logic_vector(658,11);
      WHEN "010110000" => data <= conv_std_logic_vector(657,11);
      WHEN "010110001" => data <= conv_std_logic_vector(655,11);
      WHEN "010110010" => data <= conv_std_logic_vector(654,11);
      WHEN "010110011" => data <= conv_std_logic_vector(652,11);
      WHEN "010110100" => data <= conv_std_logic_vector(651,11);
      WHEN "010110101" => data <= conv_std_logic_vector(650,11);
      WHEN "010110110" => data <= conv_std_logic_vector(648,11);
      WHEN "010110111" => data <= conv_std_logic_vector(647,11);
      WHEN "010111000" => data <= conv_std_logic_vector(645,11);
      WHEN "010111001" => data <= conv_std_logic_vector(644,11);
      WHEN "010111010" => data <= conv_std_logic_vector(643,11);
      WHEN "010111011" => data <= conv_std_logic_vector(641,11);
      WHEN "010111100" => data <= conv_std_logic_vector(640,11);
      WHEN "010111101" => data <= conv_std_logic_vector(639,11);
      WHEN "010111110" => data <= conv_std_logic_vector(637,11);
      WHEN "010111111" => data <= conv_std_logic_vector(636,11);
      WHEN "011000000" => data <= conv_std_logic_vector(634,11);
      WHEN "011000001" => data <= conv_std_logic_vector(633,11);
      WHEN "011000010" => data <= conv_std_logic_vector(632,11);
      WHEN "011000011" => data <= conv_std_logic_vector(630,11);
      WHEN "011000100" => data <= conv_std_logic_vector(629,11);
      WHEN "011000101" => data <= conv_std_logic_vector(628,11);
      WHEN "011000110" => data <= conv_std_logic_vector(626,11);
      WHEN "011000111" => data <= conv_std_logic_vector(625,11);
      WHEN "011001000" => data <= conv_std_logic_vector(624,11);
      WHEN "011001001" => data <= conv_std_logic_vector(622,11);
      WHEN "011001010" => data <= conv_std_logic_vector(621,11);
      WHEN "011001011" => data <= conv_std_logic_vector(620,11);
      WHEN "011001100" => data <= conv_std_logic_vector(619,11);
      WHEN "011001101" => data <= conv_std_logic_vector(617,11);
      WHEN "011001110" => data <= conv_std_logic_vector(616,11);
      WHEN "011001111" => data <= conv_std_logic_vector(615,11);
      WHEN "011010000" => data <= conv_std_logic_vector(613,11);
      WHEN "011010001" => data <= conv_std_logic_vector(612,11);
      WHEN "011010010" => data <= conv_std_logic_vector(611,11);
      WHEN "011010011" => data <= conv_std_logic_vector(610,11);
      WHEN "011010100" => data <= conv_std_logic_vector(608,11);
      WHEN "011010101" => data <= conv_std_logic_vector(607,11);
      WHEN "011010110" => data <= conv_std_logic_vector(606,11);
      WHEN "011010111" => data <= conv_std_logic_vector(605,11);
      WHEN "011011000" => data <= conv_std_logic_vector(603,11);
      WHEN "011011001" => data <= conv_std_logic_vector(602,11);
      WHEN "011011010" => data <= conv_std_logic_vector(601,11);
      WHEN "011011011" => data <= conv_std_logic_vector(600,11);
      WHEN "011011100" => data <= conv_std_logic_vector(598,11);
      WHEN "011011101" => data <= conv_std_logic_vector(597,11);
      WHEN "011011110" => data <= conv_std_logic_vector(596,11);
      WHEN "011011111" => data <= conv_std_logic_vector(595,11);
      WHEN "011100000" => data <= conv_std_logic_vector(594,11);
      WHEN "011100001" => data <= conv_std_logic_vector(592,11);
      WHEN "011100010" => data <= conv_std_logic_vector(591,11);
      WHEN "011100011" => data <= conv_std_logic_vector(590,11);
      WHEN "011100100" => data <= conv_std_logic_vector(589,11);
      WHEN "011100101" => data <= conv_std_logic_vector(588,11);
      WHEN "011100110" => data <= conv_std_logic_vector(586,11);
      WHEN "011100111" => data <= conv_std_logic_vector(585,11);
      WHEN "011101000" => data <= conv_std_logic_vector(584,11);
      WHEN "011101001" => data <= conv_std_logic_vector(583,11);
      WHEN "011101010" => data <= conv_std_logic_vector(582,11);
      WHEN "011101011" => data <= conv_std_logic_vector(580,11);
      WHEN "011101100" => data <= conv_std_logic_vector(579,11);
      WHEN "011101101" => data <= conv_std_logic_vector(578,11);
      WHEN "011101110" => data <= conv_std_logic_vector(577,11);
      WHEN "011101111" => data <= conv_std_logic_vector(576,11);
      WHEN "011110000" => data <= conv_std_logic_vector(575,11);
      WHEN "011110001" => data <= conv_std_logic_vector(574,11);
      WHEN "011110010" => data <= conv_std_logic_vector(572,11);
      WHEN "011110011" => data <= conv_std_logic_vector(571,11);
      WHEN "011110100" => data <= conv_std_logic_vector(570,11);
      WHEN "011110101" => data <= conv_std_logic_vector(569,11);
      WHEN "011110110" => data <= conv_std_logic_vector(568,11);
      WHEN "011110111" => data <= conv_std_logic_vector(567,11);
      WHEN "011111000" => data <= conv_std_logic_vector(566,11);
      WHEN "011111001" => data <= conv_std_logic_vector(565,11);
      WHEN "011111010" => data <= conv_std_logic_vector(563,11);
      WHEN "011111011" => data <= conv_std_logic_vector(562,11);
      WHEN "011111100" => data <= conv_std_logic_vector(561,11);
      WHEN "011111101" => data <= conv_std_logic_vector(560,11);
      WHEN "011111110" => data <= conv_std_logic_vector(559,11);
      WHEN "011111111" => data <= conv_std_logic_vector(558,11);
      WHEN "100000000" => data <= conv_std_logic_vector(557,11);
      WHEN "100000001" => data <= conv_std_logic_vector(556,11);
      WHEN "100000010" => data <= conv_std_logic_vector(555,11);
      WHEN "100000011" => data <= conv_std_logic_vector(554,11);
      WHEN "100000100" => data <= conv_std_logic_vector(553,11);
      WHEN "100000101" => data <= conv_std_logic_vector(551,11);
      WHEN "100000110" => data <= conv_std_logic_vector(550,11);
      WHEN "100000111" => data <= conv_std_logic_vector(549,11);
      WHEN "100001000" => data <= conv_std_logic_vector(548,11);
      WHEN "100001001" => data <= conv_std_logic_vector(547,11);
      WHEN "100001010" => data <= conv_std_logic_vector(546,11);
      WHEN "100001011" => data <= conv_std_logic_vector(545,11);
      WHEN "100001100" => data <= conv_std_logic_vector(544,11);
      WHEN "100001101" => data <= conv_std_logic_vector(543,11);
      WHEN "100001110" => data <= conv_std_logic_vector(542,11);
      WHEN "100001111" => data <= conv_std_logic_vector(541,11);
      WHEN "100010000" => data <= conv_std_logic_vector(540,11);
      WHEN "100010001" => data <= conv_std_logic_vector(539,11);
      WHEN "100010010" => data <= conv_std_logic_vector(538,11);
      WHEN "100010011" => data <= conv_std_logic_vector(537,11);
      WHEN "100010100" => data <= conv_std_logic_vector(536,11);
      WHEN "100010101" => data <= conv_std_logic_vector(535,11);
      WHEN "100010110" => data <= conv_std_logic_vector(534,11);
      WHEN "100010111" => data <= conv_std_logic_vector(533,11);
      WHEN "100011000" => data <= conv_std_logic_vector(532,11);
      WHEN "100011001" => data <= conv_std_logic_vector(531,11);
      WHEN "100011010" => data <= conv_std_logic_vector(530,11);
      WHEN "100011011" => data <= conv_std_logic_vector(529,11);
      WHEN "100011100" => data <= conv_std_logic_vector(528,11);
      WHEN "100011101" => data <= conv_std_logic_vector(527,11);
      WHEN "100011110" => data <= conv_std_logic_vector(526,11);
      WHEN "100011111" => data <= conv_std_logic_vector(525,11);
      WHEN "100100000" => data <= conv_std_logic_vector(524,11);
      WHEN "100100001" => data <= conv_std_logic_vector(523,11);
      WHEN "100100010" => data <= conv_std_logic_vector(522,11);
      WHEN "100100011" => data <= conv_std_logic_vector(521,11);
      WHEN "100100100" => data <= conv_std_logic_vector(520,11);
      WHEN "100100101" => data <= conv_std_logic_vector(519,11);
      WHEN "100100110" => data <= conv_std_logic_vector(518,11);
      WHEN "100100111" => data <= conv_std_logic_vector(517,11);
      WHEN "100101000" => data <= conv_std_logic_vector(516,11);
      WHEN "100101001" => data <= conv_std_logic_vector(515,11);
      WHEN "100101010" => data <= conv_std_logic_vector(514,11);
      WHEN "100101011" => data <= conv_std_logic_vector(513,11);
      WHEN "100101100" => data <= conv_std_logic_vector(512,11);
      WHEN "100101101" => data <= conv_std_logic_vector(511,11);
      WHEN "100101110" => data <= conv_std_logic_vector(510,11);
      WHEN "100101111" => data <= conv_std_logic_vector(509,11);
      WHEN "100110000" => data <= conv_std_logic_vector(508,11);
      WHEN "100110001" => data <= conv_std_logic_vector(508,11);
      WHEN "100110010" => data <= conv_std_logic_vector(507,11);
      WHEN "100110011" => data <= conv_std_logic_vector(506,11);
      WHEN "100110100" => data <= conv_std_logic_vector(505,11);
      WHEN "100110101" => data <= conv_std_logic_vector(504,11);
      WHEN "100110110" => data <= conv_std_logic_vector(503,11);
      WHEN "100110111" => data <= conv_std_logic_vector(502,11);
      WHEN "100111000" => data <= conv_std_logic_vector(501,11);
      WHEN "100111001" => data <= conv_std_logic_vector(500,11);
      WHEN "100111010" => data <= conv_std_logic_vector(499,11);
      WHEN "100111011" => data <= conv_std_logic_vector(498,11);
      WHEN "100111100" => data <= conv_std_logic_vector(497,11);
      WHEN "100111101" => data <= conv_std_logic_vector(497,11);
      WHEN "100111110" => data <= conv_std_logic_vector(496,11);
      WHEN "100111111" => data <= conv_std_logic_vector(495,11);
      WHEN "101000000" => data <= conv_std_logic_vector(494,11);
      WHEN "101000001" => data <= conv_std_logic_vector(493,11);
      WHEN "101000010" => data <= conv_std_logic_vector(492,11);
      WHEN "101000011" => data <= conv_std_logic_vector(491,11);
      WHEN "101000100" => data <= conv_std_logic_vector(490,11);
      WHEN "101000101" => data <= conv_std_logic_vector(489,11);
      WHEN "101000110" => data <= conv_std_logic_vector(489,11);
      WHEN "101000111" => data <= conv_std_logic_vector(488,11);
      WHEN "101001000" => data <= conv_std_logic_vector(487,11);
      WHEN "101001001" => data <= conv_std_logic_vector(486,11);
      WHEN "101001010" => data <= conv_std_logic_vector(485,11);
      WHEN "101001011" => data <= conv_std_logic_vector(484,11);
      WHEN "101001100" => data <= conv_std_logic_vector(483,11);
      WHEN "101001101" => data <= conv_std_logic_vector(483,11);
      WHEN "101001110" => data <= conv_std_logic_vector(482,11);
      WHEN "101001111" => data <= conv_std_logic_vector(481,11);
      WHEN "101010000" => data <= conv_std_logic_vector(480,11);
      WHEN "101010001" => data <= conv_std_logic_vector(479,11);
      WHEN "101010010" => data <= conv_std_logic_vector(478,11);
      WHEN "101010011" => data <= conv_std_logic_vector(477,11);
      WHEN "101010100" => data <= conv_std_logic_vector(477,11);
      WHEN "101010101" => data <= conv_std_logic_vector(476,11);
      WHEN "101010110" => data <= conv_std_logic_vector(475,11);
      WHEN "101010111" => data <= conv_std_logic_vector(474,11);
      WHEN "101011000" => data <= conv_std_logic_vector(473,11);
      WHEN "101011001" => data <= conv_std_logic_vector(472,11);
      WHEN "101011010" => data <= conv_std_logic_vector(472,11);
      WHEN "101011011" => data <= conv_std_logic_vector(471,11);
      WHEN "101011100" => data <= conv_std_logic_vector(470,11);
      WHEN "101011101" => data <= conv_std_logic_vector(469,11);
      WHEN "101011110" => data <= conv_std_logic_vector(468,11);
      WHEN "101011111" => data <= conv_std_logic_vector(468,11);
      WHEN "101100000" => data <= conv_std_logic_vector(467,11);
      WHEN "101100001" => data <= conv_std_logic_vector(466,11);
      WHEN "101100010" => data <= conv_std_logic_vector(465,11);
      WHEN "101100011" => data <= conv_std_logic_vector(464,11);
      WHEN "101100100" => data <= conv_std_logic_vector(464,11);
      WHEN "101100101" => data <= conv_std_logic_vector(463,11);
      WHEN "101100110" => data <= conv_std_logic_vector(462,11);
      WHEN "101100111" => data <= conv_std_logic_vector(461,11);
      WHEN "101101000" => data <= conv_std_logic_vector(460,11);
      WHEN "101101001" => data <= conv_std_logic_vector(460,11);
      WHEN "101101010" => data <= conv_std_logic_vector(459,11);
      WHEN "101101011" => data <= conv_std_logic_vector(458,11);
      WHEN "101101100" => data <= conv_std_logic_vector(457,11);
      WHEN "101101101" => data <= conv_std_logic_vector(456,11);
      WHEN "101101110" => data <= conv_std_logic_vector(456,11);
      WHEN "101101111" => data <= conv_std_logic_vector(455,11);
      WHEN "101110000" => data <= conv_std_logic_vector(454,11);
      WHEN "101110001" => data <= conv_std_logic_vector(453,11);
      WHEN "101110010" => data <= conv_std_logic_vector(453,11);
      WHEN "101110011" => data <= conv_std_logic_vector(452,11);
      WHEN "101110100" => data <= conv_std_logic_vector(451,11);
      WHEN "101110101" => data <= conv_std_logic_vector(450,11);
      WHEN "101110110" => data <= conv_std_logic_vector(449,11);
      WHEN "101110111" => data <= conv_std_logic_vector(449,11);
      WHEN "101111000" => data <= conv_std_logic_vector(448,11);
      WHEN "101111001" => data <= conv_std_logic_vector(447,11);
      WHEN "101111010" => data <= conv_std_logic_vector(446,11);
      WHEN "101111011" => data <= conv_std_logic_vector(446,11);
      WHEN "101111100" => data <= conv_std_logic_vector(445,11);
      WHEN "101111101" => data <= conv_std_logic_vector(444,11);
      WHEN "101111110" => data <= conv_std_logic_vector(443,11);
      WHEN "101111111" => data <= conv_std_logic_vector(443,11);
      WHEN "110000000" => data <= conv_std_logic_vector(442,11);
      WHEN "110000001" => data <= conv_std_logic_vector(441,11);
      WHEN "110000010" => data <= conv_std_logic_vector(440,11);
      WHEN "110000011" => data <= conv_std_logic_vector(440,11);
      WHEN "110000100" => data <= conv_std_logic_vector(439,11);
      WHEN "110000101" => data <= conv_std_logic_vector(438,11);
      WHEN "110000110" => data <= conv_std_logic_vector(438,11);
      WHEN "110000111" => data <= conv_std_logic_vector(437,11);
      WHEN "110001000" => data <= conv_std_logic_vector(436,11);
      WHEN "110001001" => data <= conv_std_logic_vector(435,11);
      WHEN "110001010" => data <= conv_std_logic_vector(435,11);
      WHEN "110001011" => data <= conv_std_logic_vector(434,11);
      WHEN "110001100" => data <= conv_std_logic_vector(433,11);
      WHEN "110001101" => data <= conv_std_logic_vector(433,11);
      WHEN "110001110" => data <= conv_std_logic_vector(432,11);
      WHEN "110001111" => data <= conv_std_logic_vector(431,11);
      WHEN "110010000" => data <= conv_std_logic_vector(430,11);
      WHEN "110010001" => data <= conv_std_logic_vector(430,11);
      WHEN "110010010" => data <= conv_std_logic_vector(429,11);
      WHEN "110010011" => data <= conv_std_logic_vector(428,11);
      WHEN "110010100" => data <= conv_std_logic_vector(428,11);
      WHEN "110010101" => data <= conv_std_logic_vector(427,11);
      WHEN "110010110" => data <= conv_std_logic_vector(426,11);
      WHEN "110010111" => data <= conv_std_logic_vector(425,11);
      WHEN "110011000" => data <= conv_std_logic_vector(425,11);
      WHEN "110011001" => data <= conv_std_logic_vector(424,11);
      WHEN "110011010" => data <= conv_std_logic_vector(423,11);
      WHEN "110011011" => data <= conv_std_logic_vector(423,11);
      WHEN "110011100" => data <= conv_std_logic_vector(422,11);
      WHEN "110011101" => data <= conv_std_logic_vector(421,11);
      WHEN "110011110" => data <= conv_std_logic_vector(421,11);
      WHEN "110011111" => data <= conv_std_logic_vector(420,11);
      WHEN "110100000" => data <= conv_std_logic_vector(419,11);
      WHEN "110100001" => data <= conv_std_logic_vector(419,11);
      WHEN "110100010" => data <= conv_std_logic_vector(418,11);
      WHEN "110100011" => data <= conv_std_logic_vector(417,11);
      WHEN "110100100" => data <= conv_std_logic_vector(417,11);
      WHEN "110100101" => data <= conv_std_logic_vector(416,11);
      WHEN "110100110" => data <= conv_std_logic_vector(415,11);
      WHEN "110100111" => data <= conv_std_logic_vector(415,11);
      WHEN "110101000" => data <= conv_std_logic_vector(414,11);
      WHEN "110101001" => data <= conv_std_logic_vector(413,11);
      WHEN "110101010" => data <= conv_std_logic_vector(413,11);
      WHEN "110101011" => data <= conv_std_logic_vector(412,11);
      WHEN "110101100" => data <= conv_std_logic_vector(411,11);
      WHEN "110101101" => data <= conv_std_logic_vector(411,11);
      WHEN "110101110" => data <= conv_std_logic_vector(410,11);
      WHEN "110101111" => data <= conv_std_logic_vector(409,11);
      WHEN "110110000" => data <= conv_std_logic_vector(409,11);
      WHEN "110110001" => data <= conv_std_logic_vector(408,11);
      WHEN "110110010" => data <= conv_std_logic_vector(407,11);
      WHEN "110110011" => data <= conv_std_logic_vector(407,11);
      WHEN "110110100" => data <= conv_std_logic_vector(406,11);
      WHEN "110110101" => data <= conv_std_logic_vector(405,11);
      WHEN "110110110" => data <= conv_std_logic_vector(405,11);
      WHEN "110110111" => data <= conv_std_logic_vector(404,11);
      WHEN "110111000" => data <= conv_std_logic_vector(404,11);
      WHEN "110111001" => data <= conv_std_logic_vector(403,11);
      WHEN "110111010" => data <= conv_std_logic_vector(402,11);
      WHEN "110111011" => data <= conv_std_logic_vector(402,11);
      WHEN "110111100" => data <= conv_std_logic_vector(401,11);
      WHEN "110111101" => data <= conv_std_logic_vector(400,11);
      WHEN "110111110" => data <= conv_std_logic_vector(400,11);
      WHEN "110111111" => data <= conv_std_logic_vector(399,11);
      WHEN "111000000" => data <= conv_std_logic_vector(399,11);
      WHEN "111000001" => data <= conv_std_logic_vector(398,11);
      WHEN "111000010" => data <= conv_std_logic_vector(397,11);
      WHEN "111000011" => data <= conv_std_logic_vector(397,11);
      WHEN "111000100" => data <= conv_std_logic_vector(396,11);
      WHEN "111000101" => data <= conv_std_logic_vector(395,11);
      WHEN "111000110" => data <= conv_std_logic_vector(395,11);
      WHEN "111000111" => data <= conv_std_logic_vector(394,11);
      WHEN "111001000" => data <= conv_std_logic_vector(394,11);
      WHEN "111001001" => data <= conv_std_logic_vector(393,11);
      WHEN "111001010" => data <= conv_std_logic_vector(392,11);
      WHEN "111001011" => data <= conv_std_logic_vector(392,11);
      WHEN "111001100" => data <= conv_std_logic_vector(391,11);
      WHEN "111001101" => data <= conv_std_logic_vector(391,11);
      WHEN "111001110" => data <= conv_std_logic_vector(390,11);
      WHEN "111001111" => data <= conv_std_logic_vector(389,11);
      WHEN "111010000" => data <= conv_std_logic_vector(389,11);
      WHEN "111010001" => data <= conv_std_logic_vector(388,11);
      WHEN "111010010" => data <= conv_std_logic_vector(388,11);
      WHEN "111010011" => data <= conv_std_logic_vector(387,11);
      WHEN "111010100" => data <= conv_std_logic_vector(386,11);
      WHEN "111010101" => data <= conv_std_logic_vector(386,11);
      WHEN "111010110" => data <= conv_std_logic_vector(385,11);
      WHEN "111010111" => data <= conv_std_logic_vector(385,11);
      WHEN "111011000" => data <= conv_std_logic_vector(384,11);
      WHEN "111011001" => data <= conv_std_logic_vector(383,11);
      WHEN "111011010" => data <= conv_std_logic_vector(383,11);
      WHEN "111011011" => data <= conv_std_logic_vector(382,11);
      WHEN "111011100" => data <= conv_std_logic_vector(382,11);
      WHEN "111011101" => data <= conv_std_logic_vector(381,11);
      WHEN "111011110" => data <= conv_std_logic_vector(381,11);
      WHEN "111011111" => data <= conv_std_logic_vector(380,11);
      WHEN "111100000" => data <= conv_std_logic_vector(379,11);
      WHEN "111100001" => data <= conv_std_logic_vector(379,11);
      WHEN "111100010" => data <= conv_std_logic_vector(378,11);
      WHEN "111100011" => data <= conv_std_logic_vector(378,11);
      WHEN "111100100" => data <= conv_std_logic_vector(377,11);
      WHEN "111100101" => data <= conv_std_logic_vector(377,11);
      WHEN "111100110" => data <= conv_std_logic_vector(376,11);
      WHEN "111100111" => data <= conv_std_logic_vector(375,11);
      WHEN "111101000" => data <= conv_std_logic_vector(375,11);
      WHEN "111101001" => data <= conv_std_logic_vector(374,11);
      WHEN "111101010" => data <= conv_std_logic_vector(374,11);
      WHEN "111101011" => data <= conv_std_logic_vector(373,11);
      WHEN "111101100" => data <= conv_std_logic_vector(373,11);
      WHEN "111101101" => data <= conv_std_logic_vector(372,11);
      WHEN "111101110" => data <= conv_std_logic_vector(372,11);
      WHEN "111101111" => data <= conv_std_logic_vector(371,11);
      WHEN "111110000" => data <= conv_std_logic_vector(370,11);
      WHEN "111110001" => data <= conv_std_logic_vector(370,11);
      WHEN "111110010" => data <= conv_std_logic_vector(369,11);
      WHEN "111110011" => data <= conv_std_logic_vector(369,11);
      WHEN "111110100" => data <= conv_std_logic_vector(368,11);
      WHEN "111110101" => data <= conv_std_logic_vector(368,11);
      WHEN "111110110" => data <= conv_std_logic_vector(367,11);
      WHEN "111110111" => data <= conv_std_logic_vector(367,11);
      WHEN "111111000" => data <= conv_std_logic_vector(366,11);
      WHEN "111111001" => data <= conv_std_logic_vector(366,11);
      WHEN "111111010" => data <= conv_std_logic_vector(365,11);
      WHEN "111111011" => data <= conv_std_logic_vector(364,11);
      WHEN "111111100" => data <= conv_std_logic_vector(364,11);
      WHEN "111111101" => data <= conv_std_logic_vector(363,11);
      WHEN "111111110" => data <= conv_std_logic_vector(363,11);
      WHEN "111111111" => data <= conv_std_logic_vector(362,11);
      WHEN others => data <= conv_std_logic_vector(0,11);
    END CASE;
  END PROCESS;

END rtl;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

-- for 36 bit mantissa for trig library

--***************************************************
--*** Notes: Latency = 17                         ***
--***************************************************

ENTITY fp_invsqr_trig1 IS 
GENERIC (synthesize : integer := 1); 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      exponentin: IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (36 DOWNTO 1);

      exponentout : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
		);
END fp_invsqr_trig1;

ARCHITECTURE rtl OF fp_invsqr_trig1 IS
  
  constant manwidth : positive := 36;
  constant expwidth : positive := 8;
  
  constant coredepth : positive := 17;
  
  type expfftype IS ARRAY (coredepth DOWNTO 1) OF STD_LOGIC_VECTOR (expwidth DOWNTO 1);

  signal expff : expfftype;
  signal radicand : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal oddexponent : STD_LOGIC;
  signal invroot : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal zerovec : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal offset : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
   
  component fp_invsqr_core IS 
  GENERIC (synthesize : integer := 1); -- 0/1 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        radicand : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
        odd : IN STD_LOGIC;

		  invroot : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
		  );
  end component;
	
BEGIN
    
  gzva: FOR k IN 1 TO manwidth GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  gxoa: FOR k IN 1 TO expwidth-1 GENERATE
    offset(k) <= '1';
  END GENERATE;
  offset(expwidth) <= '0';

  pma: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN

      FOR k IN 1 TO coredepth LOOP
        FOR j IN 1 TO expwidth LOOP
          expff(k)(j) <= '0';
        END LOOP;
      END LOOP;
  
    ELSIF (rising_edge(sysclk)) THEN
  
      expff(1)(expwidth DOWNTO 1) <= exponentin;
      expff(2)(expwidth DOWNTO 1) <= expff(1)(expwidth DOWNTO 1) - offset;
      expff(3)(expwidth DOWNTO 1) <= expff(2)(expwidth) & expff(2)(expwidth DOWNTO 2);
      expff(4)(expwidth DOWNTO 1) <= offset - expff(3)(expwidth DOWNTO 1);
      expff(5)(expwidth DOWNTO 1) <= expff(4)(expwidth DOWNTO 1) - 1;
      FOR k IN 6 TO coredepth LOOP
        expff(k)(expwidth DOWNTO 1) <= expff(k-1)(expwidth DOWNTO 1);
      END LOOP;
  
    END IF;
  
  END PROCESS;

--*******************
--*** SQUARE ROOT ***
--*******************

  radicand <= mantissain; -- already with leading '1'
  -- sub 127, so 127 (odd) = 2^0 => even
  oddexponent <= NOT(exponentin(1));

  -- does not require rounding, output of core rounded already, LSB always 0
  isqr: fp_invsqr_core
  GENERIC MAP (synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            radicand=>radicand,odd=>oddexponent,
            invroot=>invroot);
       
--***************
--*** OUTPUTS ***
--***************

  exponentout <= expff(coredepth)(expwidth DOWNTO 1);   
  mantissaout <= invroot;  

END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   ALTERA FLOATING POINT DATAPATH COMPILER   ***
--***                                             ***
--***   FP_LDEXP.VHD                              ***
--***                                             ***
--***   Function: Single Precision Load Exponent  ***
--***                                             ***
--***   ldexp(x,n) - x*2^n - IEEE in and out      ***
--***                                             ***
--***   Created 11/09/09                          ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_ldexp IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (23 DOWNTO 1);
      bb : IN STD_LOGIC_VECTOR (32 DOWNTO 1);
      
		  signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
		  satout, zeroout, nanout : OUT STD_LOGIC
		);
END fp_ldexp;

ARCHITECTURE rtl OF fp_ldexp IS
 
  signal signinff : STD_LOGIC;
  signal exponentinff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal mantissainff : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal bbff : STD_LOGIC_VECTOR (10 DOWNTO 1);
  signal signoutff : STD_LOGIC;
  signal exponentoutff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal mantissaoutff : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal satoutff, zerooutff, nanoutff : STD_LOGIC;
  signal satnode, zeronode, nannode : STD_LOGIC;
  signal expnode : STD_LOGIC_VECTOR (10 DOWNTO 1);
  signal expzeroin, expmaxin : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal expzeronode, expmaxnode : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal expzeroout, expmaxout : STD_LOGIC;
  signal manzeroin : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal manzero, mannonzero : STD_LOGIC; 

BEGIN
    
  pin: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
    
      signinff <= '0';
      signoutff <= '0';
      FOR k IN 1 TO 8 LOOP
        exponentinff(k) <= '0';
        exponentoutff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 23 LOOP
        mantissainff(k) <= '0';
        mantissaoutff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 10 LOOP
        bbff(k) <= '0';
      END LOOP;
      satoutff <= '0';
      zerooutff <= '0';
      nanoutff <= '0';
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF (enable = '1') THEN

      
        signinff <= signin;
        exponentinff <= exponentin;
        mantissainff <= mantissain;
        
        bbff <= bb(10 DOWNTO 1);
        
        signoutff <= signinff;
        FOR k IN 1 TO 8 LOOP
          exponentoutff(k) <= (expnode(k) AND NOT(zeronode)) OR satnode OR nannode;
        END LOOP;
        FOR k IN 1 TO 23 LOOP
          mantissaoutff(k) <= (mantissainff(k) AND NOT(zeronode) AND NOT(satnode)) OR nannode;
        END LOOP;
        
        satoutff <= satnode;
        zerooutff <= zeronode;
        nanoutff <= nannode;
        
      END IF;
    
    END IF;  
      
  END PROCESS;
  
  expnode <= ("00" & exponentinff) + bbff;
  
  expzeroin(1) <= exponentinff(1);
  expmaxin(1) <= exponentinff(1);
  gxa: FOR k IN 2 TO 8 GENERATE
    expzeroin(k) <= expzeroin(k-1) OR exponentinff(k);
    expmaxin(k) <= expmaxin(k-1) AND exponentinff(k);
  END GENERATE;
  
  expzeronode(1) <= expnode(1);
  expmaxnode(1) <= expnode(1);
  gxb: FOR k IN 2 TO 8 GENERATE
    expzeronode(k) <= expzeronode(k-1) OR expnode(k);
    expmaxnode(k) <= expmaxnode(k-1) AND expnode(k);
  END GENERATE;
  expzeroout <= NOT(expzeroin(8)) OR (NOT(expzeronode(8)) AND NOT(expnode(9))) OR (expnode(10));
  expmaxout <= expmaxin(8) OR (expmaxnode(8) AND NOT(expnode(9))) OR (expnode(9) AND NOT(expnode(10))); 
  
  manzeroin(1) <= mantissainff(1);
  gma: FOR k IN 2 TO 23 GENERATE
    manzeroin(k) <= manzeroin(k-1) OR mantissainff(k);
  END GENERATE;
  manzero <= NOT(manzeroin(23));
  mannonzero <= manzeroin(23);
  
  satnode <= (expmaxin(8) AND NOT(manzeroin(23))) OR expmaxout;
  zeronode <= NOT(expzeroin(8)) OR expzeroout;
  nannode <= expmaxin(8) AND manzeroin(23);
  
	signout <= signoutff;
  exponentout <= exponentoutff;
  mantissaout <= mantissaoutff;
      
  satout <= satoutff;
  zeroout <= zerooutff;
  nanout <= nanoutff;

END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   SINGLE PRECISION LOG(e) - CORE            ***
--***                                             ***
--***   FP_LN_CORE.VHD                            ***
--***                                             ***
--***   Function: Single Precision LOG (LN) Core  ***
--***                                             ***
--***   22/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** Latency = 19                                ***
--***************************************************

ENTITY fp_ln_core IS 
GENERIC (synthesize : integer := 0);
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      aaman : IN STD_LOGIC_VECTOR (23 DOWNTO 1); 
      aaexp : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      
      ccman : OUT STD_LOGIC_VECTOR (24 DOWNTO 1);
      ccexp : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
      ccsgn : OUT STD_LOGIC;
      zeroout : OUT STD_LOGIC
     );
END fp_ln_core;

ARCHITECTURE rtl OF fp_ln_core IS
    
  signal zerovec : STD_LOGIC_VECTOR (32 DOWNTO 1);
  -- input
  signal aamanff : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal aaexpff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal aaexppos, aaexpneg : STD_LOGIC_VECTOR (9 DOWNTO 1);
  signal aaexpabs, aaexpabsff : STD_LOGIC_VECTOR (7 DOWNTO 1);
  -- range reduction
  signal lutpowaddff : STD_LOGIC_VECTOR (7 DOWNTO 1);
  signal lutoneaddff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal lutpowmanff, lutonemanff : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal lutpowexpff, lutoneexpff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal lutoneinvff : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal lutpowmannode, lutonemannode : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal lutpowexpnode, lutoneexpnode : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal lutoneinvnode : STD_LOGIC_VECTOR (11 DOWNTO 1); 
  signal aanum, aanumdel : STD_LOGIC_VECTOR (24 DOWNTO 1);
  signal mulonenode : STD_LOGIC_VECTOR (35 DOWNTO 1);
  signal mulonenormff : STD_LOGIC_VECTOR (34 DOWNTO 1);    
  -- series
  signal squared : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal cubed : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal scaled : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal onethird : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal mulonedel : STD_LOGIC_VECTOR (26 DOWNTO 1);
  signal oneterm, twoterm, thrterm : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal seriesoneff, seriesonedelff, seriestwoff : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal numtwo : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal exptwo : STD_LOGIC_VECTOR (8 DOWNTO 1);
  -- addition
  signal zeroone, zeropow : STD_LOGIC;
  signal numberone, numberonedel : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal numpow, numone : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal numpowsigned : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal exppow, expone : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal numpowone, numpowonedel : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal exppowone, exppowonedel : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal numsum : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal numsumabs : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal expsum : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal ccmannode : STD_LOGIC_VECTOR (24 DOWNTO 1);
  signal ccexpnode : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal signff : STD_LOGIC_VECTOR (18 DOWNTO 1);      

  component fp_lnlutpow
  PORT (
        add : IN STD_LOGIC_VECTOR (7 DOWNTO 1);
        logman : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
        logexp : OUT STD_LOGIC_VECTOR (8 DOWNTO 1)
       );
  end component;
  
  component fp_lnlut8 
  PORT (
        add : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
        inv : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
        logman : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
        logexp : OUT STD_LOGIC_VECTOR (8 DOWNTO 1)
       );
  end component;

  component fp_del
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
  end component;
  
  component fp_fxmul
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36;
           pipes : positive := 1;
           accuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1); 
      
        result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
       );
  end component;
  
  component fp_lnadd
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aaman : IN STD_LOGIC_VECTOR (32 DOWNTO 1);
        aaexp : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
        bbman : IN STD_LOGIC_VECTOR (32 DOWNTO 1);
        bbexp : IN STD_LOGIC_VECTOR (8 DOWNTO 1);

	     ccman : OUT STD_LOGIC_VECTOR (32 DOWNTO 1);
	     ccexp : OUT STD_LOGIC_VECTOR (8 DOWNTO 1)
	   );
  end component;
  
  component fp_lnnorm
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        inman : IN STD_LOGIC_VECTOR (32 DOWNTO 1);
        inexp : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
        outman : OUT STD_LOGIC_VECTOR (24 DOWNTO 1);
        outexp : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
        zero : OUT STD_LOGIC
       );
  end component;     
                 
BEGIN
  
  gza: FOR k IN 1 TO 32 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  --*******************
  --*** INPUT BLOCK ***
  --*******************
  
  ppin: PROCESS (sysclk,reset)
  BEGIN
  
    IF (reset = '1') THEN
        
      FOR k IN 1 TO 23 LOOP
        aamanff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 8 LOOP
        aaexpff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 7 LOOP
        aaexpabsff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
     
      IF (enable = '1') THEN       
      
        aamanff <= aaman;  -- level 1
        aaexpff <= aaexp;  -- level 1
      
        aaexpabsff <= aaexpabs;  -- level 2
      
      END IF;
 
    END IF;
    
  END PROCESS;
  
  aaexppos <= ('0' & aaexpff) - "001111111";
  aaexpneg <= "001111111" - ('0' & aaexpff);
  gaba: FOR k IN 1 TO 7 GENERATE
    aaexpabs(k) <= (aaexppos(k) AND NOT(aaexppos(9))) OR (aaexpneg(k) AND aaexppos(9));
  END GENERATE;
  
  --******************************************
  --*** RANGE REDUCTION THROUGH LUT SERIES ***
  --******************************************
    
  plut: PROCESS (sysclk,reset)
  BEGIN
  
    IF (reset = '1') THEN
       
      FOR k IN 1 TO 7 LOOP 
        lutpowaddff(k) <= '0'; 
      END LOOP;
      FOR k IN 1 TO 8 LOOP
        lutoneaddff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 23 LOOP
        lutpowmanff(k) <= '0';
        lutonemanff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 8 LOOP
        lutpowexpff(k) <= '0';
        lutoneexpff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 11 LOOP
        lutoneinvff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
            
      IF (enable = '1') THEN
          
        lutpowaddff <= aaexpabsff;  -- level 3
        lutoneaddff <= aamanff(23 DOWNTO 16);  -- level 2
   
        lutpowmanff <= lutpowmannode;  -- level 4
        lutpowexpff <= lutpowexpnode; -- level 4
      
        lutoneinvff <= lutoneinvnode;  -- level 3
        lutonemanff <= lutonemannode;  -- level 3
        lutoneexpff <= lutoneexpnode; -- level 3
      
      END IF;
      
    END IF;
    
  END PROCESS;
  
  lutpow: fp_lnlutpow
  PORT MAP (add=>lutpowaddff,
            logman=>lutpowmannode,logexp=>lutpowexpnode);
              
  lutone: fp_lnlut8
  PORT MAP (add=>lutoneaddff,
            inv=>lutoneinvnode,logman=>lutonemannode,logexp=>lutoneexpnode);
  
  aanum <= '1' & aamanff;
  
  -- level 1 in, level 3 out
  delone: fp_del
  GENERIC MAP (width=>24,pipes=>2)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>aanum,cc=>aanumdel);
            
  --mulone <= aanum * invone; -- 24*11 = 35
  
  -- level 3 in, level 6 out
  mulone: fp_fxmul
  GENERIC MAP (widthaa=>24,widthbb=>11,widthcc=>35,
               pipes=>3,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>aanumdel,databb=>lutoneinvff,
            result=>mulonenode);

  pmna: PROCESS (sysclk,reset)
  BEGIN
  
    IF (reset = '1') THEN
        
      FOR k IN 1 TO 34 LOOP
        mulonenormff(k) <= '0';
      END LOOP;
   
    ELSIF (rising_edge(sysclk)) THEN
     
      IF (enable = '1') THEN
        
        -- normalize in case input is 1.000000 and inv is 0.5  
        -- level 7
        FOR k IN 1 TO 34 LOOP
          mulonenormff(k) <= (mulonenode(k+1) AND mulonenode(35)) OR 
                             (mulonenode(k) AND NOT(mulonenode(35)));
        END LOOP;
         
      END IF;       
    END IF;
    
  END PROCESS;
  
  --***********************************************************
  --*** taylor series expansion of subrange (15 bits)       ***
  --*** x - x*x/2                                           ***
  --*** 7 leading bits, so x*x 7 bits down, +1 bit for 1/2  ***
  --***********************************************************
  
  --square <= mulonenorm(25 DOWNTO 8) * mulonenorm(25 DOWNTO 8);
  --cubed <= square(36 DOWNTO 19) * mulonenorm(25 DOWNTO 8);
  --cubedscale <= cubed(36 DOWNTO 19) * onethird;
  
  onethird <= "010101010101010101";
  
  -- level 7 in, level 9 out
  multwo: fp_fxmul
  GENERIC MAP (widthaa=>18,widthbb=>18,widthcc=>36,
               pipes=>2,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>mulonenormff(26 DOWNTO 9),databb=>mulonenormff(26 DOWNTO 9),
            result=>squared);
            
  -- level 7 in, level 9 out
  multhr: fp_fxmul
  GENERIC MAP (widthaa=>18,widthbb=>18,widthcc=>36,
               pipes=>2,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>mulonenormff(26 DOWNTO 9),databb=>onethird,
            result=>scaled); 
            
  -- level 9 in, level 11 out
  mulfor: fp_fxmul
  GENERIC MAP (widthaa=>18,widthbb=>18,widthcc=>36,
               pipes=>2,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>squared(36 DOWNTO 19),databb=>scaled(36 DOWNTO 19),
            result=>cubed);
                               
  oneterm <= mulonenormff(26 DOWNTO 1) & zerovec(6 DOWNTO 1);
  twoterm <= zerovec(7 DOWNTO 1) & squared(36 DOWNTO 12);
  thrterm <= zerovec(14 DOWNTO 1) & cubed(36 DOWNTO 19);
  
  --numtwo <= '0' & ((mulonenorm(25 DOWNTO 1) & zerovec(6 DOWNTO 1)) -
  --                 (zerovec(9 DOWNTO 1) & square(36 DOWNTO 15)) +
  --                 (zerovec(16 DOWNTO 1) & cubedscale(36 DOWNTO 22)));
  
  -- level 7 in, level 9 out
  deltwo: fp_del
  GENERIC MAP (width=>26,pipes=>2)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>mulonenormff(26 DOWNTO 1),cc=>mulonedel);
            
  ptay: PROCESS (sysclk,reset)
  BEGIN
  
    IF (reset = '1') THEN
        
      FOR k IN 1 TO 32 LOOP
        seriesoneff(k) <= '0';
        seriesonedelff(k) <= '0';
        seriestwoff(k) <= '0';
      END LOOP;
   
    ELSIF (rising_edge(sysclk)) THEN
     
      IF (enable = '1') THEN
        
        -- level 10
        seriesoneff <= (mulonedel & zerovec(6 DOWNTO 1)) -
                       (zerovec(8 DOWNTO 1) & squared(36 DOWNTO 13));
        seriesonedelff <= seriesoneff;
        -- level 12          
        seriestwoff <= seriesonedelff + (zerovec(14 DOWNTO 1) & cubed(36 DOWNTO 19));
         
      END IF;       

    END IF;
    
  END PROCESS;
            
  numtwo <= '0' & seriestwoff(32 DOWNTO 2);
  -- exponent for subrange 127-8 = 119              
  exptwo <= "01110111";
  
  --***********************************************************
  --*** add logarithm values                                ***
  --***********************************************************
  
  zeroone <= lutoneexpff(8) OR lutoneexpff(7) OR lutoneexpff(6) OR lutoneexpff(5) OR 
             lutoneexpff(4) OR lutoneexpff(3) OR lutoneexpff(2) OR lutoneexpff(1);
             
  numberone <= zeroone & lutonemanff & lutoneexpff;
  
  -- level 3 in, level 4 out
  delthr: fp_del
  GENERIC MAP (width=>32,pipes=>1)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>numberone,cc=>numberonedel);
    
  numone <= '0' & numberonedel(32 DOWNTO 9) & zerovec(7 DOWNTO 1);
  expone <= numberonedel(8 DOWNTO 1);
          
  zeropow <= lutpowexpff(8) OR lutpowexpff(7) OR lutpowexpff(6) OR lutpowexpff(5) OR 
             lutpowexpff(4) OR lutpowexpff(3) OR lutpowexpff(2) OR lutpowexpff(1);
 
  numpow <= '0' & zeropow & lutpowmanff & zerovec(7 DOWNTO 1);
  exppow <= lutpowexpff;

  gmpz: FOR k IN 1 TO 32 GENERATE
    numpowsigned(k) <= numpow(k) XOR signff(3);
  END GENERATE;
  
  -- level 4 in, level 8 out
  addone: fp_lnadd
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aaman=>numpowsigned,aaexp=>exppow,
            bbman=>numone,bbexp=>expone,
            ccman=>numpowone,ccexp=>exppowone);
  
  -- level 8 in, level 12 out
  delfor: fp_del
  GENERIC MAP (width=>32,pipes=>4)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>numpowone,cc=>numpowonedel);
  delfiv: fp_del
  GENERIC MAP (width=>8,pipes=>4)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>exppowone,cc=>exppowonedel);
             
  -- level 12 in, level 16 out         
  addtwo: fp_lnadd
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aaman=>numpowonedel,aaexp=>exppowonedel,
            bbman=>numtwo,bbexp=>exptwo,
            ccman=>numsum,ccexp=>expsum);          
  
  gmsa: FOR k IN 1 TO 32 GENERATE
    numsumabs(k) <= numsum(k) XOR signff(15);
  END GENERATE;
  
  -- level 16 in, level 19 out
  norm: fp_lnnorm
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            inman=>numsumabs,inexp=>expsum,
            outman=>ccmannode,outexp=>ccexpnode,
            zero=>zeroout);
  
  psgna: PROCESS (sysclk)
  BEGIN
      
    IF (reset = '1') THEN
      FOR k IN 1 TO 18 LOOP
        signff(k) <= '0';
      END LOOP;
    ELSIF (rising_edge(sysclk)) THEN
      signff(1) <= aaexppos(9);
      FOR k IN 2 TO 18 LOOP
        signff(k) <= signff(k-1);
      END LOOP;    
    END IF;
    
  END PROCESS;
      
  ccsgn <= signff(18);
  ccman <= ccmannode;
  ccexp <= ccexpnode;
          
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_LNADD.VHD                              ***
--***                                             ***
--***   Function: Single Precision Addition of    ***
--***   LN elements                               ***
--***                                             ***
--***   22/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** Latency = 4                                 ***
--***************************************************

ENTITY fp_lnadd IS 
GENERIC (
         speed : integer := 1; -- '0' for unpiped adder, '1' for piped adder
         synthesize : integer := 1
        ); 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      aaman : IN STD_LOGIC_VECTOR (32 DOWNTO 1);
      aaexp : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      bbman : IN STD_LOGIC_VECTOR (32 DOWNTO 1);
      bbexp : IN STD_LOGIC_VECTOR (8 DOWNTO 1);

	   ccman : OUT STD_LOGIC_VECTOR (32 DOWNTO 1);
	   ccexp : OUT STD_LOGIC_VECTOR (8 DOWNTO 1)
	 );
END fp_lnadd;

ARCHITECTURE rtl OF fp_lnadd IS
  
  type expbasefftype IS ARRAY (3 DOWNTO 1) OF STD_LOGIC_VECTOR (8 DOWNTO 1);
  
  signal aamanff, bbmanff : STD_LOGIC_VECTOR (32 DOWNTO 1); 
  signal aaexpff, bbexpff : STD_LOGIC_VECTOR (8 DOWNTO 1);  
  signal manleftff, manrightff : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal aluleftff, alurightff : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal expbaseff : expbasefftype;
  signal shiftff : STD_LOGIC_VECTOR (5 DOWNTO 1);
  signal subexpone, subexptwo : STD_LOGIC_VECTOR (9 DOWNTO 1);
  signal switch : STD_LOGIC;
  signal shiftleftnode, shiftrightnode : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal aluff : STD_LOGIC_VECTOR (32 DOWNTO 1);
  
  component fp_rsft32x5 IS 
  PORT (
        inbus : IN STD_LOGIC_VECTOR (32 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (5 DOWNTO 1);
        outbus : OUT STD_LOGIC_VECTOR (32 DOWNTO 1)
      );
  end component;
     
BEGIN
     
  paa: PROCESS (sysclk, reset)
  BEGIN
      
    IF (reset = '1') THEN
       
      FOR k IN 1 TO 32 LOOP 
        aamanff(k) <= '0';
        bbmanff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 8 LOOP 
        aaexpff(k) <= '0';
        bbexpff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 32 LOOP
        manleftff(k) <= '0';
        manrightff(k) <= '0';
        aluleftff(k) <= '0';
        alurightff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 8 LOOP
        FOR j IN 1 TO 3 LOOP
          expbaseff(j)(k) <= '0';
        END LOOP;
      END LOOP;
      shiftff <= "00000";
        
    ELSIF (rising_edge(sysclk)) THEN
            
      IF (enable = '1') THEN
          
        --*** LEVEL 1 ***
        aamanff <= aaman;
        bbmanff <= bbman;
        aaexpff <= aaexp;
        bbexpff <= bbexp;
        
        --*** LEVEL 2 ***
        FOR k IN 1 TO 32 LOOP
          manleftff(k) <= (aamanff(k) AND NOT(switch)) OR (bbmanff(k) AND switch);
          manrightff(k) <= (bbmanff(k) AND NOT(switch)) OR (aamanff(k) AND switch);
        END LOOP;
          
        FOR k IN 1 TO 8 LOOP
          expbaseff(1)(k) <= (aaexpff(k) AND NOT(switch)) OR (bbexpff(k) AND switch); 
        END LOOP;
        FOR k IN 2 TO 3 LOOP
          expbaseff(k)(8 DOWNTO 1) <= expbaseff(k-1)(8 DOWNTO 1);  -- level 3 to 4
        END LOOP;
        
        FOR k IN 1 TO 5 LOOP
          shiftff(k) <= (subexpone(k) AND NOT(switch)) OR (subexptwo(k) AND switch);
        END LOOP;
        
        --*** LEVEL 3 ***
        aluleftff <= shiftleftnode;
        alurightff <= shiftrightnode;
        
        --*** LEVEL 4 ***
        aluff <= aluleftff + alurightff;
      
      END IF;
        
    END IF;
      
  END PROCESS;
  
  subexpone <= ('0' & aaexpff) - ('0' & bbexpff);
  subexptwo <= ('0' & bbexpff) - ('0' & aaexpff);

  switch <= subexpone(9);

  shifter: fp_rsft32x5
  PORT MAP (inbus=>manrightff,shift=>shiftff,
            outbus=>shiftrightnode);
              
  shiftleftnode <= manleftff;

  --*** OUTPUTS ***
  ccman <= aluff;
  ccexp <= expbaseff(3)(8 DOWNTO 1);

END rtl;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_LNCLZ.VHD                              ***
--***                                             ***
--***   Function: Single Precision CLZ            ***
--***                                             ***
--***   22/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_lnclz IS
PORT (
      mantissa : IN STD_LOGIC_VECTOR (32 DOWNTO 1);
      
      leading : OUT STD_LOGIC_VECTOR (5 DOWNTO 1)    
     );
END fp_lnclz;

ARCHITECTURE rtl of fp_lnclz IS

  type positiontype IS ARRAY (6 DOWNTO 1) OF STD_LOGIC_VECTOR (5 DOWNTO 1);
  
  signal position, positionmux : positiontype;
  signal zerogroup, firstzero : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal lastman : STD_LOGIC_VECTOR (6 DOWNTO 1);
  
  component fp_pos
  GENERIC (start: integer := 0);
  PORT 
       (
        ingroup : IN STD_LOGIC_VECTOR (6 DOWNTO 1); 
        
        position : OUT STD_LOGIC_VECTOR (5 DOWNTO 1)    
       );
  end component;
  
BEGIN
     
  zerogroup(1) <= mantissa(32) OR mantissa(31) OR mantissa(30) OR mantissa(29) OR mantissa(28) OR mantissa(27);
  zerogroup(2) <= mantissa(26) OR mantissa(25) OR mantissa(24) OR mantissa(23) OR mantissa(22) OR mantissa(21);
  zerogroup(3) <= mantissa(20) OR mantissa(19) OR mantissa(18) OR mantissa(17) OR mantissa(16) OR mantissa(15);
  zerogroup(4) <= mantissa(14) OR mantissa(13) OR mantissa(12) OR mantissa(11) OR mantissa(10) OR mantissa(9);
  zerogroup(5) <= mantissa(8) OR mantissa(7) OR mantissa(6) OR mantissa(5) OR mantissa(4) OR mantissa(3);
  zerogroup(6) <= mantissa(2) OR mantissa(1);

  pa: fp_pos 
  GENERIC MAP (start=>0) 
  PORT MAP (ingroup=>mantissa(32 DOWNTO 27),position=>position(1)(5 DOWNTO 1));
  pb: fp_pos 
  GENERIC MAP (start=>6) 
  PORT MAP (ingroup=>mantissa(26 DOWNTO 21),position=>position(2)(5 DOWNTO 1));
  pc: fp_pos 
  GENERIC MAP (start=>12) 
  PORT MAP (ingroup=>mantissa(20 DOWNTO 15),position=>position(3)(5 DOWNTO 1));
  pd: fp_pos 
  GENERIC MAP (start=>18) 
  PORT MAP (ingroup=>mantissa(14 DOWNTO 9),position=>position(4)(5 DOWNTO 1));
  pe: fp_pos 
  GENERIC MAP (start=>24) 
  PORT MAP (ingroup=>mantissa(8 DOWNTO 3),position=>position(5)(5 DOWNTO 1));
  pf: fp_pos 
  GENERIC MAP (start=>30) 
  PORT MAP (ingroup=>lastman,position=>position(6)(5 DOWNTO 1));
      
  lastman <= mantissa(2 DOWNTO 1) & "0000";

  firstzero(1) <= zerogroup(1);
  firstzero(2) <= NOT(zerogroup(1)) AND zerogroup(2);
  firstzero(3) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND zerogroup(3);
  firstzero(4) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND zerogroup(4);
  firstzero(5) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND NOT(zerogroup(4)) 
                  AND zerogroup(5);
  firstzero(6) <= NOT(zerogroup(1)) AND NOT(zerogroup(2)) AND NOT(zerogroup(3)) AND NOT(zerogroup(4)) 
                  AND NOT(zerogroup(5)) AND zerogroup(6);                
                
  gma: FOR k IN 1 TO 5 GENERATE
    positionmux(1)(k) <= position(1)(k) AND firstzero(1);
    gmb: FOR j IN 2 TO 6 GENERATE
      positionmux(j)(k) <= positionmux(j-1)(k) OR (position(j)(k) AND firstzero(j));
    END GENERATE;
  END GENERATE;
  
leading <= positionmux(6)(5 DOWNTO 1);
                                               
END rtl;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_LNLUT8.VHD                             ***
--***                                             ***
--***   Function: Look Up Table - LN()            ***
--***                                             ***
--***   Generated by MATLAB Utility               ***
--***                                             ***
--***   22/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_lnlut8 IS
PORT (
      add : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      inv : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
      logman : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
      logexp : OUT STD_LOGIC_VECTOR (8 DOWNTO 1)
     );
END fp_lnlut8;

ARCHITECTURE rtl OF fp_lnlut8 IS

BEGIN

  pca: PROCESS (add)
  BEGIN
    CASE add IS
      WHEN "00000000" =>
            inv <= conv_std_logic_vector(1024,11);
            logman <= conv_std_logic_vector(0,23);
            logexp <= conv_std_logic_vector(0,8);
      WHEN "00000001" =>
            inv <= conv_std_logic_vector(2041,11);
            logman <= conv_std_logic_vector(6316601,23);
            logexp <= conv_std_logic_vector(118,8);
      WHEN "00000010" =>
            inv <= conv_std_logic_vector(2033,11);
            logman <= conv_std_logic_vector(7397915,23);
            logexp <= conv_std_logic_vector(119,8);
      WHEN "00000011" =>
            inv <= conv_std_logic_vector(2025,11);
            logman <= conv_std_logic_vector(3738239,23);
            logexp <= conv_std_logic_vector(120,8);
      WHEN "00000100" =>
            inv <= conv_std_logic_vector(2017,11);
            logman <= conv_std_logic_vector(7988584,23);
            logexp <= conv_std_logic_vector(120,8);
      WHEN "00000101" =>
            inv <= conv_std_logic_vector(2009,11);
            logman <= conv_std_logic_vector(1933606,23);
            logexp <= conv_std_logic_vector(121,8);
      WHEN "00000110" =>
            inv <= conv_std_logic_vector(2002,11);
            logman <= conv_std_logic_vector(3807503,23);
            logexp <= conv_std_logic_vector(121,8);
      WHEN "00000111" =>
            inv <= conv_std_logic_vector(1994,11);
            logman <= conv_std_logic_vector(5957139,23);
            logexp <= conv_std_logic_vector(121,8);
      WHEN "00001000" =>
            inv <= conv_std_logic_vector(1986,11);
            logman <= conv_std_logic_vector(8115417,23);
            logexp <= conv_std_logic_vector(121,8);
      WHEN "00001001" =>
            inv <= conv_std_logic_vector(1979,11);
            logman <= conv_std_logic_vector(811223,23);
            logexp <= conv_std_logic_vector(122,8);
      WHEN "00001010" =>
            inv <= conv_std_logic_vector(1972,11);
            logman <= conv_std_logic_vector(1762400,23);
            logexp <= conv_std_logic_vector(122,8);
      WHEN "00001011" =>
            inv <= conv_std_logic_vector(1964,11);
            logman <= conv_std_logic_vector(2853602,23);
            logexp <= conv_std_logic_vector(122,8);
      WHEN "00001100" =>
            inv <= conv_std_logic_vector(1957,11);
            logman <= conv_std_logic_vector(3812057,23);
            logexp <= conv_std_logic_vector(122,8);
      WHEN "00001101" =>
            inv <= conv_std_logic_vector(1950,11);
            logman <= conv_std_logic_vector(4773946,23);
            logexp <= conv_std_logic_vector(122,8);
      WHEN "00001110" =>
            inv <= conv_std_logic_vector(1942,11);
            logman <= conv_std_logic_vector(5877485,23);
            logexp <= conv_std_logic_vector(122,8);
      WHEN "00001111" =>
            inv <= conv_std_logic_vector(1935,11);
            logman <= conv_std_logic_vector(6846817,23);
            logexp <= conv_std_logic_vector(122,8);
      WHEN "00010000" =>
            inv <= conv_std_logic_vector(1928,11);
            logman <= conv_std_logic_vector(7819662,23);
            logexp <= conv_std_logic_vector(122,8);
      WHEN "00010001" =>
            inv <= conv_std_logic_vector(1921,11);
            logman <= conv_std_logic_vector(203719,23);
            logexp <= conv_std_logic_vector(123,8);
      WHEN "00010010" =>
            inv <= conv_std_logic_vector(1914,11);
            logman <= conv_std_logic_vector(693693,23);
            logexp <= conv_std_logic_vector(123,8);
      WHEN "00010011" =>
            inv <= conv_std_logic_vector(1907,11);
            logman <= conv_std_logic_vector(1185462,23);
            logexp <= conv_std_logic_vector(123,8);
      WHEN "00010100" =>
            inv <= conv_std_logic_vector(1900,11);
            logman <= conv_std_logic_vector(1679040,23);
            logexp <= conv_std_logic_vector(123,8);
      WHEN "00010101" =>
            inv <= conv_std_logic_vector(1893,11);
            logman <= conv_std_logic_vector(2174439,23);
            logexp <= conv_std_logic_vector(123,8);
      WHEN "00010110" =>
            inv <= conv_std_logic_vector(1886,11);
            logman <= conv_std_logic_vector(2671674,23);
            logexp <= conv_std_logic_vector(123,8);
      WHEN "00010111" =>
            inv <= conv_std_logic_vector(1880,11);
            logman <= conv_std_logic_vector(3099346,23);
            logexp <= conv_std_logic_vector(123,8);
      WHEN "00011000" =>
            inv <= conv_std_logic_vector(1873,11);
            logman <= conv_std_logic_vector(3600026,23);
            logexp <= conv_std_logic_vector(123,8);
      WHEN "00011001" =>
            inv <= conv_std_logic_vector(1866,11);
            logman <= conv_std_logic_vector(4102580,23);
            logexp <= conv_std_logic_vector(123,8);
      WHEN "00011010" =>
            inv <= conv_std_logic_vector(1860,11);
            logman <= conv_std_logic_vector(4534844,23);
            logexp <= conv_std_logic_vector(123,8);
      WHEN "00011011" =>
            inv <= conv_std_logic_vector(1853,11);
            logman <= conv_std_logic_vector(5040917,23);
            logexp <= conv_std_logic_vector(123,8);
      WHEN "00011100" =>
            inv <= conv_std_logic_vector(1847,11);
            logman <= conv_std_logic_vector(5476218,23);
            logexp <= conv_std_logic_vector(123,8);
      WHEN "00011101" =>
            inv <= conv_std_logic_vector(1840,11);
            logman <= conv_std_logic_vector(5985860,23);
            logexp <= conv_std_logic_vector(123,8);
      WHEN "00011110" =>
            inv <= conv_std_logic_vector(1834,11);
            logman <= conv_std_logic_vector(6424242,23);
            logexp <= conv_std_logic_vector(123,8);
      WHEN "00011111" =>
            inv <= conv_std_logic_vector(1827,11);
            logman <= conv_std_logic_vector(6937504,23);
            logexp <= conv_std_logic_vector(123,8);
      WHEN "00100000" =>
            inv <= conv_std_logic_vector(1821,11);
            logman <= conv_std_logic_vector(7379010,23);
            logexp <= conv_std_logic_vector(123,8);
      WHEN "00100001" =>
            inv <= conv_std_logic_vector(1815,11);
            logman <= conv_std_logic_vector(7821973,23);
            logexp <= conv_std_logic_vector(123,8);
      WHEN "00100010" =>
            inv <= conv_std_logic_vector(1808,11);
            logman <= conv_std_logic_vector(8340618,23);
            logexp <= conv_std_logic_vector(123,8);
      WHEN "00100011" =>
            inv <= conv_std_logic_vector(1802,11);
            logman <= conv_std_logic_vector(199082,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00100100" =>
            inv <= conv_std_logic_vector(1796,11);
            logman <= conv_std_logic_vector(422902,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00100101" =>
            inv <= conv_std_logic_vector(1790,11);
            logman <= conv_std_logic_vector(647472,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00100110" =>
            inv <= conv_std_logic_vector(1784,11);
            logman <= conv_std_logic_vector(872796,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00100111" =>
            inv <= conv_std_logic_vector(1778,11);
            logman <= conv_std_logic_vector(1098879,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00101000" =>
            inv <= conv_std_logic_vector(1772,11);
            logman <= conv_std_logic_vector(1325726,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00101001" =>
            inv <= conv_std_logic_vector(1766,11);
            logman <= conv_std_logic_vector(1553342,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00101010" =>
            inv <= conv_std_logic_vector(1760,11);
            logman <= conv_std_logic_vector(1781734,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00101011" =>
            inv <= conv_std_logic_vector(1754,11);
            logman <= conv_std_logic_vector(2010905,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00101100" =>
            inv <= conv_std_logic_vector(1748,11);
            logman <= conv_std_logic_vector(2240861,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00101101" =>
            inv <= conv_std_logic_vector(1742,11);
            logman <= conv_std_logic_vector(2471608,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00101110" =>
            inv <= conv_std_logic_vector(1737,11);
            logman <= conv_std_logic_vector(2664505,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00101111" =>
            inv <= conv_std_logic_vector(1731,11);
            logman <= conv_std_logic_vector(2896716,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00110000" =>
            inv <= conv_std_logic_vector(1725,11);
            logman <= conv_std_logic_vector(3129733,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00110001" =>
            inv <= conv_std_logic_vector(1719,11);
            logman <= conv_std_logic_vector(3363562,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00110010" =>
            inv <= conv_std_logic_vector(1714,11);
            logman <= conv_std_logic_vector(3559044,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00110011" =>
            inv <= conv_std_logic_vector(1708,11);
            logman <= conv_std_logic_vector(3794376,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00110100" =>
            inv <= conv_std_logic_vector(1703,11);
            logman <= conv_std_logic_vector(3991119,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00110101" =>
            inv <= conv_std_logic_vector(1697,11);
            logman <= conv_std_logic_vector(4227974,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00110110" =>
            inv <= conv_std_logic_vector(1692,11);
            logman <= conv_std_logic_vector(4425994,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00110111" =>
            inv <= conv_std_logic_vector(1686,11);
            logman <= conv_std_logic_vector(4664391,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00111000" =>
            inv <= conv_std_logic_vector(1681,11);
            logman <= conv_std_logic_vector(4863705,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00111001" =>
            inv <= conv_std_logic_vector(1676,11);
            logman <= conv_std_logic_vector(5063612,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00111010" =>
            inv <= conv_std_logic_vector(1670,11);
            logman <= conv_std_logic_vector(5304290,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00111011" =>
            inv <= conv_std_logic_vector(1665,11);
            logman <= conv_std_logic_vector(5505516,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00111100" =>
            inv <= conv_std_logic_vector(1660,11);
            logman <= conv_std_logic_vector(5707347,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00111101" =>
            inv <= conv_std_logic_vector(1654,11);
            logman <= conv_std_logic_vector(5950349,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00111110" =>
            inv <= conv_std_logic_vector(1649,11);
            logman <= conv_std_logic_vector(6153525,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "00111111" =>
            inv <= conv_std_logic_vector(1644,11);
            logman <= conv_std_logic_vector(6357317,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "01000000" =>
            inv <= conv_std_logic_vector(1639,11);
            logman <= conv_std_logic_vector(6561731,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "01000001" =>
            inv <= conv_std_logic_vector(1634,11);
            logman <= conv_std_logic_vector(6766769,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "01000010" =>
            inv <= conv_std_logic_vector(1629,11);
            logman <= conv_std_logic_vector(6972435,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "01000011" =>
            inv <= conv_std_logic_vector(1624,11);
            logman <= conv_std_logic_vector(7178734,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "01000100" =>
            inv <= conv_std_logic_vector(1619,11);
            logman <= conv_std_logic_vector(7385668,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "01000101" =>
            inv <= conv_std_logic_vector(1614,11);
            logman <= conv_std_logic_vector(7593243,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "01000110" =>
            inv <= conv_std_logic_vector(1609,11);
            logman <= conv_std_logic_vector(7801462,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "01000111" =>
            inv <= conv_std_logic_vector(1604,11);
            logman <= conv_std_logic_vector(8010329,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "01001000" =>
            inv <= conv_std_logic_vector(1599,11);
            logman <= conv_std_logic_vector(8219848,23);
            logexp <= conv_std_logic_vector(124,8);
      WHEN "01001001" =>
            inv <= conv_std_logic_vector(1594,11);
            logman <= conv_std_logic_vector(20707,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01001010" =>
            inv <= conv_std_logic_vector(1589,11);
            logman <= conv_std_logic_vector(126125,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01001011" =>
            inv <= conv_std_logic_vector(1584,11);
            logman <= conv_std_logic_vector(231875,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01001100" =>
            inv <= conv_std_logic_vector(1580,11);
            logman <= conv_std_logic_vector(316716,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01001101" =>
            inv <= conv_std_logic_vector(1575,11);
            logman <= conv_std_logic_vector(423069,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01001110" =>
            inv <= conv_std_logic_vector(1570,11);
            logman <= conv_std_logic_vector(529760,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01001111" =>
            inv <= conv_std_logic_vector(1566,11);
            logman <= conv_std_logic_vector(615358,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01010000" =>
            inv <= conv_std_logic_vector(1561,11);
            logman <= conv_std_logic_vector(722664,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01010001" =>
            inv <= conv_std_logic_vector(1556,11);
            logman <= conv_std_logic_vector(830314,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01010010" =>
            inv <= conv_std_logic_vector(1552,11);
            logman <= conv_std_logic_vector(916683,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01010011" =>
            inv <= conv_std_logic_vector(1547,11);
            logman <= conv_std_logic_vector(1024958,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01010100" =>
            inv <= conv_std_logic_vector(1543,11);
            logman <= conv_std_logic_vector(1111831,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01010101" =>
            inv <= conv_std_logic_vector(1538,11);
            logman <= conv_std_logic_vector(1220738,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01010110" =>
            inv <= conv_std_logic_vector(1534,11);
            logman <= conv_std_logic_vector(1308120,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01010111" =>
            inv <= conv_std_logic_vector(1529,11);
            logman <= conv_std_logic_vector(1417667,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01011000" =>
            inv <= conv_std_logic_vector(1525,11);
            logman <= conv_std_logic_vector(1505564,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01011001" =>
            inv <= conv_std_logic_vector(1520,11);
            logman <= conv_std_logic_vector(1615759,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01011010" =>
            inv <= conv_std_logic_vector(1516,11);
            logman <= conv_std_logic_vector(1704177,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01011011" =>
            inv <= conv_std_logic_vector(1511,11);
            logman <= conv_std_logic_vector(1815027,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01011100" =>
            inv <= conv_std_logic_vector(1507,11);
            logman <= conv_std_logic_vector(1903972,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01011101" =>
            inv <= conv_std_logic_vector(1503,11);
            logman <= conv_std_logic_vector(1993153,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01011110" =>
            inv <= conv_std_logic_vector(1498,11);
            logman <= conv_std_logic_vector(2104964,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01011111" =>
            inv <= conv_std_logic_vector(1494,11);
            logman <= conv_std_logic_vector(2194682,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01100000" =>
            inv <= conv_std_logic_vector(1490,11);
            logman <= conv_std_logic_vector(2284640,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01100001" =>
            inv <= conv_std_logic_vector(1486,11);
            logman <= conv_std_logic_vector(2374840,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01100010" =>
            inv <= conv_std_logic_vector(1482,11);
            logman <= conv_std_logic_vector(2465284,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01100011" =>
            inv <= conv_std_logic_vector(1477,11);
            logman <= conv_std_logic_vector(2578682,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01100100" =>
            inv <= conv_std_logic_vector(1473,11);
            logman <= conv_std_logic_vector(2669677,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01100101" =>
            inv <= conv_std_logic_vector(1469,11);
            logman <= conv_std_logic_vector(2760919,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01100110" =>
            inv <= conv_std_logic_vector(1465,11);
            logman <= conv_std_logic_vector(2852411,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01100111" =>
            inv <= conv_std_logic_vector(1461,11);
            logman <= conv_std_logic_vector(2944152,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01101000" =>
            inv <= conv_std_logic_vector(1457,11);
            logman <= conv_std_logic_vector(3036145,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01101001" =>
            inv <= conv_std_logic_vector(1453,11);
            logman <= conv_std_logic_vector(3128391,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01101010" =>
            inv <= conv_std_logic_vector(1449,11);
            logman <= conv_std_logic_vector(3220891,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01101011" =>
            inv <= conv_std_logic_vector(1445,11);
            logman <= conv_std_logic_vector(3313647,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01101100" =>
            inv <= conv_std_logic_vector(1441,11);
            logman <= conv_std_logic_vector(3406660,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01101101" =>
            inv <= conv_std_logic_vector(1437,11);
            logman <= conv_std_logic_vector(3499932,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01101110" =>
            inv <= conv_std_logic_vector(1433,11);
            logman <= conv_std_logic_vector(3593464,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01101111" =>
            inv <= conv_std_logic_vector(1429,11);
            logman <= conv_std_logic_vector(3687257,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01110000" =>
            inv <= conv_std_logic_vector(1425,11);
            logman <= conv_std_logic_vector(3781312,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01110001" =>
            inv <= conv_std_logic_vector(1421,11);
            logman <= conv_std_logic_vector(3875633,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01110010" =>
            inv <= conv_std_logic_vector(1417,11);
            logman <= conv_std_logic_vector(3970219,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01110011" =>
            inv <= conv_std_logic_vector(1414,11);
            logman <= conv_std_logic_vector(4041334,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01110100" =>
            inv <= conv_std_logic_vector(1410,11);
            logman <= conv_std_logic_vector(4136389,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01110101" =>
            inv <= conv_std_logic_vector(1406,11);
            logman <= conv_std_logic_vector(4231714,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01110110" =>
            inv <= conv_std_logic_vector(1402,11);
            logman <= conv_std_logic_vector(4327311,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01110111" =>
            inv <= conv_std_logic_vector(1399,11);
            logman <= conv_std_logic_vector(4399188,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01111000" =>
            inv <= conv_std_logic_vector(1395,11);
            logman <= conv_std_logic_vector(4495263,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01111001" =>
            inv <= conv_std_logic_vector(1391,11);
            logman <= conv_std_logic_vector(4591615,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01111010" =>
            inv <= conv_std_logic_vector(1388,11);
            logman <= conv_std_logic_vector(4664061,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01111011" =>
            inv <= conv_std_logic_vector(1384,11);
            logman <= conv_std_logic_vector(4760899,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01111100" =>
            inv <= conv_std_logic_vector(1380,11);
            logman <= conv_std_logic_vector(4858018,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01111101" =>
            inv <= conv_std_logic_vector(1377,11);
            logman <= conv_std_logic_vector(4931041,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01111110" =>
            inv <= conv_std_logic_vector(1373,11);
            logman <= conv_std_logic_vector(5028654,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "01111111" =>
            inv <= conv_std_logic_vector(1369,11);
            logman <= conv_std_logic_vector(5126552,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10000000" =>
            inv <= conv_std_logic_vector(1366,11);
            logman <= conv_std_logic_vector(5200163,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10000001" =>
            inv <= conv_std_logic_vector(1362,11);
            logman <= conv_std_logic_vector(5298564,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10000010" =>
            inv <= conv_std_logic_vector(1359,11);
            logman <= conv_std_logic_vector(5372554,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10000011" =>
            inv <= conv_std_logic_vector(1355,11);
            logman <= conv_std_logic_vector(5471461,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10000100" =>
            inv <= conv_std_logic_vector(1352,11);
            logman <= conv_std_logic_vector(5545834,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10000101" =>
            inv <= conv_std_logic_vector(1348,11);
            logman <= conv_std_logic_vector(5645255,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10000110" =>
            inv <= conv_std_logic_vector(1345,11);
            logman <= conv_std_logic_vector(5720014,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10000111" =>
            inv <= conv_std_logic_vector(1341,11);
            logman <= conv_std_logic_vector(5819953,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10001000" =>
            inv <= conv_std_logic_vector(1338,11);
            logman <= conv_std_logic_vector(5895103,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10001001" =>
            inv <= conv_std_logic_vector(1335,11);
            logman <= conv_std_logic_vector(5970421,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10001010" =>
            inv <= conv_std_logic_vector(1331,11);
            logman <= conv_std_logic_vector(6071110,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10001011" =>
            inv <= conv_std_logic_vector(1328,11);
            logman <= conv_std_logic_vector(6146825,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10001100" =>
            inv <= conv_std_logic_vector(1324,11);
            logman <= conv_std_logic_vector(6248045,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10001101" =>
            inv <= conv_std_logic_vector(1321,11);
            logman <= conv_std_logic_vector(6324161,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10001110" =>
            inv <= conv_std_logic_vector(1318,11);
            logman <= conv_std_logic_vector(6400450,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10001111" =>
            inv <= conv_std_logic_vector(1315,11);
            logman <= conv_std_logic_vector(6476913,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10010000" =>
            inv <= conv_std_logic_vector(1311,11);
            logman <= conv_std_logic_vector(6579135,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10010001" =>
            inv <= conv_std_logic_vector(1308,11);
            logman <= conv_std_logic_vector(6656007,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10010010" =>
            inv <= conv_std_logic_vector(1305,11);
            logman <= conv_std_logic_vector(6733055,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10010011" =>
            inv <= conv_std_logic_vector(1301,11);
            logman <= conv_std_logic_vector(6836061,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10010100" =>
            inv <= conv_std_logic_vector(1298,11);
            logman <= conv_std_logic_vector(6913525,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10010101" =>
            inv <= conv_std_logic_vector(1295,11);
            logman <= conv_std_logic_vector(6991167,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10010110" =>
            inv <= conv_std_logic_vector(1292,11);
            logman <= conv_std_logic_vector(7068989,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10010111" =>
            inv <= conv_std_logic_vector(1289,11);
            logman <= conv_std_logic_vector(7146993,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10011000" =>
            inv <= conv_std_logic_vector(1286,11);
            logman <= conv_std_logic_vector(7225178,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10011001" =>
            inv <= conv_std_logic_vector(1282,11);
            logman <= conv_std_logic_vector(7329709,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10011010" =>
            inv <= conv_std_logic_vector(1279,11);
            logman <= conv_std_logic_vector(7408321,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10011011" =>
            inv <= conv_std_logic_vector(1276,11);
            logman <= conv_std_logic_vector(7487119,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10011100" =>
            inv <= conv_std_logic_vector(1273,11);
            logman <= conv_std_logic_vector(7566101,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10011101" =>
            inv <= conv_std_logic_vector(1270,11);
            logman <= conv_std_logic_vector(7645270,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10011110" =>
            inv <= conv_std_logic_vector(1267,11);
            logman <= conv_std_logic_vector(7724626,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10011111" =>
            inv <= conv_std_logic_vector(1264,11);
            logman <= conv_std_logic_vector(7804171,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10100000" =>
            inv <= conv_std_logic_vector(1261,11);
            logman <= conv_std_logic_vector(7883904,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10100001" =>
            inv <= conv_std_logic_vector(1258,11);
            logman <= conv_std_logic_vector(7963827,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10100010" =>
            inv <= conv_std_logic_vector(1255,11);
            logman <= conv_std_logic_vector(8043941,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10100011" =>
            inv <= conv_std_logic_vector(1252,11);
            logman <= conv_std_logic_vector(8124247,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10100100" =>
            inv <= conv_std_logic_vector(1249,11);
            logman <= conv_std_logic_vector(8204746,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10100101" =>
            inv <= conv_std_logic_vector(1246,11);
            logman <= conv_std_logic_vector(8285438,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10100110" =>
            inv <= conv_std_logic_vector(1243,11);
            logman <= conv_std_logic_vector(8366324,23);
            logexp <= conv_std_logic_vector(125,8);
      WHEN "10100111" =>
            inv <= conv_std_logic_vector(1240,11);
            logman <= conv_std_logic_vector(29399,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10101000" =>
            inv <= conv_std_logic_vector(1237,11);
            logman <= conv_std_logic_vector(70038,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10101001" =>
            inv <= conv_std_logic_vector(1234,11);
            logman <= conv_std_logic_vector(110776,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10101010" =>
            inv <= conv_std_logic_vector(1231,11);
            logman <= conv_std_logic_vector(151613,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10101011" =>
            inv <= conv_std_logic_vector(1228,11);
            logman <= conv_std_logic_vector(192550,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10101100" =>
            inv <= conv_std_logic_vector(1225,11);
            logman <= conv_std_logic_vector(233587,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10101101" =>
            inv <= conv_std_logic_vector(1223,11);
            logman <= conv_std_logic_vector(261001,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10101110" =>
            inv <= conv_std_logic_vector(1220,11);
            logman <= conv_std_logic_vector(302205,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10101111" =>
            inv <= conv_std_logic_vector(1217,11);
            logman <= conv_std_logic_vector(343512,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10110000" =>
            inv <= conv_std_logic_vector(1214,11);
            logman <= conv_std_logic_vector(384920,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10110001" =>
            inv <= conv_std_logic_vector(1211,11);
            logman <= conv_std_logic_vector(426431,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10110010" =>
            inv <= conv_std_logic_vector(1209,11);
            logman <= conv_std_logic_vector(454162,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10110011" =>
            inv <= conv_std_logic_vector(1206,11);
            logman <= conv_std_logic_vector(495844,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10110100" =>
            inv <= conv_std_logic_vector(1203,11);
            logman <= conv_std_logic_vector(537630,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10110101" =>
            inv <= conv_std_logic_vector(1200,11);
            logman <= conv_std_logic_vector(579521,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10110110" =>
            inv <= conv_std_logic_vector(1198,11);
            logman <= conv_std_logic_vector(607506,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10110111" =>
            inv <= conv_std_logic_vector(1195,11);
            logman <= conv_std_logic_vector(649572,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10111000" =>
            inv <= conv_std_logic_vector(1192,11);
            logman <= conv_std_logic_vector(691744,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10111001" =>
            inv <= conv_std_logic_vector(1189,11);
            logman <= conv_std_logic_vector(734021,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10111010" =>
            inv <= conv_std_logic_vector(1187,11);
            logman <= conv_std_logic_vector(762266,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10111011" =>
            inv <= conv_std_logic_vector(1184,11);
            logman <= conv_std_logic_vector(804722,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10111100" =>
            inv <= conv_std_logic_vector(1181,11);
            logman <= conv_std_logic_vector(847286,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10111101" =>
            inv <= conv_std_logic_vector(1179,11);
            logman <= conv_std_logic_vector(875722,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10111110" =>
            inv <= conv_std_logic_vector(1176,11);
            logman <= conv_std_logic_vector(918466,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "10111111" =>
            inv <= conv_std_logic_vector(1173,11);
            logman <= conv_std_logic_vector(961320,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11000000" =>
            inv <= conv_std_logic_vector(1171,11);
            logman <= conv_std_logic_vector(989950,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11000001" =>
            inv <= conv_std_logic_vector(1168,11);
            logman <= conv_std_logic_vector(1032987,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11000010" =>
            inv <= conv_std_logic_vector(1166,11);
            logman <= conv_std_logic_vector(1061740,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11000011" =>
            inv <= conv_std_logic_vector(1163,11);
            logman <= conv_std_logic_vector(1104961,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11000100" =>
            inv <= conv_std_logic_vector(1160,11);
            logman <= conv_std_logic_vector(1148295,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11000101" =>
            inv <= conv_std_logic_vector(1158,11);
            logman <= conv_std_logic_vector(1177246,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11000110" =>
            inv <= conv_std_logic_vector(1155,11);
            logman <= conv_std_logic_vector(1220767,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11000111" =>
            inv <= conv_std_logic_vector(1153,11);
            logman <= conv_std_logic_vector(1249843,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11001000" =>
            inv <= conv_std_logic_vector(1150,11);
            logman <= conv_std_logic_vector(1293553,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11001001" =>
            inv <= conv_std_logic_vector(1148,11);
            logman <= conv_std_logic_vector(1322756,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11001010" =>
            inv <= conv_std_logic_vector(1145,11);
            logman <= conv_std_logic_vector(1366656,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11001011" =>
            inv <= conv_std_logic_vector(1143,11);
            logman <= conv_std_logic_vector(1395987,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11001100" =>
            inv <= conv_std_logic_vector(1140,11);
            logman <= conv_std_logic_vector(1440080,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11001101" =>
            inv <= conv_std_logic_vector(1138,11);
            logman <= conv_std_logic_vector(1469539,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11001110" =>
            inv <= conv_std_logic_vector(1135,11);
            logman <= conv_std_logic_vector(1513826,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11001111" =>
            inv <= conv_std_logic_vector(1133,11);
            logman <= conv_std_logic_vector(1543415,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11010000" =>
            inv <= conv_std_logic_vector(1130,11);
            logman <= conv_std_logic_vector(1587898,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11010001" =>
            inv <= conv_std_logic_vector(1128,11);
            logman <= conv_std_logic_vector(1617618,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11010010" =>
            inv <= conv_std_logic_vector(1126,11);
            logman <= conv_std_logic_vector(1647391,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11010011" =>
            inv <= conv_std_logic_vector(1123,11);
            logman <= conv_std_logic_vector(1692151,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11010100" =>
            inv <= conv_std_logic_vector(1121,11);
            logman <= conv_std_logic_vector(1722056,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11010101" =>
            inv <= conv_std_logic_vector(1118,11);
            logman <= conv_std_logic_vector(1767016,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11010110" =>
            inv <= conv_std_logic_vector(1116,11);
            logman <= conv_std_logic_vector(1797055,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11010111" =>
            inv <= conv_std_logic_vector(1114,11);
            logman <= conv_std_logic_vector(1827149,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11011000" =>
            inv <= conv_std_logic_vector(1111,11);
            logman <= conv_std_logic_vector(1872391,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11011001" =>
            inv <= conv_std_logic_vector(1109,11);
            logman <= conv_std_logic_vector(1902620,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11011010" =>
            inv <= conv_std_logic_vector(1107,11);
            logman <= conv_std_logic_vector(1932904,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11011011" =>
            inv <= conv_std_logic_vector(1104,11);
            logman <= conv_std_logic_vector(1978432,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11011100" =>
            inv <= conv_std_logic_vector(1102,11);
            logman <= conv_std_logic_vector(2008853,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11011101" =>
            inv <= conv_std_logic_vector(1100,11);
            logman <= conv_std_logic_vector(2039330,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11011110" =>
            inv <= conv_std_logic_vector(1097,11);
            logman <= conv_std_logic_vector(2085148,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11011111" =>
            inv <= conv_std_logic_vector(1095,11);
            logman <= conv_std_logic_vector(2115764,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11100000" =>
            inv <= conv_std_logic_vector(1093,11);
            logman <= conv_std_logic_vector(2146435,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11100001" =>
            inv <= conv_std_logic_vector(1090,11);
            logman <= conv_std_logic_vector(2192547,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11100010" =>
            inv <= conv_std_logic_vector(1088,11);
            logman <= conv_std_logic_vector(2223360,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11100011" =>
            inv <= conv_std_logic_vector(1086,11);
            logman <= conv_std_logic_vector(2254228,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11100100" =>
            inv <= conv_std_logic_vector(1084,11);
            logman <= conv_std_logic_vector(2285154,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11100101" =>
            inv <= conv_std_logic_vector(1082,11);
            logman <= conv_std_logic_vector(2316137,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11100110" =>
            inv <= conv_std_logic_vector(1079,11);
            logman <= conv_std_logic_vector(2362719,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11100111" =>
            inv <= conv_std_logic_vector(1077,11);
            logman <= conv_std_logic_vector(2393845,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11101000" =>
            inv <= conv_std_logic_vector(1075,11);
            logman <= conv_std_logic_vector(2425030,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11101001" =>
            inv <= conv_std_logic_vector(1073,11);
            logman <= conv_std_logic_vector(2456272,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11101010" =>
            inv <= conv_std_logic_vector(1070,11);
            logman <= conv_std_logic_vector(2503245,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11101011" =>
            inv <= conv_std_logic_vector(1068,11);
            logman <= conv_std_logic_vector(2534634,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11101100" =>
            inv <= conv_std_logic_vector(1066,11);
            logman <= conv_std_logic_vector(2566082,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11101101" =>
            inv <= conv_std_logic_vector(1064,11);
            logman <= conv_std_logic_vector(2597588,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11101110" =>
            inv <= conv_std_logic_vector(1062,11);
            logman <= conv_std_logic_vector(2629154,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11101111" =>
            inv <= conv_std_logic_vector(1060,11);
            logman <= conv_std_logic_vector(2660779,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11110000" =>
            inv <= conv_std_logic_vector(1058,11);
            logman <= conv_std_logic_vector(2692464,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11110001" =>
            inv <= conv_std_logic_vector(1055,11);
            logman <= conv_std_logic_vector(2740104,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11110010" =>
            inv <= conv_std_logic_vector(1053,11);
            logman <= conv_std_logic_vector(2771940,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11110011" =>
            inv <= conv_std_logic_vector(1051,11);
            logman <= conv_std_logic_vector(2803835,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11110100" =>
            inv <= conv_std_logic_vector(1049,11);
            logman <= conv_std_logic_vector(2835792,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11110101" =>
            inv <= conv_std_logic_vector(1047,11);
            logman <= conv_std_logic_vector(2867810,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11110110" =>
            inv <= conv_std_logic_vector(1045,11);
            logman <= conv_std_logic_vector(2899888,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11110111" =>
            inv <= conv_std_logic_vector(1043,11);
            logman <= conv_std_logic_vector(2932029,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11111000" =>
            inv <= conv_std_logic_vector(1041,11);
            logman <= conv_std_logic_vector(2964231,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11111001" =>
            inv <= conv_std_logic_vector(1039,11);
            logman <= conv_std_logic_vector(2996495,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11111010" =>
            inv <= conv_std_logic_vector(1037,11);
            logman <= conv_std_logic_vector(3028821,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11111011" =>
            inv <= conv_std_logic_vector(1035,11);
            logman <= conv_std_logic_vector(3061209,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11111100" =>
            inv <= conv_std_logic_vector(1033,11);
            logman <= conv_std_logic_vector(3093660,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11111101" =>
            inv <= conv_std_logic_vector(1031,11);
            logman <= conv_std_logic_vector(3126174,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11111110" =>
            inv <= conv_std_logic_vector(1029,11);
            logman <= conv_std_logic_vector(3158751,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "11111111" =>
            inv <= conv_std_logic_vector(1027,11);
            logman <= conv_std_logic_vector(3191392,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN others =>
           inv <= conv_std_logic_vector(0,11);
           logman <= conv_std_logic_vector(0,23);
           logexp <= conv_std_logic_vector(0,8);
    END CASE;
  END PROCESS;

END rtl;
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_LNLUTPOW.VHD                           ***
--***                                             ***
--***   Function: Look Up Table - LN()            ***
--***                                             ***
--***   Generated by MATLAB Utility               ***
--***                                             ***
--***   22/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_lnlutpow IS
PORT (
      add : IN STD_LOGIC_VECTOR (7 DOWNTO 1);
      logman : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
      logexp : OUT STD_LOGIC_VECTOR (8 DOWNTO 1)
     );
END fp_lnlutpow;

ARCHITECTURE rtl OF fp_lnlutpow IS

BEGIN

  pca: PROCESS (add)
  BEGIN
    CASE add IS
      WHEN "0000000" =>
            logman <= conv_std_logic_vector(0,23);
            logexp <= conv_std_logic_vector(0,8);
      WHEN "0000001" =>
            logman <= conv_std_logic_vector(3240472,23);
            logexp <= conv_std_logic_vector(126,8);
      WHEN "0000010" =>
            logman <= conv_std_logic_vector(3240472,23);
            logexp <= conv_std_logic_vector(127,8);
      WHEN "0000011" =>
            logman <= conv_std_logic_vector(333202,23);
            logexp <= conv_std_logic_vector(128,8);
      WHEN "0000100" =>
            logman <= conv_std_logic_vector(3240472,23);
            logexp <= conv_std_logic_vector(128,8);
      WHEN "0000101" =>
            logman <= conv_std_logic_vector(6147742,23);
            logexp <= conv_std_logic_vector(128,8);
      WHEN "0000110" =>
            logman <= conv_std_logic_vector(333202,23);
            logexp <= conv_std_logic_vector(129,8);
      WHEN "0000111" =>
            logman <= conv_std_logic_vector(1786837,23);
            logexp <= conv_std_logic_vector(129,8);
      WHEN "0001000" =>
            logman <= conv_std_logic_vector(3240472,23);
            logexp <= conv_std_logic_vector(129,8);
      WHEN "0001001" =>
            logman <= conv_std_logic_vector(4694107,23);
            logexp <= conv_std_logic_vector(129,8);
      WHEN "0001010" =>
            logman <= conv_std_logic_vector(6147742,23);
            logexp <= conv_std_logic_vector(129,8);
      WHEN "0001011" =>
            logman <= conv_std_logic_vector(7601377,23);
            logexp <= conv_std_logic_vector(129,8);
      WHEN "0001100" =>
            logman <= conv_std_logic_vector(333202,23);
            logexp <= conv_std_logic_vector(130,8);
      WHEN "0001101" =>
            logman <= conv_std_logic_vector(1060019,23);
            logexp <= conv_std_logic_vector(130,8);
      WHEN "0001110" =>
            logman <= conv_std_logic_vector(1786837,23);
            logexp <= conv_std_logic_vector(130,8);
      WHEN "0001111" =>
            logman <= conv_std_logic_vector(2513654,23);
            logexp <= conv_std_logic_vector(130,8);
      WHEN "0010000" =>
            logman <= conv_std_logic_vector(3240472,23);
            logexp <= conv_std_logic_vector(130,8);
      WHEN "0010001" =>
            logman <= conv_std_logic_vector(3967289,23);
            logexp <= conv_std_logic_vector(130,8);
      WHEN "0010010" =>
            logman <= conv_std_logic_vector(4694107,23);
            logexp <= conv_std_logic_vector(130,8);
      WHEN "0010011" =>
            logman <= conv_std_logic_vector(5420924,23);
            logexp <= conv_std_logic_vector(130,8);
      WHEN "0010100" =>
            logman <= conv_std_logic_vector(6147742,23);
            logexp <= conv_std_logic_vector(130,8);
      WHEN "0010101" =>
            logman <= conv_std_logic_vector(6874559,23);
            logexp <= conv_std_logic_vector(130,8);
      WHEN "0010110" =>
            logman <= conv_std_logic_vector(7601377,23);
            logexp <= conv_std_logic_vector(130,8);
      WHEN "0010111" =>
            logman <= conv_std_logic_vector(8328194,23);
            logexp <= conv_std_logic_vector(130,8);
      WHEN "0011000" =>
            logman <= conv_std_logic_vector(333202,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0011001" =>
            logman <= conv_std_logic_vector(696611,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0011010" =>
            logman <= conv_std_logic_vector(1060019,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0011011" =>
            logman <= conv_std_logic_vector(1423428,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0011100" =>
            logman <= conv_std_logic_vector(1786837,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0011101" =>
            logman <= conv_std_logic_vector(2150246,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0011110" =>
            logman <= conv_std_logic_vector(2513654,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0011111" =>
            logman <= conv_std_logic_vector(2877063,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0100000" =>
            logman <= conv_std_logic_vector(3240472,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0100001" =>
            logman <= conv_std_logic_vector(3603881,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0100010" =>
            logman <= conv_std_logic_vector(3967289,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0100011" =>
            logman <= conv_std_logic_vector(4330698,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0100100" =>
            logman <= conv_std_logic_vector(4694107,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0100101" =>
            logman <= conv_std_logic_vector(5057516,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0100110" =>
            logman <= conv_std_logic_vector(5420924,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0100111" =>
            logman <= conv_std_logic_vector(5784333,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0101000" =>
            logman <= conv_std_logic_vector(6147742,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0101001" =>
            logman <= conv_std_logic_vector(6511151,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0101010" =>
            logman <= conv_std_logic_vector(6874559,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0101011" =>
            logman <= conv_std_logic_vector(7237968,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0101100" =>
            logman <= conv_std_logic_vector(7601377,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0101101" =>
            logman <= conv_std_logic_vector(7964786,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0101110" =>
            logman <= conv_std_logic_vector(8328194,23);
            logexp <= conv_std_logic_vector(131,8);
      WHEN "0101111" =>
            logman <= conv_std_logic_vector(151498,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "0110000" =>
            logman <= conv_std_logic_vector(333202,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "0110001" =>
            logman <= conv_std_logic_vector(514906,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "0110010" =>
            logman <= conv_std_logic_vector(696611,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "0110011" =>
            logman <= conv_std_logic_vector(878315,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "0110100" =>
            logman <= conv_std_logic_vector(1060019,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "0110101" =>
            logman <= conv_std_logic_vector(1241724,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "0110110" =>
            logman <= conv_std_logic_vector(1423428,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "0110111" =>
            logman <= conv_std_logic_vector(1605133,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "0111000" =>
            logman <= conv_std_logic_vector(1786837,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "0111001" =>
            logman <= conv_std_logic_vector(1968541,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "0111010" =>
            logman <= conv_std_logic_vector(2150246,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "0111011" =>
            logman <= conv_std_logic_vector(2331950,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "0111100" =>
            logman <= conv_std_logic_vector(2513654,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "0111101" =>
            logman <= conv_std_logic_vector(2695359,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "0111110" =>
            logman <= conv_std_logic_vector(2877063,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "0111111" =>
            logman <= conv_std_logic_vector(3058768,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1000000" =>
            logman <= conv_std_logic_vector(3240472,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1000001" =>
            logman <= conv_std_logic_vector(3422176,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1000010" =>
            logman <= conv_std_logic_vector(3603881,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1000011" =>
            logman <= conv_std_logic_vector(3785585,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1000100" =>
            logman <= conv_std_logic_vector(3967289,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1000101" =>
            logman <= conv_std_logic_vector(4148994,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1000110" =>
            logman <= conv_std_logic_vector(4330698,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1000111" =>
            logman <= conv_std_logic_vector(4512403,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1001000" =>
            logman <= conv_std_logic_vector(4694107,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1001001" =>
            logman <= conv_std_logic_vector(4875811,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1001010" =>
            logman <= conv_std_logic_vector(5057516,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1001011" =>
            logman <= conv_std_logic_vector(5239220,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1001100" =>
            logman <= conv_std_logic_vector(5420924,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1001101" =>
            logman <= conv_std_logic_vector(5602629,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1001110" =>
            logman <= conv_std_logic_vector(5784333,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1001111" =>
            logman <= conv_std_logic_vector(5966038,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1010000" =>
            logman <= conv_std_logic_vector(6147742,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1010001" =>
            logman <= conv_std_logic_vector(6329446,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1010010" =>
            logman <= conv_std_logic_vector(6511151,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1010011" =>
            logman <= conv_std_logic_vector(6692855,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1010100" =>
            logman <= conv_std_logic_vector(6874559,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1010101" =>
            logman <= conv_std_logic_vector(7056264,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1010110" =>
            logman <= conv_std_logic_vector(7237968,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1010111" =>
            logman <= conv_std_logic_vector(7419673,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1011000" =>
            logman <= conv_std_logic_vector(7601377,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1011001" =>
            logman <= conv_std_logic_vector(7783081,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1011010" =>
            logman <= conv_std_logic_vector(7964786,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1011011" =>
            logman <= conv_std_logic_vector(8146490,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1011100" =>
            logman <= conv_std_logic_vector(8328194,23);
            logexp <= conv_std_logic_vector(132,8);
      WHEN "1011101" =>
            logman <= conv_std_logic_vector(60645,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1011110" =>
            logman <= conv_std_logic_vector(151498,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1011111" =>
            logman <= conv_std_logic_vector(242350,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1100000" =>
            logman <= conv_std_logic_vector(333202,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1100001" =>
            logman <= conv_std_logic_vector(424054,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1100010" =>
            logman <= conv_std_logic_vector(514906,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1100011" =>
            logman <= conv_std_logic_vector(605759,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1100100" =>
            logman <= conv_std_logic_vector(696611,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1100101" =>
            logman <= conv_std_logic_vector(787463,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1100110" =>
            logman <= conv_std_logic_vector(878315,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1100111" =>
            logman <= conv_std_logic_vector(969167,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1101000" =>
            logman <= conv_std_logic_vector(1060019,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1101001" =>
            logman <= conv_std_logic_vector(1150872,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1101010" =>
            logman <= conv_std_logic_vector(1241724,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1101011" =>
            logman <= conv_std_logic_vector(1332576,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1101100" =>
            logman <= conv_std_logic_vector(1423428,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1101101" =>
            logman <= conv_std_logic_vector(1514280,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1101110" =>
            logman <= conv_std_logic_vector(1605133,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1101111" =>
            logman <= conv_std_logic_vector(1695985,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1110000" =>
            logman <= conv_std_logic_vector(1786837,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1110001" =>
            logman <= conv_std_logic_vector(1877689,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1110010" =>
            logman <= conv_std_logic_vector(1968541,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1110011" =>
            logman <= conv_std_logic_vector(2059394,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1110100" =>
            logman <= conv_std_logic_vector(2150246,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1110101" =>
            logman <= conv_std_logic_vector(2241098,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1110110" =>
            logman <= conv_std_logic_vector(2331950,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1110111" =>
            logman <= conv_std_logic_vector(2422802,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1111000" =>
            logman <= conv_std_logic_vector(2513654,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1111001" =>
            logman <= conv_std_logic_vector(2604507,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1111010" =>
            logman <= conv_std_logic_vector(2695359,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1111011" =>
            logman <= conv_std_logic_vector(2786211,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1111100" =>
            logman <= conv_std_logic_vector(2877063,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1111101" =>
            logman <= conv_std_logic_vector(2967915,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1111110" =>
            logman <= conv_std_logic_vector(3058768,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN "1111111" =>
            logman <= conv_std_logic_vector(3149620,23);
            logexp <= conv_std_logic_vector(133,8);
      WHEN others =>
           logman <= conv_std_logic_vector(0,23);
           logexp <= conv_std_logic_vector(0,8);
    END CASE;
  END PROCESS;

END rtl;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_LNNORM.VHD                             ***
--***                                             ***
--***   Function: Single Precision Normalization  ***
--***   of LN calculation                         ***
--***                                             ***
--***   22/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_lnnorm IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      inman : IN STD_LOGIC_VECTOR (32 DOWNTO 1);
      inexp : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      
      outman : OUT STD_LOGIC_VECTOR (24 DOWNTO 1);
      outexp : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
      zero : OUT STD_LOGIC
    );
END fp_lnnorm;

ARCHITECTURE rtl OF fp_lnnorm IS

  -- 3 latency
  
  signal shift, shiftff : STD_LOGIC_VECTOR (5 DOWNTO 1);
  signal zerochk : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal inmanff, inmandelff, outmanff : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal outmanbus : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal inexpff, expaddff, expsubff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal zeroff : STD_LOGIC_VECTOR (2 DOWNTO 1);

  component fp_lnclz
  PORT (
        mantissa : IN STD_LOGIC_VECTOR (32 DOWNTO 1);
        leading : OUT STD_LOGIC_VECTOR (5 DOWNTO 1)    
       );
  end component;
  
  component fp_lsft32x5
  PORT (
        inbus : IN STD_LOGIC_VECTOR (32 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (5 DOWNTO 1);
        outbus : OUT STD_LOGIC_VECTOR (32 DOWNTO 1)
      );
  end component;
             
BEGIN
  
  ppin: PROCESS (sysclk,reset)
  BEGIN
  
    IF (reset = '1') THEN
        
      FOR k IN 1 TO 32 LOOP
        inmanff(k) <= '0';
        inmandelff(k) <= '0';
        outmanff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 8 LOOP
        inexpff(k) <= '0';
        expaddff(k) <= '0';
        expsubff(k) <= '0';
      END LOOP;
      zeroff <= "00";
      shiftff <= "00000";
      
    ELSIF (rising_edge(sysclk)) THEN
        
      IF (enable = '1') THEN
          
        inmanff <= inman;
        inmandelff <= inmanff;
        outmanff <= outmanbus;
        
        inexpff <= inexp;
        -- add 2 - 1 for right shift to avoid overflow 
        expaddff <= inexpff + 1;
        expsubff <= expaddff - ("000" & shiftff);
        
        zeroff(1) <= zerochk(32);
        zeroff(2) <= zeroff(1);
      
        shiftff <= shift;
        
      END IF;
  
    END IF;
    
  END PROCESS;
  
  zerochk(1) <= inmanff(1);
  gza: FOR k IN 2 TO 32 GENERATE
    zerochk(k) <= zerochk(k-1) OR inmanff(k);
  END GENERATE;

  clz: fp_lnclz
  PORT MAP (mantissa=>inmanff,leading=>shift);
  
  sft: fp_lsft32x5
  PORT MAP (inbus=>inmandelff,shift=>shiftff,
            outbus=>outmanbus);

  --*** OUTPUTS ***
  outman <= outmanff(31 DOWNTO 8);
  outexp <= expsubff;
  zero <= zeroff(2);
      
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_LNRND.VHD                              ***
--***                                             ***
--***   Function: FP LOG Output Block - Rounded   ***
--***                                             ***
--***   22/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_lnrnd IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signln : IN STD_LOGIC;
      exponentln : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissaln : IN STD_LOGIC_VECTOR (24 DOWNTO 1);
      nanin : IN STD_LOGIC;
      infinityin : IN STD_LOGIC;
      zeroin : IN STD_LOGIC;
        
		signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
      --------------------------------------------------
      nanout : OUT STD_LOGIC;
      overflowout : OUT STD_LOGIC;
      zeroout : OUT STD_LOGIC
		);
END fp_lnrnd;

ARCHITECTURE rtl OF fp_lnrnd IS

  constant expwidth : positive := 8;
  constant manwidth : positive := 23;
  
  type exponentfftype IS ARRAY (2 DOWNTO 1) OF STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  
  signal zerovec : STD_LOGIC_VECTOR (manwidth-1 DOWNTO 1);
  signal nanff : STD_LOGIC_VECTOR (2 DOWNTO 1);
  signal zeroff : STD_LOGIC_VECTOR (2 DOWNTO 1);
  signal signff : STD_LOGIC_VECTOR (2 DOWNTO 1);
  signal infinityff : STD_LOGIC_VECTOR (2 DOWNTO 1);
  signal manoverflowbitff : STD_LOGIC; 
  signal roundmantissaff, mantissaff : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal exponentnode : STD_LOGIC_VECTOR (expwidth+2 DOWNTO 1);
  signal exponentoneff : STD_LOGIC_VECTOR (expwidth+2 DOWNTO 1);
  signal exponenttwoff : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
    
  signal manoverflow : STD_LOGIC_VECTOR (manwidth+1 DOWNTO 1);
  signal setmanzero, setmanmax : STD_LOGIC;
  signal setexpzero, setexpmax : STD_LOGIC;

BEGIN
    
  gzv: FOR k IN 1 TO manwidth-1 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  pra: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN
        
      nanff <= "00";
      signff <= "00";
      FOR k IN 1 TO manwidth LOOP
        roundmantissaff(k) <= '0';
        mantissaff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth+2 LOOP
        exponentoneff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        exponenttwoff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF(enable = '1') THEN 
      
        nanff(1) <= nanin;
        nanff(2) <= nanff(1);
        infinityff(1) <= infinityin;
        infinityff(2) <= infinityff(1);
        zeroff(1) <= zeroin;
        zeroff(2) <= zeroff(1);
        signff(1) <= signln;
        signff(2) <= signff(1);
       
        manoverflowbitff <= manoverflow(manwidth+1);
        
        roundmantissaff <= mantissaln(manwidth+1 DOWNTO 2) + (zerovec & mantissaln(1));
        
        FOR k IN 1 TO manwidth LOOP
          mantissaff(k) <= (roundmantissaff(k) AND NOT(setmanzero)) OR setmanmax;
        END LOOP;
        
        exponentoneff(expwidth+2 DOWNTO 1) <= "00" & exponentln;                 
        FOR k IN 1 TO expwidth LOOP
          exponenttwoff(k) <= (exponentnode(k) AND NOT(setexpzero)) OR setexpmax;
        END LOOP;
      
      END IF;
             
    END IF;
      
  END PROCESS;
  
  exponentnode <= exponentoneff(expwidth+2 DOWNTO 1) + 
                 (zerovec(expwidth+1 DOWNTO 1) & manoverflowbitff);

--*********************************
--*** PREDICT MANTISSA OVERFLOW ***   
--*********************************
     
  manoverflow(1) <= mantissaln(1);
  gmoa: FOR k IN 2 TO manwidth+1 GENERATE
    manoverflow(k) <= manoverflow(k-1) AND mantissaln(k);
  END GENERATE; 
                                                                 
--**********************************
--*** CHECK GENERATED CONDITIONS ***   
--**********************************

  -- all set to '1' when true
  
  -- set mantissa to 0 when infinity or zero condition
  setmanzero <= NOT(zeroff(1)) OR infinityff(1);
  -- setmantissa to "11..11" when nan
  setmanmax <= nanff(1);
  -- set exponent to 0 when zero condition 
  setexpzero <= NOT(zeroff(1));
  -- set exponent to "11..11" when nan or infinity
  setexpmax <= nanff(1) OR infinityff(1);
                             
--***************
--*** OUTPUTS ***
--***************
  
  signout <= signff(2);
  mantissaout <= mantissaff;
  exponentout <= exponenttwoff; 
  -----------------------------------------------
  nanout <= nanff(2);
  overflowout <= infinityff(2);
  zeroout <= zeroff(2);

END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   SINGLE PRECISION LOG(LN) - TOP LEVEL      ***
--***                                             ***
--***   FP_LOG.VHD                                ***
--***                                             ***
--***   Function: IEEE754 FP LOG()                ***
--***                                             ***
--***   21/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** Latency = 21                                ***
--***************************************************

ENTITY fp_log IS 
GENERIC (synthesize : integer := 1);
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (23 DOWNTO 1);

		  signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
      --------------------------------------------------
      nanout : OUT STD_LOGIC;
      overflowout : OUT STD_LOGIC;
      zeroout : OUT STD_LOGIC
		);
END fp_log;

ARCHITECTURE rtl OF fp_log IS
  
  constant expwidth : positive := 8;
  constant manwidth : positive := 23;
  
  constant coredepth : positive := 19;

  signal signinff : STD_LOGIC_VECTOR (2 DOWNTO 1);
  signal maninff : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal expinff : STD_LOGIC_VECTOR (expwidth DOWNTO 1);   
  signal signnode : STD_LOGIC;
  signal mantissanode : STD_LOGIC_VECTOR (24 DOWNTO 1);
  signal exponentnode : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal zeronode : STD_LOGIC;
              
  -- conditions
  signal zeroman : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal zeroexp : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal maxexp : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal zeromaninff : STD_LOGIC;
  signal zeroexpinff : STD_LOGIC;
  signal maxexpinff : STD_LOGIC;
  signal naninff : STD_LOGIC;
  signal nanff : STD_LOGIC_VECTOR (coredepth-3 DOWNTO 1);
  signal infinityinff : STD_LOGIC;
  signal infinityff : STD_LOGIC_VECTOR (coredepth-3 DOWNTO 1);
      
  component fp_ln_core 
  GENERIC (synthesize : integer := 1);
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aaman : IN STD_LOGIC_VECTOR (23 DOWNTO 1); 
        aaexp : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      
        ccman : OUT STD_LOGIC_VECTOR (24 DOWNTO 1);
        ccexp : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
        ccsgn : OUT STD_LOGIC;
        zeroout : OUT STD_LOGIC
       );
  end component;
  
  component fp_lnrnd
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        signln : IN STD_LOGIC;
        exponentln : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
        mantissaln : IN STD_LOGIC_VECTOR (24 DOWNTO 1);
        nanin : IN STD_LOGIC;
        infinityin : IN STD_LOGIC;
        zeroin : IN STD_LOGIC;

        signout : OUT STD_LOGIC;
        exponentout : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
        mantissaout : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
        --------------------------------------------------
        nanout : OUT STD_LOGIC;
        overflowout : OUT STD_LOGIC;
        zeroout : OUT STD_LOGIC
		  );
  end component;

BEGIN

  pma: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN

      FOR k IN 1 TO manwidth LOOP
        maninff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        expinff(k) <= '0';
      END LOOP;
      signinff <= "00";
    
    ELSIF (rising_edge(sysclk)) THEN

      IF (enable = '1') THEN

        maninff <= mantissain;
        expinff <= exponentin;
        signinff(1) <= signin;
        signinff(2) <= signinff(1);
                                                  
      END IF;
  
    END IF;
  
  END PROCESS;

--********************
--*** CHECK INPUTS ***
--********************

  zeroman(1) <= maninff(1);
  gca: FOR k IN 2 TO manwidth GENERATE
    zeroman(k) <= zeroman(k-1) OR maninff(k);
  END GENERATE; 
  zeroexp(1) <= expinff(1);
  gcb: FOR k IN 2 TO expwidth GENERATE
    zeroexp(k) <= zeroexp(k-1) OR expinff(k);
  END GENERATE;
  maxexp(1) <= expinff(1);
  gcc: FOR k IN 2 TO expwidth GENERATE
    maxexp(k) <= maxexp(k-1) AND expinff(k);
  END GENERATE;

  pcc: PROCESS (sysclk,reset)
  BEGIN
    
    IF (reset = '1') THEN
      
      zeromaninff <= '0';
      zeroexpinff <= '0';
      maxexpinff <= '0';  
      naninff <= '0';
      FOR k IN 1 TO coredepth-3 LOOP
        nanff(k) <= '0';
      END LOOP;
     
    ELSIF (rising_edge(sysclk)) THEN
            
      IF (enable = '1') THEN

        zeromaninff <= NOT(zeroman(manwidth));
        zeroexpinff <= NOT(zeroexp(expwidth));
        maxexpinff <= maxexp(expwidth);
    
        -- infinity when exp = zero
        -- nan when man != 0, exp = max
    
        -- all ffs '1' when condition true
        naninff <= (zeromaninff AND maxexpinff) OR signinff(2);
        infinityinff <= zeroexpinff OR maxexpinff;

        -- nan output when nan input
        nanff(1) <= naninff;
        FOR k IN 2 TO coredepth-3 LOOP
          nanff(k) <= nanff(k-1);
        END LOOP;
        
        infinityff(1) <= infinityinff;
        FOR k IN 2 TO coredepth-3 LOOP
          infinityff(k) <= infinityff(k-1);
        END LOOP;
      
      END IF;
   
    END IF;

  END PROCESS;


--***************
--*** LN CORE ***
--***************

  lncore: fp_ln_core
  GENERIC MAP (synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aaman=>mantissain,aaexp=>exponentin,
            ccman=>mantissanode,ccexp=>exponentnode,ccsgn=>signnode,
            zeroout=>zeronode);
  
--************************
--*** ROUND AND OUTPUT ***
--************************

    rndout: fp_lnrnd
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              signln=>signnode,
              exponentln=>exponentnode,
              mantissaln=>mantissanode,
              nanin=>nanff(coredepth-3),
              infinityin=>infinityff(coredepth-3),
              zeroin=>zeronode,

              signout=>signout,
              exponentout=>exponentout,
              mantissaout=>mantissaout,
              nanout=>nanout,overflowout=>overflowout,zeroout=>zeroout);

END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_LSFT23.VHD                             ***
--***                                             ***
--***   Function: 23 bit Left Shift               ***
--***                                             ***
--***   22/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_lsft23 IS 
PORT (
      inbus : IN STD_LOGIC_VECTOR (23 DOWNTO 1);
      shift : IN STD_LOGIC_VECTOR (5 DOWNTO 1);

	   outbus : OUT STD_LOGIC_VECTOR (23 DOWNTO 1)
	  );
END fp_lsft23;

ARCHITECTURE sft OF fp_lsft23 IS
  
  signal levzip, levone, levtwo, levthr : STD_LOGIC_VECTOR (23 DOWNTO 1);
    
BEGIN
        
  levzip <= inbus;
  
  -- shift by 0,1,2,3
  levone(1) <=  (levzip(1) AND NOT(shift(2)) AND NOT(shift(1)));
  levone(2) <=  (levzip(2) AND NOT(shift(2)) AND NOT(shift(1))) OR
                (levzip(1) AND NOT(shift(2)) AND     shift(1));
  levone(3) <=  (levzip(3) AND NOT(shift(2)) AND NOT(shift(1))) OR
                (levzip(2) AND NOT(shift(2)) AND     shift(1)) OR
                (levzip(1) AND     shift(2)  AND NOT(shift(1))); 
  gaa: FOR k IN 4 TO 23 GENERATE
    levone(k) <= (levzip(k)   AND NOT(shift(2)) AND NOT(shift(1))) OR
                 (levzip(k-1) AND NOT(shift(2)) AND     shift(1)) OR
                 (levzip(k-2) AND     shift(2)  AND NOT(shift(1))) OR
                 (levzip(k-3) AND     shift(2)  AND     shift(1)); 
  END GENERATE;

  -- shift by 0,4,8,12
  gba: FOR k IN 1 TO 4 GENERATE
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3)));
  END GENERATE;
  gbb: FOR k IN 5 TO 8 GENERATE
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                 (levone(k-4)  AND NOT(shift(4)) AND     shift(3));
  END GENERATE;
  gbc: FOR k IN 9 TO 12 GENERATE
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                 (levone(k-4)  AND NOT(shift(4)) AND     shift(3)) OR
                 (levone(k-8)  AND     shift(4)  AND NOT(shift(3)));
  END GENERATE;
  gbd: FOR k IN 13 TO 23 GENERATE
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                 (levone(k-4)  AND NOT(shift(4)) AND     shift(3)) OR
                 (levone(k-8)  AND     shift(4)  AND NOT(shift(3))) OR
                 (levone(k-12) AND     shift(4)  AND     shift(3)); 
  END GENERATE;

  gca: FOR k IN 1 TO 16 GENERATE
    levthr(k) <= (levtwo(k)    AND NOT(shift(5)));
  END GENERATE;
  gcb: FOR k IN 17 TO 23 GENERATE
    levthr(k) <= (levtwo(k)    AND NOT(shift(5))) OR
                 (levtwo(k-16) AND     shift(5));
  END GENERATE;

  outbus <= levthr;
  
END sft;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_LSFT32X5.VHD                           ***
--***                                             ***
--***   Function: Single Precision Left Shift     ***
--***                                             ***
--***   22/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_lsft32x5 IS 
PORT (
      inbus : IN STD_LOGIC_VECTOR (32 DOWNTO 1);
      shift : IN STD_LOGIC_VECTOR (5 DOWNTO 1);
      outbus : OUT STD_LOGIC_VECTOR (32 DOWNTO 1)
    );
END fp_lsft32x5;

ARCHITECTURE rtl OF fp_lsft32x5 IS

  signal leftone, lefttwo, leftthr : STD_LOGIC_VECTOR (32 DOWNTO 1);
            
BEGIN
  
  leftone(1) <=  inbus(1)     AND NOT(shift(2)) AND NOT(shift(1));
  leftone(2) <= (inbus(2)     AND NOT(shift(2)) AND NOT(shift(1))) OR
                (inbus(1)     AND NOT(shift(2)) AND     shift(1)); 
  leftone(3) <= (inbus(3)     AND NOT(shift(2)) AND NOT(shift(1))) OR
                (inbus(2)     AND NOT(shift(2)) AND     shift(1)) OR
                (inbus(1)     AND     shift(2)  AND NOT(shift(1))); 
  gla: FOR k IN 4 TO 32 GENERATE
    leftone(k) <= (inbus(k)   AND NOT(shift(2)) AND NOT(shift(1))) OR
                  (inbus(k-1) AND NOT(shift(2)) AND     shift(1)) OR
                  (inbus(k-2) AND     shift(2)  AND NOT(shift(1))) OR
                  (inbus(k-3) AND     shift(2)  AND     shift(1));
  END GENERATE;
             
  glb: FOR k IN 1 TO 4 GENERATE
    lefttwo(k) <=  leftone(k)    AND NOT(shift(4)) AND NOT(shift(3));
  END GENERATE;
  glc: FOR k IN 5 TO 8 GENERATE
    lefttwo(k) <= (leftone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                  (leftone(k-4)  AND NOT(shift(4)) AND     shift(3)); 
  END GENERATE;
  gld: FOR k IN 9 TO 12 GENERATE
    lefttwo(k) <= (leftone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                  (leftone(k-4)  AND NOT(shift(4)) AND     shift(3)) OR
                  (leftone(k-8)  AND     shift(4)  AND NOT(shift(3))); 
  END GENERATE;
  gle: FOR k IN 13 TO 32 GENERATE
    lefttwo(k) <= (leftone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                  (leftone(k-4)  AND NOT(shift(4)) AND     shift(3)) OR
                  (leftone(k-8)  AND     shift(4)  AND NOT(shift(3)))  OR
                  (leftone(k-12) AND     shift(4)  AND     shift(3)); 
  END GENERATE;
  
  glf: FOR k IN 1 TO 16 GENERATE
    leftthr(k) <=  lefttwo(k)    AND NOT(shift(5));
  END GENERATE;
  glg: FOR k IN 17 TO 32 GENERATE
    leftthr(k) <= (lefttwo(k)    AND NOT(shift(5))) OR
                  (lefttwo(k-16) AND     shift(5)); 
  END GENERATE;
    
  outbus <= leftthr;        
            
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_LSFT36.VHD                             ***
--***                                             ***
--***   Function: 36 bit Left Shift               ***
--***                                             ***
--***   22/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_lsft36 IS 
PORT (
      inbus : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
      shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);

	    outbus : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
	   );
END fp_lsft36;

ARCHITECTURE sft OF fp_lsft36 IS
  
  signal levzip, levone, levtwo, levthr : STD_LOGIC_VECTOR (36 DOWNTO 1);
    
BEGIN
        
  levzip <= inbus;
  
  -- shift by 0,1,2,3
  levone(1) <=  (levzip(1) AND NOT(shift(2)) AND NOT(shift(1)));
  levone(2) <=  (levzip(2) AND NOT(shift(2)) AND NOT(shift(1))) OR
                (levzip(1) AND NOT(shift(2)) AND     shift(1));
  levone(3) <=  (levzip(3) AND NOT(shift(2)) AND NOT(shift(1))) OR
                (levzip(2) AND NOT(shift(2)) AND     shift(1)) OR
                (levzip(1) AND     shift(2)  AND NOT(shift(1))); 
  gaa: FOR k IN 4 TO 36 GENERATE
    levone(k) <= (levzip(k)   AND NOT(shift(2)) AND NOT(shift(1))) OR
                 (levzip(k-1) AND NOT(shift(2)) AND     shift(1)) OR
                 (levzip(k-2) AND     shift(2)  AND NOT(shift(1))) OR
                 (levzip(k-3) AND     shift(2)  AND     shift(1)); 
  END GENERATE;

  -- shift by 0,4,8,12
  gba: FOR k IN 1 TO 4 GENERATE
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3)));
  END GENERATE;
  gbb: FOR k IN 5 TO 8 GENERATE
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                 (levone(k-4)  AND NOT(shift(4)) AND     shift(3));
  END GENERATE;
  gbc: FOR k IN 9 TO 12 GENERATE
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                 (levone(k-4)  AND NOT(shift(4)) AND     shift(3)) OR
                 (levone(k-8)  AND     shift(4)  AND NOT(shift(3)));
  END GENERATE;
  gbd: FOR k IN 13 TO 36 GENERATE
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                 (levone(k-4)  AND NOT(shift(4)) AND     shift(3)) OR
                 (levone(k-8)  AND     shift(4)  AND NOT(shift(3))) OR
                 (levone(k-12) AND     shift(4)  AND     shift(3)); 
  END GENERATE;

  -- shift by 0,16,32
  gca: FOR k IN 1 TO 16 GENERATE
    levthr(k) <= (levtwo(k)    AND NOT(shift(6)) AND NOT(shift(5)));
  END GENERATE;
  gcb: FOR k IN 17 TO 32 GENERATE
    levthr(k) <= (levtwo(k)    AND NOT(shift(6)) AND NOT(shift(5))) OR
                 (levtwo(k-16) AND NOT(shift(6)) AND     shift(5));
  END GENERATE;
  gcc: FOR k IN 33 TO 36 GENERATE
    levthr(k) <= (levtwo(k)    AND NOT(shift(6)) AND NOT(shift(5))) OR
                 (levtwo(k-16) AND NOT(shift(6)) AND     shift(5)) OR
                 (levtwo(k-32) AND     shift(6)  AND NOT(shift(5)));
  END GENERATE;

  outbus <= levthr;
  
END sft;

LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_LSFT78.VHD                             ***
--***                                             ***
--***   Function: 78 bit Left Shift               ***
--***                                             ***
--***   22/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_lsft78 IS
PORT (
      inbus : IN STD_LOGIC_VECTOR (78 DOWNTO 1); 
      shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1); 

      outbus : OUT STD_LOGIC_VECTOR (78 DOWNTO 1)
     );
END fp_lsft78;

ARCHITECTURE rtl of fp_lsft78 IS

  signal levzip, levone, levtwo : STD_LOGIC_VECTOR (78 DOWNTO 1);
  signal levthr, levfor, levfiv : STD_LOGIC_VECTOR (78 DOWNTO 1);
  signal levsix : STD_LOGIC_VECTOR (78 DOWNTO 1);
  
BEGIN

  levzip <= inbus;
  
  levone(1) <= levzip(1) AND NOT(shift(1));
  gaa: FOR k IN 2 TO 78 GENERATE
    levone(k) <= (levzip(k) AND NOT(shift(1))) OR (levzip(k-1) AND shift(1));
  END GENERATE;
  
  levtwo(1) <= levone(1) AND NOT(shift(2));
  levtwo(2) <= levone(2) AND NOT(shift(2));
  gba: FOR k IN 3 TO 78 GENERATE
    levtwo(k) <= (levone(k) AND NOT(shift(2))) OR (levone(k-2) AND shift(2));
  END GENERATE;
  
  gca: FOR k IN 1 TO 4 GENERATE
    levthr(k) <= levtwo(k) AND NOT(shift(3));
  END GENERATE;
  gcb: FOR k IN 5 TO 78 GENERATE
    levthr(k) <= (levtwo(k) AND NOT(shift(3))) OR (levtwo(k-4) AND shift(3));
  END GENERATE;
  
  gda: FOR k IN 1 TO 8 GENERATE
    levfor(k) <= levthr(k) AND NOT(shift(4));
  END GENERATE;
  gdb: FOR k IN 9 TO 78 GENERATE
    levfor(k) <= (levthr(k) AND NOT(shift(4))) OR (levthr(k-8) AND shift(4));
  END GENERATE;
  
  gea: FOR k IN 1 TO 16 GENERATE
    levfiv(k) <= levfor(k) AND NOT(shift(5));
  END GENERATE;
  geb: FOR k IN 17 TO 78 GENERATE
    levfiv(k) <= (levfor(k) AND NOT(shift(5))) OR (levfor(k-16) AND shift(5));
  END GENERATE;
  
  gfa: FOR k IN 1 TO 32 GENERATE
    levsix(k) <= levfiv(k) AND NOT(shift(6));
  END GENERATE;
  gfb: FOR k IN 33 TO 78 GENERATE
    levsix(k) <= (levfiv(k) AND NOT(shift(6))) OR (levfiv(k-32) AND shift(6));
  END GENERATE;
  
  outbus <= levsix;
  
END;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

LIBRARY altera_mf;
USE altera_mf.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_MUL23X56.VHD                           ***
--***                                             ***
--***   Function: Fixed Point Multiplier          ***
--***                                             ***
--***   23 and 56 bit inputs, 4 pipes             ***
--***                                             ***
--***   07/01/10 ML                               ***
--***                                             ***
--***   (c) 2010 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_mul23x56 IS
GENERIC (device : integer := 0);
PORT
	(
    sysclk : IN STD_LOGIC;
    reset : IN STD_LOGIC;
    enable : IN STD_LOGIC;
    dataaa : IN STD_LOGIC_VECTOR (23 DOWNTO 1);
    databb : IN STD_LOGIC_VECTOR (56 DOWNTO 1);

	 result : OUT STD_LOGIC_VECTOR (79 DOWNTO 1)
	);
END fp_mul23x56;

ARCHITECTURE SYN OF fp_mul23x56 IS
  constant AW : integer := 23;
  constant BW : integer := 56;
  constant RW : integer := AW+BW;
  
  -- use 27-bit multipliers on SV/AV/CV,
  -- use 36-bit multipliers on SIII/SIV
  -- split multiplication into two equal parts on other architectures
  function chooseMaxMulWidth(device : integer) return integer is
  begin
    if (device = 2) then
      return 27;
    elsif (device = 1) then
      return 36;
    else
      return 28;
    end if;
  end function;

  constant MAXMULWIDTH : integer := chooseMaxMulWidth(device);
  constant use_2_multipliers : boolean := BW <= 2 * MAXMULWIDTH;
  constant use_3_multipliers : boolean := not use_2_multipliers;
  
  component fp_mul2s
  GENERIC (
    widthaa : positive;
    widthbb : positive;
    widthcc : positive
  );
  PORT (
    sysclk : IN STD_LOGIC;
    reset : IN STD_LOGIC;
    enable : IN STD_LOGIC;
    dataaa : IN STD_LOGIC_VECTOR(widthaa DOWNTO 1);
    databb : IN STD_LOGIC_VECTOR(widthbb DOWNTO 1);

    result : OUT STD_LOGIC_VECTOR(widthcc DOWNTO 1)
  );
  end component;

  component fp_mul3s
  GENERIC (
    widthaa : positive;
    widthbb : positive;
    widthcc : positive
  );
  PORT (
    sysclk : IN STD_LOGIC;
    reset : IN STD_LOGIC;
    enable : IN STD_LOGIC;
    dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
    databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1);

    result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
  );
  end component; 

  signal zerovec : STD_LOGIC_VECTOR(MAXMULWIDTH DOWNTO 1);
BEGIN
  zerovec <= (others => '0');

gen2mul: IF use_2_multipliers GENERATE
  constant BLW : integer := MAXMULWIDTH;
  constant BHW : integer := BW - BLW;
  signal multiplier_low  : STD_LOGIC_VECTOR(BLW+AW DOWNTO 1);
  signal multiplier_high : STD_LOGIC_VECTOR(BHW+AW DOWNTO 1);
  signal adderff  : STD_LOGIC_VECTOR(RW DOWNTO 1);
BEGIN
  ml: fp_mul3s
  GENERIC MAP (widthaa=>AW,widthbb=>BLW,widthcc=>BLW+AW)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>dataaa,databb=>databb(BLW DOWNTO 1),
            result=>multiplier_low);

  mh: fp_mul3s
  GENERIC MAP (widthaa=>AW,widthbb=>BHW,widthcc=>BHW+AW)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>dataaa,databb=>databb(BHW+BLW DOWNTO BLW+1),
            result=>multiplier_high);

  pad: PROCESS (sysclk,reset)
  BEGIN
    IF (reset = '1') THEN
        adderff <= (others => '0');
    ELSIF (rising_edge(sysclk)) THEN
      IF (enable = '1') THEN
        adderff <= (zerovec(RW-(BLW+AW) DOWNTO 1) & multiplier_low) +
                   (multiplier_high & zerovec(RW-(BHW+AW) DOWNTO 1));
      END IF;
    END IF;
  END PROCESS;

  result <= adderff;
END GENERATE;

gen3mul: IF use_3_multipliers GENERATE
  constant BLW : integer := MAXMULWIDTH;
  constant BHW : integer := MAXMULWIDTH;
  constant BTW : integer := BW - BLW - BHW;
  signal multiplier_low :  STD_LOGIC_VECTOR(BLW+AW DOWNTO 1);
  signal multiplier_high : STD_LOGIC_VECTOR(BHW+AW DOWNTO 1);
  signal multiplier_top :  STD_LOGIC_VECTOR(BTW+AW DOWNTO 1);
  signal adderff0 : STD_LOGIC_VECTOR (RW DOWNTO 1);
  signal adderff1 : STD_LOGIC_VECTOR (RW DOWNTO 1);
BEGIN
  ml: fp_mul2s
  GENERIC MAP (widthaa=>AW,widthbb=>BLW,widthcc=>BLW+AW)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>dataaa,databb=>databb(BLW DOWNTO 1),
            result=>multiplier_low);

  mh: fp_mul2s
  GENERIC MAP (widthaa=>AW,widthbb=>BHW,widthcc=>BHW+AW)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>dataaa,databb=>databb(BHW+BLW DOWNTO BLW+1),
            result=>multiplier_high);

  mt: fp_mul2s
  GENERIC MAP (widthaa=>AW,widthbb=>BTW,widthcc=>BTW+AW)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>dataaa,databb=>databb(BTW+BHW+BLW DOWNTO BHW+BLW+1),
            result=>multiplier_top);

  pad: PROCESS (sysclk,reset)
  BEGIN
    IF (reset = '1') THEN
        adderff0 <= (others => '0');
        adderff1 <= (others => '0');
    ELSIF (rising_edge(sysclk)) THEN
      IF (enable = '1') THEN
        adderff0 <= (multiplier_top & zerovec(RW-(BTW+AW)-(BLW+AW) DOWNTO 1) & multiplier_low) +
                    (zerovec(RW-(BHW+AW)-BLW DOWNTO 1) & multiplier_high & zerovec(BLW DOWNTO 1));
        adderff1 <= adderff0;
      END IF;
    END IF;
  END PROCESS;

  result <= adderff1;
END GENERATE;

END SYN;


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_MUL2S.VHD                              ***
--***                                             ***
--***   Function: Fixed Point Multiplier          ***
--***                                             ***
--***   18-36 bit inputs, 2 pipes                 ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_mul2s IS
GENERIC (
         widthaa : positive := 18;
         widthbb : positive := 18;
         widthcc : positive := 36
        );
PORT
	(
    sysclk : IN STD_LOGIC;
    reset : IN STD_LOGIC;
    enable : IN STD_LOGIC;
    dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
    databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1);

	 result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
	);
END fp_mul2s;

ARCHITECTURE SYN OF fp_mul2s IS

	SIGNAL resultnode	: STD_LOGIC_VECTOR (widthaa+widthbb DOWNTO 1);

	COMPONENT altmult_add
	GENERIC (
		addnsub_multiplier_aclr1		: STRING;
		addnsub_multiplier_pipeline_aclr1		: STRING;
		addnsub_multiplier_pipeline_register1		: STRING;
		addnsub_multiplier_register1		: STRING;
		dedicated_multiplier_circuitry		: STRING;
		input_aclr_a0		: STRING;
		input_aclr_b0		: STRING;
		input_register_a0		: STRING;
		input_register_b0		: STRING;
		input_source_a0		: STRING;
		input_source_b0		: STRING;
		intended_device_family		: STRING;
		lpm_type		: STRING;
		multiplier1_direction		: STRING;
		multiplier_aclr0		: STRING;
		multiplier_register0		: STRING;
		number_of_multipliers		: NATURAL;
		output_register		: STRING;
		port_addnsub1		: STRING;
		port_signa		: STRING;
		port_signb		: STRING;
		representation_a		: STRING;
		representation_b		: STRING;
		signed_aclr_a		: STRING;
		signed_aclr_b		: STRING;
		signed_pipeline_aclr_a		: STRING;
		signed_pipeline_aclr_b		: STRING;
		signed_pipeline_register_a		: STRING;
		signed_pipeline_register_b		: STRING;
		signed_register_a		: STRING;
		signed_register_b		: STRING;
		width_a		: NATURAL;
		width_b		: NATURAL;
		width_result		: NATURAL
	);
	PORT (
			dataa	: IN STD_LOGIC_VECTOR (widthaa-1 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (widthbb-1 DOWNTO 0);
			clock0	: IN STD_LOGIC ;
			aclr3	: IN STD_LOGIC ;
			ena0	: IN STD_LOGIC ;
			result	: OUT STD_LOGIC_VECTOR (widthaa+widthbb-1 DOWNTO 0)
	);
	END COMPONENT;

BEGIN

	ALTMULT_ADD_component : altmult_add
	GENERIC MAP (
		addnsub_multiplier_aclr1 => "ACLR3",
		addnsub_multiplier_pipeline_aclr1 => "ACLR3",
		addnsub_multiplier_pipeline_register1 => "CLOCK0",
		addnsub_multiplier_register1 => "CLOCK0",
		dedicated_multiplier_circuitry => "AUTO",
		input_aclr_a0 => "ACLR3",
		input_aclr_b0 => "ACLR3",
		input_register_a0 => "CLOCK0",
		input_register_b0 => "CLOCK0",
		input_source_a0 => "DATAA",
		input_source_b0 => "DATAB",
		intended_device_family => "Stratix",
		lpm_type => "altmult_add",
		multiplier1_direction => "ADD",
		multiplier_aclr0 => "ACLR3",
		multiplier_register0 => "CLOCK0",
		number_of_multipliers => 1,
		output_register => "UNREGISTERED",
		port_addnsub1 => "PORT_UNUSED",
		port_signa => "PORT_UNUSED",
		port_signb => "PORT_UNUSED",
		representation_a => "UNSIGNED",
		representation_b => "UNSIGNED",
		signed_aclr_a => "ACLR3",
		signed_aclr_b => "ACLR3",
		signed_pipeline_aclr_a => "ACLR3",
		signed_pipeline_aclr_b => "ACLR3",
		signed_pipeline_register_a => "CLOCK0",
		signed_pipeline_register_b => "CLOCK0",
		signed_register_a => "CLOCK0",
		signed_register_b => "CLOCK0",
		width_a => widthaa,
		width_b => widthbb,
		width_result => widthaa+widthbb
	)
	PORT MAP (
		dataa => dataaa,
		datab => databb,
		clock0 => sysclk,
		aclr3 => reset,
		ena0 => enable,
		result => resultnode
	);

  result <= resultnode(widthaa+widthbb DOWNTO widthaa+widthbb-widthcc+1);
  
END SYN;

LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_MUL3S.VHD                              ***
--***                                             ***
--***   Function: Fixed Point Multiplier          ***
--***                                             ***
--***   18-36 bit inputs, 3 pipes                 ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_mul3s IS
GENERIC (
         widthaa : positive := 18;
         widthbb : positive := 18;
         widthcc : positive := 36
        );
PORT
	(
    sysclk : IN STD_LOGIC;
    reset : IN STD_LOGIC;
    enable : IN STD_LOGIC;
    dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
    databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1);

	 result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
	);
END fp_mul3s;

ARCHITECTURE SYN OF fp_mul3s IS

	SIGNAL resultnode	: STD_LOGIC_VECTOR (widthaa+widthbb DOWNTO 1);

  component altmult_add
	GENERIC (
		addnsub_multiplier_aclr1		: STRING;
		addnsub_multiplier_pipeline_aclr1		: STRING;
		addnsub_multiplier_pipeline_register1		: STRING;
		addnsub_multiplier_register1		: STRING;
		dedicated_multiplier_circuitry		: STRING;
		input_aclr_a0		: STRING;
		input_aclr_b0		: STRING;
		input_register_a0		: STRING;
		input_register_b0		: STRING;
		input_source_a0		: STRING;
		input_source_b0		: STRING;
		intended_device_family		: STRING;
		lpm_type		: STRING;
		multiplier1_direction		: STRING;
		multiplier_aclr0		: STRING;
		multiplier_register0		: STRING;
		number_of_multipliers		: NATURAL;
		output_aclr		: STRING;
		output_register		: STRING;
		port_addnsub1		: STRING;
		port_signa		: STRING;
		port_signb		: STRING;
		representation_a		: STRING;
		representation_b		: STRING;
		signed_aclr_a		: STRING;
		signed_aclr_b		: STRING;
		signed_pipeline_aclr_a		: STRING;
		signed_pipeline_aclr_b		: STRING;
		signed_pipeline_register_a		: STRING;
		signed_pipeline_register_b		: STRING;
		signed_register_a		: STRING;
		signed_register_b		: STRING;
		width_a		: NATURAL;
		width_b		: NATURAL;
		width_result		: NATURAL
	);
	PORT (
			dataa	: IN STD_LOGIC_VECTOR (widthaa-1 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (widthbb-1 DOWNTO 0);
			clock0	: IN STD_LOGIC ;
			aclr3	: IN STD_LOGIC ;
			ena0	: IN STD_LOGIC ;
			result	: OUT STD_LOGIC_VECTOR (widthaa+widthbb-1 DOWNTO 0)
	);
	end component;

BEGIN

  mulone : altmult_add
  GENERIC MAP (
		addnsub_multiplier_aclr1 => "ACLR3",
		addnsub_multiplier_pipeline_aclr1 => "ACLR3",
		addnsub_multiplier_pipeline_register1 => "CLOCK0",
		addnsub_multiplier_register1 => "CLOCK0",
		dedicated_multiplier_circuitry => "AUTO",
		input_aclr_a0 => "ACLR3",
		input_aclr_b0 => "ACLR3",
		input_register_a0 => "CLOCK0",
		input_register_b0 => "CLOCK0",
		input_source_a0 => "DATAA",
		input_source_b0 => "DATAB",
		intended_device_family => "Stratix II",
		lpm_type => "altmult_add",
		multiplier1_direction => "ADD",
		multiplier_aclr0 => "ACLR3",
		multiplier_register0 => "CLOCK0",
		number_of_multipliers => 1,
		output_aclr => "ACLR3",
		output_register => "CLOCK0",
		port_addnsub1 => "PORT_UNUSED",
		port_signa => "PORT_UNUSED",
		port_signb => "PORT_UNUSED",
		representation_a => "UNSIGNED",
		representation_b => "UNSIGNED",
		signed_aclr_a => "ACLR3",
		signed_aclr_b => "ACLR3",
		signed_pipeline_aclr_a => "ACLR3",
		signed_pipeline_aclr_b => "ACLR3",
		signed_pipeline_register_a => "CLOCK0",
		signed_pipeline_register_b => "CLOCK0",
		signed_register_a => "CLOCK0",
		signed_register_b => "CLOCK0",
		width_a => widthaa,
		width_b => widthbb,
		width_result => widthaa+widthbb
	)
	PORT MAP (
		dataa => dataaa,
		datab => databb,
		clock0 => sysclk,
		aclr3 => reset,
		ena0 => enable,
		result => resultnode
	);

  result <= resultnode(widthaa+widthbb DOWNTO widthaa+widthbb-widthcc+1);
  
END SYN;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_MUL5418S.VHD                           ***
--***                                             ***
--***   Function: Fixed Point Multiplier          ***
--***   54x18=54, 3 18x18 architecture,           ***
--***   Stratix II/III, 3 or 4 pipeline,          ***
--***   synthesizable                             ***
--***                                             ***
--***   09/12/07 ML                               ***
--***                                             ***
--***   (c) 2007 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***   15/01/08 - outputs up to 72 bits now      ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_mul5418s IS 
GENERIC (
         widthcc : positive := 36;
         pipes : positive := 3  --3/4
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      dataaa : IN STD_LOGIC_VECTOR (54 DOWNTO 1);
      databb : IN STD_LOGIC_VECTOR (18 DOWNTO 1);
      
		result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
		);
END fp_mul5418s;

ARCHITECTURE rtl OF fp_mul5418s IS

  signal zerovec : STD_LOGIC_VECTOR (18 DOWNTO 1);

  signal muloneout, multwoout, multhrout : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal aavec, bbvec : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal resultnode : STD_LOGIC_VECTOR (72 DOWNTO 1);
  signal lowff, lowdelff : STD_LOGIC_VECTOR (18 DOWNTO 1);
  
  component dp_fxadd IS 
  GENERIC (
           width : positive := 64;
           pipes : positive := 1;
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
        carryin : IN STD_LOGIC;
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
  end component;

  component fp_mul2s IS
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36
          );
  PORT (  
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1);

	     result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
	    ); 
  end component;
  
BEGIN
  
  gza: FOR k IN 1 TO 18 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  mulone: fp_mul2s
  GENERIC MAP (widthaa=>18,widthbb=>18,widthcc=>36)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>dataaa(18 DOWNTO 1),databb=>databb(18 DOWNTO 1),
            result=>muloneout);
            
  multwo: fp_mul2s
  GENERIC MAP (widthaa=>18,widthbb=>18,widthcc=>36)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>dataaa(36 DOWNTO 19),databb=>databb(18 DOWNTO 1),
            result=>multwoout);
            
  multhr: fp_mul2s
  GENERIC MAP (widthaa=>18,widthbb=>18,widthcc=>36)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>dataaa(54 DOWNTO 37),databb=>databb(18 DOWNTO 1),
            result=>multhrout);
  
  aavec <= multhrout & muloneout(36 DOWNTO 19);
  bbvec <= zerovec(18 DOWNTO 1) & multwoout;
  
  adder: dp_fxadd
  GENERIC MAP (width=>54,pipes=>pipes-2,synthesize=>1)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            aa=>aavec,bb=>bbvec,carryin=>'0',
            cc=>resultnode(72 DOWNTO 19));
            
  gda: IF (pipes = 3) GENERATE  
         
    pda: PROCESS (sysclk,reset)
    BEGIN
    
      IF (reset = '1') THEN
        FOR k IN 1 TO 18 LOOP
          lowff(k) <= '0';
        END LOOP;
      ELSIF (rising_edge(sysclk)) THEN
        IF (enable = '1') THEN
          lowff <= muloneout(18 DOWNTO 1);
        END IF;
      END IF;
      
    END PROCESS;
    
    resultnode(18 DOWNTO 1) <= lowff;
    
  END GENERATE;

  gdb: IF (pipes = 4) GENERATE  
         
    pdb: PROCESS (sysclk,reset)
    BEGIN
    
      IF (reset = '1') THEN
        FOR k IN 1 TO 18 LOOP
          lowff(k) <= '0';
          lowdelff(k) <= '0';
        END LOOP;
      ELSIF (rising_edge(sysclk)) THEN
        IF (enable = '1') THEN
          lowff <= muloneout(18 DOWNTO 1);
          lowdelff <= lowff;
        END IF;
      END IF;
      
    END PROCESS;
    
    resultnode(18 DOWNTO 1) <= lowdelff;
    
  END GENERATE;
  
  result <= resultnode(72 DOWNTO 73-widthcc);
              
END rtl;


LIBRARY ieee;
LIBRARY work;
LIBRARY lpm;
LIBRARY altera_mf;
USE lpm.all;
USE altera_mf.all;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   ALTERA FLOATING POINT DATAPATH COMPILER   ***
--***                                             ***
--***   FP_MUL54US_28S.VHD                        ***
--***                                             ***
--***   Function: 5/6 pipeline stage unsigned 54  ***
--***   bit multiplier                            ***
--***   28S: Stratix 2, 8 18x18, synthesizeable   ***
--***                                             ***
--***   21/04/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** 1. Identical to HCC_MUL54US_28S, except 5   ***
--*** or 6 pipeline parameter and 72 outputs      ***
--***************************************************

ENTITY fp_mul54us_28s IS
GENERIC (latency : positive := 5);
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      mulaa, mulbb : IN STD_LOGIC_VECTOR (54 DOWNTO 1);      

      mulcc : OUT STD_LOGIC_VECTOR (72 DOWNTO 1)  
     );
END fp_mul54us_28s;

ARCHITECTURE syn of fp_mul54us_28s IS

  signal muloneaa, mulonebb : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal multwoaa, multwobb, multhraa, multhrbb : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal mulforaa, mulforbb, mulfivaa, mulfivbb : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal muloneout : STD_LOGIC_VECTOR (72 DOWNTO 1);
  signal multwoout, multhrout, mulforout, mulfivout : STD_LOGIC_VECTOR (36 DOWNTO 1);

  signal vecone, vectwo, vecthr, vecfor, vecfiv : STD_LOGIC_VECTOR (58 DOWNTO 1);
  signal vecsix, vecsev : STD_LOGIC_VECTOR (58 DOWNTO 1);
  signal vecegt, vecnin, vecten : STD_LOGIC_VECTOR (72 DOWNTO 1);
  signal sumvecone, carvecone : STD_LOGIC_VECTOR (58 DOWNTO 1);
  signal sumvectwo, carvectwo : STD_LOGIC_VECTOR (58 DOWNTO 1);
  signal sumvecthr, carvecthr : STD_LOGIC_VECTOR (72 DOWNTO 1);
  signal sumoneff, caroneff : STD_LOGIC_VECTOR (58 DOWNTO 1);
  signal sumtwoff, cartwoff : STD_LOGIC_VECTOR (72 DOWNTO 1);
  signal resultnode : STD_LOGIC_VECTOR (72 DOWNTO 1);
  
  signal zerovec : STD_LOGIC_VECTOR (36 DOWNTO 1);

  component altmult_add
	GENERIC (
		addnsub_multiplier_aclr1		: STRING;
		addnsub_multiplier_pipeline_aclr1		: STRING;
		addnsub_multiplier_pipeline_register1		: STRING;
		addnsub_multiplier_register1		: STRING;
		dedicated_multiplier_circuitry		: STRING;
		input_aclr_a0		: STRING;
		input_aclr_b0		: STRING;
		input_register_a0		: STRING;
		input_register_b0		: STRING;
		input_source_a0		: STRING;
		input_source_b0		: STRING;
		intended_device_family		: STRING;
		lpm_type		: STRING;
		multiplier1_direction		: STRING;
		multiplier_aclr0		: STRING;
		multiplier_register0		: STRING;
		number_of_multipliers		: NATURAL;
		output_aclr		: STRING;
		output_register		: STRING;
		port_addnsub1		: STRING;
		port_signa		: STRING;
		port_signb		: STRING;
		representation_a		: STRING;
		representation_b		: STRING;
		signed_aclr_a		: STRING;
		signed_aclr_b		: STRING;
		signed_pipeline_aclr_a		: STRING;
		signed_pipeline_aclr_b		: STRING;
		signed_pipeline_register_a		: STRING;
		signed_pipeline_register_b		: STRING;
		signed_register_a		: STRING;
		signed_register_b		: STRING;
		width_a		: NATURAL;
		width_b		: NATURAL;
		width_result		: NATURAL
	);
	PORT (
			dataa	: IN STD_LOGIC_VECTOR (width_a-1 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (width_b-1 DOWNTO 0);
			clock0	: IN STD_LOGIC ;
			aclr3	: IN STD_LOGIC ;
			ena0	: IN STD_LOGIC ;
			result	: OUT STD_LOGIC_VECTOR (width_result-1 DOWNTO 0)
	);
	end component;
	
	-- identical component to that above, but fixed at 18x18, latency 2
	-- mul18usus generated by Quartus 
	component hcc_mul18usus
	PORT
	(
		aclr3		: IN STD_LOGIC  := '0';
		clock0		: IN STD_LOGIC  := '1';
		dataa_0		: IN STD_LOGIC_VECTOR (17 DOWNTO 0) :=  (OTHERS => '0');
		datab_0		: IN STD_LOGIC_VECTOR (17 DOWNTO 0) :=  (OTHERS => '0');
		ena0		: IN STD_LOGIC  := '1';
		result		: OUT STD_LOGIC_VECTOR (35 DOWNTO 0)
	);
	end component;

	COMPONENT lpm_add_sub
	GENERIC (
		lpm_direction		: STRING;
		lpm_hint		: STRING;
		lpm_pipeline		: NATURAL;
		lpm_type		: STRING;
		lpm_width		: NATURAL
	);
	PORT (
			dataa	: IN STD_LOGIC_VECTOR (71 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (71 DOWNTO 0);
			clken	: IN STD_LOGIC ;
			aclr	: IN STD_LOGIC ;
			clock	: IN STD_LOGIC ;
			result	: OUT STD_LOGIC_VECTOR (71 DOWNTO 0)
	);
	END COMPONENT;
		 
BEGIN

  gza: FOR k IN 1 TO 36 GENERATE
    zerovec(k) <= '0';
  END GENERATE;

  muloneaa <= mulaa(54 DOWNTO 19);
  mulonebb <= mulbb(54 DOWNTO 19);
  
  multwoaa <= mulaa(18 DOWNTO 1);
  multwobb <= mulbb(36 DOWNTO 19);
  multhraa <= mulaa(18 DOWNTO 1);
  multhrbb <= mulbb(54 DOWNTO 37);
  
  mulforaa <= mulbb(18 DOWNTO 1);
  mulforbb <= mulaa(36 DOWNTO 19);
  mulfivaa <= mulbb(18 DOWNTO 1);
  mulfivbb <= mulaa(54 DOWNTO 37);
  
  -- {A,C) * {B,D}
  -- AAC
  -- BBD
  
  -- AA*BB 36x36=72, latency 3
  mulone : altmult_add
  GENERIC MAP (
		addnsub_multiplier_aclr1 => "ACLR3",
		addnsub_multiplier_pipeline_aclr1 => "ACLR3",
		addnsub_multiplier_pipeline_register1 => "CLOCK0",
		addnsub_multiplier_register1 => "CLOCK0",
		dedicated_multiplier_circuitry => "AUTO",
		input_aclr_a0 => "ACLR3",
		input_aclr_b0 => "ACLR3",
		input_register_a0 => "CLOCK0",
		input_register_b0 => "CLOCK0",
		input_source_a0 => "DATAA",
		input_source_b0 => "DATAB",
		intended_device_family => "Stratix II",
		lpm_type => "altmult_add",
		multiplier1_direction => "ADD",
		multiplier_aclr0 => "ACLR3",
		multiplier_register0 => "CLOCK0",
		number_of_multipliers => 1,
		output_aclr => "ACLR3",
		output_register => "CLOCK0",
		port_addnsub1 => "PORT_UNUSED",
		port_signa => "PORT_UNUSED",
		port_signb => "PORT_UNUSED",
		representation_a => "UNSIGNED",
		representation_b => "UNSIGNED",
		signed_aclr_a => "ACLR3",
		signed_aclr_b => "ACLR3",
		signed_pipeline_aclr_a => "ACLR3",
		signed_pipeline_aclr_b => "ACLR3",
		signed_pipeline_register_a => "CLOCK0",
		signed_pipeline_register_b => "CLOCK0",
		signed_register_a => "CLOCK0",
		signed_register_b => "CLOCK0",
		width_a => 36,
		width_b => 36,
		width_result => 72
	)
	PORT MAP (
		dataa => muloneaa,
		datab => mulonebb,
		clock0 => sysclk,
		aclr3 => reset,
		ena0 => enable,
		result => muloneout
	);

  --	Blo*C 18*18 = 36, latency = 2
	multwo: hcc_mul18usus
	PORT MAP (
		dataa_0 => multwoaa,
		datab_0 => multwobb,
		clock0 => sysclk,
		aclr3 => reset,
		ena0 => enable,
		result => multwoout
	);
		
  --	Bhi*C 18*18 = 36, latency = 2
  multhr: hcc_mul18usus
	PORT MAP (
		dataa_0 => multhraa,
		datab_0 => multhrbb,
		clock0 => sysclk,
		aclr3 => reset,
		ena0 => enable,
		result => multhrout
	);
	
  --	Alo*D 18*18 = 36, latency = 2
  mulfor: hcc_mul18usus
	PORT MAP (
		dataa_0 => mulforaa,
		datab_0 => mulforbb,
		clock0 => sysclk,
		aclr3 => reset,
		ena0 => enable,
		result => mulforout
	);	

  --	Ahi*D 18*18 = 36, latency = 2
  mulfiv: hcc_mul18usus
	PORT MAP (
		dataa_0 => mulfivaa,
		datab_0 => mulfivbb,
		clock0 => sysclk,
		aclr3 => reset,
		ena0 => enable,
		result => mulfivout
	);

  vecone <= zerovec(22 DOWNTO 1) & multwoout;
  vectwo <= zerovec(4 DOWNTO 1) & multhrout & zerovec(18 DOWNTO 1);
  vecthr <= zerovec(22 DOWNTO 1) & mulforout;
  vecfor <= zerovec(4 DOWNTO 1) & mulfivout & zerovec(18 DOWNTO 1);

  gva: FOR k IN 1 TO 58 GENERATE
    sumvecone(k) <= vecone(k) XOR vectwo(k) XOR vecthr(k);
    carvecone(k) <= (vecone(k) AND vectwo(k)) OR 
                    (vectwo(k) AND vecthr(k)) OR 
                    (vecone(k) AND vecthr(k));
  END GENERATE;
 
  vecfiv <= vecfor;
  vecsix <= sumvecone;
  vecsev <= carvecone(57 DOWNTO 1) & '0';

  gvb: FOR k IN 1 TO 58 GENERATE
    sumvectwo(k) <= vecfiv(k) XOR vecsix(k) XOR vecsev(k);
    carvectwo(k) <= (vecfiv(k) AND vecsix(k)) OR 
                    (vecsix(k) AND vecsev(k)) OR 
                    (vecfiv(k) AND vecsev(k));
  END GENERATE;

  paa: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN

      FOR k IN 1 TO 58 LOOP
        sumoneff(k) <= '0';
        caroneff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 72 LOOP
        sumtwoff(k) <= '0';
        cartwoff(k) <= '0';
      END LOOP;
      

    ELSIF (rising_edge(sysclk)) THEN

      IF (enable = '1') THEN

        sumoneff <= sumvectwo;
        caroneff <= carvectwo(57 DOWNTO 1) & '0';
        sumtwoff <= sumvecthr;
        cartwoff <= carvecthr(71 DOWNTO 1) & '0';

      END IF;

    END IF;

  END PROCESS;
  
  vecegt <= zerovec(32 DOWNTO 1) & sumoneff(58 DOWNTO 19);
  vecnin <= zerovec(32 DOWNTO 1) & caroneff(58 DOWNTO 19);
  vecten <= muloneout(72 DOWNTO 1);
  vecten <= muloneout(72 DOWNTO 1);

  gvc: FOR k IN 1 TO 72 GENERATE
    sumvecthr(k) <= vecegt(k) XOR vecnin(k) XOR vecten(k);
    carvecthr(k) <= (vecegt(k) AND vecnin(k)) OR 
                    (vecnin(k) AND vecten(k)) OR 
                    (vecegt(k) AND vecten(k));
  END GENERATE;

	adder : lpm_add_sub
	GENERIC MAP (
		lpm_direction => "ADD",
		lpm_hint => "ONE_INPUT_IS_CONSTANT=NO,CIN_USED=NO",
		lpm_pipeline => latency-4,
		lpm_type => "LPM_ADD_SUB",
		lpm_width => 72
	)
	PORT MAP (
		dataa => sumtwoff(72 DOWNTO 1),
		datab => cartwoff(72 DOWNTO 1),
		clken => enable,
		aclr => reset,
		clock => sysclk,
		result => resultnode
	);
	
  mulcc <= resultnode;
                                  
END syn;


LIBRARY ieee;
LIBRARY work;
LIBRARY lpm;
LIBRARY altera_mf;
USE lpm.all;
USE altera_mf.all;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   ALTERA FLOATING POINT DATAPATH COMPILER   ***
--***                                             ***
--***   FP_MUL54US_29S.VHD                        ***
--***                                             ***
--***   Function: 5/6 pipeline stage unsigned 54  ***
--***   bit multiplier                            ***
--***   29S: Stratix 2, 9 18x18, synthesizeable   ***
--***                                             ***
--***   21/04/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** 1. Identical to HCC_MUL54US_29S, except 5   ***
--*** or 6 pipeline parameter and 72 outputs      ***
--***************************************************

ENTITY fp_mul54us_29s IS
GENERIC (latency : positive := 5);
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      mulaa, mulbb : IN STD_LOGIC_VECTOR (54 DOWNTO 1);      

      mulcc : OUT STD_LOGIC_VECTOR (72 DOWNTO 1)  
     );
END fp_mul54us_29s;

ARCHITECTURE syn of fp_mul54us_29s IS

  signal muloneaa, mulonebb : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal multwoaa, multwobb, multhraa, multhrbb : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal mulforaa, mulforbb, mulfivaa, mulfivbb : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal mulsixaa, mulsixbb : STD_LOGIC_VECTOR (18 DOWNTO 1);
  signal muloneout : STD_LOGIC_VECTOR (72 DOWNTO 1);
  signal multwoout, multhrout, mulforout, mulfivout, mulsixout : STD_LOGIC_VECTOR (36 DOWNTO 1);

  signal vecone, vectwo, vecthr, vecfor, vecfiv : STD_LOGIC_VECTOR (72 DOWNTO 1);
  signal vecsix, vecsev, vecegt, vecnin, vecten : STD_LOGIC_VECTOR (72 DOWNTO 1);
  signal sumvecone, carvecone : STD_LOGIC_VECTOR (72 DOWNTO 1);
  signal sumvectwo, carvectwo : STD_LOGIC_VECTOR (72 DOWNTO 1);
  signal sumvecthr, carvecthr : STD_LOGIC_VECTOR (72 DOWNTO 1);
  signal sumoneff, caroneff : STD_LOGIC_VECTOR (72 DOWNTO 1);
  signal sumtwoff, cartwoff : STD_LOGIC_VECTOR (72 DOWNTO 1);
  signal resultnode : STD_LOGIC_VECTOR (72 DOWNTO 1);
  
  signal zerovec : STD_LOGIC_VECTOR (36 DOWNTO 1);

  component altmult_add
	GENERIC (
		addnsub_multiplier_aclr1		: STRING;
		addnsub_multiplier_pipeline_aclr1		: STRING;
		addnsub_multiplier_pipeline_register1		: STRING;
		addnsub_multiplier_register1		: STRING;
		dedicated_multiplier_circuitry		: STRING;
		input_aclr_a0		: STRING;
		input_aclr_b0		: STRING;
		input_register_a0		: STRING;
		input_register_b0		: STRING;
		input_source_a0		: STRING;
		input_source_b0		: STRING;
		intended_device_family		: STRING;
		lpm_type		: STRING;
		multiplier1_direction		: STRING;
		multiplier_aclr0		: STRING;
		multiplier_register0		: STRING;
		number_of_multipliers		: NATURAL;
		output_aclr		: STRING;
		output_register		: STRING;
		port_addnsub1		: STRING;
		port_signa		: STRING;
		port_signb		: STRING;
		representation_a		: STRING;
		representation_b		: STRING;
		signed_aclr_a		: STRING;
		signed_aclr_b		: STRING;
		signed_pipeline_aclr_a		: STRING;
		signed_pipeline_aclr_b		: STRING;
		signed_pipeline_register_a		: STRING;
		signed_pipeline_register_b		: STRING;
		signed_register_a		: STRING;
		signed_register_b		: STRING;
		width_a		: NATURAL;
		width_b		: NATURAL;
		width_result		: NATURAL
	);
	PORT (
			dataa	: IN STD_LOGIC_VECTOR (width_a-1 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (width_b-1 DOWNTO 0);
			clock0	: IN STD_LOGIC ;
			aclr3	: IN STD_LOGIC ;
			ena0	: IN STD_LOGIC ;
			result	: OUT STD_LOGIC_VECTOR (width_result-1 DOWNTO 0)
	);
	end component;
	
	-- identical component to that above, but fixed at 18x18, latency 2
	-- mul18usus generated by Quartus 
	component hcc_mul18usus
	PORT
	(
		aclr3		: IN STD_LOGIC  := '0';
		clock0		: IN STD_LOGIC  := '1';
		dataa_0		: IN STD_LOGIC_VECTOR (17 DOWNTO 0) :=  (OTHERS => '0');
		datab_0		: IN STD_LOGIC_VECTOR (17 DOWNTO 0) :=  (OTHERS => '0');
		ena0		: IN STD_LOGIC  := '1';
		result		: OUT STD_LOGIC_VECTOR (35 DOWNTO 0)
	);
	end component;

	COMPONENT lpm_add_sub
	GENERIC (
		lpm_direction		: STRING;
		lpm_hint		: STRING;
		lpm_pipeline		: NATURAL;
		lpm_type		: STRING;
		lpm_width		: NATURAL
	);
	PORT (
			dataa	: IN STD_LOGIC_VECTOR (71 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (71 DOWNTO 0);
			clken	: IN STD_LOGIC ;
			aclr	: IN STD_LOGIC ;
			clock	: IN STD_LOGIC ;
			result	: OUT STD_LOGIC_VECTOR (71 DOWNTO 0)
	);
	END COMPONENT;
		 
BEGIN

  gza: FOR k IN 1 TO 36 GENERATE
    zerovec(k) <= '0';
  END GENERATE;

  muloneaa <= mulaa(36 DOWNTO 1);
  mulonebb <= mulbb(36 DOWNTO 1);
  
  multwoaa <= mulaa(54 DOWNTO 37);
  multwobb <= mulbb(18 DOWNTO 1);
  multhraa <= mulaa(54 DOWNTO 37);
  multhrbb <= mulbb(36 DOWNTO 19);
  
  mulforaa <= mulbb(54 DOWNTO 37);
  mulforbb <= mulaa(18 DOWNTO 1);
  mulfivaa <= mulbb(54 DOWNTO 37);
  mulfivbb <= mulaa(36 DOWNTO 19);
  
  mulsixaa <= mulbb(54 DOWNTO 37);
  mulsixbb <= mulaa(54 DOWNTO 37);
  
  -- {C,A) * {D,B}
  -- CAA
  -- DBB
  
  -- AA*BB 36x36=72, latency 3
  mulone : altmult_add
  GENERIC MAP (
		addnsub_multiplier_aclr1 => "ACLR3",
		addnsub_multiplier_pipeline_aclr1 => "ACLR3",
		addnsub_multiplier_pipeline_register1 => "CLOCK0",
		addnsub_multiplier_register1 => "CLOCK0",
		dedicated_multiplier_circuitry => "AUTO",
		input_aclr_a0 => "ACLR3",
		input_aclr_b0 => "ACLR3",
		input_register_a0 => "CLOCK0",
		input_register_b0 => "CLOCK0",
		input_source_a0 => "DATAA",
		input_source_b0 => "DATAB",
		intended_device_family => "Stratix II",
		lpm_type => "altmult_add",
		multiplier1_direction => "ADD",
		multiplier_aclr0 => "ACLR3",
		multiplier_register0 => "CLOCK0",
		number_of_multipliers => 1,
		output_aclr => "ACLR3",
		output_register => "CLOCK0",
		port_addnsub1 => "PORT_UNUSED",
		port_signa => "PORT_UNUSED",
		port_signb => "PORT_UNUSED",
		representation_a => "UNSIGNED",
		representation_b => "UNSIGNED",
		signed_aclr_a => "ACLR3",
		signed_aclr_b => "ACLR3",
		signed_pipeline_aclr_a => "ACLR3",
		signed_pipeline_aclr_b => "ACLR3",
		signed_pipeline_register_a => "CLOCK0",
		signed_pipeline_register_b => "CLOCK0",
		signed_register_a => "CLOCK0",
		signed_register_b => "CLOCK0",
		width_a => 36,
		width_b => 36,
		width_result => 72
	)
	PORT MAP (
		dataa => muloneaa,
		datab => mulonebb,
		clock0 => sysclk,
		aclr3 => reset,
		ena0 => enable,
		result => muloneout
	);

  --	Blo*C 18*18 = 36, latency = 2
	multwo: hcc_mul18usus
	PORT MAP (
		dataa_0 => multwoaa,
		datab_0 => multwobb,
		clock0 => sysclk,
		aclr3 => reset,
		ena0 => enable,
		result => multwoout
	);
		
  --	Bhi*C 18*18 = 36, latency = 2
  multhr: hcc_mul18usus
	PORT MAP (
		dataa_0 => multhraa,
		datab_0 => multhrbb,
		clock0 => sysclk,
		aclr3 => reset,
		ena0 => enable,
		result => multhrout
	);
	
  --	Alo*D 18*18 = 36, latency = 2
  mulfor: hcc_mul18usus
	PORT MAP (
		dataa_0 => mulforaa,
		datab_0 => mulforbb,
		clock0 => sysclk,
		aclr3 => reset,
		ena0 => enable,
		result => mulforout
	);	

  --	Ahi*D 18*18 = 36, latency = 2
  mulfiv: hcc_mul18usus
	PORT MAP (
		dataa_0 => mulfivaa,
		datab_0 => mulfivbb,
		clock0 => sysclk,
		aclr3 => reset,
		ena0 => enable,
		result => mulfivout
	);

  --	C*D 18*18 = 36, latency = 3
  mulsix : altmult_add
  GENERIC MAP (
		addnsub_multiplier_aclr1 => "ACLR3",
		addnsub_multiplier_pipeline_aclr1 => "ACLR3",
		addnsub_multiplier_pipeline_register1 => "CLOCK0",
		addnsub_multiplier_register1 => "CLOCK0",
		dedicated_multiplier_circuitry => "AUTO",
		input_aclr_a0 => "ACLR3",
		input_aclr_b0 => "ACLR3",
		input_register_a0 => "CLOCK0",
		input_register_b0 => "CLOCK0",
		input_source_a0 => "DATAA",
		input_source_b0 => "DATAB",
		intended_device_family => "Stratix II",
		lpm_type => "altmult_add",
		multiplier1_direction => "ADD",
		multiplier_aclr0 => "ACLR3",
		multiplier_register0 => "CLOCK0",
		number_of_multipliers => 1,
		output_aclr => "ACLR3",
		output_register => "CLOCK0",
		port_addnsub1 => "PORT_UNUSED",
		port_signa => "PORT_UNUSED",
		port_signb => "PORT_UNUSED",
		representation_a => "UNSIGNED",
		representation_b => "UNSIGNED",
		signed_aclr_a => "ACLR3",
		signed_aclr_b => "ACLR3",
		signed_pipeline_aclr_a => "ACLR3",
		signed_pipeline_aclr_b => "ACLR3",
		signed_pipeline_register_a => "CLOCK0",
		signed_pipeline_register_b => "CLOCK0",
		signed_register_a => "CLOCK0",
		signed_register_b => "CLOCK0",
		width_a => 18,
		width_b => 18,
		width_result => 36
	)
	PORT MAP (
		dataa => mulsixaa,
		datab => mulsixbb,
		clock0 => sysclk,
		aclr3 => reset,
		ena0 => enable,
		result => mulsixout
	);
	
  vecone <= zerovec(36 DOWNTO 1) & multwoout;
  vectwo <= zerovec(18 DOWNTO 1) & multhrout & zerovec(18 DOWNTO 1);
  vecthr <= zerovec(36 DOWNTO 1) & mulforout;
  vecfor <= zerovec(18 DOWNTO 1) & mulfivout & zerovec(18 DOWNTO 1);

  gva: FOR k IN 1 TO 72 GENERATE
    sumvecone(k) <= vecone(k) XOR vectwo(k) XOR vecthr(k);
    carvecone(k) <= (vecone(k) AND vectwo(k)) OR 
                    (vectwo(k) AND vecthr(k)) OR 
                    (vecone(k) AND vecthr(k));
  END GENERATE;
 
  vecfiv <= vecfor;
  vecsix <= sumvecone;
  vecsev <= carvecone(71 DOWNTO 1) & '0';

  gvb: FOR k IN 1 TO 72 GENERATE
    sumvectwo(k) <= vecfiv(k) XOR vecsix(k) XOR vecsev(k);
    carvectwo(k) <= (vecfiv(k) AND vecsix(k)) OR 
                    (vecsix(k) AND vecsev(k)) OR 
                    (vecfiv(k) AND vecsev(k));
  END GENERATE;

  paa: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN

      FOR k IN 1 TO 72 LOOP
        sumoneff(k) <= '0';
        caroneff(k) <= '0';
        sumtwoff(k) <= '0';
        cartwoff(k) <= '0';
      END LOOP;

    ELSIF (rising_edge(sysclk)) THEN

      IF (enable = '1') THEN

        sumoneff <= sumvectwo;
        caroneff <= carvectwo(71 DOWNTO 1) & '0';
        sumtwoff <= sumvecthr;
        cartwoff <= carvecthr(71 DOWNTO 1) & '0';

      END IF;

    END IF;

  END PROCESS;

  vecegt <= sumoneff;
  vecnin <= caroneff;
  vecten <= mulsixout & muloneout(72 DOWNTO 37);

  gvc: FOR k IN 1 TO 72 GENERATE
    sumvecthr(k) <= vecegt(k) XOR vecnin(k) XOR vecten(k);
    carvecthr(k) <= (vecegt(k) AND vecnin(k)) OR 
                    (vecnin(k) AND vecten(k)) OR 
                    (vecegt(k) AND vecten(k));
  END GENERATE;

  -- according to marcel, 2 pipes = 1 pipe in middle, on on output
	adder : lpm_add_sub
	GENERIC MAP (
		lpm_direction => "ADD",
		lpm_hint => "ONE_INPUT_IS_CONSTANT=NO,CIN_USED=NO",
		lpm_pipeline => latency-4,
		lpm_type => "LPM_ADD_SUB",
		lpm_width => 72
	)
	PORT MAP (
		dataa => sumtwoff(72 DOWNTO 1),
		datab => cartwoff(72 DOWNTO 1),
		clken => enable,
		aclr => reset,
		clock => sysclk,
		result => resultnode
	);
	
  mulcc <= resultnode;
                                  
END syn;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   ALTERA FLOATING POINT DATAPATH COMPILER   ***
--***                                             ***
--***   FP_MUL54US_38S.VHD                        ***
--***                                             ***
--***   Function: 4 pipeline stage unsigned 54    ***
--***   bit multiplier                            ***
--***   38S: Stratix 3, 8 18x18, synthesizeable   ***
--***                                             ***
--***   20/08/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** Build explicitlyout of two SIII/SIV         ***
--*** DSP Blocks                                  ***
--***************************************************

ENTITY fp_mul54us_38s IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      mulaa : IN STD_LOGIC_VECTOR (54 DOWNTO 1);
      mulbb : IN STD_LOGIC_VECTOR (54 DOWNTO 1);
      
		  mulcc : OUT STD_LOGIC_VECTOR (72 DOWNTO 1)
		);
END fp_mul54us_38s;

ARCHITECTURE rtl OF fp_mul54us_38s IS

  signal zerovec : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal multone : STD_LOGIC_VECTOR (72 DOWNTO 1);
  signal multtwo : STD_LOGIC_VECTOR (55 DOWNTO 1);
  signal addmultff : STD_LOGIC_VECTOR (72 DOWNTO 1);
  
  component fp_mul3s
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1);

	      result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
	     );
  end component;

  component fp_sum36x18
	PORT (
		    aclr3		: IN STD_LOGIC  := '0';
		    clock0		: IN STD_LOGIC  := '1';
		    dataa_0		: IN STD_LOGIC_VECTOR (17 DOWNTO 0) :=  (OTHERS => '0');
		    dataa_1		: IN STD_LOGIC_VECTOR (17 DOWNTO 0) :=  (OTHERS => '0');
		    datab_0		: IN STD_LOGIC_VECTOR (35 DOWNTO 0) :=  (OTHERS => '0');
		    datab_1		: IN STD_LOGIC_VECTOR (35 DOWNTO 0) :=  (OTHERS => '0');
		    ena0		: IN STD_LOGIC  := '1';
		    result		: OUT STD_LOGIC_VECTOR (54 DOWNTO 0)
	    );
	end component;
	
BEGIN
  
  gza: FOR k IN 1 TO 36 GENERATE
    zerovec(k) <= '0';
  END GENERATE;

  mone: fp_mul3s
  GENERIC MAP (widthaa=>36,widthbb=>36,widthcc=>72)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dataaa=>mulaa(54 DOWNTO 19),databb=>mulbb(54 DOWNTO 19),
            result=>multone);
      
  mtwo: fp_sum36x18
  PORT MAP (aclr3=>reset,clock0=>sysclk,
            dataa_0=>mulaa(18 DOWNTO 1),
            dataa_1=>mulbb(18 DOWNTO 1),
            datab_0=>mulbb(54 DOWNTO 19),
            datab_1=>mulaa(54 DOWNTO 19),
            ena0=>enable,
            result=>multtwo);
            
  paa: PROCESS (sysclk,reset)
  BEGIN
    
    IF (reset = '1') THEN
      FOR k IN 1 TO 72 LOOP
        addmultff(k) <= '0';
      END LOOP;
    ELSIF (rising_edge(sysclk)) THEN
      IF (enable = '1') THEN
        addmultff <= multone + (zerovec(35 DOWNTO 1) & multtwo(55 DOWNTO 19));
      END IF;
    END IF;
    
  END PROCESS;
        
  mulcc <= addmultff;
         
END rtl;


	
LIBRARY ieee;
LIBRARY work;
LIBRARY lpm;
LIBRARY altera_mf;
USE lpm.all;
USE altera_mf.all;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   ALTERA FLOATING POINT DATAPATH COMPILER   ***
--***                                             ***
--***   FP_MUL54US_3XS.VHD                        ***
--***                                             ***
--***   Function: 4 pipeline stage unsigned 54    ***
--***   bit multiplier                            ***
--***   3XS: Stratix 3, 10 18x18, synthesizeable  ***
--***                                             ***
--***   21/04/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** 1. For QII8.0 LPM_MULT always creates a 10  ***
--*** 18x18 multiplier 54x54 core                 ***
--*** 2. Identical to HCC_MUL54US_3XS, but 72     ***
--*** outputs                                     ***
--***                                             ***
--***************************************************

ENTITY fp_mul54us_3xs IS
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      mulaa, mulbb : IN STD_LOGIC_VECTOR (54 DOWNTO 1);      

      mulcc : OUT STD_LOGIC_VECTOR (72 DOWNTO 1)  
     );
END fp_mul54us_3xs;

ARCHITECTURE syn of fp_mul54us_3xs IS

  component lpm_mult
  GENERIC (
		     lpm_hint		: STRING;
		     lpm_pipeline		: NATURAL;
		     lpm_representation		: STRING;
		     lpm_type		: STRING;
		     lpm_widtha		: NATURAL;
		     lpm_widthb		: NATURAL;
		     lpm_widthp		: NATURAL
	      );
	PORT (
			dataa	: IN STD_LOGIC_VECTOR (53 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (53 DOWNTO 0);
			clken	: IN STD_LOGIC ;
			aclr	: IN STD_LOGIC ;
			clock	: IN STD_LOGIC ;
			result	: OUT STD_LOGIC_VECTOR (71 DOWNTO 0)
	);
	end component;
 
BEGIN

 	lpm_mult_component : lpm_mult
	GENERIC MAP (
		lpm_hint => "MAXIMIZE_SPEED=5",
		lpm_pipeline => 4,
		lpm_representation => "UNSIGNED",
		lpm_type => "LPM_MULT",
		lpm_widtha => 54,
		lpm_widthb => 54,
		lpm_widthp => 72
	)
	PORT MAP (
		dataa => mulaa,
		datab => mulbb,
		clken => enable,
		aclr => reset,
		clock => sysclk,
		result => mulcc
	);
                                  
END syn;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   ALTERA FLOATING POINT DATAPATH COMPILER   ***
--***                                             ***
--***   FP_MUL54USB.VHD                           ***
--***                                             ***
--***   Function: 4/5/6 pipeline stage unsigned   ***
--***             54 bit multiplier (behavioral)  ***
--***                                             ***
--***   24/04/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***   31/01/08 ML see below                     ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_mul54usb IS 

 GENERIC (
          latency : positive := 5; -- 4/5/6
          device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
          prune : integer := 0 -- 0 = pruned multiplier, 1 = normal multiplier
         );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      aa, bb : IN STD_LOGIC_VECTOR (54 DOWNTO 1);
      
	cc : OUT STD_LOGIC_VECTOR (72 DOWNTO 1)
	);
END fp_mul54usb;

ARCHITECTURE rtl OF fp_mul54usb IS
 
  constant delaydepth : integer := latency - 2;
  
  type muldelfftype IS ARRAY (delaydepth DOWNTO 1) OF STD_LOGIC_VECTOR (72 DOWNTO 1);
  
  signal zerovec : STD_LOGIC_VECTOR (72 DOWNTO 1);
  
  signal aaff, bbff : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal mulff : STD_LOGIC_VECTOR (108 DOWNTO 1);
  signal muldelff : muldelfftype;
  
  signal mulnode : STD_LOGIC_VECTOR (108 DOWNTO 1);
  signal mulonenode, multwonode : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal multhrnode : STD_LOGIC_VECTOR (72 DOWNTO 1);
    
BEGIN
    
  gza: FOR k IN 1 TO 72 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  pma: PROCESS (sysclk, reset)
  BEGIN
  
    IF (reset = '1') THEN
        
      FOR k IN 1 TO 54 LOOP
        mulff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 108 LOOP
        mulff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO delaydepth LOOP
        FOR j IN 1 TO 72 LOOP
          muldelff(k)(j) <= '0';
        END LOOP;
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
        
      IF (enable = '1') THEN

        aaff <= aa; 
        bbff <= bb;
        mulff <= mulnode;
        muldelff(1)(72 DOWNTO 1) <= mulff(108 DOWNTO 37);
        FOR k IN 2 TO delaydepth LOOP
          muldelff(k)(72 DOWNTO 1) <= muldelff(k-1)(72 DOWNTO 1);
        END LOOP;
         
      END IF;
                 
    END IF;
  
  END PROCESS;
  
  -- full multiplier
  gpa: IF (prune = 1) GENERATE
    mulonenode <= zerovec(54 DOWNTO 1);
    multwonode <= zerovec(54 DOWNTO 1);
    multhrnode <= zerovec(72 DOWNTO 1);
    mulnode <= aaff * bbff;
  END GENERATE;
    
  -- pruned multiplier (18x18 LSB contribution missing)
  gpb: IF (prune = 0) GENERATE
    mulonenode <= aaff(18 DOWNTO 1) * bbff(54 DOWNTO 19);
    multwonode <= bbff(18 DOWNTO 1) * aaff(54 DOWNTO 19);
    multhrnode <= aaff(54 DOWNTO 19) * bbff(54 DOWNTO 19);
    mulnode <= (multhrnode & zerovec(36 DOWNTO 1)) +  
               (zerovec(36 DOWNTO 1) & mulonenode & zerovec(18 DOWNTO 1)) + 
               (zerovec(36 DOWNTO 1) & multwonode & zerovec(18 DOWNTO 1));
  END GENERATE; 
                               
  cc <= muldelff(delaydepth)(72 DOWNTO 1); 
  
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   ALTERA FLOATING POINT DATAPATH COMPILER   ***
--***                                             ***
--***   FP_NEG.VHD                                ***
--***                                             ***
--***   Function: Single Precision Negative Value ***
--***                                             ***
--***   Created 11/09/09                          ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_neg IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (23 DOWNTO 1);

		  signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
		  satout, zeroout, nanout : OUT STD_LOGIC
		);
END fp_neg;

ARCHITECTURE rtl OF fp_neg IS
 
  signal signff : STD_LOGIC;
  signal exponentff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal mantissaff : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal expnode : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal expzerochk, expmaxchk : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal expzero, expmax : STD_LOGIC;
  signal manzerochk : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal manzero, mannonzero : STD_LOGIC; 

BEGIN
    
  pin: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
    
      signff <= '0';
      FOR k IN 1 TO 8 LOOP
        exponentff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 23 LOOP
        mantissaff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF (enable = '1') THEN
          
        signff <= NOT(signin);
        exponentff <= exponentin;
        mantissaff <= mantissain;
        
      END IF;
    
    END IF;  
      
  END PROCESS;

  expzerochk(1) <= exponentff(1);
  expmaxchk(1) <= exponentff(1);
  gxa: FOR k IN 2 TO 8 GENERATE
    expzerochk(k) <= expzerochk(k-1) OR exponentff(k);
    expmaxchk(k) <= expmaxchk(k-1) AND exponentff(k);
  END GENERATE;
  expzero <= NOT(expzerochk(8));
  expmax <= expmaxchk(8);
  
  manzerochk(1) <= mantissaff(1);
  gma: FOR k IN 2 TO 23 GENERATE
    manzerochk(k) <= manzerochk(k-1) OR mantissaff(k);
  END GENERATE;
  manzero <= NOT(manzerochk(23));
  mannonzero <= manzerochk(23);
  
  signout <= signff;
  exponentout <= exponentff;
  mantissaout <= mantissaff;
  satout <= expmax AND manzero;
  zeroout <= expzero;
  nanout <= expmax AND mannonzero;

END rtl;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT LIBRARY                    ***
--***                                             ***
--***   FP_POS.VHD                                ***
--***                                             ***
--***   Function: Local Count Leading Zeroes      ***
--***                                             ***
--***   22/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_pos IS
GENERIC (start : integer := 10);
PORT (
      ingroup : IN STD_LOGIC_VECTOR (6 DOWNTO 1);
      
      position : OUT STD_LOGIC_VECTOR (5 DOWNTO 1)   
     );
END fp_pos;

ARCHITECTURE rtl of fp_pos IS
  
BEGIN

ptab: PROCESS (ingroup)
BEGIN

  CASE ingroup IS
      
      WHEN "000000" => position <= conv_std_logic_vector(0,5);
          
      WHEN "000001" => position <= conv_std_logic_vector(start+5,5);
          
      WHEN "000010" => position <= conv_std_logic_vector(start+4,5);
      WHEN "000011" => position <= conv_std_logic_vector(start+4,5); 
          
      WHEN "000100" => position <= conv_std_logic_vector(start+3,5);
      WHEN "000101" => position <= conv_std_logic_vector(start+3,5);
      WHEN "000110" => position <= conv_std_logic_vector(start+3,5);
      WHEN "000111" => position <= conv_std_logic_vector(start+3,5);
       
      WHEN "001000" => position <= conv_std_logic_vector(start+2,5); 
      WHEN "001001" => position <= conv_std_logic_vector(start+2,5);
      WHEN "001010" => position <= conv_std_logic_vector(start+2,5);
      WHEN "001011" => position <= conv_std_logic_vector(start+2,5);
      WHEN "001100" => position <= conv_std_logic_vector(start+2,5);
      WHEN "001101" => position <= conv_std_logic_vector(start+2,5);
      WHEN "001110" => position <= conv_std_logic_vector(start+2,5);
      WHEN "001111" => position <= conv_std_logic_vector(start+2,5); 
              
      WHEN "010000" => position <= conv_std_logic_vector(start+1,5);
      WHEN "010001" => position <= conv_std_logic_vector(start+1,5);
      WHEN "010010" => position <= conv_std_logic_vector(start+1,5);
      WHEN "010011" => position <= conv_std_logic_vector(start+1,5);
      WHEN "010100" => position <= conv_std_logic_vector(start+1,5);
      WHEN "010101" => position <= conv_std_logic_vector(start+1,5);
      WHEN "010110" => position <= conv_std_logic_vector(start+1,5);
      WHEN "010111" => position <= conv_std_logic_vector(start+1,5);
      WHEN "011000" => position <= conv_std_logic_vector(start+1,5);
      WHEN "011001" => position <= conv_std_logic_vector(start+1,5);
      WHEN "011010" => position <= conv_std_logic_vector(start+1,5);
      WHEN "011011" => position <= conv_std_logic_vector(start+1,5);
      WHEN "011100" => position <= conv_std_logic_vector(start+1,5);
      WHEN "011101" => position <= conv_std_logic_vector(start+1,5);
      WHEN "011110" => position <= conv_std_logic_vector(start+1,5); 
      WHEN "011111" => position <= conv_std_logic_vector(start+1,5);  
 
      WHEN "100000" => position <= conv_std_logic_vector(start,5);
      WHEN "100001" => position <= conv_std_logic_vector(start,5);
      WHEN "100010" => position <= conv_std_logic_vector(start,5);
      WHEN "100011" => position <= conv_std_logic_vector(start,5);
      WHEN "100100" => position <= conv_std_logic_vector(start,5);
      WHEN "100101" => position <= conv_std_logic_vector(start,5);
      WHEN "100110" => position <= conv_std_logic_vector(start,5);
      WHEN "100111" => position <= conv_std_logic_vector(start,5);
      WHEN "101000" => position <= conv_std_logic_vector(start,5);
      WHEN "101001" => position <= conv_std_logic_vector(start,5);
      WHEN "101010" => position <= conv_std_logic_vector(start,5);
      WHEN "101011" => position <= conv_std_logic_vector(start,5);
      WHEN "101100" => position <= conv_std_logic_vector(start,5);
      WHEN "101101" => position <= conv_std_logic_vector(start,5);
      WHEN "101110" => position <= conv_std_logic_vector(start,5); 
      WHEN "101111" => position <= conv_std_logic_vector(start,5);      
      WHEN "110000" => position <= conv_std_logic_vector(start,5);
      WHEN "110001" => position <= conv_std_logic_vector(start,5);
      WHEN "110010" => position <= conv_std_logic_vector(start,5);
      WHEN "110011" => position <= conv_std_logic_vector(start,5);
      WHEN "110100" => position <= conv_std_logic_vector(start,5);
      WHEN "110101" => position <= conv_std_logic_vector(start,5);
      WHEN "110110" => position <= conv_std_logic_vector(start,5);
      WHEN "110111" => position <= conv_std_logic_vector(start,5);
      WHEN "111000" => position <= conv_std_logic_vector(start,5);
      WHEN "111001" => position <= conv_std_logic_vector(start,5);
      WHEN "111010" => position <= conv_std_logic_vector(start,5);
      WHEN "111011" => position <= conv_std_logic_vector(start,5);
      WHEN "111100" => position <= conv_std_logic_vector(start,5);
      WHEN "111101" => position <= conv_std_logic_vector(start,5);
      WHEN "111110" => position <= conv_std_logic_vector(start,5); 
      WHEN "111111" => position <= conv_std_logic_vector(start,5);
          
      WHEN others => position <= conv_std_logic_vector(0,5);
          
  END CASE;
               
END PROCESS;    
    
END rtl;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_POS51.VHD                              ***
--***                                             ***
--***   Function: 5 Bit Count Leading Zeros       ***
--***   Component                                 ***
--***                                             ***
--***   22/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_pos51 IS
GENERIC (start : integer := 10);
PORT (
      ingroup : IN STD_LOGIC_VECTOR (6 DOWNTO 1);
      
      position : OUT STD_LOGIC_VECTOR (5 DOWNTO 1)   
     );
END fp_pos51;

ARCHITECTURE sss of fp_pos51 IS
  
BEGIN

ptab: PROCESS (ingroup)
BEGIN

  CASE ingroup IS
      
      WHEN "000000" => position <= conv_std_logic_vector(0,5);
          
      WHEN "000001" => position <= conv_std_logic_vector(start+5,5);
          
      WHEN "000010" => position <= conv_std_logic_vector(start+4,5);
      WHEN "000011" => position <= conv_std_logic_vector(start+4,5); 
          
      WHEN "000100" => position <= conv_std_logic_vector(start+3,5);
      WHEN "000101" => position <= conv_std_logic_vector(start+3,5);
      WHEN "000110" => position <= conv_std_logic_vector(start+3,5);
      WHEN "000111" => position <= conv_std_logic_vector(start+3,5);
       
      WHEN "001000" => position <= conv_std_logic_vector(start+2,5); 
      WHEN "001001" => position <= conv_std_logic_vector(start+2,5);
      WHEN "001010" => position <= conv_std_logic_vector(start+2,5);
      WHEN "001011" => position <= conv_std_logic_vector(start+2,5);
      WHEN "001100" => position <= conv_std_logic_vector(start+2,5);
      WHEN "001101" => position <= conv_std_logic_vector(start+2,5);
      WHEN "001110" => position <= conv_std_logic_vector(start+2,5);
      WHEN "001111" => position <= conv_std_logic_vector(start+2,5); 
              
      WHEN "010000" => position <= conv_std_logic_vector(start+1,5);
      WHEN "010001" => position <= conv_std_logic_vector(start+1,5);
      WHEN "010010" => position <= conv_std_logic_vector(start+1,5);
      WHEN "010011" => position <= conv_std_logic_vector(start+1,5);
      WHEN "010100" => position <= conv_std_logic_vector(start+1,5);
      WHEN "010101" => position <= conv_std_logic_vector(start+1,5);
      WHEN "010110" => position <= conv_std_logic_vector(start+1,5);
      WHEN "010111" => position <= conv_std_logic_vector(start+1,5);
      WHEN "011000" => position <= conv_std_logic_vector(start+1,5);
      WHEN "011001" => position <= conv_std_logic_vector(start+1,5);
      WHEN "011010" => position <= conv_std_logic_vector(start+1,5);
      WHEN "011011" => position <= conv_std_logic_vector(start+1,5);
      WHEN "011100" => position <= conv_std_logic_vector(start+1,5);
      WHEN "011101" => position <= conv_std_logic_vector(start+1,5);
      WHEN "011110" => position <= conv_std_logic_vector(start+1,5); 
      WHEN "011111" => position <= conv_std_logic_vector(start+1,5);  

      WHEN "100000" => position <= conv_std_logic_vector(start,5);
      WHEN "100001" => position <= conv_std_logic_vector(start,5);
      WHEN "100010" => position <= conv_std_logic_vector(start,5);
      WHEN "100011" => position <= conv_std_logic_vector(start,5);
      WHEN "100100" => position <= conv_std_logic_vector(start,5);
      WHEN "100101" => position <= conv_std_logic_vector(start,5);
      WHEN "100110" => position <= conv_std_logic_vector(start,5);
      WHEN "100111" => position <= conv_std_logic_vector(start,5);
      WHEN "101000" => position <= conv_std_logic_vector(start,5);
      WHEN "101001" => position <= conv_std_logic_vector(start,5);
      WHEN "101010" => position <= conv_std_logic_vector(start,5);
      WHEN "101011" => position <= conv_std_logic_vector(start,5);
      WHEN "101100" => position <= conv_std_logic_vector(start,5);
      WHEN "101101" => position <= conv_std_logic_vector(start,5);
      WHEN "101110" => position <= conv_std_logic_vector(start,5); 
      WHEN "101111" => position <= conv_std_logic_vector(start,5);      
      WHEN "110000" => position <= conv_std_logic_vector(start,5);
      WHEN "110001" => position <= conv_std_logic_vector(start,5);
      WHEN "110010" => position <= conv_std_logic_vector(start,5);
      WHEN "110011" => position <= conv_std_logic_vector(start,5);
      WHEN "110100" => position <= conv_std_logic_vector(start,5);
      WHEN "110101" => position <= conv_std_logic_vector(start,5);
      WHEN "110110" => position <= conv_std_logic_vector(start,5);
      WHEN "110111" => position <= conv_std_logic_vector(start,5);
      WHEN "111000" => position <= conv_std_logic_vector(start,5);
      WHEN "111001" => position <= conv_std_logic_vector(start,5);
      WHEN "111010" => position <= conv_std_logic_vector(start,5);
      WHEN "111011" => position <= conv_std_logic_vector(start,5);
      WHEN "111100" => position <= conv_std_logic_vector(start,5);
      WHEN "111101" => position <= conv_std_logic_vector(start,5);
      WHEN "111110" => position <= conv_std_logic_vector(start,5); 
      WHEN "111111" => position <= conv_std_logic_vector(start,5);
          
      WHEN others => position <= conv_std_logic_vector(0,5);
          
  END CASE;
               
END PROCESS;    
    
END sss;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_POS52.VHD                              ***
--***                                             ***
--***   Function: 6 Bit Count Leading Zeros       ***
--***   Component                                 ***
--***                                             ***
--***   22/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_pos52 IS
GENERIC (start : integer := 10);
PORT (
      ingroup : IN STD_LOGIC_VECTOR (6 DOWNTO 1);
      
      position : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)   
     );
END fp_pos52;

ARCHITECTURE sss of fp_pos52 IS
  
BEGIN

ptab: PROCESS (ingroup)
BEGIN

  CASE ingroup IS
      
      WHEN "000000" => position <= conv_std_logic_vector(0,6);
          
      WHEN "000001" => position <= conv_std_logic_vector(start+5,6);
          
      WHEN "000010" => position <= conv_std_logic_vector(start+4,6);
      WHEN "000011" => position <= conv_std_logic_vector(start+4,6); 
          
      WHEN "000100" => position <= conv_std_logic_vector(start+3,6);
      WHEN "000101" => position <= conv_std_logic_vector(start+3,6);
      WHEN "000110" => position <= conv_std_logic_vector(start+3,6);
      WHEN "000111" => position <= conv_std_logic_vector(start+3,6);
       
      WHEN "001000" => position <= conv_std_logic_vector(start+2,6); 
      WHEN "001001" => position <= conv_std_logic_vector(start+2,6);
      WHEN "001010" => position <= conv_std_logic_vector(start+2,6);
      WHEN "001011" => position <= conv_std_logic_vector(start+2,6);
      WHEN "001100" => position <= conv_std_logic_vector(start+2,6);
      WHEN "001101" => position <= conv_std_logic_vector(start+2,6);
      WHEN "001110" => position <= conv_std_logic_vector(start+2,6);
      WHEN "001111" => position <= conv_std_logic_vector(start+2,6); 
              
      WHEN "010000" => position <= conv_std_logic_vector(start+1,6);
      WHEN "010001" => position <= conv_std_logic_vector(start+1,6);
      WHEN "010010" => position <= conv_std_logic_vector(start+1,6);
      WHEN "010011" => position <= conv_std_logic_vector(start+1,6);
      WHEN "010100" => position <= conv_std_logic_vector(start+1,6);
      WHEN "010101" => position <= conv_std_logic_vector(start+1,6);
      WHEN "010110" => position <= conv_std_logic_vector(start+1,6);
      WHEN "010111" => position <= conv_std_logic_vector(start+1,6);
      WHEN "011000" => position <= conv_std_logic_vector(start+1,6);
      WHEN "011001" => position <= conv_std_logic_vector(start+1,6);
      WHEN "011010" => position <= conv_std_logic_vector(start+1,6);
      WHEN "011011" => position <= conv_std_logic_vector(start+1,6);
      WHEN "011100" => position <= conv_std_logic_vector(start+1,6);
      WHEN "011101" => position <= conv_std_logic_vector(start+1,6);
      WHEN "011110" => position <= conv_std_logic_vector(start+1,6); 
      WHEN "011111" => position <= conv_std_logic_vector(start+1,6);  

      WHEN "100000" => position <= conv_std_logic_vector(start,6);
      WHEN "100001" => position <= conv_std_logic_vector(start,6);
      WHEN "100010" => position <= conv_std_logic_vector(start,6);
      WHEN "100011" => position <= conv_std_logic_vector(start,6);
      WHEN "100100" => position <= conv_std_logic_vector(start,6);
      WHEN "100101" => position <= conv_std_logic_vector(start,6);
      WHEN "100110" => position <= conv_std_logic_vector(start,6);
      WHEN "100111" => position <= conv_std_logic_vector(start,6);
      WHEN "101000" => position <= conv_std_logic_vector(start,6);
      WHEN "101001" => position <= conv_std_logic_vector(start,6);
      WHEN "101010" => position <= conv_std_logic_vector(start,6);
      WHEN "101011" => position <= conv_std_logic_vector(start,6);
      WHEN "101100" => position <= conv_std_logic_vector(start,6);
      WHEN "101101" => position <= conv_std_logic_vector(start,6);
      WHEN "101110" => position <= conv_std_logic_vector(start,6); 
      WHEN "101111" => position <= conv_std_logic_vector(start,6);      
      WHEN "110000" => position <= conv_std_logic_vector(start,6);
      WHEN "110001" => position <= conv_std_logic_vector(start,6);
      WHEN "110010" => position <= conv_std_logic_vector(start,6);
      WHEN "110011" => position <= conv_std_logic_vector(start,6);
      WHEN "110100" => position <= conv_std_logic_vector(start,6);
      WHEN "110101" => position <= conv_std_logic_vector(start,6);
      WHEN "110110" => position <= conv_std_logic_vector(start,6);
      WHEN "110111" => position <= conv_std_logic_vector(start,6);
      WHEN "111000" => position <= conv_std_logic_vector(start,6);
      WHEN "111001" => position <= conv_std_logic_vector(start,6);
      WHEN "111010" => position <= conv_std_logic_vector(start,6);
      WHEN "111011" => position <= conv_std_logic_vector(start,6);
      WHEN "111100" => position <= conv_std_logic_vector(start,6);
      WHEN "111101" => position <= conv_std_logic_vector(start,6);
      WHEN "111110" => position <= conv_std_logic_vector(start,6); 
      WHEN "111111" => position <= conv_std_logic_vector(start,6);
          
      WHEN others => position <= conv_std_logic_vector(0,6);
          
  END CASE;
               
END PROCESS;    
    
END sss;


LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_RANGE1.VHD                             ***
--***                                             ***
--***   Function: Single Precision Range Reduction***
--***   Core. Output as a fraction of 2PI.        ***
--***                                             ***
--***   22/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_range1 IS
GENERIC (device : integer := 0);
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (8 DOWNTO 1); 
      mantissain : IN STD_LOGIC_VECTOR (23 DOWNTO 1); 

      circle : OUT STD_LOGIC_VECTOR (36 DOWNTO 1);
      negcircle : OUT STD_LOGIC_VECTOR (36 DOWNTO 1) 
     );
END fp_range1;

ARCHITECTURE rtl of fp_range1 IS

  type rangeexponentfftype IS ARRAY (6 DOWNTO 1) OF STD_LOGIC_VECTOR (9 DOWNTO 1);
 
  signal mantissaff : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal mantissadelff : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal mantissamultipliernode : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal mantissamultiplierff : STD_LOGIC_VECTOR (23 DOWNTO 1);
  
  signal exponentff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal mantissaexponentnode : STD_LOGIC_VECTOR (9 DOWNTO 1);
 
  signal leadnode, leadff : STD_LOGIC_VECTOR (5 DOWNTO 1);
  
  signal rangeexponentff : rangeexponentfftype;
  signal negrangeexponentff : STD_LOGIC_VECTOR (9 DOWNTO 1);
  
  signal tableaddressff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal basefractionnode, basefractionff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal incmantissanode, incmantissaff : STD_LOGIC_VECTOR (56 DOWNTO 1);
  signal incexponentnode, incexponentff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal basefractiondelnode, basefractiondelff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  
  signal multipliernode : STD_LOGIC_VECTOR (79 DOWNTO 1);
  signal multipliernormnode : STD_LOGIC_VECTOR (78 DOWNTO 1);
  signal multipliernormff : STD_LOGIC_VECTOR (78 DOWNTO 1);
  
  signal leftrotatenode, rightrotatenode : STD_LOGIC_VECTOR (78 DOWNTO 1);
  signal leftrotateff, rightrotateff : STD_LOGIC_VECTOR (78 DOWNTO 1);
  signal rotatenode : STD_LOGIC_VECTOR (78 DOWNTO 1);
  signal rotateff : STD_LOGIC_VECTOR (78 DOWNTO 1);
  signal selectrotateff : STD_LOGIC;
  signal circlenode : STD_LOGIC_VECTOR (37 DOWNTO 1);
  signal circleff : STD_LOGIC_VECTOR (37 DOWNTO 1);
  
  signal negbasefractiondelnode : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal negbasefractiondelff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal negrotatenode : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal negcirclenode : STD_LOGIC_VECTOR (37 DOWNTO 1);
  signal negcircleff : STD_LOGIC_VECTOR (37 DOWNTO 1);
 
  component fp_clz23 
  PORT (
        mantissa : IN STD_LOGIC_VECTOR (23 DOWNTO 1);
       
        leading : OUT STD_LOGIC_VECTOR (5 DOWNTO 1)    
      );
  end component;
  
  component fp_lsft23  
  PORT (
        inbus : IN STD_LOGIC_VECTOR (23 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (5 DOWNTO 1);

	      outbus : OUT STD_LOGIC_VECTOR (23 DOWNTO 1)
	     );
  end component;
  
  component fp_lsft78  
  PORT (
        inbus : IN STD_LOGIC_VECTOR (78 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);

	      outbus : OUT STD_LOGIC_VECTOR (78 DOWNTO 1)
	     );
  end component;
  
  component fp_rsft78  
  PORT (
        inbus : IN STD_LOGIC_VECTOR (78 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);

	     outbus : OUT STD_LOGIC_VECTOR (78 DOWNTO 1)
	    );
  end component;
 
  component fp_range_table1 
  PORT (
        address : IN STD_LOGIC_VECTOR (8 DOWNTO 1); 
 
        basefraction : OUT STD_LOGIC_VECTOR (36 DOWNTO 1);  
        incmantissa : OUT STD_LOGIC_VECTOR (56 DOWNTO 1);
        incexponent : OUT STD_LOGIC_VECTOR (8 DOWNTO 1)
     );
  end component;

  component fp_mul23x56 IS
  GENERIC (device : integer);
  PORT (  
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (23 DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (56 DOWNTO 1);

        result : OUT STD_LOGIC_VECTOR (79 DOWNTO 1)
  );
  end component;

  component fp_del IS 
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
   end component;
     
BEGIN

    pca: PROCESS (sysclk,reset)
    BEGIN
        
      IF (reset = '1') THEN
      
        FOR k IN 1 TO 23 LOOP
          mantissaff(k) <= '0';
          mantissadelff(k) <= '0';
          mantissamultiplierff(k) <= '0';
        END LOOP;
        exponentff <= "00000000";
        FOR k IN 1 TO 6 LOOP
          rangeexponentff(k)(9 DOWNTO 1) <= "000000000";
        END LOOP;
        negrangeexponentff(9 DOWNTO 1) <= "000000000";
        leadff <= "00000";
        tableaddressff <= "00000000";
        FOR k IN 1 TO 36 LOOP
          basefractionff(k) <= '0';
        END LOOP;
        FOR k IN 1 TO 56 LOOP
          incmantissaff(k) <= '0';
        END LOOP;
        incexponentff <= "00000000";
        FOR k IN 1 TO 78 LOOP
          multipliernormff(k) <= '0';
          leftrotateff(k) <= '0';
          rightrotateff(k) <= '0';
        END LOOP;
        selectrotateff <= '0';
        FOR k IN 1 TO 37 LOOP
          circleff(k) <= '0';
          negcircleff(k) <= '0';
        END LOOP;

      ELSIF (rising_edge(sysclk)) THEN
      
        IF (enable = '1') THEN
            
          mantissaff <= mantissain; -- level 1
          mantissadelff <= mantissaff; -- level 2
          exponentff <= exponentin;  -- level 1
          
          leadff <= leadnode; -- level 2
          mantissamultiplierff <= mantissamultipliernode; -- level 3
          
          tableaddressff <= exponentff; -- level 2
          basefractionff <= basefractionnode; -- level 3
          incmantissaff <= incmantissanode; -- level 3
          incexponentff <= incexponentnode; -- level 3
          
          rangeexponentff(1)(9 DOWNTO 1) <= mantissaexponentnode; -- levels 3,4,5,6,7, and 8
          rangeexponentff(2)(9 DOWNTO 1) <= rangeexponentff(1)(9 DOWNTO 1) - ('0' & incexponentff);
          rangeexponentff(3)(9 DOWNTO 1) <= rangeexponentff(2)(9 DOWNTO 1);
          rangeexponentff(4)(9 DOWNTO 1) <= rangeexponentff(3)(9 DOWNTO 1);
          rangeexponentff(5)(9 DOWNTO 1) <= rangeexponentff(4)(9 DOWNTO 1);
          rangeexponentff(6)(9 DOWNTO 1) <= rangeexponentff(5)(9 DOWNTO 1) - ("00000000" & NOT(multipliernode(79)));
          
          negrangeexponentff <= "100000000" - 
                                (rangeexponentff(5)(9 DOWNTO 1) - 
                                ("00000000" & NOT(multipliernode(79)))); -- level 8
          
          multipliernormff <= multipliernormnode;
          
          leftrotateff <= leftrotatenode;
          rightrotateff <= rightrotatenode;
          rotateff <= rotatenode;
          selectrotateff <= negrangeexponentff(9);
          
          basefractiondelff <= basefractiondelnode;
          negbasefractiondelff <= negbasefractiondelnode;
            
          circleff <= circlenode;
          negcircleff <= negcirclenode;
                
        END IF;
      
      END IF;    
        
    END PROCESS;

    cbfd: fp_del  
    GENERIC MAP (width=>36,pipes=>6)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>basefractionff,
              cc=>basefractiondelnode);

    --turn mantissa fractional part into floating point number
    -- level 1 in
    cclzin: fp_clz23
    PORT MAP (mantissa=>mantissaff,leading=>leadnode);
    
    -- need to do this shift so that both mult inputs normalized, so we can see
    -- if 1 bit mult output normalization required
    -- level 2 in
    csftin: fp_lsft23
    PORT MAP (inbus=>mantissadelff,shift=>leadff,
              outbus=>mantissamultipliernode);
           
    -- exponents (expin, baseexp, incexp) reversed
    -- exponents show shift from 0.9999 posisition
    -- ex: 0.111e3 = 0.000111, 0.111e5 = 0.00000111
    -- if no shift, expin = 23
    -- ex: mantissain = 123, after shift = 0.1111011 (0.96), same as 7
    -- level 2 in
    mantissaexponentnode <= "000010111" - ("0000" & leadff); -- 23 - shift
    
    -- level 2 in
    clut: fp_range_table1 
    PORT MAP (address=>tableaddressff,
              basefraction=>basefractionnode,
              incmantissa=>incmantissanode,
              incexponent=>incexponentnode);
    
    -- 23 x 56 = 79 bits
    -- mantissamulin, incman both in range 0.5 to 0.9999, so result is range 0.25 to 0.999
    -- if < 0.5, shift left and add 1 to exponent
    -- levels 4,5,6,7 
    cmul: fp_mul23x56
    GENERIC MAP(device=>device) 
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              dataaa=>mantissamultiplierff,databb=>incmantissaff,
              result=>multipliernode);  
    
    -- level 7 in
    gma: FOR k IN 1 TO 78 GENERATE
      multipliernormnode(k) <= (multipliernode(k+1) AND multipliernode(79)) OR 
                               (multipliernode(k) AND NOT(multipliernode(79))); 
    END GENERATE;
    
    lftsft: fp_lsft78
    PORT MAP (inbus=>multipliernormff,shift=>rangeexponentff(6)(6 DOWNTO 1),
              outbus=>leftrotatenode);
              
    rgtsft: fp_rsft78
    PORT MAP (inbus=>multipliernormff,shift=>negrangeexponentff(6 DOWNTO 1),
              outbus=>rightrotatenode);
              
    gra: FOR k IN 1 TO 78 GENERATE
      rotatenode(k) <= (leftrotateff(k) AND NOT(selectrotateff)) OR 
                       (rightrotateff(k) AND selectrotateff);
    END GENERATE;
    
    -- use 3-1 adder to round as well?
    
    -- max will be 1.9999, but only interested in fractional part          
    circlenode <= ('0' & basefractiondelff) + ('0' & rotateff(78 DOWNTO 43));
    
    negbasefractiondelnode <= 0 - (basefractiondelnode(36 DOWNTO 1));
    gnra: FOR k IN 1 TO 36 GENERATE
      negrotatenode(k) <= NOT(rotateff(k+42));
    END GENERATE;
    negcirclenode <= ('1' & negbasefractiondelff) + ('1' & negrotatenode) + 1;
    
    -- fractional part of 2pi will be circle(36 DOWNTO 1)
    circle <= circleff(36 DOWNTO 1);
    negcircle <= negcircleff(36 DOWNTO 1);
 
  END rtl;
  
    LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_RANGE_TABLE1.VHD                       ***
--***                                             ***
--***   Function: Single Precision Range Reduction***
--***   Component                                 ***
--***                                             ***
--***   22/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_range_table1 IS
PORT (
      address : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      basefraction : OUT STD_LOGIC_VECTOR (36 DOWNTO 1);
      incmantissa : OUT STD_LOGIC_VECTOR (56 DOWNTO 1);
		  incexponent : OUT STD_LOGIC_VECTOR (8 DOWNTO 1)
     );
END fp_range_table1;

ARCHITECTURE rtl OF fp_range_table1 IS

BEGIN

  pca: PROCESS (address)
  BEGIN
    CASE address IS
      WHEN "01101110" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(0,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(83443,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(42,8);
      WHEN "01101111" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(0,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(166886,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(41,8);
      WHEN "01110000" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(0,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(333772,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(40,8);
      WHEN "01110001" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(0,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(667544,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(39,8);
      WHEN "01110010" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(0,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(1335088,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(38,8);
      WHEN "01110011" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(0,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(2670177,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(37,8);
      WHEN "01110100" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(0,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(5340354,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(36,8);
      WHEN "01110101" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(0,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(10680707,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(35,8);
      WHEN "01110110" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(0,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(21361415,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(34,8);
      WHEN "01110111" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(0,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(42722830,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(33,8);
      WHEN "01111000" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(0,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(85445659,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(32,8);
      WHEN "01111001" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(0,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(170891319,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(31,8);
      WHEN "01111010" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(1,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(73347182,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(30,8);
      WHEN "01111011" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(2,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(146694364,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(29,8);
      WHEN "01111100" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(5,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(24953271,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(28,8);
      WHEN "01111101" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(10,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(49906542,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(27,8);
      WHEN "01111110" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(20,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(99813085,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(26,8);
      WHEN "01111111" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(40,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(199626169,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(25,8);
      WHEN "10000000" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(81,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(130816882,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891319,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(14297640,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(24,8);
      WHEN "10000001" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(162,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(261633765,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(23,8);
      WHEN "10000010" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(69,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(254832074,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(22,8);
      WHEN "10000011" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(139,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(241228692,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(21,8);
      WHEN "10000100" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(23,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(214021927,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(20,8);
      WHEN "10000101" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(47,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(159608398,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(241345352,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(19,8);
      WHEN "10000110" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(95,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(50781341,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(18,8);
      WHEN "10000111" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(190,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(101562681,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(237340088,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(17,8);
      WHEN "10001000" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(124,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(203125362,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(16,8);
      WHEN "10001001" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(249,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(137815268,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(15,8);
      WHEN "10001010" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(243,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(7195081,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(14,8);
      WHEN "10001011" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(230,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(14390161,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(13,8);
      WHEN "10001100" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(204,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(28780322,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(12,8);
      WHEN "10001101" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(152,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(57560644,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(11,8);
      WHEN "10001110" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(48,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(115121288,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(10,8);
      WHEN "10001111" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(96,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(230242576,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(9,8);
      WHEN "10010000" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(193,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(192049697,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240015480,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(8,8);
      WHEN "10010001" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(131,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(115663937,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(7,8);
      WHEN "10010010" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(6,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(231327875,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(6,8);
      WHEN "10010011" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(13,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(194220293,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(5,8);
      WHEN "10010100" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(27,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(120005131,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(4,8);
      WHEN "10010101" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(54,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(240010261,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(3,8);
      WHEN "10010110" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(109,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(211585066,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(2,8);
      WHEN "10010111" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(219,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(154734677,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "10011000" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(183,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(41033897,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(170891318,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(240010256,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "10011001" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(110,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(82067795,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(146694363,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(154734672,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "10011010" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(220,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(164135589,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(146694363,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(154734680,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "10011011" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(185,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(59835722,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(199626169,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(59835760,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(3,8);
      WHEN "10011100" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(114,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(119671445,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(199626169,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(59835712,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(2,8);
      WHEN "10011101" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(228,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(239342890,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(199626169,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(59835736,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "10011110" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(201,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(210250324,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(199626169,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(59835728,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "10011111" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(147,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(152065192,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(261633764,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(239342888,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "10100000" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(39,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(35694928,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(261633764,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(239342888,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "10100001" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(78,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(71389856,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(254832073,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(210250312,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "10100010" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(156,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(142779712,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(241228691,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(152065192,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "10100011" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(57,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(17123967,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(214021927,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(35694928,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "10100100" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(114,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(34247934,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(159608398,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(71389856,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "10100101" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(228,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(68495868,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(203125362,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(34247944,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(2,8);
      WHEN "10100110" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(200,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(136991736,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(203125362,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(34247920,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "10100111" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(145,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(5548017,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(203125362,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(34247944,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "10101000" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(34,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(11096033,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(137815268,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(68495872,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "10101001" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(68,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(22192066,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(230242576,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(88768104,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(5,8);
      WHEN "10101010" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(136,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(44384133,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(230242576,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(88768184,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(4,8);
      WHEN "10101011" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(16,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(88768266,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(230242576,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(88768288,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(3,8);
      WHEN "10101100" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(32,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(177536532,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(230242576,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(88768264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(2,8);
      WHEN "10101101" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(65,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(86637607,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(230242576,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(88768248,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "10101110" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(130,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(173275215,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(230242576,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(88768264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "10101111" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(5,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(78114973,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(192049696,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(177536536,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "10110000" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(10,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(156229947,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(231327874,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(173275224,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "10110001" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(21,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(44024437,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(231327874,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(173275224,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "10110010" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(42,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(88048875,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(194220293,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(78114968,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "10110011" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(84,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(176097750,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(240010261,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(44024424,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "10110100" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(169,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(83760044,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(240010261,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(44024440,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "10110101" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(82,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(167520088,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(211585066,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(88048872,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "10110110" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(165,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(66604720,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(154734676,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(176097752,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "10110111" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(74,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(133209439,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(164135589,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(66604720,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(2,8);
      WHEN "10111000" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(148,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(266418879,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(164135589,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(66604728,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "10111001" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(41,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(264402301,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(164135589,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(66604728,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "10111010" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(83,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(260369146,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(239342889,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(264402312,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(2,8);
      WHEN "10111011" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(167,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(252302836,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(239342889,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(264402288,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "10111100" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(79,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(236170217,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(239342889,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(264402296,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "10111101" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(159,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(203904978,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(210250323,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(260369144,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "10111110" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(63,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(139374500,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(152065191,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(252302864,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "10111111" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(127,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(10313544,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(142779711,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(139374496,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(2,8);
      WHEN "11000000" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(254,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(20627088,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(142779711,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(139374496,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "11000001" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(252,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(41254175,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(142779711,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(139374496,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11000010" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(248,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(82508351,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(136991736,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(82508384,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(3,8);
      WHEN "11000011" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(240,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(165016701,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(136991736,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(82508344,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(2,8);
      WHEN "11000100" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(225,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(61597947,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(136991736,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(82508368,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "11000101" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(194,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(123195893,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(136991736,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(82508360,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11000110" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(132,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(246391786,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(177536531,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(180260912,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(5,8);
      WHEN "11000111" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(9,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(224348117,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(177536531,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(180260792,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(4,8);
      WHEN "11001000" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(19,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(180260778,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(177536531,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(180260792,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(3,8);
      WHEN "11001001" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(39,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(92086099,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(177536531,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(180260792,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(2,8);
      WHEN "11001010" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(78,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(184172199,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(177536531,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(180260792,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "11001011" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(157,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(99908941,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(177536531,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(180260776,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11001100" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(58,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(199817882,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(173275214,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(184172200,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "11001101" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(117,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(131200309,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(173275214,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(184172200,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11001110" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(234,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(262400618,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(156229946,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(199817896,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "11001111" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(213,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(256365779,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(156229946,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(199817880,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11010000" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(171,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(244296103,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(176097749,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(256365776,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(2,8);
      WHEN "11010001" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(87,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(220156750,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(176097749,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(256365792,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "11010010" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(175,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(171878044,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(176097749,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(256365776,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11010011" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(95,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(75320631,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(167520087,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(220156768,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "11010100" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(190,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(150641263,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(167520087,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(220156760,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11010101" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(125,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(32847070,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(266418878,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(150641264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(2,8);
      WHEN "11010110" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(250,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(65694140,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(266418878,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(150641280,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "11010111" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(244,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(131388279,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(266418878,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(150641264,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11011000" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(232,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(262776558,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(264402301,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(32847064,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11011001" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(209,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(257117660,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(260369146,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(65694136,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11011010" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(163,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(245799864,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(252302836,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(131388288,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11011011" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(71,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(223164272,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(236170216,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(262776560,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11011100" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(143,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(177893088,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(203904977,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(257117656,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11011101" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(31,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(87350721,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(139374499,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(245799872,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11011110" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(62,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(174701442,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(165016701,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(80967568,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(4,8);
      WHEN "11011111" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(125,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(80967427,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(165016701,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(80967448,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(3,8);
      WHEN "11100000" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(250,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(161934855,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(165016701,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(80967448,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(2,8);
      WHEN "11100001" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(245,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(55434254,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(165016701,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(80967448,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "11100010" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(234,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(110868507,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(165016701,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(80967424,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11100011" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(212,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(221737015,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(246391786,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(110868472,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(2,8);
      WHEN "11100100" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(169,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(175038574,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(246391786,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(110868512,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "11100101" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(83,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(81641691,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(246391786,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(110868528,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11100110" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(166,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(163283383,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(224348116,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(221737016,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11100111" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(77,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(58131310,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(180260777,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(175038576,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11101000" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(154,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(116262619,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(184172198,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(163283376,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "11101001" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(52,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(232525238,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(184172198,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(163283384,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11101010" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(105,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(196615020,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(199817882,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(116262632,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "11101011" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(211,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(124794585,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(199817882,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(116262624,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11101100" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(166,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(249589169,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(262400617,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(196615040,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "11101101" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(77,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(230742883,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(262400617,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(196615016,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11101110" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(155,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(193050309,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(256365779,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(124794584,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11101111" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(55,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(117665162,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(244296102,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(249589176,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11110000" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(110,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(235330325,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(220156749,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(230742864,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11110001" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(221,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(202225193,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(171878043,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(193050312,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11110010" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(187,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(136014931,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(150641262,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(235330336,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "11110011" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(119,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(3594405,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(150641262,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(235330328,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11110100" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(238,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(7188811,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(262776558,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(7188776,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(3,8);
      WHEN "11110101" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(220,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(14377622,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(262776558,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(7188816,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(2,8);
      WHEN "11110110" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(184,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(28755243,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(262776558,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(7188816,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "11110111" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(112,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(57510486,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(262776558,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(7188816,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11111000" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(224,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(115020973,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(257117660,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(14377624,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11111001" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(192,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(230041946,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(245799864,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(28755224,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11111010" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(129,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(191648435,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(223164272,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(57510496,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11111011" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(3,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(114861414,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(177893088,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(115020976,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11111100" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(6,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(229722829,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(174701441,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(191648432,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "11111101" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(13,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(191010201,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(174701441,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(191648440,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN "11111110" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(27,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(113584946,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(161934854,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(229722832,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(1,8);
      WHEN "11111111" => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(54,8);
                         basefraction(28 DOWNTO 1) <= conv_std_logic_vector(227169893,28);
                         incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(161934854,28);
                         incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(229722824,28);
                         incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
      WHEN others => basefraction(36 DOWNTO 29) <= conv_std_logic_vector(0,8);
                     basefraction(28 DOWNTO 1) <= conv_std_logic_vector(0,28);
                     incmantissa(56 DOWNTO 29) <= conv_std_logic_vector(0,28);
                     incmantissa(28 DOWNTO 1) <= conv_std_logic_vector(0,28);
                     incexponent(8 DOWNTO 1) <= conv_std_logic_vector(0,8);
    END CASE;
  END PROCESS;

END rtl;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_RSFT32X5.VHD                           ***
--***                                             ***
--***   Function: Single Precision Right Shift    ***
--***                                             ***
--***   22/02/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_rsft32x5 IS 
PORT (
      inbus : IN STD_LOGIC_VECTOR (32 DOWNTO 1);
      shift : IN STD_LOGIC_VECTOR (5 DOWNTO 1);
      outbus : OUT STD_LOGIC_VECTOR (32 DOWNTO 1)
    );
END fp_rsft32x5;

ARCHITECTURE rtl OF fp_rsft32x5 IS

  signal rightone, righttwo, rightthr : STD_LOGIC_VECTOR (32 DOWNTO 1);
            
BEGIN

  gra: FOR k IN 1 TO 29 GENERATE
    rightone(k) <= (inbus(k)   AND NOT(shift(2)) AND NOT(shift(1))) OR
                   (inbus(k+1) AND NOT(shift(2)) AND     shift(1)) OR
                   (inbus(k+2) AND     shift(2)  AND NOT(shift(1))) OR
                   (inbus(k+3) AND     shift(2)  AND     shift(1));
  END GENERATE;
  rightone(30) <= (inbus(30) AND NOT(shift(2)) AND NOT(shift(1))) OR
                  (inbus(31) AND NOT(shift(2)) AND     shift(1)) OR
                  (inbus(32) AND     shift(2)  AND NOT(shift(1))); 
  rightone(31) <= (inbus(31) AND NOT(shift(2)) AND NOT(shift(1))) OR
                  (inbus(32) AND NOT(shift(2)) AND     shift(1));
  rightone(32) <=  inbus(32) AND NOT(shift(2)) AND NOT(shift(1));
  
  grb: FOR k IN 1 TO 20 GENERATE
    righttwo(k) <= (rightone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                   (rightone(k+4)  AND NOT(shift(4)) AND     shift(3)) OR
                   (rightone(k+8)  AND     shift(4)  AND NOT(shift(3))) OR
                   (rightone(k+12) AND     shift(4)  AND     shift(3)); 
  END GENERATE;
  grc: FOR k IN 21 TO 24 GENERATE
    righttwo(k) <= (rightone(k)   AND NOT(shift(4)) AND NOT(shift(3))) OR
                   (rightone(k+4) AND NOT(shift(4)) AND     shift(3)) OR
                   (rightone(k+8) AND     shift(4)  AND NOT(shift(3))); 
  END GENERATE; 
  grd: FOR k IN 25 TO 28 GENERATE
    righttwo(k) <= (rightone(k)   AND NOT(shift(4)) AND NOT(shift(3))) OR
                   (rightone(k+4) AND NOT(shift(4)) AND     shift(3));
  END GENERATE; 
  gre: FOR k IN 29 TO 32 GENERATE
    righttwo(k) <= (rightone(k)   AND NOT(shift(4)) AND NOT(shift(3)));
  END GENERATE;  
  
  grf: FOR k IN 1 TO 16 GENERATE
    rightthr(k) <= (righttwo(k)    AND NOT(shift(5))) OR 
                   (righttwo(k+16) AND shift(5));
  END GENERATE;
  grg: FOR k IN 17 TO 32 GENERATE
    rightthr(k) <= (righttwo(k)    AND NOT(shift(5)));
  END GENERATE;
  
  outbus <= rightthr;        
            
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_RSFT36.VHD                             ***
--***                                             ***
--***   Function: 36 bit Unsigned Right Shift     ***
--***                                             ***
--***   22/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_rsft36 IS 
PORT (
      inbus : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
      shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);

	   outbus : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
	  );
END fp_rsft36;

ARCHITECTURE rtl OF fp_rsft36 IS
  
  signal levzip, levone, levtwo, levthr : STD_LOGIC_VECTOR (36 DOWNTO 1);
    
BEGIN
        
  levzip <= inbus;
  
  -- shift by 0,1,2,3
  gaa: FOR k IN 1 TO 33 GENERATE
    levone(k) <= (levzip(k)   AND NOT(shift(2)) AND NOT(shift(1))) OR
                 (levzip(k+1) AND NOT(shift(2)) AND     shift(1)) OR
                 (levzip(k+2) AND     shift(2)  AND NOT(shift(1))) OR
                 (levzip(k+3) AND     shift(2)  AND     shift(1)); 
  END GENERATE;
  levone(34) <=  (levzip(34) AND NOT(shift(2)) AND NOT(shift(1))) OR
                 (levzip(35) AND NOT(shift(2)) AND     shift(1)) OR
                 (levzip(36) AND     shift(2)  AND NOT(shift(1)));
  levone(35) <=  (levzip(35) AND NOT(shift(2)) AND NOT(shift(1))) OR
                 (levzip(36) AND NOT(shift(2)) AND     shift(1));
  levone(36) <= levzip(36)   AND NOT(shift(2)) AND NOT(shift(1));
                              
  -- shift by 0,4,8,12
  gba: FOR k IN 1 TO 24 GENERATE
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                 (levone(k+4)  AND NOT(shift(4)) AND     shift(3)) OR
                 (levone(k+8)  AND     shift(4)  AND NOT(shift(3))) OR
                 (levone(k+12) AND     shift(4)  AND     shift(3)); 
  END GENERATE;
  gbb: FOR k IN 25 TO 28 GENERATE
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                 (levone(k+4)  AND NOT(shift(4)) AND     shift(3)) OR
                 (levone(k+8)  AND     shift(4)  AND NOT(shift(3)));
  END GENERATE;
  gbc: FOR k IN 29 TO 32 GENERATE
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                 (levone(k+4)  AND NOT(shift(4)) AND     shift(3));
  END GENERATE;
  gbd: FOR k IN 33 TO 36 GENERATE
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3)));
  END GENERATE;
  
  gca: FOR k IN 1 TO 4 GENERATE
    levthr(k) <= (levtwo(k)    AND NOT(shift(6)) AND NOT(shift(5))) OR
                 (levtwo(k+16) AND NOT(shift(6)) AND     shift(5)) OR
                 (levtwo(k+32) AND     shift(6));
  END GENERATE;
  gcb: FOR k IN 5 TO 20 GENERATE
    levthr(k) <= (levtwo(k)    AND NOT(shift(6)) AND NOT(shift(5))) OR
                 (levtwo(k+16) AND NOT(shift(6)) AND     shift(5));
  END GENERATE;
  gcc: FOR k IN 21 TO 36 GENERATE
    levthr(k) <= (levtwo(k)    AND NOT(shift(6)) AND NOT(shift(5)));
  END GENERATE;

  outbus <= levthr;
  
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_RSFT56X20.VHD                          ***
--***                                             ***
--***   Function: 56 bit Unsigned Right Shift     ***
--***   (Maximum 20 bit Shift)                    ***
--***                                             ***
--***   22/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_rsft56x20 IS 
PORT (
      inbus : IN STD_LOGIC_VECTOR (56 DOWNTO 1);
      shift : IN STD_LOGIC_VECTOR (5 DOWNTO 1);

	   outbus : OUT STD_LOGIC_VECTOR (56 DOWNTO 1)
	  );
END fp_rsft56x20;

ARCHITECTURE rtl OF fp_rsft56x20 IS
  
  signal levzip, levone, levtwo, levthr : STD_LOGIC_VECTOR (56 DOWNTO 1);
    
BEGIN
        
  levzip <= inbus;
  
  -- shift by 0,1,2,3
  gaa: FOR k IN 1 TO 53 GENERATE
    levone(k) <= (levzip(k)   AND NOT(shift(2)) AND NOT(shift(1))) OR
                 (levzip(k+1) AND NOT(shift(2)) AND     shift(1)) OR
                 (levzip(k+2) AND     shift(2)  AND NOT(shift(1))) OR
                 (levzip(k+3) AND     shift(2)  AND     shift(1)); 
  END GENERATE;
  levone(54) <=  (levzip(54) AND NOT(shift(2)) AND NOT(shift(1))) OR
                 (levzip(55) AND NOT(shift(2)) AND     shift(1)) OR
                 (levzip(56) AND     shift(2)  AND NOT(shift(1)));
  levone(55) <=  (levzip(55) AND NOT(shift(2)) AND NOT(shift(1))) OR
                 (levzip(56) AND NOT(shift(2)) AND     shift(1));
  levone(56) <= levzip(56)   AND NOT(shift(2)) AND NOT(shift(1));
                              
  -- shift by 0,4,8,12
  gba: FOR k IN 1 TO 44 GENERATE
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                 (levone(k+4)  AND NOT(shift(4)) AND     shift(3)) OR
                 (levone(k+8)  AND     shift(4)  AND NOT(shift(3))) OR
                 (levone(k+12) AND     shift(4)  AND     shift(3)); 
  END GENERATE;
  gbb: FOR k IN 45 TO 48 GENERATE
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                 (levone(k+4)  AND NOT(shift(4)) AND     shift(3)) OR
                 (levone(k+8)  AND     shift(4)  AND NOT(shift(3)));
  END GENERATE;
  gbc: FOR k IN 49 TO 52 GENERATE
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3))) OR
                 (levone(k+4)  AND NOT(shift(4)) AND     shift(3));
  END GENERATE;
  gbd: FOR k IN 53 TO 56 GENERATE
    levtwo(k) <= (levone(k)    AND NOT(shift(4)) AND NOT(shift(3)));
  END GENERATE;
  
  gca: FOR k IN 1 TO 40 GENERATE
    levthr(k) <= (levtwo(k)    AND NOT(shift(5))) OR
                 (levtwo(k+16) AND     shift(5));
  END GENERATE;
  gcc: FOR k IN 41 TO 56 GENERATE
    levthr(k) <= (levtwo(k)    AND NOT(shift(5)));
  END GENERATE;

  outbus <= levthr;
  
END rtl;

LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_RSFT78.VHD                             ***
--***                                             ***
--***   Function: 78 bit Arithmetic Right Shift   ***
--***                                             ***
--***   22/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_rsft78 IS
PORT (
      inbus : IN STD_LOGIC_VECTOR (78 DOWNTO 1); 
      shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1); 

      outbus : OUT STD_LOGIC_VECTOR (78 DOWNTO 1)
     );
END fp_rsft78;

ARCHITECTURE rtl of fp_rsft78 IS

  signal levzip, levone, levtwo : STD_LOGIC_VECTOR (78 DOWNTO 1);
  signal levthr, levfor, levfiv : STD_LOGIC_VECTOR (78 DOWNTO 1);
  signal levsix : STD_LOGIC_VECTOR (78 DOWNTO 1);
  
BEGIN

  levzip <= inbus;
 
  gaa: FOR k IN 1 TO 77 GENERATE
    levone(k) <= (levzip(k) AND NOT(shift(1))) OR (levzip(k+1) AND shift(1));
  END GENERATE;
  levone(78) <= levzip(78) AND NOT(shift(1));
  
  gba: FOR k IN 1 TO 76 GENERATE
    levtwo(k) <= (levone(k) AND NOT(shift(2))) OR (levone(k+2) AND shift(2));
  END GENERATE;
  levtwo(77) <= levone(77) AND NOT(shift(2));
  levtwo(78) <= levone(78) AND NOT(shift(2));
  
  gca: FOR k IN 1 TO 74 GENERATE
    levthr(k) <= (levtwo(k) AND NOT(shift(3))) OR (levtwo(k+4) AND shift(3));
  END GENERATE;
  gcb: FOR k IN 75 TO 78 GENERATE
    levthr(k) <= levtwo(k) AND NOT(shift(3));
  END GENERATE;
  
  gda: FOR k IN 1 TO 70 GENERATE
    levfor(k) <= (levthr(k) AND NOT(shift(4))) OR (levthr(k+8) AND shift(4));
  END GENERATE;
  gdb: FOR k IN 71 TO 78 GENERATE
    levfor(k) <= levthr(k) AND NOT(shift(4));
  END GENERATE;
 
  gea: FOR k IN 1 TO 62 GENERATE
    levfiv(k) <= (levfor(k) AND NOT(shift(5))) OR (levfor(k+16) AND shift(5));
  END GENERATE;
  geb: FOR k IN 63 TO 78 GENERATE
    levfiv(k) <= levfor(k) AND NOT(shift(5));
  END GENERATE;
   
  gfa: FOR k IN 1 TO 46 GENERATE
    levsix(k) <= (levfiv(k) AND NOT(shift(6))) OR (levfiv(k+32) AND shift(6));
  END GENERATE;
  gfb: FOR k IN 47 TO 78 GENERATE
    levsix(k) <= levfiv(k) AND NOT(shift(6));
  END GENERATE;
    
  outbus <= levsix;
  
END;


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_SGN_MUL3S.VHD                          ***
--***                                             ***
--***   Function: Signed Multiplier - 3 Pipe      ***
--***   Stages                                    ***
--***                                             ***
--***   22/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_sgn_mul3s IS
GENERIC (
         widthaa : positive := 18;
         widthbb : positive := 18;
         widthcc : positive := 36
        );
PORT
	(
    sysclk : IN STD_LOGIC;
    reset : IN STD_LOGIC;
    enable : IN STD_LOGIC;
    dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
    databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1);

	 result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
	);
END fp_sgn_mul3s;

ARCHITECTURE SYN OF fp_sgn_mul3s IS

	SIGNAL resultnode	: STD_LOGIC_VECTOR (widthaa+widthbb DOWNTO 1);

  component altmult_add
	GENERIC (
		addnsub_multiplier_aclr1		: STRING;
		addnsub_multiplier_pipeline_aclr1		: STRING;
		addnsub_multiplier_pipeline_register1		: STRING;
		addnsub_multiplier_register1		: STRING;
		dedicated_multiplier_circuitry		: STRING;
		input_aclr_a0		: STRING;
		input_aclr_b0		: STRING;
		input_register_a0		: STRING;
		input_register_b0		: STRING;
		input_source_a0		: STRING;
		input_source_b0		: STRING;
		intended_device_family		: STRING;
		lpm_type		: STRING;
		multiplier1_direction		: STRING;
		multiplier_aclr0		: STRING;
		multiplier_register0		: STRING;
		number_of_multipliers		: NATURAL;
		output_aclr		: STRING;
		output_register		: STRING;
		port_addnsub1		: STRING;
		port_signa		: STRING;
		port_signb		: STRING;
		representation_a		: STRING;
		representation_b		: STRING;
		signed_aclr_a		: STRING;
		signed_aclr_b		: STRING;
		signed_pipeline_aclr_a		: STRING;
		signed_pipeline_aclr_b		: STRING;
		signed_pipeline_register_a		: STRING;
		signed_pipeline_register_b		: STRING;
		signed_register_a		: STRING;
		signed_register_b		: STRING;
		width_a		: NATURAL;
		width_b		: NATURAL;
		width_result		: NATURAL
	);
	PORT (
			dataa	: IN STD_LOGIC_VECTOR (widthaa-1 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (widthbb-1 DOWNTO 0);
			clock0	: IN STD_LOGIC ;
			aclr3	: IN STD_LOGIC ;
			ena0	: IN STD_LOGIC ;
			result	: OUT STD_LOGIC_VECTOR (widthaa+widthbb-1 DOWNTO 0)
	);
	end component;

BEGIN

  mulone : altmult_add
  GENERIC MAP (
		addnsub_multiplier_aclr1 => "ACLR3",
		addnsub_multiplier_pipeline_aclr1 => "ACLR3",
		addnsub_multiplier_pipeline_register1 => "CLOCK0",
		addnsub_multiplier_register1 => "CLOCK0",
		dedicated_multiplier_circuitry => "AUTO",
		input_aclr_a0 => "ACLR3",
		input_aclr_b0 => "ACLR3",
		input_register_a0 => "CLOCK0",
		input_register_b0 => "CLOCK0",
		input_source_a0 => "DATAA",
		input_source_b0 => "DATAB",
		intended_device_family => "Stratix II",
		lpm_type => "altmult_add",
		multiplier1_direction => "ADD",
		multiplier_aclr0 => "ACLR3",
		multiplier_register0 => "CLOCK0",
		number_of_multipliers => 1,
		output_aclr => "ACLR3",
		output_register => "CLOCK0",
		port_addnsub1 => "PORT_UNUSED",
		port_signa => "PORT_UNUSED",
		port_signb => "PORT_UNUSED",
		representation_a => "SIGNED",
		representation_b => "SIGNED",
		signed_aclr_a => "ACLR3",
		signed_aclr_b => "ACLR3",
		signed_pipeline_aclr_a => "ACLR3",
		signed_pipeline_aclr_b => "ACLR3",
		signed_pipeline_register_a => "CLOCK0",
		signed_pipeline_register_b => "CLOCK0",
		signed_register_a => "CLOCK0",
		signed_register_b => "CLOCK0",
		width_a => widthaa,
		width_b => widthbb,
		width_result => widthaa+widthbb
	)
	PORT MAP (
		dataa => dataaa,
		datab => databb,
		clock0 => sysclk,
		aclr3 => reset,
		ena0 => enable,
		result => resultnode
	);

  result <= resultnode(widthaa+widthbb DOWNTO widthaa+widthbb-widthcc+1);
  
END SYN;

LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_SIN.VHD                               ***
--***                                             ***
--***   Function: Single Precision SIN Core       ***
--***                                             ***
--***   10/01/10 ML                               ***
--***                                             ***
--***   (c) 2010 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** 1. Input < 0.5 radians, take cos(pi/2-input)***
--*** 2. latency = depth + range_depth (11) + 7   ***
--*** (1 more than cos)                           ***
--***************************************************

ENTITY fp_sin IS
GENERIC (
          device : integer := 0;
          width : positive := 30;
          depth : positive := 18;
          indexpoint : positive := 2
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (8 DOWNTO 1); 
      mantissain : IN STD_LOGIC_VECTOR (23 DOWNTO 1); 

      signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (8 DOWNTO 1); 
      mantissaout : OUT STD_LOGIC_VECTOR (23 DOWNTO 1) 
     );
END fp_sin;

ARCHITECTURE rtl of fp_sin IS

  constant cordic_width : positive := width;
  constant cordic_depth : positive := depth;
  constant range_depth : positive := 11;

  signal piovertwo : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal zerovec : STD_LOGIC_VECTOR (36 DOWNTO 1);

  signal input_number : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal input_number_delay : STD_LOGIC_VECTOR (32 DOWNTO 1);
  signal exponentinff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal exponentcheck : STD_LOGIC_VECTOR (9 DOWNTO 1);
  
  -- range reduction
  signal circle : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal negcircle : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal quadrantsign, quadrantselect : STD_LOGIC;
  signal positive_quadrant, negative_quadrant : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal fraction_quadrant : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal one_term : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal quadrant : STD_LOGIC_VECTOR (34 DOWNTO 1);
  
  -- circle to radians mult
  signal radiansnode : STD_LOGIC_VECTOR (cordic_width DOWNTO 1);
  signal indexcheck : STD_LOGIC_VECTOR (16 DOWNTO 1);
  signal indexbit : STD_LOGIC;
  
  signal signinff : STD_LOGIC_VECTOR (range_depth DOWNTO 1);
  signal selectoutputff : STD_LOGIC_VECTOR (range_depth+cordic_depth+5 DOWNTO 1);
  signal signcalcff : STD_LOGIC_VECTOR (cordic_depth+6 DOWNTO 1);
  signal quadrant_sumff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal select_sincosff : STD_LOGIC_VECTOR (4 DOWNTO 1);

  signal fixed_sincos : STD_LOGIC_VECTOR (cordic_width DOWNTO 1);
  signal fixed_sincosnode : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal fixed_sincosff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  
  signal countnode : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal countff : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal mantissanormnode : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal mantissanormff : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal exponentnormnode : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal exponentnormff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal overflownode : STD_LOGIC_VECTOR (24 DOWNTO 1);
  signal mantissaoutff : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal exponentoutff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal signoutff : STD_LOGIC;
  
  component fp_range1
  GENERIC (device : integer);
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        signin : IN STD_LOGIC;
        exponentin : IN STD_LOGIC_VECTOR (8 DOWNTO 1); 
        mantissain : IN STD_LOGIC_VECTOR (23 DOWNTO 1); 

        circle : OUT STD_LOGIC_VECTOR (36 DOWNTO 1);
        negcircle : OUT STD_LOGIC_VECTOR (36 DOWNTO 1) 
  );
  end component;
   
  component fp_cordic_m1
  GENERIC (
         width : positive := 36;
         depth : positive := 20;
         indexpoint : positive := 2
        );  
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        radians : IN STD_LOGIC_VECTOR (width DOWNTO 1); --'0'&[width-1:1]   
        indexbit : IN STD_LOGIC;   
        sincosbit : IN STD_LOGIC;

        sincos : OUT STD_LOGIC_VECTOR (width DOWNTO 1)     
       );
  end component;

  component fp_clz36 IS
  PORT (
        mantissa : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
      
        leading : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
       );
  end component;

  component fp_lsft36 IS 
  PORT (
        inbus : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);

        outbus : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
  );
  end component;

  component fp_fxmul
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36;
           pipes : positive := 1;
           accuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 0
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1); 
      
        result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
       );
  end component;
   
  component fp_del IS
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
   end component;
   
  BEGIN
    
    -- pi/2 = 1.57
    piovertwo <= x"c90fdaa22";
  
    zerovec <= x"000000000";
    
    --*** SIN(X) = X when exponent < 115 ***
    input_number <= signin & exponentin & mantissain; 
    
    -- level 1 in, level range_depth+cordic_depth+7 out
    cdin: fp_del 
    GENERIC MAP (width=>32,pipes=>range_depth+cordic_depth+6)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>input_number,
              cc=>input_number_delay);
              
    --*** RANGE REDUCTION ***
    crr: fp_range1
    GENERIC MAP(device=>device)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              signin=>signin,exponentin=>exponentin,mantissain=>mantissain,
              circle=>circle,negcircle=>negcircle); 

    quadrantsign <= circle(36); -- sin negative in quadrants 3&4
    quadrantselect <= circle(35); -- sin (1-x) in quadants 2&4

    gra: FOR k IN 1 TO 34 GENERATE
      quadrant(k) <= (circle(k) AND NOT(quadrantselect)) OR
                     (negcircle(k) AND quadrantselect);
    END GENERATE;   
    
    -- if quadrant >0.5 (when quadrant(34) = 1), use quadrant, else use 1-quadrant, and take cos rather than sin
    positive_quadrant <= '0' & quadrant & '0';
    gnqa: FOR k IN 1 TO 36 GENERATE
      negative_quadrant(k) <= NOT(positive_quadrant(k));
      fraction_quadrant(k) <= (positive_quadrant(k) AND quadrant(34)) OR
                              (negative_quadrant(k) AND NOT(quadrant(34)));
    END GENERATE;

    one_term <= NOT(quadrant(34)) & zerovec(35 DOWNTO 1); -- 0 if positive quadrant
      
    pfa: PROCESS (sysclk,reset)
    BEGIN        
      IF (reset = '1') THEN
          
        FOR k IN 1 TO range_depth LOOP
          signinff(k) <= '0';
        END LOOP;
        FOR k IN 1 TO cordic_depth+6 LOOP
          signcalcff(k) <= '0';
        END LOOP;
        FOR k IN 1 TO 8 LOOP
          exponentinff(k) <= '0';
        END LOOP;
        FOR k IN 1 TO range_depth+cordic_depth+5 LOOP
          selectoutputff(k) <= '0';
        END LOOP;
        FOR k IN 1 TO 36 LOOP
          quadrant_sumff(k) <= '0';
        END LOOP;
        FOR k IN 1 TO 4 LOOP
          select_sincosff(k) <= '0';
        END LOOP;
 
      ELSIF (rising_edge(sysclk)) THEN
         
        IF (enable = '1') THEN
        
          signinff(1) <= signin;
          FOR k IN 2 TO range_depth LOOP
            signinff(k) <= signinff(k-1);
          END LOOP;
          -- level range_depth+1 to range_depth+cordic_depth+6
          signcalcff(1) <= quadrantsign XOR signinff(range_depth); 
          FOR k IN 2 TO cordic_depth+6 LOOP
            signcalcff(k) <= signcalcff(k-1);
          END LOOP;
          
          exponentinff <= exponentin; -- level 1
          selectoutputff(1) <= exponentcheck(9); -- level 2 to range_depth+cordic_depth+6
          FOR k IN 2 TO range_depth+cordic_depth+5 LOOP
            selectoutputff(k) <= selectoutputff(k-1);
          END LOOP;
          
          -- range 0-0.9999
          quadrant_sumff <= one_term + fraction_quadrant + NOT(quadrant(34)); -- level range_depth+1
          
          -- level range depth+1 to range_depth+4 
          select_sincosff(1) <= quadrant(34);
          FOR k IN 2 TO 4 LOOP
            select_sincosff(k) <= select_sincosff(k-1);
          END LOOP;
   
        END IF;
         
      END IF;
        
    END PROCESS;
    
    -- if exponent < 115, sin = input
    exponentcheck <= ('0' & exponentinff) - ('0' & x"73");

    -- levels range_depth+2,3,4
    cmul: fp_fxmul  
    GENERIC MAP (widthaa=>36,widthbb=>36,widthcc=>cordic_width,
                 pipes=>3,synthesize=>1)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              dataaa=>quadrant_sumff,databb=>piovertwo,
              result=>radiansnode);
                    
    indexcheck(1) <= radiansnode(cordic_width-1);
    gica: FOR k IN 2 TO 16 GENERATE
      indexcheck(k) <= indexcheck(k-1) OR radiansnode(cordic_width-k);
    END GENERATE;
    -- for safety, give an extra bit of space
    indexbit <= NOT(indexcheck(indexpoint+1));
   
    ccc: fp_cordic_m1
    GENERIC MAP (width=>cordic_width,depth=>cordic_depth,indexpoint=>indexpoint)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              radians=>radiansnode,
              indexbit=>indexbit,
              sincosbit=>select_sincosff(4),
              sincos=>fixed_sincos);
   
    gfxa: IF (width < 36) GENERATE
      fixed_sincosnode <= fixed_sincos & zerovec(36-width DOWNTO 1);
    END GENERATE;
    gfxb: IF (width = 36) GENERATE
      fixed_sincosnode <= fixed_sincos;
    END GENERATE;
    
    clz: fp_clz36
    PORT MAP (mantissa=>fixed_sincosnode,leading=>countnode);
        
    sft: fp_lsft36  
    PORT MAP (inbus=>fixed_sincosff,shift=>countff,
              outbus=>mantissanormnode);
    
    -- maximum sin or cos = 1.0 = 1.0e127 single precision
    -- 1e128 - 1 (leading one) gives correct number
    exponentnormnode <= "10000000" - ("00" & countff); 
    
    overflownode(1) <= mantissanormnode(12);
    gova: FOR k IN 2 TO 24 GENERATE
      overflownode(k) <= mantissanormnode(k+11) AND overflownode(k-1);
    END GENERATE;
    
    -- OUTPUT
    poa: PROCESS (sysclk,reset)
    BEGIN
        
      IF (reset = '1') THEN
          
        FOR k IN 1 TO 36 LOOP
          fixed_sincosff(k) <= '0';
        END LOOP;
        countff <= "000000";
        FOR k IN 1 TO 23 LOOP
          mantissanormff(k) <= '0';
          mantissaoutff(k) <= '0';
        END LOOP;
        FOR k IN 1 TO 8 LOOP
          exponentnormff(k) <= '0';
          exponentoutff(k) <= '0';
        END LOOP;
        signoutff <= '0';

      ELSIF (rising_edge(sysclk)) THEN
          
        IF (enable = '1') THEN
           
          fixed_sincosff <= fixed_sincosnode; -- level range_depth+cordic_depth+5
          countff <= countnode; -- level range_depth+4+cordic_depth+5

          -- level range_depth+cordic_depth+6
          mantissanormff <= mantissanormnode(35 DOWNTO 13) + mantissanormnode(12);
          exponentnormff <= exponentnormnode(8 DOWNTO 1) + overflownode(24);
          
          -- level range_depth+cordic_depth+7         
          FOR k IN 1 TO 23 LOOP
            mantissaoutff(k) <= (mantissanormff(k) AND NOT(selectoutputff(range_depth+cordic_depth+5))) OR
                                (input_number_delay(k) AND selectoutputff(range_depth+cordic_depth+5));
          END LOOP;
          FOR k IN 1 TO 8 LOOP
            exponentoutff(k) <= (exponentnormff(k) AND NOT(selectoutputff(range_depth+cordic_depth+5))) OR
                                (input_number_delay(k+23) AND selectoutputff(range_depth+cordic_depth+5));
          END LOOP;
          signoutff <= (signcalcff(cordic_depth+6) AND NOT(selectoutputff(range_depth+cordic_depth+5))) OR
                       (input_number_delay(32) AND selectoutputff(range_depth+cordic_depth+5));
          
        END IF;
        
      END IF;
      
    END PROCESS;
    
    mantissaout <= mantissaoutff; 
    exponentout <= exponentoutff;
    signout <= signoutff;    
    
  END rtl;
  
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   SINGLE PRECISION SQUARE ROOT - TOP LEVEL  ***
--***                                             ***
--***   FP_SQR.VHD                                ***
--***                                             ***
--***   Function: IEEE754 FP Square Root          ***
--***                                             ***
--***   31/01/08 ML                               ***
--***                                             ***
--***   (c) 2008 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** Latency = 28                                ***
--*** Based on FPROOT1.VHD (12/06)                ***
--***************************************************

ENTITY fp_sqr IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (23 DOWNTO 1);

		  signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (8 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (23 DOWNTO 1);
      --------------------------------------------------
      nanout : OUT STD_LOGIC;
      invalidout : OUT STD_LOGIC
		);
END fp_sqr;

ARCHITECTURE rtl OF fp_sqr IS
  
  constant manwidth : positive := 23;
  constant expwidth : positive := 8;
  
  type expfftype IS ARRAY (manwidth+4 DOWNTO 1) OF STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  
  signal signinff : STD_LOGIC;
  signal maninff : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal expinff : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal signff : STD_LOGIC_VECTOR (manwidth+4 DOWNTO 1);
  signal expnode, expdiv : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal expff : expfftype;
  signal radicand : STD_LOGIC_VECTOR (manwidth+3 DOWNTO 1);
  signal squareroot : STD_LOGIC_VECTOR (manwidth+2 DOWNTO 1);
  signal roundff, manff : STD_LOGIC_VECTOR (manwidth DOWNTO 1); 
  signal roundbit : STD_LOGIC;
  signal preadjust : STD_LOGIC;
  signal zerovec : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal offset : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
    
  -- conditions
  signal nanmanff, nanexpff : STD_LOGIC_VECTOR (manwidth+4 DOWNTO 1);
  signal zeroexpff, zeromanff : STD_LOGIC_VECTOR (manwidth+3 DOWNTO 1); 
  signal expinzero, expinmax : STD_LOGIC_VECTOR (expwidth DOWNTO 1);
  signal maninzero : STD_LOGIC_VECTOR (manwidth DOWNTO 1);
  signal expzero, expmax, manzero : STD_LOGIC;
  signal infinitycondition, nancondition : STD_LOGIC;

  component fp_sqrroot IS 
  GENERIC (width : positive := 52);
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        rad : IN STD_LOGIC_VECTOR (width+1 DOWNTO 1);

		  root : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
		  );
	end component;
		
BEGIN
    
  gzva: FOR k IN 1 TO manwidth GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  gxoa: FOR k IN 1 TO expwidth-1 GENERATE
    offset(k) <= '1';
  END GENERATE;
  offset(expwidth) <= '0';

  pma: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
      
      signinff <= '0';
      FOR k IN 1 TO manwidth LOOP
        maninff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        expinff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO manwidth+4 LOOP
        signff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO manwidth+4 LOOP
        FOR j IN 1 TO expwidth LOOP
          expff(k)(j) <= '0';
        END LOOP;
      END LOOP;
      FOR k IN 1 TO manwidth LOOP
        roundff(k) <= '0';
        manff(k) <= '0';
      END LOOP;
  
    ELSIF (rising_edge(sysclk)) THEN

      signinff <= signin;
      maninff <= mantissain;
      expinff <= exponentin;
    
      signff(1) <= signinff;
      FOR k IN 2 TO manwidth+4 LOOP
        signff(k) <= signff(k-1);
      END LOOP;
      
      expff(1)(expwidth DOWNTO 1) <= expdiv;
      expff(2)(expwidth DOWNTO 1) <= expff(1)(expwidth DOWNTO 1) + offset;
      FOR k IN 3 TO manwidth+3 LOOP
        expff(k)(expwidth DOWNTO 1) <= expff(k-1)(expwidth DOWNTO 1);
      END LOOP;
      FOR k IN 1 TO expwidth LOOP
        expff(manwidth+4)(k) <= (expff(manwidth+3)(k) AND zeroexpff(manwidth+3)) OR nanexpff(manwidth+3);
      END LOOP;
    
      roundff <= squareroot(manwidth+1 DOWNTO 2) + (zerovec(manwidth-1 DOWNTO 1) & roundbit);
    
      FOR k IN 1 TO manwidth LOOP
        manff(k) <= (roundff(k) AND zeromanff(manwidth+3)) OR nanmanff(manwidth+3);
      END LOOP;
  
    END IF;
  
  END PROCESS;

--*******************
--*** CONDITIONS ***
--*******************

  pcc: PROCESS (sysclk,reset)
  BEGIN

    IF (reset = '1') THEN
      
      FOR k IN 1 TO manwidth+4 LOOP
        nanmanff(k) <= '0';
        nanexpff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO manwidth+3 LOOP
        zeroexpff(k) <= '0';
        zeromanff(k) <= '0';
      END LOOP;
    
    ELSIF (rising_edge(sysclk)) THEN
      
      nanmanff(1) <= nancondition; -- level 1
      nanexpff(1) <= nancondition OR infinitycondition; -- also max exp when infinity
      FOR k IN 2 TO manwidth+4 LOOP
        nanmanff(k) <= nanmanff(k-1);
        nanexpff(k) <= nanexpff(k-1);
      END LOOP;

      zeromanff(1) <= expzero AND NOT(infinitycondition); -- level 1
      zeroexpff(1) <= expzero; -- level 1
      FOR k IN 2 TO manwidth+3 LOOP
        zeromanff(k) <= zeromanff(k-1);
        zeroexpff(k) <= zeroexpff(k-1);
      END LOOP;
    
    END IF;
  
  END PROCESS;

--*******************
--*** SQUARE ROOT ***
--*******************

  -- if exponent is odd, double mantissa and adjust exponent
  -- core latency manwidth+2 = 25
  -- top latency = core + 1 (input) + 2 (output) = 28
  sqr: fp_sqrroot
  GENERIC MAP (width=>manwidth+2)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            rad=>radicand,
            root=>squareroot);

  radicand(1) <= '0';
  radicand(2) <= maninff(1) AND NOT(preadjust);
  gra: FOR k IN 3 TO manwidth+1 GENERATE
    radicand(k) <= (maninff(k-1) AND NOT(preadjust)) OR (maninff(k-2) AND preadjust);
  END GENERATE; 
  radicand(manwidth+2) <= NOT(preadjust) OR (maninff(manwidth) AND preadjust);
  radicand(manwidth+3) <= preadjust;   

--****************
--*** EXPONENT ***
--****************

  -- subtract 1023, divide result/2, if odd - preadjust
  -- if zero input, zero exponent and mantissa
  expnode <= expinff - offset;

  preadjust <= expnode(1);

  expdiv <= expnode(expwidth) & expnode(expwidth DOWNTO 2);

--*************
--*** ROUND ***
--*************

  -- only need to round up, round to nearest not possible out of root
  roundbit <= squareroot(1);

--*********************
--*** SPECIAL CASES ***
--*********************
-- 1. if negative input, invalid operation, NAN  (unless -0)
-- 2. -0 in -0 out
-- 3. infinity in, invalid operation, infinity out
-- 4. NAN in, invalid operation, NAN

  -- '0' if 0 
  expinzero(1) <= expinff(1);
  gxza: FOR k IN 2 TO expwidth GENERATE
    expinzero(k) <= expinzero(k-1) OR expinff(k);
  END GENERATE;
  expzero <= expinzero(expwidth); -- '0' when zero
                 
  -- '1' if nan or infinity
  expinmax(1) <= expinff(1);
  gxia: FOR k IN 2 TO expwidth GENERATE
    expinmax(k) <= expinmax(k-1) AND expinff(k);
  END GENERATE;
  expmax <= expinmax(expwidth); -- '1' when true
          
  -- '1' if not zero or infinity
  maninzero(1) <= maninff(1);
  gmza: FOR k IN 2 TO manwidth GENERATE
    maninzero(k) <= maninzero(k-1) OR maninff(k);
  END GENERATE;
  manzero <= maninzero(manwidth); 
    
  infinitycondition <= NOT(manzero) AND expmax; 

  nancondition <= (signinff AND expzero) OR (expmax AND manzero);
                
--***************
--*** OUTPUTS ***
--***************

  signout <= signff(manwidth+4);
  exponentout <= expff(manwidth+4)(expwidth DOWNTO 1);   
  mantissaout <= manff;
  -----------------------------------------------
  nanout <= nanmanff(manwidth+4);
  invalidout <= nanmanff(manwidth+4);

END rtl;



LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--********************************************************************
--***                                                              ***
--***  FP_SQRROOT.VHD                                              ***
--***                                                              ***
--***  Fixed Point Square Root Core - Restoring                    ***
--***                                                              ***
--***  21/12/06  ML                                                ***
--***                                                              ***
--***  Copyright Altera 2006                                       ***
--***                                                              ***
--***                                                              ***
--********************************************************************

ENTITY fp_sqrroot IS 
GENERIC (width : positive := 52);
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      rad : IN STD_LOGIC_VECTOR (width+1 DOWNTO 1);

		root : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
		);
END fp_sqrroot;

ARCHITECTURE rtl OF fp_sqrroot IS
  
  type nodetype IS ARRAY (width DOWNTO 1) OF STD_LOGIC_VECTOR (width+2 DOWNTO 1);
  type qfftype IS ARRAY (width-1 DOWNTO 1) OF STD_LOGIC_VECTOR (width-1 DOWNTO 1);
  
  signal zerovec : STD_LOGIC_VECTOR (width DOWNTO 1);
  signal onevec : STD_LOGIC_VECTOR (width+1 DOWNTO 1);
  signal subnode, slevel, qlevel, radff : nodetype;
  signal qff : qfftype;
    
BEGIN

gza: FOR k IN 1 TO width GENERATE
  zerovec(k) <= '0';
END GENERATE;
  
onevec <= "01" & zerovec(width-1 DOWNTO 1);

-- 1 <= input range < 4, therefore 1 <= root < 2
-- input may be shifted left by 1, therefore first subtract "001" not "01" 
slevel(1)(width+2 DOWNTO 1) <= '0' & rad;
qlevel(1)(width+2 DOWNTO 1) <= "001" & zerovec(width-1  DOWNTO 1);
subnode(1)(width+2 DOWNTO width) <= slevel(1)(width+2 DOWNTO width) - qlevel(1)(width+2 DOWNTO width);
subnode(1)(width-1 DOWNTO 1) <= slevel(1)(width-1  DOWNTO 1);

slevel(2)(width+2 DOWNTO 1) <= radff(1)(width+1 DOWNTO 1) & '0';
qlevel(2)(width+2 DOWNTO 1) <= "0101" & zerovec(width-2 DOWNTO 1); 
subnode(2)(width+2 DOWNTO width-1) <= slevel(2)(width+2 DOWNTO width-1) - qlevel(2)(width+2 DOWNTO width-1);
subnode(2)(width-2 DOWNTO 1) <= slevel(2)(width-2 DOWNTO 1);

gla: FOR k IN 3 TO width GENERATE
  glb: FOR j IN 1 TO k-2 GENERATE
    qlevel(k)(width+1-j) <= qff(width-j)(k-1-j);
  END GENERATE;
END GENERATE;

gsa: FOR k IN 3 TO width-1 GENERATE
  slevel(k)(width+2 DOWNTO 1) <= radff(k-1)(width+1 DOWNTO 1) & '0';
  qlevel(k)(width+2 DOWNTO width+1) <= "01";
  qlevel(k)(width+2-k DOWNTO 1) <= "01" & zerovec(width-k DOWNTO 1);
  subnode(k)(width+2 DOWNTO width+1-k) <= slevel(k)(width+2 DOWNTO width+1-k) - 
                                          qlevel(k)(width+2 DOWNTO width+1-k);
  subnode(k)(width-k DOWNTO 1) <= slevel(k)(width-k DOWNTO 1);
END GENERATE;

slevel(width)(width+2 DOWNTO 1) <= radff(width-1)(width+1 DOWNTO 1) & '0';
qlevel(width)(width+2 DOWNTO width+1) <= "01";
qlevel(width)(2 DOWNTO 1) <= "01";
subnode(width)(width+2 DOWNTO 1) <= slevel(width)(width+2 DOWNTO 1) - qlevel(width)(width+2 DOWNTO 1);
  
pma: PROCESS (sysclk,reset)
BEGIN

  IF (reset = '1') THEN
      
    FOR k IN 1 TO width LOOP
      FOR j IN 1 TO width+2 LOOP
        radff(k)(j) <= '0';
      END LOOP;
    END LOOP;
    FOR k IN 1 TO width-1 LOOP
      FOR j IN 1 TO width-1 LOOP
        qff(k)(j) <= '0';
      END LOOP;
    END LOOP;
      
  ELSIF (rising_edge(sysclk)) THEN
     
    IF (enable = '1') THEN
        
      radff(1)(width+2 DOWNTO 1) <= subnode(1)(width+2 DOWNTO 1); 
      FOR k IN 2 TO width LOOP
        FOR j IN 1 TO width+2 LOOP
          radff(k)(j) <= (slevel(k)(j) AND subnode(k)(width+2)) OR 
                         (subnode(k)(j) AND NOT(subnode(k)(width+2))); 
        END LOOP;
      END LOOP;
    
      FOR k IN 1 TO width-1 LOOP
        qff(width-k)(1) <= NOT(subnode(k+1)(width+2));
        FOR j IN 2 TO width-1 LOOP
          qff(k)(j) <= qff(k)(j-1);
        END LOOP;
      END LOOP;
    
    END IF;
 
  END IF;

END PROCESS;

fro: FOR k IN 1 TO width-1 GENERATE
  root(k) <= qff(k)(k);
END GENERATE;
root(width) <= '1';

END rtl;

-- megafunction wizard: %ALTMULT_ADD%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTMULT_ADD 

-- ============================================================
-- File Name: sum36x18.vhd
-- Megafunction Name(s):
-- 			ALTMULT_ADD
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 8.1 Build 163 10/28/2008 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2008 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

ENTITY fp_sum36x18 IS
	PORT
	(
		aclr3		: IN STD_LOGIC  := '0';
		clock0		: IN STD_LOGIC  := '1';
		dataa_0		: IN STD_LOGIC_VECTOR (17 DOWNTO 0) :=  (OTHERS => '0');
		dataa_1		: IN STD_LOGIC_VECTOR (17 DOWNTO 0) :=  (OTHERS => '0');
		datab_0		: IN STD_LOGIC_VECTOR (35 DOWNTO 0) :=  (OTHERS => '0');
		datab_1		: IN STD_LOGIC_VECTOR (35 DOWNTO 0) :=  (OTHERS => '0');
		ena0		: IN STD_LOGIC  := '1';
		result		: OUT STD_LOGIC_VECTOR (54 DOWNTO 0)
	);
END fp_sum36x18;


ARCHITECTURE SYN OF fp_sum36x18 IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (54 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (17 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (35 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (17 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (35 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (71 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (35 DOWNTO 0);



	COMPONENT altmult_add
	GENERIC (
		accumulator		: STRING;
		addnsub_multiplier_aclr1		: STRING;
		addnsub_multiplier_pipeline_aclr1		: STRING;
		addnsub_multiplier_pipeline_register1		: STRING;
		addnsub_multiplier_register1		: STRING;
		chainout_adder		: STRING;
		chainout_register		: STRING;
		dedicated_multiplier_circuitry		: STRING;
		input_aclr_a0		: STRING;
		input_aclr_a1		: STRING;
		input_aclr_b0		: STRING;
		input_aclr_b1		: STRING;
		input_register_a0		: STRING;
		input_register_a1		: STRING;
		input_register_b0		: STRING;
		input_register_b1		: STRING;
		input_source_a0		: STRING;
		input_source_a1		: STRING;
		input_source_b0		: STRING;
		input_source_b1		: STRING;
		intended_device_family		: STRING;
		lpm_type		: STRING;
		multiplier1_direction		: STRING;
		multiplier_aclr0		: STRING;
		multiplier_aclr1		: STRING;
		multiplier_register0		: STRING;
		multiplier_register1		: STRING;
		number_of_multipliers		: NATURAL;
		output_aclr		: STRING;
		output_register		: STRING;
		port_addnsub1		: STRING;
		port_signa		: STRING;
		port_signb		: STRING;
		representation_a		: STRING;
		representation_b		: STRING;
		signed_aclr_a		: STRING;
		signed_aclr_b		: STRING;
		signed_pipeline_aclr_a		: STRING;
		signed_pipeline_aclr_b		: STRING;
		signed_pipeline_register_a		: STRING;
		signed_pipeline_register_b		: STRING;
		signed_register_a		: STRING;
		signed_register_b		: STRING;
		width_a		: NATURAL;
		width_b		: NATURAL;
		width_chainin		: NATURAL;
		width_result		: NATURAL;
		zero_chainout_output_aclr		: STRING;
		zero_chainout_output_register		: STRING;
		zero_loopback_aclr		: STRING;
		zero_loopback_output_aclr		: STRING;
		zero_loopback_output_register		: STRING;
		zero_loopback_pipeline_aclr		: STRING;
		zero_loopback_pipeline_register		: STRING;
		zero_loopback_register		: STRING
	);
	PORT (
			dataa	: IN STD_LOGIC_VECTOR (35 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (71 DOWNTO 0);
			clock0	: IN STD_LOGIC ;
			aclr3	: IN STD_LOGIC ;
			ena0	: IN STD_LOGIC ;
			result	: OUT STD_LOGIC_VECTOR (54 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	sub_wire6    <= datab_1(35 DOWNTO 0);
	sub_wire3    <= dataa_1(17 DOWNTO 0);
	result    <= sub_wire0(54 DOWNTO 0);
	sub_wire1    <= dataa_0(17 DOWNTO 0);
	sub_wire2    <= sub_wire3(17 DOWNTO 0) & sub_wire1(17 DOWNTO 0);
	sub_wire4    <= datab_0(35 DOWNTO 0);
	sub_wire5    <= sub_wire6(35 DOWNTO 0) & sub_wire4(35 DOWNTO 0);

	ALTMULT_ADD_component : ALTMULT_ADD
	GENERIC MAP (
		accumulator => "NO",
		addnsub_multiplier_aclr1 => "ACLR3",
		addnsub_multiplier_pipeline_aclr1 => "ACLR3",
		addnsub_multiplier_pipeline_register1 => "CLOCK0",
		addnsub_multiplier_register1 => "CLOCK0",
		chainout_adder => "NO",
		chainout_register => "UNREGISTERED",
		dedicated_multiplier_circuitry => "AUTO",
		input_aclr_a0 => "ACLR3",
		input_aclr_a1 => "ACLR3",
		input_aclr_b0 => "ACLR3",
		input_aclr_b1 => "ACLR3",
		input_register_a0 => "CLOCK0",
		input_register_a1 => "CLOCK0",
		input_register_b0 => "CLOCK0",
		input_register_b1 => "CLOCK0",
		input_source_a0 => "DATAA",
		input_source_a1 => "DATAA",
		input_source_b0 => "DATAB",
		input_source_b1 => "DATAB",
		intended_device_family => "Stratix III",
		lpm_type => "altmult_add",
		multiplier1_direction => "ADD",
		multiplier_aclr0 => "ACLR3",
		multiplier_aclr1 => "ACLR3",
		multiplier_register0 => "CLOCK0",
		multiplier_register1 => "CLOCK0",
		number_of_multipliers => 2,
		output_aclr => "ACLR3",
		output_register => "CLOCK0",
		port_addnsub1 => "PORT_UNUSED",
		port_signa => "PORT_UNUSED",
		port_signb => "PORT_UNUSED",
		representation_a => "UNSIGNED",
		representation_b => "UNSIGNED",
		signed_aclr_a => "ACLR3",
		signed_aclr_b => "ACLR3",
		signed_pipeline_aclr_a => "ACLR3",
		signed_pipeline_aclr_b => "ACLR3",
		signed_pipeline_register_a => "CLOCK0",
		signed_pipeline_register_b => "CLOCK0",
		signed_register_a => "CLOCK0",
		signed_register_b => "CLOCK0",
		width_a => 18,
		width_b => 36,
		width_chainin => 1,
		width_result => 55,
		zero_chainout_output_aclr => "ACLR3",
		zero_chainout_output_register => "CLOCK0",
		zero_loopback_aclr => "ACLR3",
		zero_loopback_output_aclr => "ACLR3",
		zero_loopback_output_register => "CLOCK0",
		zero_loopback_pipeline_aclr => "ACLR3",
		zero_loopback_pipeline_register => "CLOCK0",
		zero_loopback_register => "CLOCK0"
	)
	PORT MAP (
		dataa => sub_wire2,
		datab => sub_wire5,
		clock0 => clock0,
		aclr3 => aclr3,
		ena0 => ena0,
		result => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ACCUM_DIRECTION STRING "Add"
-- Retrieval info: PRIVATE: ACCUM_SLOAD_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ACCUM_SLOAD_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ACCUM_SLOAD_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ACCUM_SLOAD_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ACCUM_SLOAD_PIPE_REG STRING "1"
-- Retrieval info: PRIVATE: ACCUM_SLOAD_REG STRING "1"
-- Retrieval info: PRIVATE: ADDNSUB1_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADDNSUB1_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB1_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADDNSUB1_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB1_PIPE_REG STRING "1"
-- Retrieval info: PRIVATE: ADDNSUB1_REG STRING "1"
-- Retrieval info: PRIVATE: ADDNSUB3_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADDNSUB3_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB3_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADDNSUB3_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB3_PIPE_REG STRING "1"
-- Retrieval info: PRIVATE: ADDNSUB3_REG STRING "1"
-- Retrieval info: PRIVATE: ADD_ENABLE NUMERIC "1"
-- Retrieval info: PRIVATE: ALL_REG_ACLR NUMERIC "1"
-- Retrieval info: PRIVATE: A_ACLR_SRC_MULT0 NUMERIC "3"
-- Retrieval info: PRIVATE: A_CLK_SRC_MULT0 NUMERIC "0"
-- Retrieval info: PRIVATE: B_ACLR_SRC_MULT0 NUMERIC "3"
-- Retrieval info: PRIVATE: B_CLK_SRC_MULT0 NUMERIC "0"
-- Retrieval info: PRIVATE: CHAINOUT_OUTPUT_ACLR NUMERIC "3"
-- Retrieval info: PRIVATE: CHAINOUT_OUTPUT_REG STRING "0"
-- Retrieval info: PRIVATE: CHAINOUT_OUTPUT_REGISTER NUMERIC "0"
-- Retrieval info: PRIVATE: CHAINOUT_OUTPUT_REGISTERED NUMERIC "0"
-- Retrieval info: PRIVATE: CHAS_ZERO_CHAINOUT NUMERIC "1"
-- Retrieval info: PRIVATE: HAS_ACCUMULATOR NUMERIC "0"
-- Retrieval info: PRIVATE: HAS_ACUMM_SLOAD NUMERIC "0"
-- Retrieval info: PRIVATE: HAS_CHAININ_PORT NUMERIC "0"
-- Retrieval info: PRIVATE: HAS_CHAINOUT_ADDER NUMERIC "0"
-- Retrieval info: PRIVATE: HAS_LOOPBACK NUMERIC "0"
-- Retrieval info: PRIVATE: HAS_MAC STRING "0"
-- Retrieval info: PRIVATE: HAS_SAT_ROUND STRING "0"
-- Retrieval info: PRIVATE: HAS_ZERO_LOOPBACK NUMERIC "0"
-- Retrieval info: PRIVATE: IMPL_STYLE_DEDICATED NUMERIC "0"
-- Retrieval info: PRIVATE: IMPL_STYLE_DEFAULT NUMERIC "1"
-- Retrieval info: PRIVATE: IMPL_STYLE_LCELL NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix III"
-- Retrieval info: PRIVATE: MULT_REGA0 NUMERIC "1"
-- Retrieval info: PRIVATE: MULT_REGB0 NUMERIC "1"
-- Retrieval info: PRIVATE: MULT_REGOUT0 NUMERIC "1"
-- Retrieval info: PRIVATE: NUM_MULT STRING "2"
-- Retrieval info: PRIVATE: OP1 STRING "Add"
-- Retrieval info: PRIVATE: OP3 STRING "Add"
-- Retrieval info: PRIVATE: OUTPUT_EXTRA_LAT NUMERIC "0"
-- Retrieval info: PRIVATE: OUTPUT_REG_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: OUTPUT_REG_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: Q_ACLR_SRC_MULT0 NUMERIC "3"
-- Retrieval info: PRIVATE: Q_CLK_SRC_MULT0 NUMERIC "0"
-- Retrieval info: PRIVATE: REG_OUT NUMERIC "1"
-- Retrieval info: PRIVATE: RNFORMAT STRING "55"
-- Retrieval info: PRIVATE: ROTATE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ROTATE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ROTATE_OUT_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ROTATE_OUT_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ROTATE_OUT_REG STRING "1"
-- Retrieval info: PRIVATE: ROTATE_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ROTATE_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ROTATE_PIPE_REG STRING "1"
-- Retrieval info: PRIVATE: ROTATE_REG STRING "1"
-- Retrieval info: PRIVATE: RQFORMAT STRING "Q1.15"
-- Retrieval info: PRIVATE: RTS_WIDTH STRING "55"
-- Retrieval info: PRIVATE: SAME_CONFIG NUMERIC "1"
-- Retrieval info: PRIVATE: SAME_CONTROL_SRC_A0 NUMERIC "1"
-- Retrieval info: PRIVATE: SAME_CONTROL_SRC_B0 NUMERIC "1"
-- Retrieval info: PRIVATE: SCANOUTA NUMERIC "0"
-- Retrieval info: PRIVATE: SCANOUTB NUMERIC "0"
-- Retrieval info: PRIVATE: SHIFTOUTA_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: SHIFTOUTA_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SHIFTOUTA_REG STRING "0"
-- Retrieval info: PRIVATE: SHIFT_RIGHT_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: SHIFT_RIGHT_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SHIFT_RIGHT_OUT_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: SHIFT_RIGHT_OUT_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SHIFT_RIGHT_OUT_REG STRING "1"
-- Retrieval info: PRIVATE: SHIFT_RIGHT_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: SHIFT_RIGHT_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SHIFT_RIGHT_PIPE_REG STRING "1"
-- Retrieval info: PRIVATE: SHIFT_RIGHT_REG STRING "1"
-- Retrieval info: PRIVATE: SHIFT_ROTATE_MODE STRING "None"
-- Retrieval info: PRIVATE: SIGNA STRING "Unsigned"
-- Retrieval info: PRIVATE: SIGNA_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: SIGNA_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SIGNA_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: SIGNA_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SIGNA_PIPE_REG STRING "1"
-- Retrieval info: PRIVATE: SIGNA_REG STRING "1"
-- Retrieval info: PRIVATE: SIGNB STRING "Unsigned"
-- Retrieval info: PRIVATE: SIGNB_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: SIGNB_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SIGNB_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: SIGNB_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SIGNB_PIPE_REG STRING "1"
-- Retrieval info: PRIVATE: SIGNB_REG STRING "1"
-- Retrieval info: PRIVATE: SRCA0 STRING "Multiplier input"
-- Retrieval info: PRIVATE: SRCB0 STRING "Multiplier input"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: WIDTHA STRING "18"
-- Retrieval info: PRIVATE: WIDTHB STRING "36"
-- Retrieval info: PRIVATE: ZERO_CHAINOUT_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ZERO_CHAINOUT_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ZERO_CHAINOUT_REG STRING "1"
-- Retrieval info: PRIVATE: ZERO_LOOPBACK_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ZERO_LOOPBACK_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ZERO_LOOPBACK_OUT_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ZERO_LOOPBACK_OUT_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ZERO_LOOPBACK_OUT_REG STRING "1"
-- Retrieval info: PRIVATE: ZERO_LOOPBACK_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ZERO_LOOPBACK_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ZERO_LOOPBACK_PIPE_REG STRING "1"
-- Retrieval info: PRIVATE: ZERO_LOOPBACK_REG STRING "1"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: ACCUMULATOR STRING "NO"
-- Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_ACLR1 STRING "ACLR3"
-- Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_PIPELINE_ACLR1 STRING "ACLR3"
-- Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_PIPELINE_REGISTER1 STRING "CLOCK0"
-- Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_REGISTER1 STRING "CLOCK0"
-- Retrieval info: CONSTANT: CHAINOUT_ADDER STRING "NO"
-- Retrieval info: CONSTANT: CHAINOUT_REGISTER STRING "UNREGISTERED"
-- Retrieval info: CONSTANT: DEDICATED_MULTIPLIER_CIRCUITRY STRING "AUTO"
-- Retrieval info: CONSTANT: INPUT_ACLR_A0 STRING "ACLR3"
-- Retrieval info: CONSTANT: INPUT_ACLR_A1 STRING "ACLR3"
-- Retrieval info: CONSTANT: INPUT_ACLR_B0 STRING "ACLR3"
-- Retrieval info: CONSTANT: INPUT_ACLR_B1 STRING "ACLR3"
-- Retrieval info: CONSTANT: INPUT_REGISTER_A0 STRING "CLOCK0"
-- Retrieval info: CONSTANT: INPUT_REGISTER_A1 STRING "CLOCK0"
-- Retrieval info: CONSTANT: INPUT_REGISTER_B0 STRING "CLOCK0"
-- Retrieval info: CONSTANT: INPUT_REGISTER_B1 STRING "CLOCK0"
-- Retrieval info: CONSTANT: INPUT_SOURCE_A0 STRING "DATAA"
-- Retrieval info: CONSTANT: INPUT_SOURCE_A1 STRING "DATAA"
-- Retrieval info: CONSTANT: INPUT_SOURCE_B0 STRING "DATAB"
-- Retrieval info: CONSTANT: INPUT_SOURCE_B1 STRING "DATAB"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix III"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altmult_add"
-- Retrieval info: CONSTANT: MULTIPLIER1_DIRECTION STRING "ADD"
-- Retrieval info: CONSTANT: MULTIPLIER_ACLR0 STRING "ACLR3"
-- Retrieval info: CONSTANT: MULTIPLIER_ACLR1 STRING "ACLR3"
-- Retrieval info: CONSTANT: MULTIPLIER_REGISTER0 STRING "CLOCK0"
-- Retrieval info: CONSTANT: MULTIPLIER_REGISTER1 STRING "CLOCK0"
-- Retrieval info: CONSTANT: NUMBER_OF_MULTIPLIERS NUMERIC "2"
-- Retrieval info: CONSTANT: OUTPUT_ACLR STRING "ACLR3"
-- Retrieval info: CONSTANT: OUTPUT_REGISTER STRING "CLOCK0"
-- Retrieval info: CONSTANT: PORT_ADDNSUB1 STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SIGNA STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SIGNB STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: REPRESENTATION_A STRING "UNSIGNED"
-- Retrieval info: CONSTANT: REPRESENTATION_B STRING "UNSIGNED"
-- Retrieval info: CONSTANT: SIGNED_ACLR_A STRING "ACLR3"
-- Retrieval info: CONSTANT: SIGNED_ACLR_B STRING "ACLR3"
-- Retrieval info: CONSTANT: SIGNED_PIPELINE_ACLR_A STRING "ACLR3"
-- Retrieval info: CONSTANT: SIGNED_PIPELINE_ACLR_B STRING "ACLR3"
-- Retrieval info: CONSTANT: SIGNED_PIPELINE_REGISTER_A STRING "CLOCK0"
-- Retrieval info: CONSTANT: SIGNED_PIPELINE_REGISTER_B STRING "CLOCK0"
-- Retrieval info: CONSTANT: SIGNED_REGISTER_A STRING "CLOCK0"
-- Retrieval info: CONSTANT: SIGNED_REGISTER_B STRING "CLOCK0"
-- Retrieval info: CONSTANT: WIDTH_A NUMERIC "18"
-- Retrieval info: CONSTANT: WIDTH_B NUMERIC "36"
-- Retrieval info: CONSTANT: WIDTH_CHAININ NUMERIC "1"
-- Retrieval info: CONSTANT: WIDTH_RESULT NUMERIC "55"
-- Retrieval info: CONSTANT: ZERO_CHAINOUT_OUTPUT_ACLR STRING "ACLR3"
-- Retrieval info: CONSTANT: ZERO_CHAINOUT_OUTPUT_REGISTER STRING "CLOCK0"
-- Retrieval info: CONSTANT: ZERO_LOOPBACK_ACLR STRING "ACLR3"
-- Retrieval info: CONSTANT: ZERO_LOOPBACK_OUTPUT_ACLR STRING "ACLR3"
-- Retrieval info: CONSTANT: ZERO_LOOPBACK_OUTPUT_REGISTER STRING "CLOCK0"
-- Retrieval info: CONSTANT: ZERO_LOOPBACK_PIPELINE_ACLR STRING "ACLR3"
-- Retrieval info: CONSTANT: ZERO_LOOPBACK_PIPELINE_REGISTER STRING "CLOCK0"
-- Retrieval info: CONSTANT: ZERO_LOOPBACK_REGISTER STRING "CLOCK0"
-- Retrieval info: USED_PORT: aclr3 0 0 0 0 INPUT GND "aclr3"
-- Retrieval info: USED_PORT: clock0 0 0 0 0 INPUT VCC "clock0"
-- Retrieval info: USED_PORT: dataa_0 0 0 18 0 INPUT GND "dataa_0[17..0]"
-- Retrieval info: USED_PORT: dataa_1 0 0 18 0 INPUT GND "dataa_1[17..0]"
-- Retrieval info: USED_PORT: datab_0 0 0 36 0 INPUT GND "datab_0[35..0]"
-- Retrieval info: USED_PORT: datab_1 0 0 36 0 INPUT GND "datab_1[35..0]"
-- Retrieval info: USED_PORT: ena0 0 0 0 0 INPUT VCC "ena0"
-- Retrieval info: USED_PORT: result 0 0 55 0 OUTPUT GND "result[54..0]"
-- Retrieval info: CONNECT: @datab 0 0 36 36 datab_1 0 0 36 0
-- Retrieval info: CONNECT: @aclr3 0 0 0 0 aclr3 0 0 0 0
-- Retrieval info: CONNECT: @clock0 0 0 0 0 clock0 0 0 0 0
-- Retrieval info: CONNECT: result 0 0 55 0 @result 0 0 55 0
-- Retrieval info: CONNECT: @dataa 0 0 18 0 dataa_0 0 0 18 0
-- Retrieval info: CONNECT: @dataa 0 0 18 18 dataa_1 0 0 18 0
-- Retrieval info: CONNECT: @ena0 0 0 0 0 ena0 0 0 0 0
-- Retrieval info: CONNECT: @datab 0 0 36 0 datab_0 0 0 36 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL sum36x18.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL sum36x18.inc FALSE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL sum36x18.cmp TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL sum36x18.bsf FALSE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL sum36x18_inst.vhd FALSE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL sum36x18_waveforms.html TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL sum36x18_wave*.jpg FALSE FALSE
-- Retrieval info: LIB_FILE: altera_mf

LIBRARY ieee;
LIBRARY work;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_TAN1.VHD                               ***
--***                                             ***
--***   Function: Single Precision Floating Point ***
--***   Tangent                                   ***
--***                                             ***
--***   23/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** NOTES                                       ***
--***************************************************

--*** 1. for very top of range (last 256 mantissa lsbs before pi/2), use seperate ROM, not  
--*** calculation
--*** 2. if round up starting when X.49999, errors reduce about 25%, need to tweak this, still getting
--*** all -1 errors with bX.111111111. less errors with less tail bits for smaller exponents (like 122)
--*** more for exponent = 126

ENTITY fp_tan IS
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      mantissain : IN STD_LOGIC_VECTOR (23 DOWNTO 1); 
      exponentin : IN STD_LOGIC_VECTOR (8 DOWNTO 1);

      signout : OUT STD_LOGIC;
      mantissaout : OUT STD_LOGIC_VECTOR (23 DOWNTO 1); 
      exponentout : OUT STD_LOGIC_VECTOR (8 DOWNTO 1)  
     );
END fp_tan;

ARCHITECTURE rtl of fp_tan IS

  -- input section
  signal zerovec : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal mantissainff : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal exponentinff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal argumentff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal topargumentff : STD_LOGIC_VECTOR (9 DOWNTO 1);
  signal middleargumentff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal tanhighmantissaff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal tanmiddleff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal tanhighexponentff : STD_LOGIC_VECTOR (5 DOWNTO 1);
  signal tanlowsumff : STD_LOGIC_VECTOR (37 DOWNTO 1);
  signal shiftin : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal shiftinbus : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal argumentbus : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal tanhighmantissa : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal tanhighexponent : STD_LOGIC_VECTOR (5 DOWNTO 1);
  signal tanmiddle : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal deltwo_tailnode : STD_LOGIC_VECTOR (19 DOWNTO 1);
  signal tantailnode : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal tanlowsumnode : STD_LOGIC_VECTOR (37 DOWNTO 1);
  signal tanlowmantissabus : STD_LOGIC_VECTOR (56 DOWNTO 1);
  
  -- numerator section
  signal tanlowff : STD_LOGIC_VECTOR (56 DOWNTO 1);
  signal numeratorsumff : STD_LOGIC_VECTOR (57 DOWNTO 1);
  signal tanlowshift : STD_LOGIC_VECTOR (5 DOWNTO 1);
  signal numeratormantissaff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal numeratorexponentff : STD_LOGIC_VECTOR (5 DOWNTO 1);
  signal delone_tanhighexponent : STD_LOGIC_VECTOR (5 DOWNTO 1);
  signal delthr_tanhighexponent : STD_LOGIC_VECTOR (5 DOWNTO 1);
  signal deltwo_tanhighmantissa : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal tanlowbus : STD_LOGIC_VECTOR (56 DOWNTO 1);
  signal numeratorsum : STD_LOGIC_VECTOR (57 DOWNTO 1);
  signal numeratorlead, numeratorleadnode : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal numeratormantissa : STD_LOGIC_VECTOR (36 DOWNTO 1); 
  signal numeratorexponent : STD_LOGIC_VECTOR (5 DOWNTO 1);
  
  -- denominator section
  signal lowleadff : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal denominatorleadff : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal multshiftff : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal denominatorproductff : STD_LOGIC_VECTOR (36 DOWNTO 1); 
  signal denominatorff : STD_LOGIC_VECTOR (36 DOWNTO 1); 
  signal denominatormantissaff : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal inverseexponentff : STD_LOGIC_VECTOR (6 DOWNTO 1); 
  signal lowleadnode : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal multshiftnode : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal denominatorproductbus : STD_LOGIC_VECTOR (36 DOWNTO 1); 
  signal denominator : STD_LOGIC_VECTOR (36 DOWNTO 1); 
  signal delone_denominator : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal denominatorlead : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal denominatormantissa : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal delone_tanlowsum : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal lowmantissabus : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal delthr_tanhighmantissa : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal multipliernode : STD_LOGIC_VECTOR (72 DOWNTO 1);
  signal delfor_tanhighexponent : STD_LOGIC_VECTOR (5 DOWNTO 1);
  signal deltwo_lowlead : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal multexponent : STD_LOGIC_VECTOR (6 DOWNTO 1);         
  signal denominatorexponent : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal inverseexponent : STD_LOGIC_VECTOR (6 DOWNTO 1);

  -- divider section
  signal tanexponentff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal tanexponentnormff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal tanexponentoutff : STD_LOGIC_VECTOR (8 DOWNTO 1); 
  signal tanmantissanormff : STD_LOGIC_VECTOR (24 DOWNTO 1);
  signal roundbitff : STD_LOGIC;
  signal mantissaoutff : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal exponentoutff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal overff : STD_LOGIC;
  signal denominatorinverse : STD_LOGIC_VECTOR (36 DOWNTO 1); 
  signal del_numeratormantissa : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal multiplier_tan : STD_LOGIC_VECTOR (72 DOWNTO 1);
  signal tanmantissa : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal tanmantissanorm : STD_LOGIC_VECTOR (24 DOWNTO 1);
  signal tanmantissatail : STD_LOGIC_VECTOR (9 DOWNTO 1);
  signal overcheck : STD_LOGIC_VECTOR (24 DOWNTO 1);
  signal del_inverseexponent : STD_LOGIC_VECTOR (6 DOWNTO 1);
  signal del_numeratorexponent : STD_LOGIC_VECTOR (5 DOWNTO 1);
  signal tanexponent, tanexponentnorm : STD_LOGIC_VECTOR (8 DOWNTO 1); 
  signal exponentoutnode : STD_LOGIC_VECTOR (8 DOWNTO 1); 
  signal mantissaoutnode : STD_LOGIC_VECTOR (23 DOWNTO 1);

  -- small inputs
  signal signff : STD_LOGIC_VECTOR (30 DOWNTO 1);
  signal small_mantissa : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal small_exponent : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal exponentcheck : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal small_inputff : STD_LOGIC_VECTOR (28 DOWNTO 1);
  signal mantissabase : STD_LOGIC_VECTOR (24 DOWNTO 1);
  signal exponentbase : STD_LOGIC_VECTOR (8 DOWNTO 1);
   
  component fp_tanlut1 
  PORT (
        add : IN STD_LOGIC_VECTOR (9 DOWNTO 1);
        mantissa : OUT STD_LOGIC_VECTOR (36 DOWNTO 1);
        exponent : OUT STD_LOGIC_VECTOR (5 DOWNTO 1)
       );
   end component;
 
   component fp_tanlut2 
   PORT (
         add : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
         tanfraction : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
        );
   end component;
  
  component fp_clz36
  PORT (
        mantissa : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
      
        leading : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
     );
  end component;

  component fp_clz36x6
  PORT (
        mantissa : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
      
        leading : OUT STD_LOGIC_VECTOR (6 DOWNTO 1)    
     );
  end component;
      
  component fp_lsft36 
  PORT (
        inbus : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);

	     outbus : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
	    );
	end component;

  component fp_rsft36 
  PORT (
        inbus : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (6 DOWNTO 1);

	     outbus : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
	    );
	end component;

  component fp_rsft56x20  
  PORT (
        inbus : IN STD_LOGIC_VECTOR (56 DOWNTO 1);
        shift : IN STD_LOGIC_VECTOR (5 DOWNTO 1);

	     outbus : OUT STD_LOGIC_VECTOR (56 DOWNTO 1)
	    );	 
	end component;

  component fp_inv_core 
  GENERIC (synthesize : integer := 1); 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        divisor : IN STD_LOGIC_VECTOR (36 DOWNTO 1);

		    quotient : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
		    );
  end component;
	
	component fp_del 
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
   end component;

  component fp_fxmul
  GENERIC (
           widthaa : positive := 18;
           widthbb : positive := 18;
           widthcc : positive := 36;
           pipes : positive := 1;
           accuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
           device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
           synthesize : integer := 0
          );
   PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dataaa : IN STD_LOGIC_VECTOR (widthaa DOWNTO 1);
        databb : IN STD_LOGIC_VECTOR (widthbb DOWNTO 1); 
      
        result : OUT STD_LOGIC_VECTOR (widthcc DOWNTO 1)
       );
  end component;
   	       
BEGIN
    
  gza: FOR k IN 1 TO 36 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  -- convert to fixed point
  pin: PROCESS (sysclk,reset)
  BEGIN
    
    IF  (reset = '1') THEN
      
      FOR k IN 1 TO 23 LOOP
        mantissainff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 8 LOOP
        exponentinff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 36 LOOP
        argumentff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 9 LOOP
        topargumentff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 8 LOOP
        middleargumentff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 36 LOOP
        tanhighmantissaff(k) <= '0';
        tanmiddleff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 5 LOOP
        tanhighexponentff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 5 LOOP
        tanlowsumff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN
      
        mantissainff <= mantissain;
        exponentinff <= exponentin;
        
        argumentff <= argumentbus;
        topargumentff <= argumentff(36 DOWNTO 28);
        middleargumentff <= argumentff(27 DOWNTO 20);
  
        tanhighmantissaff <= tanhighmantissa;
        tanhighexponentff <= tanhighexponent;
        tanmiddleff <= tanmiddle;  
        
        tanlowsumff <= tanlowsumnode;  
           
      END IF;
      
    END IF;
    
  END PROCESS;
  
  shiftin <= 127 - exponentinff;
  shiftinbus <= '1' & mantissainff & zerovec(12 DOWNTO 1);
  
  csftin: fp_rsft36 
  PORT MAP (inbus=>shiftinbus,shift=>shiftin(6 DOWNTO 1),
            outbus=>argumentbus);

  chtt: fp_tanlut1
  PORT MAP (add=>topargumentff,
            mantissa=>tanhighmantissa,
            exponent=>tanhighexponent);
            
  cltt: fp_tanlut2
  PORT MAP (add=>middleargumentff,
           tanfraction=>tanmiddle);
   
  -- in level 2, out level 4        
  dtail: fp_del 
  GENERIC MAP (width=>19,pipes=>2)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable, -- use reset to force to ffs here
            aa=>argumentff(19 DOWNTO 1),
            cc=>deltwo_tailnode); 
                   
  tantailnode <= zerovec(8 DOWNTO 1) & deltwo_tailnode & zerovec(9 DOWNTO 1);
  
  tanlowsumnode <= ('0' & tanmiddleff(36 DOWNTO 1)) + ('0' & tantailnode);
  
  tanlowmantissabus <= tanlowsumff & zerovec(19 DOWNTO 1);
  
  --*********************************************
  --*** Align two tangent values for addition ***
  --*********************************************
 
  padd: PROCESS (sysclk,reset)
  BEGIN
    
    IF  (reset = '1') THEN
      
      FOR k IN 1 TO 56 LOOP
        tanlowff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 57 LOOP
        numeratorsumff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 36 LOOP
        numeratormantissaff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 5 LOOP
        numeratorexponentff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN
      
        tanlowff <= tanlowbus;
        numeratorsumff <= numeratorsum;
        numeratormantissaff <= numeratormantissa;
        numeratorexponentff <= numeratorexponent;
          
      END IF;
      
    END IF;
    
  END PROCESS;
  
  -- in level 4, out level 5        
  dhxa: fp_del 
  GENERIC MAP (width=>5,pipes=>1)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable, -- use reset to force to ffs here
            aa=>tanhighexponentff,
            cc=>delone_tanhighexponent); 

  -- in level 5, out level 7        
  dhxb: fp_del 
  GENERIC MAP (width=>5,pipes=>2)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable, -- use reset to force to ffs here
            aa=>delone_tanhighexponent,
            cc=>delthr_tanhighexponent); 
              
  -- in level 4, out level 6        
  dhm: fp_del 
  GENERIC MAP (width=>36,pipes=>2)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable, -- use reset to force to ffs here
            aa=>tanhighmantissaff,
            cc=>deltwo_tanhighmantissa); 
              
  -- tan high mantissa format 1.XXX, tan low mantissa format 0.XXXXX 
  -- tan high exponent base is 119 (top of middle range)
  tanlowshift <= delone_tanhighexponent;
  
  crsadd: fp_rsft56x20
  PORT MAP (inbus=>tanlowmantissabus,
            shift=>tanlowshift,
            outbus=>tanlowbus);
  
  numeratorsum <= ('0' & deltwo_tanhighmantissa & zerovec(20 DOWNTO 1)) + ('0' & tanlowff);
  
  -- level 8
  -- no pipe between clz and shift as only 6 bit shift 
  -- middle exponent is 119, and 2 overflow bits in numerator sum, so this will
  -- cover downto (119+2-6) = 115 exponent
  -- below 115 exponent, output mantissa = input mantissa
  clznuma: fp_clz36x6
  PORT MAP (mantissa=>numeratorsumff(57 DOWNTO 22),
            leading=>numeratorlead);
 
  numeratorleadnode <= "000" & numeratorlead(3 DOWNTO 1); -- force [6:4] to 0 to optimize away logic in LSFT
  clsnuma: fp_lsft36 
  PORT MAP (inbus=>numeratorsumff(57 DOWNTO 22),shift=>numeratorleadnode,
            outbus=>numeratormantissa);
   
  numeratorexponent <= delthr_tanhighexponent - numeratorlead(5 DOWNTO 1) + 1;
            
  --gnnadd: FOR k IN 1 TO 36 GENERATE
  --  numeratormantissa(k) <= (numeratorsumff(k+20) AND NOT(numeratorsumff(57))) OR 
  --                          (numeratorsumff(k+21) AND numeratorsumff(57));
  --END GENERATE;
  --numeratorexponent <= delthr_tanhighexponent + ("0000" & numeratorsumff(57));
  
  --***************************************************
  --*** Align two tangent values for multiplication ***
  --***************************************************  

  pmul: PROCESS (sysclk,reset)
  BEGIN
    
    IF  (reset = '1') THEN

      FOR k IN 1 TO 6 LOOP
        lowleadff(k) <= '0';
        denominatorleadff(k) <= '0';
        inverseexponentff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 6 LOOP
        multshiftff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 36 LOOP
        denominatorproductff(k) <= '0';
        denominatorff(k) <= '0';
        denominatormantissaff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN
      
        lowleadff <= lowleadnode;
        multshiftff <= multshiftnode;
        denominatorproductff <= denominatorproductbus;
        denominatorff <= denominator;
        denominatorleadff <= denominatorlead;
        denominatormantissaff <= denominatormantissa;
        inverseexponentff <= inverseexponent;
        
      END IF;
      
    END IF;
    
  END PROCESS;
  
  clzmula: fp_clz36
  PORT MAP (mantissa=>tanlowsumff(37 DOWNTO 2),
            leading=>lowleadnode);
  
  -- in level 5, out level 6       
  dlm: fp_del 
  GENERIC MAP (width=>36,pipes=>1)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable, -- use reset to force to ffs here
            aa=>tanlowsumff(37 DOWNTO 2),
            cc=>delone_tanlowsum); 
                      
  clsmula: fp_lsft36 
  PORT MAP (inbus=>delone_tanlowsum,shift=>lowleadff,
            outbus=>lowmantissabus);
            
  cma: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>36,widthcc=>72,
               pipes=>3,synthesize=>0)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,  
            dataaa=>deltwo_tanhighmantissa,
            databb=>lowmantissabus,
            result=>multipliernode);

  -- in level 5, out level 8        
  dhxc: fp_del 
  GENERIC MAP (width=>5,pipes=>3)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable, -- use reset to force to ffs here
            aa=>delone_tanhighexponent,
            cc=>delfor_tanhighexponent); 
  
  -- in level 6, out level 8        
  dlla: fp_del 
  GENERIC MAP (width=>6,pipes=>2)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable, -- use reset to force to ffs here
            aa=>lowleadff,
            cc=>deltwo_lowlead); 
                      
  -- msb of lowmantissa(37) is at exponent 0 for highmantissa
  multexponent <= ('0' & delfor_tanhighexponent);
  
  --multshiftnode <= "001000" - multexponent + 8 - 1 + lowlead;
  multshiftnode <= "001111" - multexponent + deltwo_lowlead;
  
  -- '1.0' is at exponent 8 compared to highmantissa 
  crsmul: fp_rsft36 
  PORT MAP (inbus=>multipliernode(72 DOWNTO 37),shift=>multshiftff,
            outbus=>denominatorproductbus);
                
  denominator <= ('1' & zerovec(35 DOWNTO 1)) - denominatorproductff;
  
  -- in level 11, out level 12        
  dda: fp_del 
  GENERIC MAP (width=>36,pipes=>1)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable, -- use reset to force to ffs here
            aa=>denominatorff,
            cc=>delone_denominator); 
            
  clzmulb: fp_clz36
  PORT MAP (mantissa=>denominatorff,
            leading=>denominatorlead);
            
  -- denominatormantissa level 12, (denominatormantissaff level 13)
  clsmulb: fp_lsft36 
  PORT MAP (inbus=>delone_denominator,shift=>denominatorleadff,
            outbus=>denominatormantissa); 
            
  denominatorexponent <= denominatorleadff; -- actually inverse of exponent i.e. 4 => -4, so sign does not have to change after inverting
  -- inverseexponentff level 13
  inverseexponent <= denominatorexponent - 1;
 
  --****************************   
  --*** main divider section ***
  --****************************
  
  pdiv: PROCESS (sysclk,reset)
  BEGIN
    
    IF  (reset = '1') THEN

      FOR k IN 1 TO 8 LOOP
        tanexponentff(k) <= '0';
        tanexponentnormff(k) <= '0';
        exponentoutff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 24 LOOP
        tanmantissanormff(k) <= '0';
      END LOOP;
      roundbitff <= '0';
      FOR k IN 1 TO 23 LOOP
        mantissaoutff(k) <= '0';
      END LOOP;
      overff <= '0';
      
    ELSIF (rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN
      
        tanexponentff <= tanexponent; 
        tanmantissanormff <= tanmantissanorm; -- level 29
        tanexponentnormff <= tanexponentnorm;  -- level 29
        overff <= overcheck(24);
        -- round up if 0.4999
        roundbitff <= tanmantissanorm(1) OR 
                     (tanmantissatail(9) AND
                      tanmantissatail(8) AND tanmantissatail(7) AND 
                      tanmantissatail(6) AND tanmantissatail(5) AND
                      tanmantissatail(4) AND tanmantissatail(3) AND 
                      tanmantissatail(2) AND tanmantissatail(1));
         
        mantissaoutff <= mantissaoutnode; -- level 30
        exponentoutff <= exponentoutnode; -- level 30
        
      END IF;
      
    END IF;
    
  END PROCESS;
  
  -- latency 12
  -- will give output between 0.5 and 0.99999...
  -- will always need to be normalized
  -- level 13 in, level 25 out
  cinv: fp_inv_core 
  GENERIC MAP (synthesize=>0) 
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            divisor=>denominatormantissaff,
            quotient=>denominatorinverse);
   
  -- level 8 in, level 25 out         
	dnuma: fp_del 
  GENERIC MAP (width=>36,pipes=>17)
  PORT MAP (sysclk=>sysclk,reset=>'0',enable=>enable, -- no resets for memory
            aa=>numeratormantissaff,
            cc=>del_numeratormantissa);
   
  -- level 25 in, level 28 out
  cmt: fp_fxmul
  GENERIC MAP (widthaa=>36,widthbb=>36,widthcc=>72,
               pipes=>3,synthesize=>0)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,  
            dataaa=>del_numeratormantissa,
            databb=>denominatorinverse,
            result=>multiplier_tan);
 
  tanmantissa <= multiplier_tan(72 DOWNTO 37);
  
  gmna: FOR k IN 1 TO 24 GENERATE
    tanmantissanorm(k) <= (tanmantissa(k+9) AND NOT(tanmantissa(35))) OR
                          (tanmantissa(k+10) AND tanmantissa(35));
  END GENERATE;
  gmnb: FOR k IN 1 TO 9 GENERATE
    tanmantissatail(k) <= (tanmantissa(k) AND NOT(tanmantissa(35))) OR
                          (tanmantissa(k+1) AND tanmantissa(35));
  END GENERATE;
  
  overcheck(1) <= tanmantissanorm(1);
  gova: FOR k IN 2 TO 24 GENERATE
    overcheck(k) <= overcheck(k-1) AND tanmantissanorm(k); 
  END GENERATE;
    
  -- level 13 in, level 27 out
  ddena: fp_del 
  GENERIC MAP (width=>6,pipes=>14)
  PORT MAP (sysclk=>sysclk,reset=>'0',enable=>enable, -- no resets for memory
            aa=>inverseexponentff,
            cc=>del_inverseexponent); 
  
  -- level 8 in, level 27 out         
	dnumb: fp_del 
  GENERIC MAP (width=>5,pipes=>19)
  PORT MAP (sysclk=>sysclk,reset=>'0',enable=>enable, -- no resets for memory
            aa=>numeratorexponentff,
            cc=>del_numeratorexponent); 
                      
  tanexponent <= "01110111" + 
                (del_numeratorexponent(5) & del_numeratorexponent(5) & del_numeratorexponent(5) & del_numeratorexponent) + 
                (del_inverseexponent(6) & del_inverseexponent(6) & del_inverseexponent); -- 119 + exponent
  
  tanexponentnorm <= tanexponentff + tanmantissa(35);
  
  --*** handle small inputs ****
  dsma: fp_del
  GENERIC MAP (width=>23,pipes=>29)
  PORT MAP (sysclk=>sysclk,reset=>'0',enable=>enable, -- no resets for memory
            aa=>mantissain,
            cc=>small_mantissa); 
  dsxa: fp_del
  GENERIC MAP (width=>8,pipes=>29)
  PORT MAP (sysclk=>sysclk,reset=>'0',enable=>enable, -- no resets for memory
            aa=>exponentin,
            cc=>small_exponent); 
        
  exponentcheck <= exponentinff - 115;
                
  psa: PROCESS (sysclk,reset)
  BEGIN
  
    IF (reset = '1') THEN
      
      FOR k IN 1 TO 30 LOOP
        signff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 28 LOOP
        small_inputff(k) <= '0';
      END LOOP;
    
    ELSIF(rising_edge(sysclk)) THEN
      
      IF (enable = '1') THEN
         
        signff(1) <= signin;
        FOR k IN 2 TO 30 LOOP
          signff(k) <= signff(k-1);
        END LOOP;
           
        small_inputff(1) <= exponentcheck(8);
        FOR k IN 2 TO 28 LOOP
          small_inputff(k) <= small_inputff(k-1);
        END LOOP;
        
      END IF;
    
    END IF;
  
  END PROCESS;
  
  --mantissabase(1) <= (tanmantissanormff(1) AND NOT(small_inputff(28)));
  mantissabase(1) <= (roundbitff AND NOT(small_inputff(28)));
  gmba: FOR k IN 2 TO 24 GENERATE
    mantissabase(k) <= (small_mantissa(k-1) AND small_inputff(28)) OR
                       (tanmantissanormff(k) AND NOT(small_inputff(28)));
  END GENERATE;
  gxba: FOR k IN 1 TO 8 GENERATE
    exponentbase(k) <= (small_exponent(k) AND small_inputff(28)) OR
                       (tanexponentnormff(k) AND NOT(small_inputff(28)));
  END GENERATE;

  mantissaoutnode <= mantissabase(24 DOWNTO 2) + mantissabase(1);  

  exponentoutnode <= exponentbase + (overff AND NOT(small_inputff(28)));
  
  --***************
  --*** OUTPUTS ***
  --***************
  
  signout <= signff(30);
  mantissaout <= mantissaoutff;
  exponentout <= exponentoutff;
  
END rtl;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_TANLUT1.VHD                            ***
--***                                             ***
--***   Function: Tangent Look Up Table           ***
--***   (Generated by MATLAB Utility)             ***
--***                                             ***
--***   22/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_tanlut1 IS
PORT (
      add : IN STD_LOGIC_VECTOR (9 DOWNTO 1);
      mantissa : OUT STD_LOGIC_VECTOR (36 DOWNTO 1);
      exponent : OUT STD_LOGIC_VECTOR (5 DOWNTO 1)
     );
END fp_tanlut1;

ARCHITECTURE rtl OF fp_tanlut1 IS

BEGIN

  pca: PROCESS (add)
  BEGIN
    CASE add IS
      WHEN "000000000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(0,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(0,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(0,5);
      WHEN "000000001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(131072,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(174764,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(0,5);
      WHEN "000000010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(131074,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(174780,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(1,5);
      WHEN "000000011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(196617,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(130,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(1,5);
      WHEN "000000100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(131082,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(175036,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(2,5);
      WHEN "000000101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(163860,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(219287,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(2,5);
      WHEN "000000110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(196644,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(2074,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(2,5);
      WHEN "000000111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(229433,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(48174,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(2,5);
      WHEN "000001000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(131114,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(179133,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(3,5);
      WHEN "000001001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(147516,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(204485,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(3,5);
      WHEN "000001010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(163923,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(100723,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(3,5);
      WHEN "000001011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(180334,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(261788,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(3,5);
      WHEN "000001100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(196752,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(33207,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(3,5);
      WHEN "000001101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(213175,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(71403,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(3,5);
      WHEN "000001110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(229604,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(246559,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(3,5);
      WHEN "000001111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(246041,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(166927,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(3,5);
      WHEN "000010000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(131242,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(244778,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(4,5);
      WHEN "000010001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(139469,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(18368,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(4,5);
      WHEN "000010010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(147699,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(126224,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(4,5);
      WHEN "000010011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(155934,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(110829,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(4,5);
      WHEN "000010100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(164174,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(39099,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(4,5);
      WHEN "000010101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(172418,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(240249,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(4,5);
      WHEN "000010110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(180668,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(257224,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(4,5);
      WHEN "000010111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(188924,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(157429,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(4,5);
      WHEN "000011000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(197186,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(8449,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(4,5);
      WHEN "000011001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(205453,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(140199,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(4,5);
      WHEN "000011010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(213727,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(96362,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(4,5);
      WHEN "000011011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(222007,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(207256,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(4,5);
      WHEN "000011100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(230295,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(16983,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(4,5);
      WHEN "000011101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(238589,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(118443,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(4,5);
      WHEN "000011110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(246891,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(56191,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(4,5);
      WHEN "000011111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(255200,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(161457,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(4,5);
      WHEN "000100000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(131758,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(251787,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000100001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(135921,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(182851,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000100010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(140088,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(170994,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000100011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(144259,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(251287,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000100100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(148435,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(196795,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000100101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(152616,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(42877,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000100110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(156801,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(87190,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000100111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(160991,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(103258,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000101000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(165186,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(126910,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000101001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(169386,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(194144,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000101010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(173592,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(78984,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000101011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(177803,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(79918,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000101100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(182019,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(233473,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000101101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(186242,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(52073,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000101110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(190470,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(96910,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000101111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(194704,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(142940,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000110000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(198944,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(227466,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000110001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(203191,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(125851,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000110010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(207444,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(137961,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000110011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(211704,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(39590,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000110100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(215970,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(131044,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000110101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(220243,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(188568,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000110110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(224523,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(250786,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000110111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(228811,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(94417,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000111000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(233106,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(20713,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000111001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(237408,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(69033,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000111010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(241718,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(16848,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000111011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(246035,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(166180,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000111100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(250361,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(32888,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000111101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(254694,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(181681,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000111110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(259036,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(128971,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(5,5);
      WHEN "000111111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(131693,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(88946,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001000000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(133872,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(184862,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001000001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(136056,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(110880,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001000010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(138244,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(150087,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001000011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(140437,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(61438,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001000100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(142634,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(128336,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001000101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(144836,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(110058,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001000110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(147043,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(28193,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001000111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(149254,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(166641,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001001000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(151471,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(23046,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001001001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(153692,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(143802,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001001010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(155919,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(26909,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001001011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(158150,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(219127,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001001100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(160387,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(218828,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001001101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(162630,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(48862,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001001110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(164877,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(256563,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001001111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(167131,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(78745,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001010000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(169390,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(63145,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001010001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(171654,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(233418,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001010010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(173925,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(89145,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001010011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(176201,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(178694,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001010100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(178484,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(2082,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001010101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(180772,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(108121,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001010110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(183066,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(259423,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001010111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(185367,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(218831,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001011000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(187675,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(11570,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001011001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(189988,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(187394,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001011010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(192308,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(247729,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001011011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(194635,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(218538,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001011100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(196969,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(126042,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001011101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(199309,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(258866,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001011110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(201657,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(119470,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001011111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(204011,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(259160,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001100000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(206373,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(180942,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001100001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(208742,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(174537,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001100010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(211119,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(5664,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001100011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(213502,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(226767,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001100100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(215894,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(79866,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001100101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(218293,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(118006,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001100110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(220700,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(108111,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001100111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(223115,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(79560,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001101000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(225538,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(62056,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001101001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(227969,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(85630,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001101010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(230408,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(180644,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001101011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(232856,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(115658,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001101100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(235312,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(183865,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001101101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(237777,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(154523,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001101110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(240251,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(59395,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001101111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(242733,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(192751,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001110000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(245225,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(62806,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001110001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(247725,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(226729,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001110010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(250235,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(193502,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001110011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(252754,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(258933,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001110100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(255283,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(194946,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001110101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(257822,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(36018,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001110110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(260370,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(79189,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(6,5);
      WHEN "001110111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(131464,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(48818,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "001111000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(132748,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(63557,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "001111001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(134037,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(101912,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "001111010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(135331,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(182207,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "001111011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(136631,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(60853,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "001111100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(137936,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(18783,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "001111101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(139246,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(75024,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "001111110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(140561,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(248849,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "001111111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(141883,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(35488,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010000000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(143209,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(241146,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010000001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(144542,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(99421,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010000010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(145880,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(154894,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010000011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(147224,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(165983,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010000100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(148574,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(153522,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010000101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(149930,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(138624,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010000110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(151292,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(142687,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010000111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(152660,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(187397,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010001000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(154035,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(32592,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010001001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(155415,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(224845,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010001010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(156803,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(313,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010001011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(158196,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(168333,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010001100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(159596,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(227841,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010001101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(161003,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(202385,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010001110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(162417,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(115847,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010001111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(163837,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(254593,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010010000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(165265,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(118901,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010010001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(166699,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(257978,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010010010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(168141,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(172818,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010010011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(169590,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(151210,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010010100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(171046,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(219176,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010010101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(172510,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(140977,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010010110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(173981,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(205552,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010010111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(175460,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(177949,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010011000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(176947,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(85768,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010011001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(178441,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(219166,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010011010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(179944,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(82294,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010011011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(181454,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(228309,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010011100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(182973,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(162236,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010011101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(184500,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(175979,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010011110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(186036,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(37616,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010011111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(187580,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(39982,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010100000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(189132,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(214250,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010100001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(190694,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(67791,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010100010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(192264,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(157055,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010100011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(193843,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(252568,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010100100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(195432,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(125382,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010100101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(197030,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(71365,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010100110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(198637,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(124791,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010100111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(200254,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(58341,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010101000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(201880,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(169556,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010101001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(203516,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(232268,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010101010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(205163,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(20904,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010101011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(206819,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(96928,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010101100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(208485,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(235993,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010101101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(210162,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(214385,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010101110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(211850,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(71183,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010101111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(213548,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(108271,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010110000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(215257,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(103923,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010110001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(216977,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(99249,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010110010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(218708,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(136066,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010110011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(220450,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(256917,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010110100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(222204,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(242940,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010110101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(223970,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(138174,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010110110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(225747,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(249580,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010110111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(227537,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(98477,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010111000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(229338,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(255571,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010111001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(231152,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(243824,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010111010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(232979,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(111333,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010111011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(234818,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(169210,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010111100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(236670,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(205169,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010111101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(238536,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(7833,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010111110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(240414,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(153192,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "010111111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(242306,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(169612,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "011000000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(244212,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(110728,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "011000001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(246132,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(31174,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "011000010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(248065,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(248754,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "011000011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(250014,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(33745,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "011000100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(251976,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(230368,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "011000101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(253954,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(111078,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "011000110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(255946,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(260182,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "011000111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(257954,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(214570,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "011001000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(259978,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(36603,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "011001001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(262017,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(52004,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(7,5);
      WHEN "011001010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(132036,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(31728,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011001011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(133071,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(199603,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011001100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(134115,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(170119,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011001101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(135167,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(239798,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011001110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(136228,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(181565,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011001111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(137298,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(31195,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011010000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(138376,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(87334,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011010001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(139463,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(125082,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011010010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(140559,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(182447,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011010011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(141665,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(36078,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011010100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(142779,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(249858,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011010101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(143904,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(77779,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011010110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(145038,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(85397,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011010111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(146182,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(52708,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011011000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(147336,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(22748,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011011001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(148500,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(39467,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011011010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(149674,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(147762,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011011011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(150859,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(131351,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011011100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(152055,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(37096,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011011101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(153261,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(175023,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011011110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(154479,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(69779,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011011111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(155708,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(33524,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011100000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(156948,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(117385,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011100001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(158200,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(111488,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011100010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(159464,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(69279,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011100011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(160740,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(45413,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011100100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(162028,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(95789,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011100101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(163329,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(15442,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011100110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(164642,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(125012,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011100111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(165968,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(222206,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011101000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(167308,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(106129,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011101001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(168661,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(101608,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011101010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(170028,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(10664,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011101011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(171408,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(161129,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011101100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(172803,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(95974,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011101101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(174212,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(146219,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011101110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(175636,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(120264,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011101111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(177075,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(90370,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011110000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(178529,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(130571,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011110001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(179999,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(54581,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011110010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(181484,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(202287,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011110011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(182986,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(129087,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011110100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(184504,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(178815,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011110101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(186039,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(173083,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011110110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(187591,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(197786,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011110111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(189161,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(78873,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011111000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(190748,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(168858,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011111001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(192354,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(36174,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011111010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(193978,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(38109,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011111011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(195621,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(10173,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011111100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(197283,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(52606,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011111101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(198965,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(6187,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011111110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(200666,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(238745,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "011111111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(202389,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(72398,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100000000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(204132,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(142943,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100000001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(205897,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(40664,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100000010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(207683,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(145442,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100000011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(209492,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(54008,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100000100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(211323,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(152917,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100000101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(213178,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(45809,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100000110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(215056,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(126393,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100000111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(216959,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(5720,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100001000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(218886,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(85177,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100001001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(220838,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(245917,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100001010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(222817,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(111146,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100001011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(224822,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(94854,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100001100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(226854,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(91265,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100001101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(228913,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(261427,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100001110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(231001,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(246970,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100001111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(233118,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(218857,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100010000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(235265,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(91152,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100010001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(237442,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(45510,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100010010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(239650,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(7099,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100010011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(241889,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(169116,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100010100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(244161,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(206583,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100010101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(246467,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(63025,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100010110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(248806,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(212871,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100010111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(251181,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(88861,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100011000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(253591,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(179473,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100011001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(256038,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(194218,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100011010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(258523,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(112522,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100011011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(261046,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(184058,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(8,5);
      WHEN "100011100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(131804,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(202396,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100011101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(133106,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(127604,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100011110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(134429,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(5700,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100011111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(135772,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(241668,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100100000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(137138,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(196914,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100100001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(138527,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(24498,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100100010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(139938,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(145076,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100100011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(141373,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(198575,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100100100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(142833,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(93021,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100100101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(144318,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(4818,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100100110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(145828,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(116886,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100100111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(147365,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(94683,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100101000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(148929,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(135102,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100101001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(150521,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(180373,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100101010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(152142,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(180573,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100101011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(153793,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(94005,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100101100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(155474,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(149742,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100101101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(157187,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(61623,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100101110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(158932,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(77284,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100101111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(160710,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(192200,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100110000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(162523,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(150199,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100110001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(164371,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(230433,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100110010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(166256,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(199372,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100110011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(168179,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(97853,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100110100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(170140,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(241724,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100110101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(172142,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(173961,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100110110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(174185,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(238269,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100110111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(176272,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(6999,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100111000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(178402,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(116996,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100111001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(180578,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(173338,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100111010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(182802,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(61011,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100111011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(185074,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(208074,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100111100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(187398,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(13879,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100111101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(189773,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(209544,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100111110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(192203,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(237754,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "100111111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(194690,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(89118,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "101000000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(197235,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(41457,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "101000001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(199840,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(137068,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "101000010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(202508,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(184378,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "101000011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(205242,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(21881,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "101000100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(208043,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(44347,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "101000101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(210914,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(156319,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "101000110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(213859,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(36498,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "101000111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(216879,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(188732,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "101001000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(219979,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(109619,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "101001001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(223161,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(126346,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "101001010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(226429,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(89021,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "101001011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(229786,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(160435,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "101001100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(233237,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(33224,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "101001101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(236784,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(244509,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "101001110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(240434,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(83006,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "101001111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(244189,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(215105,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "101010000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(248056,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(68494,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "101010001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(252038,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(196984,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "101010010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(256142,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(189406,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "101010011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(260373,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(249093,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(9,5);
      WHEN "101010100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(132369,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(76283,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101010101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(134621,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(153043,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101010110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(136947,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(90777,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101010111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(139350,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(80594,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101011000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(141834,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(118724,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101011001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(144404,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(12410,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101011010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(147063,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(172855,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101011011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(149818,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(49588,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101011100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(152672,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(235640,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101011101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(155633,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(117182,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101011110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(158705,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(242792,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101011111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(161896,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(237423,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101100000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(165213,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(125600,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101100001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(168663,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(83253,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101100010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(172254,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(191313,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101100011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(175996,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(191297,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101100100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(179899,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(29637,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101100101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(183972,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(142533,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101100110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(188228,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(171026,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101100111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(192680,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(38953,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101101000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(197340,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(248662,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101101001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(202226,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(84469,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101101010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(207353,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(16170,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101101011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(212739,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(177173,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101101100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(218406,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(161382,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101101101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(224376,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(140334,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101101110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(230674,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(156722,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101101111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(237328,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(218000,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101110000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(244370,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(144312,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101110001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(251834,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(222783,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101110010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(259761,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(51093,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(10,5);
      WHEN "101110011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(134097,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(16112,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(11,5);
      WHEN "101110100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(138592,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(11144,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(11,5);
      WHEN "101110101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(143394,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(60483,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(11,5);
      WHEN "101110110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(148536,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(104003,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(11,5);
      WHEN "101110111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(154056,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(37731,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(11,5);
      WHEN "101111000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(159996,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(218457,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(11,5);
      WHEN "101111001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(166408,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(191255,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(11,5);
      WHEN "101111010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(173350,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(113148,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(11,5);
      WHEN "101111011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(180890,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(176944,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(11,5);
      WHEN "101111100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(189110,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(163200,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(11,5);
      WHEN "101111101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(198106,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(211327,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(11,5);
      WHEN "101111110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(207994,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(247747,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(11,5);
      WHEN "101111111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(218914,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(252397,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(11,5);
      WHEN "110000000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(231037,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(174172,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(11,5);
      WHEN "110000001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(244573,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(197553,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(11,5);
      WHEN "110000010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(259786,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(53842,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(11,5);
      WHEN "110000011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(138503,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(202780,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(12,5);
      WHEN "110000100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(148332,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(62994,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(12,5);
      WHEN "110000101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(159656,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(230897,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(12,5);
      WHEN "110000110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(172847,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(240508,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(12,5);
      WHEN "110000111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(188408,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(183509,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(12,5);
      WHEN "110001000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(207041,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(119228,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(12,5);
      WHEN "110001001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(229756,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(71260,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(12,5);
      WHEN "110001010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(258060,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(153597,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(12,5);
      WHEN "110001011" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(147154,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(32322,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(13,5);
      WHEN "110001100" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(171195,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(78299,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(13,5);
      WHEN "110001101" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(204618,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(105365,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(13,5);
      WHEN "110001110" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(254248,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(141622,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(13,5);
      WHEN "110001111" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(167825,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(19278,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(14,5);
      WHEN "110010000" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(246850,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(149873,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(14,5);
      WHEN "110010001" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(233251,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(216105,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(15,5);
      WHEN "110010010" =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(132278,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(191927,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(19,5);
      WHEN others =>
           mantissa(36 DOWNTO 19) <= conv_std_logic_vector(0,18);
           mantissa(18 DOWNTO 1) <= conv_std_logic_vector(0,18);
           exponent(5 DOWNTO 1) <= conv_std_logic_vector(0,5);
    END CASE;
  END PROCESS;

END rtl;
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all;

--***************************************************
--***                                             ***
--***   FLOATING POINT CORE LIBRARY               ***
--***                                             ***
--***   FP_TANLUT2.VHD                            ***
--***                                             ***
--***   Function: Tangent Look Up Table           ***
--***   (Generated by MATLAB Utility)             ***
--***                                             ***
--***   22/12/09 ML                               ***
--***                                             ***
--***   (c) 2009 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***                                             ***
--***                                             ***
--***************************************************

ENTITY fp_tanlut2 IS
PORT (
      add : IN STD_LOGIC_VECTOR (8 DOWNTO 1);
      tanfraction : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
     );
END fp_tanlut2;

ARCHITECTURE rtl OF fp_tanlut2 IS

BEGIN

  pca: PROCESS (add)
  BEGIN
    CASE add IS
      WHEN "00000000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(0,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(0,18);
      WHEN "00000001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(1024,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(0,18);
      WHEN "00000010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(2048,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(0,18);
      WHEN "00000011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(3072,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(1,18);
      WHEN "00000100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(4096,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(1,18);
      WHEN "00000101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(5120,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(3,18);
      WHEN "00000110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(6144,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(5,18);
      WHEN "00000111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(7168,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(7,18);
      WHEN "00001000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(8192,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(11,18);
      WHEN "00001001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(9216,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(15,18);
      WHEN "00001010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(10240,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(21,18);
      WHEN "00001011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(11264,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(28,18);
      WHEN "00001100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(12288,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(36,18);
      WHEN "00001101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(13312,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(46,18);
      WHEN "00001110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(14336,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(57,18);
      WHEN "00001111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(15360,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(70,18);
      WHEN "00010000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(16384,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(85,18);
      WHEN "00010001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(17408,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(102,18);
      WHEN "00010010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(18432,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(122,18);
      WHEN "00010011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(19456,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(143,18);
      WHEN "00010100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(20480,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(167,18);
      WHEN "00010101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(21504,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(193,18);
      WHEN "00010110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(22528,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(222,18);
      WHEN "00010111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(23552,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(253,18);
      WHEN "00011000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(24576,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(288,18);
      WHEN "00011001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(25600,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(326,18);
      WHEN "00011010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(26624,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(366,18);
      WHEN "00011011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(27648,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(410,18);
      WHEN "00011100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(28672,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(457,18);
      WHEN "00011101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(29696,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(508,18);
      WHEN "00011110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(30720,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(563,18);
      WHEN "00011111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(31744,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(621,18);
      WHEN "00100000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(32768,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(683,18);
      WHEN "00100001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(33792,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(749,18);
      WHEN "00100010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(34816,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(819,18);
      WHEN "00100011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(35840,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(893,18);
      WHEN "00100100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(36864,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(972,18);
      WHEN "00100101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(37888,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(1055,18);
      WHEN "00100110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(38912,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(1143,18);
      WHEN "00100111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(39936,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(1236,18);
      WHEN "00101000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(40960,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(1333,18);
      WHEN "00101001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(41984,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(1436,18);
      WHEN "00101010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(43008,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(1544,18);
      WHEN "00101011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(44032,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(1656,18);
      WHEN "00101100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(45056,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(1775,18);
      WHEN "00101101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(46080,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(1898,18);
      WHEN "00101110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(47104,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(2028,18);
      WHEN "00101111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(48128,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(2163,18);
      WHEN "00110000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(49152,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(2304,18);
      WHEN "00110001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(50176,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(2451,18);
      WHEN "00110010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(51200,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(2604,18);
      WHEN "00110011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(52224,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(2764,18);
      WHEN "00110100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(53248,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(2929,18);
      WHEN "00110101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(54272,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(3102,18);
      WHEN "00110110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(55296,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(3281,18);
      WHEN "00110111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(56320,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(3466,18);
      WHEN "00111000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(57344,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(3659,18);
      WHEN "00111001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(58368,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(3858,18);
      WHEN "00111010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(59392,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(4065,18);
      WHEN "00111011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(60416,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(4279,18);
      WHEN "00111100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(61440,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(4500,18);
      WHEN "00111101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(62464,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(4729,18);
      WHEN "00111110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(63488,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(4965,18);
      WHEN "00111111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(64512,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(5209,18);
      WHEN "01000000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(65536,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(5461,18);
      WHEN "01000001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(66560,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(5721,18);
      WHEN "01000010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(67584,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(5990,18);
      WHEN "01000011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(68608,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(6266,18);
      WHEN "01000100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(69632,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(6551,18);
      WHEN "01000101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(70656,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(6844,18);
      WHEN "01000110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(71680,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(7146,18);
      WHEN "01000111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(72704,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(7456,18);
      WHEN "01001000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(73728,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(7776,18);
      WHEN "01001001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(74752,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(8105,18);
      WHEN "01001010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(75776,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(8442,18);
      WHEN "01001011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(76800,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(8789,18);
      WHEN "01001100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(77824,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(9145,18);
      WHEN "01001101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(78848,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(9511,18);
      WHEN "01001110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(79872,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(9887,18);
      WHEN "01001111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(80896,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(10272,18);
      WHEN "01010000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(81920,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(10667,18);
      WHEN "01010001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(82944,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(11072,18);
      WHEN "01010010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(83968,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(11487,18);
      WHEN "01010011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(84992,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(11912,18);
      WHEN "01010100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(86016,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(12348,18);
      WHEN "01010101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(87040,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(12794,18);
      WHEN "01010110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(88064,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(13251,18);
      WHEN "01010111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(89088,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(13719,18);
      WHEN "01011000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(90112,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(14197,18);
      WHEN "01011001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(91136,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(14687,18);
      WHEN "01011010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(92160,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(15188,18);
      WHEN "01011011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(93184,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(15699,18);
      WHEN "01011100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(94208,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(16223,18);
      WHEN "01011101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(95232,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(16757,18);
      WHEN "01011110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(96256,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(17304,18);
      WHEN "01011111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(97280,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(17862,18);
      WHEN "01100000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(98304,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(18432,18);
      WHEN "01100001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(99328,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(19014,18);
      WHEN "01100010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(100352,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(19608,18);
      WHEN "01100011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(101376,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(20215,18);
      WHEN "01100100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(102400,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(20833,18);
      WHEN "01100101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(103424,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(21465,18);
      WHEN "01100110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(104448,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(22109,18);
      WHEN "01100111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(105472,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(22765,18);
      WHEN "01101000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(106496,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(23435,18);
      WHEN "01101001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(107520,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(24117,18);
      WHEN "01101010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(108544,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(24813,18);
      WHEN "01101011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(109568,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(25522,18);
      WHEN "01101100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(110592,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(26244,18);
      WHEN "01101101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(111616,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(26980,18);
      WHEN "01101110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(112640,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(27729,18);
      WHEN "01101111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(113664,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(28492,18);
      WHEN "01110000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(114688,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(29269,18);
      WHEN "01110001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(115712,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(30060,18);
      WHEN "01110010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(116736,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(30866,18);
      WHEN "01110011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(117760,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(31685,18);
      WHEN "01110100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(118784,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(32519,18);
      WHEN "01110101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(119808,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(33367,18);
      WHEN "01110110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(120832,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(34230,18);
      WHEN "01110111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(121856,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(35108,18);
      WHEN "01111000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(122880,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(36000,18);
      WHEN "01111001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(123904,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(36908,18);
      WHEN "01111010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(124928,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(37830,18);
      WHEN "01111011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(125952,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(38768,18);
      WHEN "01111100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(126976,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(39721,18);
      WHEN "01111101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(128000,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(40690,18);
      WHEN "01111110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(129024,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(41675,18);
      WHEN "01111111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(130048,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(42675,18);
      WHEN "10000000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(131072,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(43691,18);
      WHEN "10000001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(132096,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(44723,18);
      WHEN "10000010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(133120,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(45771,18);
      WHEN "10000011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(134144,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(46835,18);
      WHEN "10000100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(135168,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(47916,18);
      WHEN "10000101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(136192,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(49013,18);
      WHEN "10000110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(137216,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(50127,18);
      WHEN "10000111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(138240,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(51258,18);
      WHEN "10001000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(139264,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(52405,18);
      WHEN "10001001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(140288,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(53570,18);
      WHEN "10001010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(141312,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(54752,18);
      WHEN "10001011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(142336,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(55950,18);
      WHEN "10001100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(143360,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(57167,18);
      WHEN "10001101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(144384,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(58401,18);
      WHEN "10001110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(145408,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(59652,18);
      WHEN "10001111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(146432,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(60921,18);
      WHEN "10010000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(147456,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(62208,18);
      WHEN "10010001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(148480,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(63513,18);
      WHEN "10010010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(149504,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(64836,18);
      WHEN "10010011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(150528,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(66178,18);
      WHEN "10010100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(151552,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(67537,18);
      WHEN "10010101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(152576,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(68916,18);
      WHEN "10010110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(153600,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(70313,18);
      WHEN "10010111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(154624,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(71728,18);
      WHEN "10011000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(155648,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(73163,18);
      WHEN "10011001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(156672,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(74616,18);
      WHEN "10011010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(157696,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(76089,18);
      WHEN "10011011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(158720,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(77581,18);
      WHEN "10011100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(159744,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(79092,18);
      WHEN "10011101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(160768,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(80623,18);
      WHEN "10011110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(161792,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(82173,18);
      WHEN "10011111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(162816,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(83744,18);
      WHEN "10100000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(163840,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(85334,18);
      WHEN "10100001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(164864,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(86944,18);
      WHEN "10100010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(165888,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(88574,18);
      WHEN "10100011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(166912,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(90224,18);
      WHEN "10100100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(167936,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(91895,18);
      WHEN "10100101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(168960,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(93586,18);
      WHEN "10100110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(169984,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(95298,18);
      WHEN "10100111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(171008,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(97031,18);
      WHEN "10101000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(172032,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(98784,18);
      WHEN "10101001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(173056,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(100559,18);
      WHEN "10101010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(174080,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(102354,18);
      WHEN "10101011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(175104,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(104171,18);
      WHEN "10101100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(176128,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(106010,18);
      WHEN "10101101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(177152,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(107869,18);
      WHEN "10101110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(178176,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(109751,18);
      WHEN "10101111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(179200,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(111654,18);
      WHEN "10110000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(180224,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(113579,18);
      WHEN "10110001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(181248,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(115526,18);
      WHEN "10110010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(182272,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(117495,18);
      WHEN "10110011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(183296,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(119487,18);
      WHEN "10110100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(184320,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(121500,18);
      WHEN "10110101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(185344,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(123537,18);
      WHEN "10110110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(186368,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(125596,18);
      WHEN "10110111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(187392,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(127677,18);
      WHEN "10111000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(188416,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(129782,18);
      WHEN "10111001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(189440,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(131909,18);
      WHEN "10111010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(190464,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(134060,18);
      WHEN "10111011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(191488,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(136234,18);
      WHEN "10111100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(192512,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(138431,18);
      WHEN "10111101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(193536,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(140652,18);
      WHEN "10111110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(194560,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(142896,18);
      WHEN "10111111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(195584,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(145164,18);
      WHEN "11000000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(196608,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(147457,18);
      WHEN "11000001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(197632,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(149773,18);
      WHEN "11000010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(198656,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(152113,18);
      WHEN "11000011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(199680,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(154477,18);
      WHEN "11000100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(200704,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(156866,18);
      WHEN "11000101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(201728,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(159279,18);
      WHEN "11000110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(202752,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(161717,18);
      WHEN "11000111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(203776,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(164180,18);
      WHEN "11001000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(204800,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(166667,18);
      WHEN "11001001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(205824,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(169180,18);
      WHEN "11001010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(206848,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(171717,18);
      WHEN "11001011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(207872,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(174280,18);
      WHEN "11001100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(208896,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(176869,18);
      WHEN "11001101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(209920,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(179482,18);
      WHEN "11001110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(210944,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(182122,18);
      WHEN "11001111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(211968,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(184787,18);
      WHEN "11010000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(212992,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(187478,18);
      WHEN "11010001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(214016,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(190195,18);
      WHEN "11010010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(215040,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(192938,18);
      WHEN "11010011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(216064,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(195708,18);
      WHEN "11010100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(217088,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(198503,18);
      WHEN "11010101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(218112,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(201326,18);
      WHEN "11010110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(219136,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(204175,18);
      WHEN "11010111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(220160,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(207050,18);
      WHEN "11011000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(221184,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(209953,18);
      WHEN "11011001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(222208,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(212882,18);
      WHEN "11011010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(223232,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(215839,18);
      WHEN "11011011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(224256,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(218823,18);
      WHEN "11011100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(225280,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(221834,18);
      WHEN "11011101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(226304,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(224873,18);
      WHEN "11011110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(227328,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(227940,18);
      WHEN "11011111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(228352,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(231034,18);
      WHEN "11100000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(229376,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(234156,18);
      WHEN "11100001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(230400,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(237306,18);
      WHEN "11100010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(231424,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(240484,18);
      WHEN "11100011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(232448,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(243690,18);
      WHEN "11100100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(233472,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(246925,18);
      WHEN "11100101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(234496,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(250188,18);
      WHEN "11100110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(235520,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(253480,18);
      WHEN "11100111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(236544,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(256801,18);
      WHEN "11101000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(237568,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(260151,18);
      WHEN "11101001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(238593,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(1385,18);
      WHEN "11101010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(239617,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(4793,18);
      WHEN "11101011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(240641,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(8230,18);
      WHEN "11101100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(241665,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(11696,18);
      WHEN "11101101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(242689,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(15192,18);
      WHEN "11101110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(243713,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(18717,18);
      WHEN "11101111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(244737,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(22272,18);
      WHEN "11110000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(245761,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(25858,18);
      WHEN "11110001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(246785,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(29473,18);
      WHEN "11110010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(247809,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(33118,18);
      WHEN "11110011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(248833,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(36793,18);
      WHEN "11110100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(249857,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(40499,18);
      WHEN "11110101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(250881,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(44235,18);
      WHEN "11110110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(251905,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(48002,18);
      WHEN "11110111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(252929,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(51800,18);
      WHEN "11111000" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(253953,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(55628,18);
      WHEN "11111001" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(254977,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(59488,18);
      WHEN "11111010" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(256001,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(63379,18);
      WHEN "11111011" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(257025,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(67301,18);
      WHEN "11111100" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(258049,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(71254,18);
      WHEN "11111101" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(259073,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(75239,18);
      WHEN "11111110" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(260097,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(79255,18);
      WHEN "11111111" =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(261121,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(83303,18);
      WHEN others =>
           tanfraction(36 DOWNTO 19) <= conv_std_logic_vector(0,18);
           tanfraction(18 DOWNTO 1) <= conv_std_logic_vector(0,18);
    END CASE;
  END PROCESS;

END rtl;

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   ALTERA FLOATING POINT DATAPATH COMPILER   ***
--***                                             ***
--***   HCC_DIVFP1X.VHD                           ***
--***                                             ***
--***   Function: Internal format single divide - ***
--***              unsigned mantissa              ***
--***                                             ***
--***   Uses new multiplier based divider core    ***
--***   from floating point library               ***
--***                                             ***
--***   24/12/07 ML                               ***
--***                                             ***
--***   (c) 2007 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***   22/04/09 - added NAN support, IEEE NAN    ***
--***   output, sign bug                          ***
--***   11/08/09 - add divider interface output   ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--*** Latency = 13 (X)                            ***
--*** Latency = 13 (M)                            ***
--*** Latency = 13 (D)                            ***
--*** Latency = 13 + roundconvert (ieee)          ***
--***************************************************

ENTITY hcc_divfp1x IS 
GENERIC (
         mantissa : positive := 32; -- 32/36 mantissa
         ieeeoutput : integer := 1; -- 1 = ieee754 (1/u23/8)
         xoutput : integer := 0; -- 1 = single x format (s32/13)
         multoutput : integer := 0; -- 1 = to another single muliplier (s/1/34/10) - signed
         divoutput : integer := 0; -- 1 = to a single divider (s/1/34/10) - signed magnitude
         roundconvert : integer := 0;
         synthesize : integer := 0
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      aa : IN STD_LOGIC_VECTOR (mantissa+10 DOWNTO 1);
      aasat, aazip, aanan : IN STD_LOGIC; 
      bb : IN STD_LOGIC_VECTOR (mantissa+10 DOWNTO 1);
      bbsat, bbzip, bbnan : IN STD_LOGIC;
      
		  cc : OUT STD_LOGIC_VECTOR (32*ieeeoutput+(mantissa+10)*(xoutput+multoutput+divoutput) DOWNTO 1);
		  ccsat, cczip, ccnan : OUT STD_LOGIC
		);
END hcc_divfp1x;

ARCHITECTURE rtl OF hcc_divfp1x IS
    
  -- latency = 13 + ieeeoutput*roundconvert

  type divexpfftype IS ARRAY (11 DOWNTO 1) OF STD_LOGIC_VECTOR (10 DOWNTO 1);

  signal zerovec : STD_LOGIC_VECTOR (24 DOWNTO 1);
        
  -- multiplier core interface
  signal divinaaman, divinbbman : STD_LOGIC_VECTOR(mantissa DOWNTO 1);
  signal divinaaexp, divinbbexp : STD_LOGIC_VECTOR(10 DOWNTO 1);
  signal divinaaexpff, divinbbexpff : STD_LOGIC_VECTOR(10 DOWNTO 1);
  signal divinaasat, divinaazip, divinaanan : STD_LOGIC;
  signal divinbbsat, divinbbzip, divinbbnan : STD_LOGIC;
  signal divinaasatff, divinaazipff, divinaananff : STD_LOGIC;
  signal divinbbsatff, divinbbzipff, divinbbnanff : STD_LOGIC;
  signal divinaasign, divinbbsign : STD_LOGIC;
  signal divinaasignff, divinbbsignff : STD_LOGIC;
  signal divsignff : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal divsatff, divzipff, divnanff : STD_LOGIC_VECTOR (11 DOWNTO 1);
  signal divexpff : divexpfftype;
  signal dividend, divisor : STD_LOGIC_VECTOR (36 DOWNTO 1);
  signal divmannode : STD_LOGIC_VECTOR (36 DOWNTO 1);

  -- output section (x out)
  signal signeddivmannode : STD_LOGIC_VECTOR (mantissa DOWNTO 1);
  signal divxmanff : STD_LOGIC_VECTOR (mantissa DOWNTO 1);
  signal divxexpff : STD_LOGIC_VECTOR (10 DOWNTO 1);
  signal divxsatff, divxzipff, divxnanff : STD_LOGIC;

  -- output section (mult out)
  signal normalizemult : STD_LOGIC;
  signal normmultnode : STD_LOGIC_VECTOR (mantissa DOWNTO 1);
  signal signedmultnode : STD_LOGIC_VECTOR (mantissa DOWNTO 1);
  signal divmultmanff : STD_LOGIC_VECTOR (mantissa DOWNTO 1);
  signal divmultexpff : STD_LOGIC_VECTOR (10 DOWNTO 1);
  signal divmultsatff, divmultzipff, divmultnanff : STD_LOGIC;
      
  -- output section (div out)
  signal normalizediv : STD_LOGIC;
  signal normdivnode : STD_LOGIC_VECTOR (mantissa-1 DOWNTO 1);
  signal divdivsignff : STD_LOGIC;
  signal divdivmanff : STD_LOGIC_VECTOR (mantissa-1 DOWNTO 1);
  signal divdivexpff : STD_LOGIC_VECTOR (10 DOWNTO 1);
  signal divdivsatff, divdivzipff, divdivnanff : STD_LOGIC;  

  -- output section (ieeeout)  
  signal normalize : STD_LOGIC;
  signal normmannode : STD_LOGIC_VECTOR (25 DOWNTO 1);
  signal manoverflow : STD_LOGIC_VECTOR (24 DOWNTO 1);
  signal ccmanff : STD_LOGIC_VECTOR (24 DOWNTO 1);
  signal ccexpff : STD_LOGIC_VECTOR (10 DOWNTO 1);
  signal divexpminus : STD_LOGIC_VECTOR (10 DOWNTO 1);
  signal ccsignff, ccsatff, cczipff, ccnanff, ccoverff : STD_LOGIC;
  signal manoutff : STD_LOGIC_VECTOR (23 DOWNTO 1);
  signal expoutff : STD_LOGIC_VECTOR (8 DOWNTO 1);
  signal signoutff : STD_LOGIC;
  signal ccexpplus : STD_LOGIC_VECTOR (10 DOWNTO 1);
  signal expmax, expzero : STD_LOGIC;
  signal manoutzero, manoutmax, expoutzero, expoutmax : STD_LOGIC;
     
  -- Signals to convert division format to mult format
  signal aaxor : STD_LOGIC_VECTOR (mantissa DOWNTO 1);
  signal bbxor : STD_LOGIC_VECTOR (mantissa DOWNTO 1);

  -- 12 latency
  component fp_div_core IS 
  GENERIC (synthesize : integer := 1);
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dividend : IN STD_LOGIC_VECTOR (36 DOWNTO 1);
        divisor : IN STD_LOGIC_VECTOR (36 DOWNTO 1);

		  quotient : OUT STD_LOGIC_VECTOR (36 DOWNTO 1)
		  );
  end component;
  
BEGIN
 
  gza: IF (ieeeoutput = 1) GENERATE
    gzb: FOR k IN 1 TO 24 GENERATE
      zerovec(k) <= '0';
    END GENERATE;
  END GENERATE;

  --**************************************************
  --***                                            ***
  --*** Input Section                              *** 
  --***                                            ***
  --**************************************************

  --********************************************************
  --*** NOTE THAT THE SIGN BIT IS PACKED IN THE MSB OF   ***
  --*** THE MANTISSA                                     ***
  --********************************************************

  aaxor <= (others => aa(mantissa+10));
  bbxor <= (others => bb(mantissa+10));

  divinaaman <= (aa(mantissa+9 DOWNTO 11) & '0') XOR aaxor;
  divinaaexp <= aa(10 DOWNTO 1);
  divinbbman <= (bb(mantissa+9 DOWNTO 11) & '0') XOR bbxor;
  divinbbexp <= bb(10 DOWNTO 1);
  divinaasat <= aasat;
  divinbbsat <= bbsat;
  divinaazip <= aazip;
  divinbbzip <= bbzip;
  divinaanan <= aanan;
  divinbbnan <= bbnan;
  -- signbits packed in MSB of mantissas
  divinaasign <= aa(mantissa+10);
  divinbbsign <= bb(mantissa+10);

  --**************************************************
  --***                                            ***
  --*** Divider Section                            *** 
  --***                                            ***
  --**************************************************

  gdda: IF (mantissa = 32) GENERATE
    dividend <= divinaaman & "0000";
    divisor <= divinbbman & "0000";
  END GENERATE;
  gddb: IF (mantissa = 36) GENERATE
    dividend <= divinaaman;
    divisor <= divinbbman;
  END GENERATE;

  -- 12 latency
  div: fp_div_core
  GENERIC MAP (synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dividend=>dividend,divisor=>divisor,
            quotient=>divmannode);

  -- 12 pipes here : 1 input stage, so 11 stages left 
  pda: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN
        
      FOR k IN 1 TO 10 LOOP
        divinaaexpff(k) <= '0';
        divinbbexpff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 11 LOOP
        FOR j IN 1 TO 10 LOOP
          divexpff(k)(j) <= '0';
        END LOOP;
      END LOOP;
      divinaasignff <= '0';
      divinbbsignff <= '0';
      divinaasatff <= '0';
      divinbbsatff <= '0';
      divinaazipff <= '0';
      divinbbzipff <= '0';
      divinaananff <= '0';
      divinbbnanff <= '0';
      FOR k IN 1 TO 11 LOOP
        divsignff(k) <= '0';
        divsatff(k) <= '0';
        divzipff(k) <= '0';
        divnanff(k) <= '0';
      END LOOP;
         
    ELSIF (rising_edge(sysclk)) THEN
        
      IF (enable = '1') THEN
          
        divinaaexpff <= divinaaexp;
        divinbbexpff <= divinbbexp;
        divexpff(1)(10 DOWNTO 1) <= divinaaexpff - divinbbexpff;
        divexpff(2)(10 DOWNTO 1) <= divexpff(1)(10 DOWNTO 1) + "0001111111";
        FOR k IN 3 TO 11 LOOP
          divexpff(k)(10 DOWNTO 1) <= divexpff(k-1)(10 DOWNTO 1);
        END LOOP; 
        
        divinaasignff <= divinaasign;
        divinbbsignff <= divinbbsign;
        divsignff(1) <= divinaasignff XOR divinbbsignff;
        FOR k IN 2 TO 11 LOOP
          divsignff(k) <= divsignff(k-1);
        END LOOP;
     
        divinaasatff <= divinaasat;
        divinbbsatff <= divinbbsat;
        divinaazipff <= divinaazip;
        divinbbzipff <= divinbbzip;
        divinaananff <= divinaanan;
        divinbbnanff <= divinbbnan;
        -- special condition: infinity = x/0
        divsatff(1) <= (divinaasatff OR divinbbsatff) OR
                       (NOT(divinaazipff) AND divinbbzipff);
        divzipff(1) <= divinaazipff;
        -- 0/0 or infinity/infinity is invalid OP, NAN out
        divnanff(1) <= divinaananff OR divinbbnanff OR 
                      (divinaazipff AND divinbbzipff) OR
                      (divinaasatff AND divinbbsatff);
        FOR k IN 2 TO 11 LOOP
          divsatff(k) <= divsatff(k-1);
          divzipff(k) <= divzipff(k-1);
          divnanff(k) <= divnanff(k-1);
        END LOOP;
         
      END IF;
        
    END IF;
      
  END PROCESS;
       
  --**************************************************
  --***                                            ***
  --*** Output Section                             *** 
  --***                                            ***
  --**************************************************

  --********************************************************
  --*** internal format output, convert back to signed   ***
  --*** no need for fine normalization                   ***
  --********************************************************    
   
  goxa: IF (xoutput = 1) GENERATE 
    
    goxb: FOR k IN 1 TO mantissa-5 GENERATE
      signeddivmannode(k) <= divmannode(36-mantissa+5+k) XOR divsignff(11);
    END GENERATE;
    goxc: FOR k IN mantissa-4 TO mantissa GENERATE
      signeddivmannode(k) <= divsignff(11);
    END GENERATE;

    pox: PROCESS (sysclk,reset)
    BEGIN
        
      IF (reset = '1') THEN
          
        FOR k IN 1 TO mantissa LOOP
          divxmanff(k) <= '0';
        END LOOP;
        divxexpff <= "0000000000";
        divxsatff <= '0';
        divxzipff <= '0';
        divxnanff <= '0';
      
      ELSIF (rising_edge(sysclk)) THEN
      
        IF (enable = '1') THEN
            
          divxmanff <= signeddivmannode;
          
          divxexpff(10 DOWNTO 1) <= divexpff(11)(10 DOWNTO 1);
          
          divxsatff <= divsatff(11);
          divxzipff <= divzipff(11);
          divxnanff <= divnanff(11);

        END IF;        
              
      END IF;
        
    END PROCESS;
       
    cc(mantissa+10 DOWNTO 11) <= divxmanff;
    cc(10 DOWNTO 1) <= divxexpff(10 DOWNTO 1);
    ccsat <= divxsatff;
    cczip <= divxzipff;
    ccnan <= divxnanff;
    
  END GENERATE;

  --*********************************
  --*** multiplier format output  ***
  --*********************************  
   
  gofa: IF (multoutput = 1) GENERATE 
  
    -- output either "01XXX" (0.5 < x < 1) or "1XXX" (1 < x < 2), normalize to "01XXX"
    -- this is opposite direction to divider normalization
    normalizemult <= NOT(divmannode(36));
    goeb: FOR k IN 1 TO mantissa-1 GENERATE -- includes leading '1' and round bit
      normmultnode(k) <= (divmannode(36-mantissa+k) AND     normalizemult) OR
                         (divmannode(37-mantissa+k) AND NOT(normalizemult));
    END GENERATE;
    normmultnode(mantissa) <= '0';
    goec: FOR k IN 1 TO mantissa GENERATE
      signedmultnode(k) <= normmultnode(k) XOR divsignff(11);
    END GENERATE;
    
    pof: PROCESS (sysclk,reset)
    BEGIN
        
      IF (reset = '1') THEN
          
        FOR k IN 1 TO mantissa LOOP
          divmultmanff(k) <= '0';
        END LOOP;
        divmultexpff <= "0000000000";
        divmultsatff <= '0';
        divmultzipff <= '0';
        divmultnanff <= '0';
      
      ELSIF (rising_edge(sysclk)) THEN
      
        IF (enable = '1') THEN

          divmultmanff <= signedmultnode + divsignff(11);
          
          divmultexpff(10 DOWNTO 1) <= divexpff(11)(10 DOWNTO 1) - normalizemult;
          
          divmultsatff <= divsatff(11);
          divmultzipff <= divzipff(11);
          divmultnanff <= divnanff(11);

        END IF;        
              
      END IF;
        
    END PROCESS;

    cc(mantissa+10 DOWNTO 11) <= divmultmanff;
    cc(10 DOWNTO 1) <= divmultexpff(10 DOWNTO 1);
    ccsat <= divmultsatff;
    cczip <= divmultzipff;
    ccnan <= divmultnanff;
    
  END GENERATE; 
   
  --******************************
  --*** divider format output  ***
  --******************************  
   
  goda: IF (divoutput = 1) GENERATE 
  
    -- output either "01XXX" (0.5 < x < 1) or "1XXX" (1 < x < 2), normalize to "1XXX"
    normalizediv <= NOT(divmannode(36));
    godb: FOR k IN 1 TO mantissa-1 GENERATE -- includes leading '1' and round bit
      normdivnode(k) <= (divmannode(36-mantissa+k) AND     normalizediv) OR
                        (divmannode(37-mantissa+k) AND NOT(normalizediv));
    END GENERATE;
    
    pof: PROCESS (sysclk,reset)
    BEGIN
        
      IF (reset = '1') THEN
          
        divdivsignff <= '0';
        FOR k IN 1 TO mantissa-1 LOOP
          divdivmanff(k) <= '0';
        END LOOP;
        divdivexpff <= "0000000000";
        divdivsatff <= '0';
        divdivzipff <= '0';
        divdivnanff <= '0';
      
      ELSIF (rising_edge(sysclk)) THEN
      
        IF (enable = '1') THEN
            
          divdivsignff <= divsignff(11);
           
          divdivmanff <= normdivnode;
          
          divdivexpff(10 DOWNTO 1) <= divexpff(11)(10 DOWNTO 1) - normalizediv;
          
          divdivsatff <= divsatff(11);
          divdivzipff <= divzipff(11);
          divdivnanff <= divnanff(11);

        END IF;        
              
      END IF;
        
    END PROCESS;
    
    cc(mantissa+10) <= divdivsignff;
    cc(mantissa+9 DOWNTO 11) <= divdivmanff;
    cc(10 DOWNTO 1) <= divdivexpff(10 DOWNTO 1);
    ccsat <= divdivsatff;
    cczip <= divdivzipff;
    ccnan <= divdivnanff;
    
  END GENERATE;
  
  --********************************************************
  --*** if output directly out of datapath, convert here ***
  --********************************************************
  goea: IF (ieeeoutput = 1) GENERATE -- ieee754 out of datapath, do conversion
     
    -- output either "01XXX" (0.5 < x < 1) or "1XXX" (1 < x < 2), normalize to "1XXX"
    normalize <= NOT(divmannode(36));
    goeb: FOR k IN 1 TO 25 GENERATE -- includes leading '1' and round bit
      normmannode(k) <= (divmannode(k+11) AND NOT(normalize)) OR
                        (divmannode(k+10) AND normalize);
    END GENERATE;
                  
    -- always round, need 
    goec: IF (roundconvert = 0) GENERATE

      poea: PROCESS (sysclk,reset)
      BEGIN
    
        IF (reset = '1') THEN
        
          FOR k IN 1 TO 23 LOOP
            manoutff(k) <= '0';  
          END LOOP; 
          FOR k IN 1 TO 8 LOOP
            expoutff(k) <= '0';  
          END LOOP; 
          signoutff <= '0';
          
        ELSIF (rising_edge(sysclk)) THEN
           
          IF (enable = '1') THEN  
            FOR k IN 1 TO 23 LOOP
              manoutff(k) <= (normmannode(k+1) AND NOT(manoutzero)) OR manoutmax;
            END LOOP;
            FOR k IN 1 TO 8 LOOP
              expoutff(k) <= (divexpminus(k) AND NOT(expoutzero)) OR expoutmax;
            END LOOP;
            signoutff <= divsignff(11);
          END IF;
                
        END IF;
        
      END PROCESS;

      divexpminus <= divexpff(11)(10 DOWNTO 1) - ("000000000" & normalize);
      
      -- both '1' when true
      expmax <= divexpminus(8) AND divexpminus(7) AND divexpminus(6) AND divexpminus(5) AND 
                divexpminus(4) AND divexpminus(3) AND divexpminus(2) AND divexpminus(1);
      expzero <= NOT(divexpminus(8) OR divexpminus(7) OR divexpminus(6) OR divexpminus(5) OR 
                     divexpminus(4) OR divexpminus(3) OR divexpminus(2) OR divexpminus(1));      
                     
      -- any special condition turns mantissa zero
      manoutzero <= divsatff(11) OR divzipff(11) OR expmax OR expzero OR 
                    divexpminus(10) OR divexpminus(9);
      manoutmax <= divnanff(11);
      expoutzero <= divzipff(11) OR expzero OR divexpminus(10);
      -- 12/05/09 - make sure ccexpminus = -1 doesnt create infinity
      expoutmax <= (expmax AND NOT(divexpminus(9)) AND NOT(divexpminus(10))) OR 
                   (divexpminus(9) AND NOT(divexpminus(10))) OR divnanff(11);  
      
    END GENERATE;
  
    goed: IF (roundconvert = 1) GENERATE
            
      manoverflow(1) <= normmannode(1);
      gva: FOR k IN 2 TO 24 GENERATE
        manoverflow(k) <= manoverflow(k-1) AND normmannode(k);
      END GENERATE;
  
      poeb: PROCESS (sysclk,reset)
      BEGIN
    
        IF (reset = '1') THEN
          
          FOR k IN 1 TO 24 LOOP
            ccmanff(k) <= '0';
          END LOOP;
          FOR k IN 1 TO 10 LOOP
            ccexpff(k) <= '0';
          END LOOP;
          ccsignff <= '0';
          ccsatff <= '0';
          cczipff <= '0';
          ccnanff <= '0';
          ccoverff <= '0';
          FOR k IN 1 TO 23 LOOP
            manoutff(k) <= '0';
          END LOOP;
          FOR k IN 1 TO 8 LOOP
            expoutff(k) <= '0';
          END LOOP;
          signoutff <= '0';
        
        ELSIF (rising_edge(sysclk)) THEN
        
          IF (enable = '1') THEN   
           
            ccmanff <= normmannode(25 DOWNTO 2) + (zerovec(23 DOWNTO 1) & normmannode(1));
            ccexpff(10 DOWNTO 1) <= divexpff(11)(10 DOWNTO 1) - ("000000000" & normalize);
            ccsignff <= divsignff(11);
            ccsatff <= divsatff(11);
            cczipff <= divzipff(11);
            ccnanff <= divnanff(11);
            ccoverff <= manoverflow(23);
          
            FOR k IN 1 TO 23 LOOP
              manoutff(k) <= (ccmanff(k) AND NOT(manoutzero)) OR manoutmax; 
            END LOOP;
            FOR k IN 1 TO 8 LOOP
              expoutff(k) <= (ccexpplus(k) AND NOT(expoutzero)) OR expoutmax;
            END LOOP;
            signoutff <= ccsignff;
      
          END IF;
          
        END IF;
        
      END PROCESS;

      ccexpplus <= ccexpff + ("000000000" & ccoverff);
      
       -- both '1' when true
      expmax <= ccexpplus(8) AND ccexpplus(7) AND ccexpplus(6) AND ccexpplus(5) AND 
                ccexpplus(4) AND ccexpplus(3) AND ccexpplus(2) AND ccexpplus(1);
      expzero <= NOT(ccexpplus(8) OR ccexpplus(7) OR ccexpplus(6) OR ccexpplus(5) OR 
                     ccexpplus(4) OR ccexpplus(3) OR ccexpplus(2) OR ccexpplus(1));      
                     
      -- any special condition turns mantissa zero
      manoutzero <= ccsatff OR cczipff OR expmax OR expzero OR 
                    ccexpplus(10) OR ccexpplus(9);
      manoutmax <= ccnanff;
      expoutzero <= cczipff OR expzero OR ccexpplus(10);
      -- 12/05/09 - make sure ccexpplus = -1 doesnt create infinity
      expoutmax <= (expmax AND NOT(ccexpplus(9)) AND NOT(ccexpplus(10))) OR 
                   (ccexpplus(9) AND NOT(ccexpplus(10))) OR ccnanff;  
    
    END GENERATE;
    
    cc(32) <= signoutff;
    cc(31 DOWNTO 24) <= expoutff;
    cc(23 DOWNTO 1) <= manoutff;
    -- dummy only
    ccsat <= '0';
    cczip <= '0';   
    ccnan <= '0';
      
  END GENERATE;
    
END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   ALTERA FLOATING POINT DATAPATH COMPILER   ***
--***                                             ***
--***   HCC_DIVFP2X.VHD                           ***
--***                                             ***
--***   Function: Internal format double divide - ***
--***              unsigned mantissa              ***
--***                                             ***
--***   Uses new multiplier based divider core    ***
--***   from floating point library               ***
--***                                             ***
--***   24/12/07 ML                               ***
--***                                             ***
--***   (c) 2007 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***   23/04/09 - added NAN support              ***
--***   27/04/09 - added SIII/SIV support         ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes:                                      ***
--***                                             ***
--*** Stratix II                                  ***
--*** Latency = 20 + 4*doublespeed +              ***
--*** doublespeed*roundconvert (Y)                ***
--*** Latency = 20 + 4*doublespeed (F)            ***
--*** Latency = 20 + 4*doublespeed +              ***
--*** roundconvert*(1+doublespeed) (ieee)         ***
--***                                             ***
--*** Stratix III/IV                              ***
--*** Latency = 19 + 2*doublespeed +              ***
--*** doublespeed*roundconvert (Y)                ***
--*** Latency = 19 + 2*doublespeed (F)            ***
--*** Latency = 19 + 2*doublespeed +              ***
--*** roundconvert*(1+doublespeed) (ieee)         ***
--***************************************************

ENTITY hcc_divfp2x IS 
GENERIC (
         ieeeoutput : integer := 0; -- 1 = ieee754 (1/u52/11)
         xoutput : integer := 1; -- 1 = double x format (s64/13)
         divoutput : integer := 1; -- output to another multiplier or divider (S'1'u54/13)
         roundconvert : integer := 1; -- global switch - round all ieee<=>x conversion when '1'
         doublespeed : integer := 0; -- global switch - '0' unpiped adders, '1' piped adders for doubles
         doubleaccuracy : integer := 0; -- 0 = pruned multiplier, 1 = normal multiplier
         device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
         synthesize : integer := 1
        );
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      aa : IN STD_LOGIC_VECTOR (67 DOWNTO 1);
      aasat, aazip, aanan : IN STD_LOGIC; 
      bb : IN STD_LOGIC_VECTOR (67 DOWNTO 1);
      bbsat, bbzip, bbnan : IN STD_LOGIC;
      
		cc : OUT STD_LOGIC_VECTOR (64+13*xoutput+3*divoutput DOWNTO 1);
		ccsat, cczip, ccnan : OUT STD_LOGIC
		);
END hcc_divfp2x;

ARCHITECTURE rtl OF hcc_divfp2x IS

  -- SII: div_core latency 19+4*doublespeed 
  -- SIII/IV: div_core latency 18+2*doublespeed 
  constant midlatency : positive := 18+4*doublespeed - device - 2*device*doublespeed;
  
  type divinexpfftype IS ARRAY (midlatency DOWNTO 1) OF STD_LOGIC_VECTOR (13 DOWNTO 1);
  type divexpdelfftype IS ARRAY (2 DOWNTO 1) OF STD_LOGIC_VECTOR (13 DOWNTO 1);
  
  signal zerovec : STD_LOGIC_VECTOR (64 DOWNTO 1);
        
  -- divider core interface
  signal divinaaman, divinbbman : STD_LOGIC_VECTOR(53 DOWNTO 1);
  signal divinaaexp, divinbbexp : STD_LOGIC_VECTOR(13 DOWNTO 1);
  signal divinaaexpff, divinbbexpff : STD_LOGIC_VECTOR(13 DOWNTO 1);
  signal divinaasat, divinaazip, divinaanan : STD_LOGIC;
  signal divinbbsat, divinbbzip, divinbbnan : STD_LOGIC;
  signal divinaasatff, divinaazipff, divinaananff : STD_LOGIC;
  signal divinbbsatff, divinbbzipff, divinbbnanff : STD_LOGIC;
  signal divinaasign, divinbbsign : STD_LOGIC;
  signal divinaasignff, divinbbsignff : STD_LOGIC;
  signal divinexpff : divinexpfftype;
  signal divinsignff : STD_LOGIC_VECTOR (midlatency DOWNTO 1);
  signal divinsatff, divinzipff, divinnanff : STD_LOGIC_VECTOR (midlatency DOWNTO 1);
  signal dividend, divisor : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal divmannode : STD_LOGIC_VECTOR (55 DOWNTO 1);

  -- output section (x out)
  signal signeddivmannode : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal divroundnode : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal divmanout : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal divymanff : STD_LOGIC_VECTOR (64 DOWNTO 1);
  signal divyexpff : STD_LOGIC_VECTOR (13 DOWNTO 1);
  signal divysatbitff, divyzipbitff, divynanbitff : STD_LOGIC;
  signal divexpplus : STD_LOGIC_VECTOR (13 DOWNTO 1);
  signal divyexpdelff : divexpdelfftype;
  signal divysatdelff, divyzipdelff, divynandelff : STD_LOGIC_VECTOR (2 DOWNTO 1);
  signal divsatbase, divzipbase : STD_LOGIC;
  
  -- output section (divout)
  signal normmannode : STD_LOGIC_VECTOR (53 DOWNTO 1);
  signal divdivmanff : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal divdivexpff : STD_LOGIC_VECTOR (13 DOWNTO 1);
  signal divdivsatff, divdivzipff, divdivnanff : STD_LOGIC;
        
  -- output section (ieeeout)  
  signal normsignff, normsatff, normzipff, normnanff : STD_LOGIC;
  signal normalize : STD_LOGIC;
  signal normalnode : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal normalff : STD_LOGIC_VECTOR (54 DOWNTO 1);
  signal normalexpff : STD_LOGIC_VECTOR (13 DOWNTO 1);
                                
  component hcc_addpipeb
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
        carryin : IN STD_LOGIC;
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
  end component;

  component hcc_addpipes
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
        carryin : IN STD_LOGIC;
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
  end component;

  -- SII: latency 19+4*doublespeed 
  -- SIII/IV: latency 18+2*doublespeed 
  component dp_div_core IS 
  GENERIC (
         doublespeed : integer := 0; -- 0/1
         doubleaccuracy : integer := 0;  -- 0 = pruned multiplier, 1 = normal multiplier
         device : integer := 0; -- 0 = "Stratix II", 1 = "Stratix III" (also 4)
         synthesize : integer := 1      -- 0/1      
        ); 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        dividend : IN STD_LOGIC_VECTOR (54 DOWNTO 1);
        divisor : IN STD_LOGIC_VECTOR (54 DOWNTO 1);

		  quotient : OUT STD_LOGIC_VECTOR (55 DOWNTO 1)
		  );
  end component;

  -- latency 1
  component hcc_divnornd 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        signin : IN STD_LOGIC;
        exponentin : IN STD_LOGIC_VECTOR (13 DOWNTO 1);
        mantissain : IN STD_LOGIC_VECTOR (53 DOWNTO 1); -- includes roundbit
        satin, zipin, nanin : IN STD_LOGIC;

		  signout : OUT STD_LOGIC;
        exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
        mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1)
		 );
  end component;
  
  -- latency 2
  component hcc_divrnd
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        signin : IN STD_LOGIC;
        exponentin : IN STD_LOGIC_VECTOR (13 DOWNTO 1);
        mantissain : IN STD_LOGIC_VECTOR (53 DOWNTO 1); -- includes roundbit
        satin, zipin, nanin : IN STD_LOGIC;

		  signout : OUT STD_LOGIC;
        exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
        mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1)
		 );
  end component; 
  
  -- latency 3
  component hcc_divrndpipe 
  GENERIC (synthesize : integer := 1); 
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        signin : IN STD_LOGIC;
        exponentin : IN STD_LOGIC_VECTOR (13 DOWNTO 1);
        mantissain : IN STD_LOGIC_VECTOR (53 DOWNTO 1); -- includes roundbit
        satin, zipin, nanin : IN STD_LOGIC;

		  signout : OUT STD_LOGIC;
        exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
        mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1)
		 );
  end component;
    
BEGIN
 
  gza: FOR k IN 1 TO 64 GENERATE
    zerovec(k) <= '0';
  END GENERATE;

  --**************************************************
  --***                                            ***
  --*** Input Section                              *** 
  --***                                            ***
  --**************************************************

  --********************************************************
  --*** NOTE THAT THE SIGN BIT IS PACKED IN THE MSB OF   ***
  --*** THE MANTISSA                                     ***
  --********************************************************

  divinaaman <= aa(66 DOWNTO 14);
  divinaaexp <= aa(13 DOWNTO 1);
  divinbbman <= bb(66 DOWNTO 14);
  divinbbexp <= bb(13 DOWNTO 1);
  divinaasat <= aasat;
  divinbbsat <= bbsat;
  divinaazip <= aazip;
  divinbbzip <= bbzip;
  divinaanan <= aanan;
  divinbbnan <= bbnan;
  -- signbits packed in MSB of mantissas
  divinaasign <= aa(67);
  divinbbsign <= bb(67);

  --**************************************************
  --***                                            ***
  --*** Divider Section                            *** 
  --***                                            ***
  --**************************************************
  
  dividend <= divinaaman & '0';
  divisor <= divinbbman & '0';
  
  -- SII: latency 19+4*doublespeed 
  -- SIII/IV: latency 18+2*doublespeed 
  div: dp_div_core
  GENERIC MAP (doublespeed=>doublespeed,doubleaccuracy=>doubleaccuracy,
               device=>device,synthesize=>synthesize)
  PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
            dividend=>dividend,divisor=>divisor,
            quotient=>divmannode);
        
  pda: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN
        
      FOR k IN 1 TO 13 LOOP
        divinaaexpff(k) <= '0';
        divinbbexpff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO midlatency LOOP
        FOR j IN 1 TO 13 LOOP
          divinexpff(k)(j) <= '0';
        END LOOP;
      END LOOP;
      divinaasignff <= '0';
      divinbbsignff <= '0';
      divinaasatff <= '0';
      divinbbsatff <= '0';
      divinaazipff <= '0';
      divinbbzipff <= '0';
      divinaananff <= '0';
      divinbbnanff <= '0';
      FOR k IN 1 TO midlatency LOOP
        divinsignff(k) <= '0';
        divinsatff(k) <= '0';
        divinzipff(k) <= '0';
        divinnanff(k) <= '0';
      END LOOP;
         
    ELSIF (rising_edge(sysclk)) THEN
        
      IF (enable = '1') THEN
          
        divinaaexpff <= divinaaexp;
        divinbbexpff <= divinbbexp;
        divinexpff(1)(13 DOWNTO 1) <= divinaaexpff - divinbbexpff;
        divinexpff(2)(13 DOWNTO 1) <= divinexpff(1)(13 DOWNTO 1) + "0001111111111";
        FOR k IN 3 TO midlatency LOOP
          divinexpff(k)(13 DOWNTO 1) <= divinexpff(k-1)(13 DOWNTO 1);
        END LOOP; 
        
        divinaasignff <= divinaasign;
        divinbbsignff <= divinbbsign;
        divinsignff(1) <= divinaasignff XOR divinbbsignff;
        FOR k IN 2 TO midlatency LOOP
          divinsignff(k) <= divinsignff(k-1);
        END LOOP;
     
        divinaasatff <= divinaasat;
        divinbbsatff <= divinbbsat;
        divinaazipff <= divinaazip;
        divinbbzipff <= divinbbzip;
        divinaananff <= divinaanan;
        divinbbnanff <= divinbbnan;
        -- special condition: infinity = x/0
        divinsatff(1) <= (divinaasatff OR divinbbsatff) OR
                         (NOT(divinaazipff) AND divinbbzipff);
        divinzipff(1) <= divinaazipff;
        -- 0/0 or infinity/infinity is invalid OP, NAN out
        divinnanff(1) <= divinaananff OR divinbbnanff OR 
                        (divinaazipff AND divinbbzipff) OR
                        (divinaasatff AND divinbbsatff);      
        FOR k IN 2 TO midlatency LOOP
          divinsatff(k) <= divinsatff(k-1);
          divinzipff(k) <= divinzipff(k-1);
          divinnanff(k) <= divinnanff(k-1);
        END LOOP;
         
      END IF;
        
    END IF;
      
  END PROCESS;
       
  --**************************************************
  --***                                            ***
  --*** Output Section                             *** 
  --***                                            ***
  --**************************************************

  --********************************************************
  --*** internal format output, convert back to signed   ***
  --*** no need for fine normalization                   ***
  --********************************************************     
  goya: IF (xoutput = 1) GENERATE 
  
    -- output either "01XXXX..RR" (<1) or "1XXXX..RR" (>=1)
    -- if <1, SSSSSS1'manSSSSS
    -- if >1, SSSSS1'manSSSS
    goyb: FOR k IN 1 TO 4 GENERATE
      signeddivmannode(k) <= divinsignff(midlatency);
    END GENERATE;
    goyc: FOR k IN 1 TO 55 GENERATE
      signeddivmannode(k+4) <= divmannode(k) XOR divinsignff(midlatency);
    END GENERATE;
    goyd: FOR k IN 60 TO 64 GENERATE
      signeddivmannode(k) <= divinsignff(midlatency);
    END GENERATE;

    goye: IF ((roundconvert = 0) OR
              (roundconvert = 1 AND doublespeed = 0)) GENERATE

      goyf: IF (roundconvert = 0) GENERATE
        divroundnode <= signeddivmannode;
      END GENERATE;

      goyg: IF (roundconvert = 1) GENERATE
        divroundnode <= signeddivmannode + (zerovec(63 DOWNTO 1) & divinsignff(midlatency));
      END GENERATE;

      poxa: PROCESS (sysclk,reset)
      BEGIN
        
        IF (reset = '1') THEN
          
          FOR k IN 1 TO 64 LOOP
            divymanff(k) <= '0';
          END LOOP;
          FOR j IN 1 TO 13 LOOP
            divyexpff(j) <= '0';
          END LOOP;
          divysatbitff <= '0';
          divyzipbitff <= '0';
          divynanbitff <= '0';
      
        ELSIF (rising_edge(sysclk)) THEN
      
          IF (enable = '1') THEN
            
            divymanff <= divroundnode;
            divyexpff <= divinexpff(midlatency)(13 DOWNTO 1);
            divysatbitff <= divinsatff(midlatency);
            divyzipbitff <= divinzipff(midlatency);
            divynanbitff <= divinnanff(midlatency);
          
          END IF;        
              
        END IF;
        
      END PROCESS;

      cc(77 DOWNTO 14) <= divymanff;
      cc(13 DOWNTO 1) <= divyexpff;
      ccsat <= divysatbitff;
      cczip <= divyzipbitff;
      ccnan <= divynanbitff;

    END GENERATE;

    goyh: IF (roundconvert = 1 AND doublespeed = 1) GENERATE

      goyi: IF (synthesize = 0) GENERATE
        rndaddone: hcc_addpipeb 
        GENERIC MAP (width=>64,pipes=>2)
        PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
                  aa=>signeddivmannode,bb=>zerovec(64 DOWNTO 1),carryin=>divinsignff(midlatency),
                  cc=>divmanout);
      END GENERATE;

      goyj: IF (synthesize = 1) GENERATE
        rndaddtwo: hcc_addpipes 
        GENERIC MAP (width=>64,pipes=>2)
        PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
                  aa=>signeddivmannode,bb=>zerovec(64 DOWNTO 1),carryin=>divinsignff(midlatency),
                  cc=>divmanout);
      END GENERATE;

      poxb: PROCESS (sysclk,reset)
      BEGIN
        
        IF (reset = '1') THEN
          
          FOR j IN 1 TO 13 LOOP
            divyexpdelff(1)(j) <= '0';
            divyexpdelff(2)(j) <= '0';
          END LOOP;
          divysatdelff <= "00";
          divyzipdelff <= "00";
          divynandelff <= "00";
      
        ELSIF (rising_edge(sysclk)) THEN
      
          IF (enable = '1') THEN

            divyexpdelff(1)(13 DOWNTO 1) <= divinexpff(midlatency)(13 DOWNTO 1);
            divyexpdelff(2)(13 DOWNTO 1) <= divyexpdelff(1)(13 DOWNTO 1);
            divysatdelff(1) <= divinsatff(midlatency);
            divysatdelff(2) <= divysatdelff(1);
            divyzipdelff(1) <= divinzipff(midlatency);
            divyzipdelff(2) <= divyzipdelff(1);
            divynandelff(1) <= divinnanff(midlatency);
            divynandelff(2) <= divynandelff(1);

          END IF;        
              
        END IF;
        
      END PROCESS;

      cc(77 DOWNTO 14) <= divmanout;
      cc(13 DOWNTO 1) <= divyexpdelff(2)(13 DOWNTO 1);
      ccsat <= divysatdelff(2);
      cczip <= divyzipdelff(2);
      ccnan <= divynandelff(2);

    END GENERATE;
           
  END GENERATE;
  
  --**************************************************
  --*** if output to another multiplier or divider *** 
  --*** use output directly                        ***
  --**************************************************
  
  --*** NOTE: roundconvert options must still be added
  
  gofa: IF (divoutput = 1) GENERATE
  
    -- [55:1] output either "01XXXX..RR" (<1) or "1XXXX..RR" (>=1)
    normalize <= NOT(divmannode(55));
    gofb: FOR k IN 1 TO 53 GENERATE
      normmannode(k) <= (divmannode(k+1) AND normalize) OR
                        (divmannode(k+2) AND NOT(normalize));
    END GENERATE;    
        
    -- exp[54:1] always '1'manR
    poda: PROCESS (sysclk,reset)
    BEGIN
        
      IF (reset = '1') THEN
          
        FOR k IN 1 TO 54 LOOP
          divdivmanff(k) <= '0';
        END LOOP;
        FOR j IN 1 TO 13 LOOP
          divdivexpff(j) <= '0';
        END LOOP;
        divdivsatff <= '0';
        divdivzipff <= '0';
        divdivnanff <= '0';
        
      ELSIF (rising_edge(sysclk)) THEN
          
        divdivmanff <= divinsignff(midlatency) & normmannode;
         -- 20/05/09 add normalize adjustement
        divdivexpff <= divinexpff(midlatency)(13 DOWNTO 1) - (zerovec(12 DOWNTO 1) & normalize); 
        divdivsatff <= divinsatff(midlatency);
        divdivzipff <= divinzipff(midlatency);
        divdivnanff <= divinnanff(midlatency);
        
      END IF;
           
    END PROCESS;

    cc(67 DOWNTO 14) <= divdivmanff;
    cc(13 DOWNTO 1) <= divdivexpff;
    ccsat <= divdivsatff;
    cczip <= divdivzipff;
    ccnan <= divdivnanff;
  
  END GENERATE;
  
  --********************************************************
  --*** if output directly out of datapath, convert here ***
  --*** input to multiplier always "01XXX" format, so    ***
  --*** just 1 bit normalization required                ***
  --********************************************************
  goea: IF (ieeeoutput = 1) GENERATE -- ieee754 out of datapath, do conversion
  
    -- output either "01XXXX..RR" (<2) or "1XXXX..RR" (>=2), need to make output
    -- 01XXXX
    normalize <= NOT(divmannode(55));
    goeb: FOR k IN 1 TO 54 GENERATE -- format "01"[52..1]R
      normalnode(k) <= (divmannode(k+1) AND NOT(normalize)) OR 
                       (divmannode(k) AND normalize); 
    END GENERATE;
    
    poea: PROCESS (sysclk,reset)
    BEGIN
    
      IF (reset = '1') THEN
          
        normsignff <= '0';
        normsatff <= '0';
        normzipff <= '0';
        normnanff <= '0';
        FOR k IN 1 TO 54 LOOP
          normalff(k) <= '0';
        END LOOP;
        FOR k IN 1 TO 13 LOOP
          normalexpff(k) <= '0';
        END LOOP;
        
      ELSIF (rising_edge(sysclk)) THEN
        
        IF (enable = '1') THEN
            
          normsignff <= divinsignff(midlatency);
          normsatff <= divinsatff(midlatency);
          normzipff <= divinzipff(midlatency);
          normnanff <= divinnanff(midlatency);
          
          normalff <= normalnode;
          
          normalexpff <= divinexpff(midlatency)(13 DOWNTO 1) -
                         (zerovec(12 DOWNTO 1) & normalize);
                         
        END IF;      
              
      END IF;
      
    END PROCESS;

    goec: IF (roundconvert = 0) GENERATE

      norndout: hcc_divnornd
      PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
                signin=>normsignff,
                exponentin=>normalexpff,
                mantissain=>normalff(53 DOWNTO 1),
                satin=>normsatff,
                zipin=>normzipff,
                nanin=>normnanff,

                signout=>cc(64),exponentout=>cc(63 DOWNTO 53),mantissaout=>cc(52 DOWNTO 1));
                
      -- dummy only
      ccsat <= '0';
      cczip <= '0';
      ccnan <= '0';    
            
    END GENERATE;
    
    goed: IF ((roundconvert = 1) AND (doublespeed = 0)) GENERATE

      rndout: hcc_divrnd
      PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
                signin=>normsignff,
                exponentin=>normalexpff,
                mantissain=>normalff(53 DOWNTO 1),
                satin=>normsatff,
                zipin=>normzipff,
                nanin=>normnanff,

                signout=>cc(64),exponentout=>cc(63 DOWNTO 53),mantissaout=>cc(52 DOWNTO 1));
                
      -- dummy only
      ccsat <= '0';
      cczip <= '0';
      ccnan <= '0';    
            
    END GENERATE;
    
    goee: IF ((roundconvert = 1) AND (doublespeed = 1)) GENERATE

      rndpipout: hcc_divrndpipe
      GENERIC MAP (synthesize=>synthesize)
      PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
                signin=>normsignff,
                exponentin=>normalexpff,
                mantissain=>normalff(53 DOWNTO 1),
                satin=>normsatff,
                zipin=>normzipff,
                nanin=>normnanff,

                signout=>cc(64),exponentout=>cc(63 DOWNTO 53),mantissaout=>cc(52 DOWNTO 1));
                
      -- dummy only
      ccsat <= '0';
      cczip <= '0';    
      ccnan <= '0';
            
    END GENERATE;
    
  END GENERATE;

END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   ALTERA FLOATING POINT DATAPATH COMPILER   ***
--***                                             ***
--***   HCC_DIVNORND.VHD                          ***
--***                                             ***
--***   Function: Output Stage, No Rounding       ***
--***                                             ***
--***                                             ***
--***   24/12/07 ML                               ***
--***                                             ***
--***   (c) 2007 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***   22/04/09 - added NAN support, IEEE NAN    ***
--***   output                                    ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes: Latency = 1                          ***
--***************************************************

ENTITY hcc_divnornd IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (13 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (53 DOWNTO 1); -- includes roundbit
      satin, zipin, nanin : IN STD_LOGIC;

		signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1)
		);
END hcc_divnornd;

ARCHITECTURE rtl OF hcc_divnornd IS

  type exponentfftype IS ARRAY (2 DOWNTO 1) OF STD_LOGIC_VECTOR (13 DOWNTO 1);
  
  signal zerovec : STD_LOGIC_VECTOR (51 DOWNTO 1);
  signal signff : STD_LOGIC;
  signal nanff : STD_LOGIC;
  signal dividebyzeroff : STD_LOGIC;  
  signal mantissaff : STD_LOGIC_VECTOR (52 DOWNTO 1);
  signal exponentff : STD_LOGIC_VECTOR (11 DOWNTO 1);
  
  signal infinitygen : STD_LOGIC_VECTOR (12 DOWNTO 1);
  signal zerogen : STD_LOGIC_VECTOR (12 DOWNTO 1);  
  signal setmanzero, setmanmax : STD_LOGIC;
  signal setexpzero, setexpmax : STD_LOGIC;

BEGIN
    
  gzv: FOR k IN 1 TO 51 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  pra: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN
        
      signff <= '0';
      FOR k IN 1 TO 52 LOOP
        mantissaff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 11 LOOP
        exponentff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF(enable = '1') THEN 
      
        signff <= signin;
  
        FOR k IN 1 TO 52 LOOP
          mantissaff(k) <= (mantissain(k+1) AND NOT(setmanzero)) OR setmanmax;
        END LOOP;
               
        FOR k IN 1 TO 11 LOOP
          exponentff(k) <= (exponentin(k) AND NOT(setexpzero)) OR setexpmax;
        END LOOP;
      
      END IF;
             
    END IF;
      
  END PROCESS;
                                                  
--**********************************
--*** CHECK GENERATED CONDITIONS ***   
--**********************************

  -- '1' when true for all cases
  
  -- infinity if exponent >= 255
  infinitygen(1) <= exponentin(1);
  gia: FOR k IN 2 TO 11 GENERATE
    infinitygen(k) <= infinitygen(k-1) AND exponentin(k);
  END GENERATE;
  -- 12/05/09 - make sure exponentin = -1 doesnt make infinity
  infinitygen(12) <= (infinitygen(11) AND NOT(exponentin(12)) AND NOT(exponentin(13))) OR 
                     satin OR (exponentin(12) AND NOT(exponentin(13))); -- '1' if infinity
                         
  -- zero if exponent <= 0
  zerogen(1) <= exponentin(1);
  gza: FOR k IN 2 TO 11 GENERATE
    zerogen(k) <= zerogen(k-1) OR exponentin(k);
  END GENERATE;
  zerogen(12) <= NOT(zerogen(11)) OR zipin OR exponentin(13); -- '1' if zero
                    
  -- set mantissa to 0 when infinity or zero condition
  setmanzero <= infinitygen(12) OR zerogen(12);
  setmanmax <= nanin;
  -- set exponent to 0 when zero condition 
  setexpzero <= zerogen(12);
  -- set exponent to "11..11" infinity
  setexpmax <= infinitygen(12) OR nanin;
                             
--***************
--*** OUTPUTS ***
--***************

  signout <= signff;   
  mantissaout <= mantissaff;
  exponentout <= exponentff; 

END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   ALTERA FLOATING POINT DATAPATH COMPILER   ***
--***                                             ***
--***   HCC_DIVRND.VHD                            ***
--***                                             ***
--***   Function: Output Stage, Rounding          ***
--***                                             ***
--***   24/12/07 ML                               ***
--***                                             ***
--***   (c) 2007 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***   22/04/09 - added NAN support, IEEE NAN    ***
--***   output                                    ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes: Latency = 2                          ***
--***************************************************

ENTITY hcc_divrnd IS 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (13 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (53 DOWNTO 1); -- includes roundbit
      satin, zipin, nanin : IN STD_LOGIC;

		signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1)
		);
END hcc_divrnd;

ARCHITECTURE rtl OF hcc_divrnd IS

  signal zerovec : STD_LOGIC_VECTOR (51 DOWNTO 1);
  signal signff : STD_LOGIC_VECTOR (2 DOWNTO 1);
  signal satinff, zipinff, naninff : STD_LOGIC;
  signal overflowbitff : STD_LOGIC; 
  signal roundmantissaff, mantissaff : STD_LOGIC_VECTOR (52 DOWNTO 1);
  signal exponentnode : STD_LOGIC_VECTOR (13 DOWNTO 1);
  signal exponentoneff : STD_LOGIC_VECTOR (13 DOWNTO 1);
  signal exponenttwoff : STD_LOGIC_VECTOR (11 DOWNTO 1);
  
  signal manoverflow : STD_LOGIC_VECTOR (53 DOWNTO 1);
  signal infinitygen : STD_LOGIC_VECTOR (12 DOWNTO 1);
  signal zerogen : STD_LOGIC_VECTOR (12 DOWNTO 1);  
  signal setmanzero, setmanmax : STD_LOGIC;
  signal setexpzero, setexpmax : STD_LOGIC;

BEGIN
    
  gzv: FOR k IN 1 TO 51 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  pra: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN
        
      signff <= "00";
      satinff <= '0';
      zipinff <= '0';
      naninff <= '0';
      overflowbitff <= '0';
      FOR k IN 1 TO 52 LOOP
        roundmantissaff(k) <= '0';
        mantissaff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 13 LOOP
        exponentoneff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 11 LOOP
        exponenttwoff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF(enable = '1') THEN 
      
        signff(1) <= signin;
        signff(2) <= signff(1);
        satinff <= satin;
        zipinff <= zipin;
        naninff <= nanin;
        
        overflowbitff <= manoverflow(53);
        
        roundmantissaff <= mantissain(53 DOWNTO 2) + (zerovec & mantissain(1));

        FOR k IN 1 TO 52 LOOP
          mantissaff(k) <= (roundmantissaff(k) AND NOT(setmanzero)) OR setmanmax;
        END LOOP;
        
        exponentoneff(13 DOWNTO 1) <= exponentin(13 DOWNTO 1);                 
        FOR k IN 1 TO 11 LOOP
          exponenttwoff(k) <= (exponentnode(k) AND NOT(setexpzero)) OR setexpmax;
        END LOOP;
      
      END IF;
             
    END IF;
      
  END PROCESS;
  
  exponentnode <= exponentoneff(13 DOWNTO 1) + 
                 (zerovec(12 DOWNTO 1) & overflowbitff);

--*********************************
--*** PREDICT MANTISSA OVERFLOW ***   
--*********************************
     
  manoverflow(1) <= mantissain(1);
  gmoa: FOR k IN 2 TO 53 GENERATE
    manoverflow(k) <= manoverflow(k-1) AND mantissain(k);
  END GENERATE; 
                                                                 
--**********************************
--*** CHECK GENERATED CONDITIONS ***   
--**********************************

  -- '1' when true for all cases
  
  -- infinity if exponent >= 255
  infinitygen(1) <= exponentnode(1);
  gia: FOR k IN 2 TO 11 GENERATE
    infinitygen(k) <= infinitygen(k-1) AND exponentnode(k);
  END GENERATE;
  -- 12/05/09 - make sure exponentnode = -1 doesnt make infinity
  infinitygen(12) <= (infinitygen(11) AND NOT(exponentnode(12)) AND NOT(exponentnode(13))) OR 
                      satinff OR (exponentnode(12) AND NOT(exponentnode(13))); -- '1' if infinity
                         
  -- zero if exponent <= 0
  zerogen(1) <= exponentnode(1);
  gza: FOR k IN 2 TO 11 GENERATE
    zerogen(k) <= zerogen(k-1) OR exponentnode(k);
  END GENERATE;
  zerogen(12) <= NOT(zerogen(11)) OR zipinff OR exponentnode(13); -- '1' if zero
                    
  -- set mantissa to 0 when infinity or zero condition
  setmanzero <= infinitygen(12) OR zerogen(12);
  setmanmax <= naninff;
  -- set exponent to 0 when zero condition 
  setexpzero <= zerogen(12);
  -- set exponent to "11..11" infinity
  setexpmax <= infinitygen(12) OR naninff;
                        
--***************
--*** OUTPUTS ***
--***************

  signout <= signff(2);   
  mantissaout <= mantissaff;
  exponentout <= exponenttwoff;

END rtl;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_arith.all; 

--***************************************************
--***                                             ***
--***   ALTERA FLOATING POINT DATAPATH COMPILER   ***
--***                                             ***
--***   HCC_DIVRNDPIPE.VHD                        ***
--***                                             ***
--***   Function: Output Stage, Pipelined Round   ***
--***                                             ***
--***   24/12/07 ML                               ***
--***                                             ***
--***   (c) 2007 Altera Corporation               ***
--***                                             ***
--***   Change History                            ***
--***                                             ***
--***   22/04/09 - added NAN support, IEEE NAN    ***
--***   output                                    ***
--***                                             ***
--***                                             ***
--***************************************************

--***************************************************
--*** Notes: Latency = 3                          ***
--***************************************************

ENTITY hcc_divrndpipe IS 
GENERIC (synthesize : integer := 1); 
PORT (
      sysclk : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      enable : IN STD_LOGIC;
      signin : IN STD_LOGIC;
      exponentin : IN STD_LOGIC_VECTOR (13 DOWNTO 1);
      mantissain : IN STD_LOGIC_VECTOR (53 DOWNTO 1); -- includes roundbit
      satin, zipin, nanin : IN STD_LOGIC;

		signout : OUT STD_LOGIC;
      exponentout : OUT STD_LOGIC_VECTOR (11 DOWNTO 1);
      mantissaout : OUT STD_LOGIC_VECTOR (52 DOWNTO 1)
		);
END hcc_divrndpipe;

ARCHITECTURE rtl OF hcc_divrndpipe IS

  signal zerovec : STD_LOGIC_VECTOR (53 DOWNTO 1);
  signal signff : STD_LOGIC_VECTOR (3 DOWNTO 1);
  signal satinff, zipinff, naninff : STD_LOGIC_VECTOR (2 DOWNTO 1);  
  signal roundmantissanode : STD_LOGIC_VECTOR (52 DOWNTO 1);
  signal mantissaff : STD_LOGIC_VECTOR (52 DOWNTO 1);
  signal exponentoneff, exponenttwoff : STD_LOGIC_VECTOR (13 DOWNTO 1);
  signal exponentff : STD_LOGIC_VECTOR (11 DOWNTO 1);
  
  signal manoverflow : STD_LOGIC_VECTOR (53 DOWNTO 1);
  signal manoverflowff : STD_LOGIC;
  signal infinitygen : STD_LOGIC_VECTOR (12 DOWNTO 1);
  signal zerogen : STD_LOGIC_VECTOR (12 DOWNTO 1);  
  signal setmanzero, setmanmax : STD_LOGIC;
  signal setexpzero, setexpmax : STD_LOGIC;

  component hcc_addpipeb
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
        carryin : IN STD_LOGIC;
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
  end component;

  component hcc_addpipes
  GENERIC (
           width : positive := 64;
           pipes : positive := 1
          );
  PORT (
        sysclk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        enable : IN STD_LOGIC;
        aa, bb : IN STD_LOGIC_VECTOR (width DOWNTO 1); 
        carryin : IN STD_LOGIC;
      
        cc : OUT STD_LOGIC_VECTOR (width DOWNTO 1)
       );
  end component;
  
BEGIN
    
  gzv: FOR k IN 1 TO 53 GENERATE
    zerovec(k) <= '0';
  END GENERATE;
  
  pra: PROCESS (sysclk,reset)
  BEGIN
      
    IF (reset = '1') THEN
        
      signff <= "000";
      satinff <= "00";
      zipinff <= "00";
      naninff <= "00";
      manoverflowff <= '0';
      FOR k IN 1 TO 52 LOOP
        mantissaff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 13 LOOP
        exponentoneff(k) <= '0';
        exponenttwoff(k) <= '0';
      END LOOP;
      FOR k IN 1 TO 11 LOOP
        exponentff(k) <= '0';
      END LOOP;
      
    ELSIF (rising_edge(sysclk)) THEN
    
      IF(enable = '1') THEN 
      
        signff(1) <= signin;
        signff(2) <= signff(1);
        signff(3) <= signff(2);
        
        satinff(1) <= satin;
        satinff(2) <= satinff(1);
        zipinff(1) <= zipin;
        zipinff(2) <= zipinff(1);
        naninff(1) <= nanin;
        naninff(2) <= naninff(1);
         
        FOR k IN 1 TO 52 LOOP
          mantissaff(k) <= (roundmantissanode(k) AND NOT(setmanzero)) OR setmanmax;
        END LOOP;
        
        exponentoneff(13 DOWNTO 1) <= exponentin;
        exponenttwoff(13 DOWNTO 1) <= exponentoneff(13 DOWNTO 1) + 
                                      (zerovec(12 DOWNTO 1) & manoverflowff);                 
        FOR k IN 1 TO 11 LOOP
          exponentff(k) <= (exponenttwoff(k) AND NOT(setexpzero)) OR setexpmax;
        END LOOP;
      
      END IF;
             
    END IF;
      
  END PROCESS;

  gaa: IF (synthesize = 0) GENERATE
    addb: hcc_addpipeb
    GENERIC MAP (width=>52,pipes=>2)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>mantissain(53 DOWNTO 2),bb=>zerovec(52 DOWNTO 1),
              carryin=>mantissain(1),
              cc=>roundmantissanode);
  END GENERATE;
         
  gab: IF (synthesize = 1) GENERATE
    addb: hcc_addpipes
    GENERIC MAP (width=>52,pipes=>2)
    PORT MAP (sysclk=>sysclk,reset=>reset,enable=>enable,
              aa=>mantissain(53 DOWNTO 2),bb=>zerovec(52 DOWNTO 1),
              carryin=>mantissain(1),
              cc=>roundmantissanode);
  END GENERATE;
  
--*********************************
--*** PREDICT MANTISSA OVERFLOW ***   
--*********************************
     
  manoverflow(1) <= mantissain(1);
  gmoa: FOR k IN 2 TO 53 GENERATE
    manoverflow(k) <= manoverflow(k-1) AND mantissain(k);
  END GENERATE;                                           
    
--**********************************
--*** CHECK GENERATED CONDITIONS ***   
--**********************************

  -- infinity if exponent >= 255
  infinitygen(1) <= exponenttwoff(1);
  gia: FOR k IN 2 TO 11 GENERATE
    infinitygen(k) <= infinitygen(k-1) AND exponenttwoff(k);
  END GENERATE;
  -- 12/05/09 - make sure exponent = -1 doesnt make infinity
  infinitygen(12) <= (infinitygen(11) AND NOT(exponenttwoff(12)) AND NOT(exponenttwoff(13))) OR 
                      satinff(2) OR (exponenttwoff(12) AND NOT(exponenttwoff(13))); -- '1' if infinity
                         
  -- zero if exponent <= 0
  zerogen(1) <= exponenttwoff(1);
  gza: FOR k IN 2 TO 11 GENERATE
    zerogen(k) <= zerogen(k-1) OR exponenttwoff(k);
  END GENERATE;
  zerogen(12) <= NOT(zerogen(11)) OR zipinff(2) OR exponenttwoff(13); -- '1' if zero
                    
  -- set mantissa to 0 when infinity or zero condition
  setmanzero <= infinitygen(12) OR zerogen(12);
  setmanmax <= naninff(2);
  -- set exponent to 0 when zero condition 
  setexpzero <= zerogen(12);
  -- set exponent to "11..11" infinity
  setexpmax <= infinitygen(12) OR naninff(2);
                             
--***************
--*** OUTPUTS ***
--***************

  signout <= signff(3);   
  mantissaout <= mantissaff;
  exponentout <= exponentff; 

END rtl;

