
library ieee;
use ieee.std_logic_1164.all;

entity DECODER is
generic(
 WIDTH : integer := 32);
port(	I:	in std_logic_vector(WIDTH-1 downto 0);
	    O:	out std_logic_vector(WIDTH-1 downto 0)
);
end DECODER;

architecture when_else of DECODER is
begin

    O <= 	"11111111111111111111111111111110" when I = "00000000000000000000000000000000" else
		    "11111111111111111111111111111101" when I = "00000000000000000000000000000001" else
		    "11111111111111111111111111111011" when I = "00000000000000000000000000000010" else
		    "11111111111111111111111111110111" when I = "00000000000000000000000000000011" else
		    "11111111111111111111111111101111" when I = "00000000000000000000000000000100" else
            "11111111111111111111111111011111" when I = "00000000000000000000000000000101" else
            "11111111111111111111111110111111" when I = "00000000000000000000000000000110" else
            "11111111111111111111111101111111" when I = "00000000000000000000000000000111" else
            "11111111111111111111111011111111" when I = "00000000000000000000000000001000" else
            "11111111111111111111110111111111" when I = "00000000000000000000000000001001" else
            "11111111111111111111101111111111" when I = "00000000000000000000000000001010" else
            "11111111111111111111011111111111" when I = "00000000000000000000000000001011" else
            "11111111111111111110111111111111" when I = "00000000000000000000000000001100" else
            "11111111111111111101111111111111" when I = "00000000000000000000000000001101" else
            "11111111111111111011111111111111" when I = "00000000000000000000000000001110" else
            "11111111111111110111111111111111" when I = "00000000000000000000000000001111" else
            "11111111111111101111111111111111" when I = "00000000000000000000000000010000" else
            "11111111111111011111111111111111" when I = "00000000000000000000000000010001" else
            "11111111111110111111111111111111" when I = "00000000000000000000000000010010" else
            "11111111111101111111111111111111" when I = "00000000000000000000000000010011" else
            "11111111111011111111111111111111" when I = "00000000000000000000000000010100" else
            "11111111110111111111111111111111" when I = "00000000000000000000000000010101" else
            "11111111101111111111111111111111" when I = "00000000000000000000000000010110" else
            "11111111011111111111111111111111" when I = "00000000000000000000000000010111" else
            "11111110111111111111111111111111" when I = "00000000000000000000000000011000" else
            "11111101111111111111111111111111" when I = "00000000000000000000000000011001" else
            "11111011111111111111111111111111" when I = "00000000000000000000000000011010" else
            "11110111111111111111111111111111" when I = "00000000000000000000000000011011" else
            "11101111111111111111111111111111" when I = "00000000000000000000000000011100" else
            "11011111111111111111111111111111" when I = "00000000000000000000000000011101" else
            "10111111111111111111111111111111" when I = "00000000000000000000000000011110" else
            "01111111111111111111111111111111" when I = "00000000000000000000000000011111" else
		    "11111111111111111111111111111111";

end when_else;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity decoder_top_vhd is
generic(
 WIDTH : integer := 32);
port(
    data_in: in std_logic_vector(WIDTH-1 downto 0);
    clk: in std_logic;
    rst: in std_logic;
    data_out: out std_logic_vector(WIDTH-1 downto 0));
end decoder_top_vhd;

architecture rtl of decoder_top_vhd is
    signal data_out_tmp: std_logic_vector(WIDTH-1 downto 0);
    
begin
    process(clk,rst)
    begin
        if rst = '0' then
            data_out<=(data_out_tmp'range=>'0');
        elsif (clk'event and clk='1') then
            data_out<=data_out_tmp;
        end if;   
    end process;
    
DEC : entity work.DECODER(when_else)
    generic map (
    WIDTH => WIDTH)
    port map(
    I => data_in(WIDTH-1 downto 0),
    O  => data_out_tmp(WIDTH-1 downto 0)
);
    
end rtl;