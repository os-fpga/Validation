// `include "encoder.v"
// `include "invertion.v"
// `include "large_mux.v"
// `include "register.v"
module design21_20_30_top #(parameter WIDTH=32,CHANNEL=20) (clk, rst, in, out);

	localparam OUT_BUS=CHANNEL*WIDTH;
	input clk,rst;
	input [WIDTH-1:0] in;
	output [WIDTH-1:0] out;

	reg [WIDTH-1:0] d_in0;
	reg [WIDTH-1:0] d_in1;
	reg [WIDTH-1:0] d_in2;
	reg [WIDTH-1:0] d_in3;
	reg [WIDTH-1:0] d_in4;
	reg [WIDTH-1:0] d_in5;
	reg [WIDTH-1:0] d_in6;
	reg [WIDTH-1:0] d_in7;
	reg [WIDTH-1:0] d_in8;
	reg [WIDTH-1:0] d_in9;
	reg [WIDTH-1:0] d_in10;
	reg [WIDTH-1:0] d_in11;
	reg [WIDTH-1:0] d_in12;
	reg [WIDTH-1:0] d_in13;
	reg [WIDTH-1:0] d_in14;
	reg [WIDTH-1:0] d_in15;
	reg [WIDTH-1:0] d_in16;
	reg [WIDTH-1:0] d_in17;
	reg [WIDTH-1:0] d_in18;
	reg [WIDTH-1:0] d_in19;
	wire [WIDTH-1:0] d_out0;
	wire [WIDTH-1:0] d_out1;
	wire [WIDTH-1:0] d_out2;
	wire [WIDTH-1:0] d_out3;
	wire [WIDTH-1:0] d_out4;
	wire [WIDTH-1:0] d_out5;
	wire [WIDTH-1:0] d_out6;
	wire [WIDTH-1:0] d_out7;
	wire [WIDTH-1:0] d_out8;
	wire [WIDTH-1:0] d_out9;
	wire [WIDTH-1:0] d_out10;
	wire [WIDTH-1:0] d_out11;
	wire [WIDTH-1:0] d_out12;
	wire [WIDTH-1:0] d_out13;
	wire [WIDTH-1:0] d_out14;
	wire [WIDTH-1:0] d_out15;
	wire [WIDTH-1:0] d_out16;
	wire [WIDTH-1:0] d_out17;
	wire [WIDTH-1:0] d_out18;
	wire [WIDTH-1:0] d_out19;

	reg [OUT_BUS-1:0] tmp;

	always @ (posedge clk or posedge rst) begin
		if (rst)
			tmp <= 0;
		else
			tmp <= {tmp[OUT_BUS-(WIDTH-1):0],in};
	end

	always @ (posedge clk) begin
		d_in0 <= tmp[WIDTH-1:0];
		d_in1 <= tmp[(WIDTH*2)-1:WIDTH*1];
		d_in2 <= tmp[(WIDTH*3)-1:WIDTH*2];
		d_in3 <= tmp[(WIDTH*4)-1:WIDTH*3];
		d_in4 <= tmp[(WIDTH*5)-1:WIDTH*4];
		d_in5 <= tmp[(WIDTH*6)-1:WIDTH*5];
		d_in6 <= tmp[(WIDTH*7)-1:WIDTH*6];
		d_in7 <= tmp[(WIDTH*8)-1:WIDTH*7];
		d_in8 <= tmp[(WIDTH*9)-1:WIDTH*8];
		d_in9 <= tmp[(WIDTH*10)-1:WIDTH*9];
		d_in10 <= tmp[(WIDTH*11)-1:WIDTH*10];
		d_in11 <= tmp[(WIDTH*12)-1:WIDTH*11];
		d_in12 <= tmp[(WIDTH*13)-1:WIDTH*12];
		d_in13 <= tmp[(WIDTH*14)-1:WIDTH*13];
		d_in14 <= tmp[(WIDTH*15)-1:WIDTH*14];
		d_in15 <= tmp[(WIDTH*16)-1:WIDTH*15];
		d_in16 <= tmp[(WIDTH*17)-1:WIDTH*16];
		d_in17 <= tmp[(WIDTH*18)-1:WIDTH*17];
		d_in18 <= tmp[(WIDTH*19)-1:WIDTH*18];
		d_in19 <= tmp[(WIDTH*20)-1:WIDTH*19];
	end

	design21_20_30 #(.WIDTH(WIDTH)) design21_20_30_inst(.d_in0(d_in0),.d_in1(d_in1),.d_in2(d_in2),.d_in3(d_in3),.d_in4(d_in4),.d_in5(d_in5),.d_in6(d_in6),.d_in7(d_in7),.d_in8(d_in8),.d_in9(d_in9),.d_in10(d_in10),.d_in11(d_in11),.d_in12(d_in12),.d_in13(d_in13),.d_in14(d_in14),.d_in15(d_in15),.d_in16(d_in16),.d_in17(d_in17),.d_in18(d_in18),.d_in19(d_in19),.d_out0(d_out0),.d_out1(d_out1),.d_out2(d_out2),.d_out3(d_out3),.d_out4(d_out4),.d_out5(d_out5),.d_out6(d_out6),.d_out7(d_out7),.d_out8(d_out8),.d_out9(d_out9),.d_out10(d_out10),.d_out11(d_out11),.d_out12(d_out12),.d_out13(d_out13),.d_out14(d_out14),.d_out15(d_out15),.d_out16(d_out16),.d_out17(d_out17),.d_out18(d_out18),.d_out19(d_out19),.clk(clk),.rst(rst));

	assign out = d_out0^d_out1^d_out2^d_out3^d_out4^d_out5^d_out6^d_out7^d_out8^d_out9^d_out10^d_out11^d_out12^d_out13^d_out14^d_out15^d_out16^d_out17^d_out18^d_out19;

endmodule

module design21_20_30 #(parameter WIDTH=32) (d_in0, d_in1, d_in2, d_in3, d_in4, d_in5, d_in6, d_in7, d_in8, d_in9, d_in10, d_in11, d_in12, d_in13, d_in14, d_in15, d_in16, d_in17, d_in18, d_in19, d_out0, d_out1, d_out2, d_out3, d_out4, d_out5, d_out6, d_out7, d_out8, d_out9, d_out10, d_out11, d_out12, d_out13, d_out14, d_out15, d_out16, d_out17, d_out18, d_out19, clk, rst);
	input clk;
	input rst;
	input [WIDTH-1:0] d_in0; 
	input [WIDTH-1:0] d_in1; 
	input [WIDTH-1:0] d_in2; 
	input [WIDTH-1:0] d_in3; 
	input [WIDTH-1:0] d_in4; 
	input [WIDTH-1:0] d_in5; 
	input [WIDTH-1:0] d_in6; 
	input [WIDTH-1:0] d_in7; 
	input [WIDTH-1:0] d_in8; 
	input [WIDTH-1:0] d_in9; 
	input [WIDTH-1:0] d_in10; 
	input [WIDTH-1:0] d_in11; 
	input [WIDTH-1:0] d_in12; 
	input [WIDTH-1:0] d_in13; 
	input [WIDTH-1:0] d_in14; 
	input [WIDTH-1:0] d_in15; 
	input [WIDTH-1:0] d_in16; 
	input [WIDTH-1:0] d_in17; 
	input [WIDTH-1:0] d_in18; 
	input [WIDTH-1:0] d_in19; 
	output [WIDTH-1:0] d_out0; 
	output [WIDTH-1:0] d_out1; 
	output [WIDTH-1:0] d_out2; 
	output [WIDTH-1:0] d_out3; 
	output [WIDTH-1:0] d_out4; 
	output [WIDTH-1:0] d_out5; 
	output [WIDTH-1:0] d_out6; 
	output [WIDTH-1:0] d_out7; 
	output [WIDTH-1:0] d_out8; 
	output [WIDTH-1:0] d_out9; 
	output [WIDTH-1:0] d_out10; 
	output [WIDTH-1:0] d_out11; 
	output [WIDTH-1:0] d_out12; 
	output [WIDTH-1:0] d_out13; 
	output [WIDTH-1:0] d_out14; 
	output [WIDTH-1:0] d_out15; 
	output [WIDTH-1:0] d_out16; 
	output [WIDTH-1:0] d_out17; 
	output [WIDTH-1:0] d_out18; 
	output [WIDTH-1:0] d_out19; 

	wire [WIDTH-1:0] wire_d0_0;
	wire [WIDTH-1:0] wire_d0_1;
	wire [WIDTH-1:0] wire_d0_2;
	wire [WIDTH-1:0] wire_d0_3;
	wire [WIDTH-1:0] wire_d0_4;
	wire [WIDTH-1:0] wire_d0_5;
	wire [WIDTH-1:0] wire_d0_6;
	wire [WIDTH-1:0] wire_d0_7;
	wire [WIDTH-1:0] wire_d0_8;
	wire [WIDTH-1:0] wire_d0_9;
	wire [WIDTH-1:0] wire_d0_10;
	wire [WIDTH-1:0] wire_d0_11;
	wire [WIDTH-1:0] wire_d0_12;
	wire [WIDTH-1:0] wire_d0_13;
	wire [WIDTH-1:0] wire_d0_14;
	wire [WIDTH-1:0] wire_d0_15;
	wire [WIDTH-1:0] wire_d0_16;
	wire [WIDTH-1:0] wire_d0_17;
	wire [WIDTH-1:0] wire_d0_18;
	wire [WIDTH-1:0] wire_d0_19;
	wire [WIDTH-1:0] wire_d0_20;
	wire [WIDTH-1:0] wire_d0_21;
	wire [WIDTH-1:0] wire_d0_22;
	wire [WIDTH-1:0] wire_d0_23;
	wire [WIDTH-1:0] wire_d0_24;
	wire [WIDTH-1:0] wire_d0_25;
	wire [WIDTH-1:0] wire_d0_26;
	wire [WIDTH-1:0] wire_d0_27;
	wire [WIDTH-1:0] wire_d0_28;
	wire [WIDTH-1:0] wire_d1_0;
	wire [WIDTH-1:0] wire_d1_1;
	wire [WIDTH-1:0] wire_d1_2;
	wire [WIDTH-1:0] wire_d1_3;
	wire [WIDTH-1:0] wire_d1_4;
	wire [WIDTH-1:0] wire_d1_5;
	wire [WIDTH-1:0] wire_d1_6;
	wire [WIDTH-1:0] wire_d1_7;
	wire [WIDTH-1:0] wire_d1_8;
	wire [WIDTH-1:0] wire_d1_9;
	wire [WIDTH-1:0] wire_d1_10;
	wire [WIDTH-1:0] wire_d1_11;
	wire [WIDTH-1:0] wire_d1_12;
	wire [WIDTH-1:0] wire_d1_13;
	wire [WIDTH-1:0] wire_d1_14;
	wire [WIDTH-1:0] wire_d1_15;
	wire [WIDTH-1:0] wire_d1_16;
	wire [WIDTH-1:0] wire_d1_17;
	wire [WIDTH-1:0] wire_d1_18;
	wire [WIDTH-1:0] wire_d1_19;
	wire [WIDTH-1:0] wire_d1_20;
	wire [WIDTH-1:0] wire_d1_21;
	wire [WIDTH-1:0] wire_d1_22;
	wire [WIDTH-1:0] wire_d1_23;
	wire [WIDTH-1:0] wire_d1_24;
	wire [WIDTH-1:0] wire_d1_25;
	wire [WIDTH-1:0] wire_d1_26;
	wire [WIDTH-1:0] wire_d1_27;
	wire [WIDTH-1:0] wire_d1_28;
	wire [WIDTH-1:0] wire_d2_0;
	wire [WIDTH-1:0] wire_d2_1;
	wire [WIDTH-1:0] wire_d2_2;
	wire [WIDTH-1:0] wire_d2_3;
	wire [WIDTH-1:0] wire_d2_4;
	wire [WIDTH-1:0] wire_d2_5;
	wire [WIDTH-1:0] wire_d2_6;
	wire [WIDTH-1:0] wire_d2_7;
	wire [WIDTH-1:0] wire_d2_8;
	wire [WIDTH-1:0] wire_d2_9;
	wire [WIDTH-1:0] wire_d2_10;
	wire [WIDTH-1:0] wire_d2_11;
	wire [WIDTH-1:0] wire_d2_12;
	wire [WIDTH-1:0] wire_d2_13;
	wire [WIDTH-1:0] wire_d2_14;
	wire [WIDTH-1:0] wire_d2_15;
	wire [WIDTH-1:0] wire_d2_16;
	wire [WIDTH-1:0] wire_d2_17;
	wire [WIDTH-1:0] wire_d2_18;
	wire [WIDTH-1:0] wire_d2_19;
	wire [WIDTH-1:0] wire_d2_20;
	wire [WIDTH-1:0] wire_d2_21;
	wire [WIDTH-1:0] wire_d2_22;
	wire [WIDTH-1:0] wire_d2_23;
	wire [WIDTH-1:0] wire_d2_24;
	wire [WIDTH-1:0] wire_d2_25;
	wire [WIDTH-1:0] wire_d2_26;
	wire [WIDTH-1:0] wire_d2_27;
	wire [WIDTH-1:0] wire_d2_28;
	wire [WIDTH-1:0] wire_d3_0;
	wire [WIDTH-1:0] wire_d3_1;
	wire [WIDTH-1:0] wire_d3_2;
	wire [WIDTH-1:0] wire_d3_3;
	wire [WIDTH-1:0] wire_d3_4;
	wire [WIDTH-1:0] wire_d3_5;
	wire [WIDTH-1:0] wire_d3_6;
	wire [WIDTH-1:0] wire_d3_7;
	wire [WIDTH-1:0] wire_d3_8;
	wire [WIDTH-1:0] wire_d3_9;
	wire [WIDTH-1:0] wire_d3_10;
	wire [WIDTH-1:0] wire_d3_11;
	wire [WIDTH-1:0] wire_d3_12;
	wire [WIDTH-1:0] wire_d3_13;
	wire [WIDTH-1:0] wire_d3_14;
	wire [WIDTH-1:0] wire_d3_15;
	wire [WIDTH-1:0] wire_d3_16;
	wire [WIDTH-1:0] wire_d3_17;
	wire [WIDTH-1:0] wire_d3_18;
	wire [WIDTH-1:0] wire_d3_19;
	wire [WIDTH-1:0] wire_d3_20;
	wire [WIDTH-1:0] wire_d3_21;
	wire [WIDTH-1:0] wire_d3_22;
	wire [WIDTH-1:0] wire_d3_23;
	wire [WIDTH-1:0] wire_d3_24;
	wire [WIDTH-1:0] wire_d3_25;
	wire [WIDTH-1:0] wire_d3_26;
	wire [WIDTH-1:0] wire_d3_27;
	wire [WIDTH-1:0] wire_d3_28;
	wire [WIDTH-1:0] wire_d4_0;
	wire [WIDTH-1:0] wire_d4_1;
	wire [WIDTH-1:0] wire_d4_2;
	wire [WIDTH-1:0] wire_d4_3;
	wire [WIDTH-1:0] wire_d4_4;
	wire [WIDTH-1:0] wire_d4_5;
	wire [WIDTH-1:0] wire_d4_6;
	wire [WIDTH-1:0] wire_d4_7;
	wire [WIDTH-1:0] wire_d4_8;
	wire [WIDTH-1:0] wire_d4_9;
	wire [WIDTH-1:0] wire_d4_10;
	wire [WIDTH-1:0] wire_d4_11;
	wire [WIDTH-1:0] wire_d4_12;
	wire [WIDTH-1:0] wire_d4_13;
	wire [WIDTH-1:0] wire_d4_14;
	wire [WIDTH-1:0] wire_d4_15;
	wire [WIDTH-1:0] wire_d4_16;
	wire [WIDTH-1:0] wire_d4_17;
	wire [WIDTH-1:0] wire_d4_18;
	wire [WIDTH-1:0] wire_d4_19;
	wire [WIDTH-1:0] wire_d4_20;
	wire [WIDTH-1:0] wire_d4_21;
	wire [WIDTH-1:0] wire_d4_22;
	wire [WIDTH-1:0] wire_d4_23;
	wire [WIDTH-1:0] wire_d4_24;
	wire [WIDTH-1:0] wire_d4_25;
	wire [WIDTH-1:0] wire_d4_26;
	wire [WIDTH-1:0] wire_d4_27;
	wire [WIDTH-1:0] wire_d4_28;
	wire [WIDTH-1:0] wire_d5_0;
	wire [WIDTH-1:0] wire_d5_1;
	wire [WIDTH-1:0] wire_d5_2;
	wire [WIDTH-1:0] wire_d5_3;
	wire [WIDTH-1:0] wire_d5_4;
	wire [WIDTH-1:0] wire_d5_5;
	wire [WIDTH-1:0] wire_d5_6;
	wire [WIDTH-1:0] wire_d5_7;
	wire [WIDTH-1:0] wire_d5_8;
	wire [WIDTH-1:0] wire_d5_9;
	wire [WIDTH-1:0] wire_d5_10;
	wire [WIDTH-1:0] wire_d5_11;
	wire [WIDTH-1:0] wire_d5_12;
	wire [WIDTH-1:0] wire_d5_13;
	wire [WIDTH-1:0] wire_d5_14;
	wire [WIDTH-1:0] wire_d5_15;
	wire [WIDTH-1:0] wire_d5_16;
	wire [WIDTH-1:0] wire_d5_17;
	wire [WIDTH-1:0] wire_d5_18;
	wire [WIDTH-1:0] wire_d5_19;
	wire [WIDTH-1:0] wire_d5_20;
	wire [WIDTH-1:0] wire_d5_21;
	wire [WIDTH-1:0] wire_d5_22;
	wire [WIDTH-1:0] wire_d5_23;
	wire [WIDTH-1:0] wire_d5_24;
	wire [WIDTH-1:0] wire_d5_25;
	wire [WIDTH-1:0] wire_d5_26;
	wire [WIDTH-1:0] wire_d5_27;
	wire [WIDTH-1:0] wire_d5_28;
	wire [WIDTH-1:0] wire_d6_0;
	wire [WIDTH-1:0] wire_d6_1;
	wire [WIDTH-1:0] wire_d6_2;
	wire [WIDTH-1:0] wire_d6_3;
	wire [WIDTH-1:0] wire_d6_4;
	wire [WIDTH-1:0] wire_d6_5;
	wire [WIDTH-1:0] wire_d6_6;
	wire [WIDTH-1:0] wire_d6_7;
	wire [WIDTH-1:0] wire_d6_8;
	wire [WIDTH-1:0] wire_d6_9;
	wire [WIDTH-1:0] wire_d6_10;
	wire [WIDTH-1:0] wire_d6_11;
	wire [WIDTH-1:0] wire_d6_12;
	wire [WIDTH-1:0] wire_d6_13;
	wire [WIDTH-1:0] wire_d6_14;
	wire [WIDTH-1:0] wire_d6_15;
	wire [WIDTH-1:0] wire_d6_16;
	wire [WIDTH-1:0] wire_d6_17;
	wire [WIDTH-1:0] wire_d6_18;
	wire [WIDTH-1:0] wire_d6_19;
	wire [WIDTH-1:0] wire_d6_20;
	wire [WIDTH-1:0] wire_d6_21;
	wire [WIDTH-1:0] wire_d6_22;
	wire [WIDTH-1:0] wire_d6_23;
	wire [WIDTH-1:0] wire_d6_24;
	wire [WIDTH-1:0] wire_d6_25;
	wire [WIDTH-1:0] wire_d6_26;
	wire [WIDTH-1:0] wire_d6_27;
	wire [WIDTH-1:0] wire_d6_28;
	wire [WIDTH-1:0] wire_d7_0;
	wire [WIDTH-1:0] wire_d7_1;
	wire [WIDTH-1:0] wire_d7_2;
	wire [WIDTH-1:0] wire_d7_3;
	wire [WIDTH-1:0] wire_d7_4;
	wire [WIDTH-1:0] wire_d7_5;
	wire [WIDTH-1:0] wire_d7_6;
	wire [WIDTH-1:0] wire_d7_7;
	wire [WIDTH-1:0] wire_d7_8;
	wire [WIDTH-1:0] wire_d7_9;
	wire [WIDTH-1:0] wire_d7_10;
	wire [WIDTH-1:0] wire_d7_11;
	wire [WIDTH-1:0] wire_d7_12;
	wire [WIDTH-1:0] wire_d7_13;
	wire [WIDTH-1:0] wire_d7_14;
	wire [WIDTH-1:0] wire_d7_15;
	wire [WIDTH-1:0] wire_d7_16;
	wire [WIDTH-1:0] wire_d7_17;
	wire [WIDTH-1:0] wire_d7_18;
	wire [WIDTH-1:0] wire_d7_19;
	wire [WIDTH-1:0] wire_d7_20;
	wire [WIDTH-1:0] wire_d7_21;
	wire [WIDTH-1:0] wire_d7_22;
	wire [WIDTH-1:0] wire_d7_23;
	wire [WIDTH-1:0] wire_d7_24;
	wire [WIDTH-1:0] wire_d7_25;
	wire [WIDTH-1:0] wire_d7_26;
	wire [WIDTH-1:0] wire_d7_27;
	wire [WIDTH-1:0] wire_d7_28;
	wire [WIDTH-1:0] wire_d8_0;
	wire [WIDTH-1:0] wire_d8_1;
	wire [WIDTH-1:0] wire_d8_2;
	wire [WIDTH-1:0] wire_d8_3;
	wire [WIDTH-1:0] wire_d8_4;
	wire [WIDTH-1:0] wire_d8_5;
	wire [WIDTH-1:0] wire_d8_6;
	wire [WIDTH-1:0] wire_d8_7;
	wire [WIDTH-1:0] wire_d8_8;
	wire [WIDTH-1:0] wire_d8_9;
	wire [WIDTH-1:0] wire_d8_10;
	wire [WIDTH-1:0] wire_d8_11;
	wire [WIDTH-1:0] wire_d8_12;
	wire [WIDTH-1:0] wire_d8_13;
	wire [WIDTH-1:0] wire_d8_14;
	wire [WIDTH-1:0] wire_d8_15;
	wire [WIDTH-1:0] wire_d8_16;
	wire [WIDTH-1:0] wire_d8_17;
	wire [WIDTH-1:0] wire_d8_18;
	wire [WIDTH-1:0] wire_d8_19;
	wire [WIDTH-1:0] wire_d8_20;
	wire [WIDTH-1:0] wire_d8_21;
	wire [WIDTH-1:0] wire_d8_22;
	wire [WIDTH-1:0] wire_d8_23;
	wire [WIDTH-1:0] wire_d8_24;
	wire [WIDTH-1:0] wire_d8_25;
	wire [WIDTH-1:0] wire_d8_26;
	wire [WIDTH-1:0] wire_d8_27;
	wire [WIDTH-1:0] wire_d8_28;
	wire [WIDTH-1:0] wire_d9_0;
	wire [WIDTH-1:0] wire_d9_1;
	wire [WIDTH-1:0] wire_d9_2;
	wire [WIDTH-1:0] wire_d9_3;
	wire [WIDTH-1:0] wire_d9_4;
	wire [WIDTH-1:0] wire_d9_5;
	wire [WIDTH-1:0] wire_d9_6;
	wire [WIDTH-1:0] wire_d9_7;
	wire [WIDTH-1:0] wire_d9_8;
	wire [WIDTH-1:0] wire_d9_9;
	wire [WIDTH-1:0] wire_d9_10;
	wire [WIDTH-1:0] wire_d9_11;
	wire [WIDTH-1:0] wire_d9_12;
	wire [WIDTH-1:0] wire_d9_13;
	wire [WIDTH-1:0] wire_d9_14;
	wire [WIDTH-1:0] wire_d9_15;
	wire [WIDTH-1:0] wire_d9_16;
	wire [WIDTH-1:0] wire_d9_17;
	wire [WIDTH-1:0] wire_d9_18;
	wire [WIDTH-1:0] wire_d9_19;
	wire [WIDTH-1:0] wire_d9_20;
	wire [WIDTH-1:0] wire_d9_21;
	wire [WIDTH-1:0] wire_d9_22;
	wire [WIDTH-1:0] wire_d9_23;
	wire [WIDTH-1:0] wire_d9_24;
	wire [WIDTH-1:0] wire_d9_25;
	wire [WIDTH-1:0] wire_d9_26;
	wire [WIDTH-1:0] wire_d9_27;
	wire [WIDTH-1:0] wire_d9_28;
	wire [WIDTH-1:0] wire_d10_0;
	wire [WIDTH-1:0] wire_d10_1;
	wire [WIDTH-1:0] wire_d10_2;
	wire [WIDTH-1:0] wire_d10_3;
	wire [WIDTH-1:0] wire_d10_4;
	wire [WIDTH-1:0] wire_d10_5;
	wire [WIDTH-1:0] wire_d10_6;
	wire [WIDTH-1:0] wire_d10_7;
	wire [WIDTH-1:0] wire_d10_8;
	wire [WIDTH-1:0] wire_d10_9;
	wire [WIDTH-1:0] wire_d10_10;
	wire [WIDTH-1:0] wire_d10_11;
	wire [WIDTH-1:0] wire_d10_12;
	wire [WIDTH-1:0] wire_d10_13;
	wire [WIDTH-1:0] wire_d10_14;
	wire [WIDTH-1:0] wire_d10_15;
	wire [WIDTH-1:0] wire_d10_16;
	wire [WIDTH-1:0] wire_d10_17;
	wire [WIDTH-1:0] wire_d10_18;
	wire [WIDTH-1:0] wire_d10_19;
	wire [WIDTH-1:0] wire_d10_20;
	wire [WIDTH-1:0] wire_d10_21;
	wire [WIDTH-1:0] wire_d10_22;
	wire [WIDTH-1:0] wire_d10_23;
	wire [WIDTH-1:0] wire_d10_24;
	wire [WIDTH-1:0] wire_d10_25;
	wire [WIDTH-1:0] wire_d10_26;
	wire [WIDTH-1:0] wire_d10_27;
	wire [WIDTH-1:0] wire_d10_28;
	wire [WIDTH-1:0] wire_d11_0;
	wire [WIDTH-1:0] wire_d11_1;
	wire [WIDTH-1:0] wire_d11_2;
	wire [WIDTH-1:0] wire_d11_3;
	wire [WIDTH-1:0] wire_d11_4;
	wire [WIDTH-1:0] wire_d11_5;
	wire [WIDTH-1:0] wire_d11_6;
	wire [WIDTH-1:0] wire_d11_7;
	wire [WIDTH-1:0] wire_d11_8;
	wire [WIDTH-1:0] wire_d11_9;
	wire [WIDTH-1:0] wire_d11_10;
	wire [WIDTH-1:0] wire_d11_11;
	wire [WIDTH-1:0] wire_d11_12;
	wire [WIDTH-1:0] wire_d11_13;
	wire [WIDTH-1:0] wire_d11_14;
	wire [WIDTH-1:0] wire_d11_15;
	wire [WIDTH-1:0] wire_d11_16;
	wire [WIDTH-1:0] wire_d11_17;
	wire [WIDTH-1:0] wire_d11_18;
	wire [WIDTH-1:0] wire_d11_19;
	wire [WIDTH-1:0] wire_d11_20;
	wire [WIDTH-1:0] wire_d11_21;
	wire [WIDTH-1:0] wire_d11_22;
	wire [WIDTH-1:0] wire_d11_23;
	wire [WIDTH-1:0] wire_d11_24;
	wire [WIDTH-1:0] wire_d11_25;
	wire [WIDTH-1:0] wire_d11_26;
	wire [WIDTH-1:0] wire_d11_27;
	wire [WIDTH-1:0] wire_d11_28;
	wire [WIDTH-1:0] wire_d12_0;
	wire [WIDTH-1:0] wire_d12_1;
	wire [WIDTH-1:0] wire_d12_2;
	wire [WIDTH-1:0] wire_d12_3;
	wire [WIDTH-1:0] wire_d12_4;
	wire [WIDTH-1:0] wire_d12_5;
	wire [WIDTH-1:0] wire_d12_6;
	wire [WIDTH-1:0] wire_d12_7;
	wire [WIDTH-1:0] wire_d12_8;
	wire [WIDTH-1:0] wire_d12_9;
	wire [WIDTH-1:0] wire_d12_10;
	wire [WIDTH-1:0] wire_d12_11;
	wire [WIDTH-1:0] wire_d12_12;
	wire [WIDTH-1:0] wire_d12_13;
	wire [WIDTH-1:0] wire_d12_14;
	wire [WIDTH-1:0] wire_d12_15;
	wire [WIDTH-1:0] wire_d12_16;
	wire [WIDTH-1:0] wire_d12_17;
	wire [WIDTH-1:0] wire_d12_18;
	wire [WIDTH-1:0] wire_d12_19;
	wire [WIDTH-1:0] wire_d12_20;
	wire [WIDTH-1:0] wire_d12_21;
	wire [WIDTH-1:0] wire_d12_22;
	wire [WIDTH-1:0] wire_d12_23;
	wire [WIDTH-1:0] wire_d12_24;
	wire [WIDTH-1:0] wire_d12_25;
	wire [WIDTH-1:0] wire_d12_26;
	wire [WIDTH-1:0] wire_d12_27;
	wire [WIDTH-1:0] wire_d12_28;
	wire [WIDTH-1:0] wire_d13_0;
	wire [WIDTH-1:0] wire_d13_1;
	wire [WIDTH-1:0] wire_d13_2;
	wire [WIDTH-1:0] wire_d13_3;
	wire [WIDTH-1:0] wire_d13_4;
	wire [WIDTH-1:0] wire_d13_5;
	wire [WIDTH-1:0] wire_d13_6;
	wire [WIDTH-1:0] wire_d13_7;
	wire [WIDTH-1:0] wire_d13_8;
	wire [WIDTH-1:0] wire_d13_9;
	wire [WIDTH-1:0] wire_d13_10;
	wire [WIDTH-1:0] wire_d13_11;
	wire [WIDTH-1:0] wire_d13_12;
	wire [WIDTH-1:0] wire_d13_13;
	wire [WIDTH-1:0] wire_d13_14;
	wire [WIDTH-1:0] wire_d13_15;
	wire [WIDTH-1:0] wire_d13_16;
	wire [WIDTH-1:0] wire_d13_17;
	wire [WIDTH-1:0] wire_d13_18;
	wire [WIDTH-1:0] wire_d13_19;
	wire [WIDTH-1:0] wire_d13_20;
	wire [WIDTH-1:0] wire_d13_21;
	wire [WIDTH-1:0] wire_d13_22;
	wire [WIDTH-1:0] wire_d13_23;
	wire [WIDTH-1:0] wire_d13_24;
	wire [WIDTH-1:0] wire_d13_25;
	wire [WIDTH-1:0] wire_d13_26;
	wire [WIDTH-1:0] wire_d13_27;
	wire [WIDTH-1:0] wire_d13_28;
	wire [WIDTH-1:0] wire_d14_0;
	wire [WIDTH-1:0] wire_d14_1;
	wire [WIDTH-1:0] wire_d14_2;
	wire [WIDTH-1:0] wire_d14_3;
	wire [WIDTH-1:0] wire_d14_4;
	wire [WIDTH-1:0] wire_d14_5;
	wire [WIDTH-1:0] wire_d14_6;
	wire [WIDTH-1:0] wire_d14_7;
	wire [WIDTH-1:0] wire_d14_8;
	wire [WIDTH-1:0] wire_d14_9;
	wire [WIDTH-1:0] wire_d14_10;
	wire [WIDTH-1:0] wire_d14_11;
	wire [WIDTH-1:0] wire_d14_12;
	wire [WIDTH-1:0] wire_d14_13;
	wire [WIDTH-1:0] wire_d14_14;
	wire [WIDTH-1:0] wire_d14_15;
	wire [WIDTH-1:0] wire_d14_16;
	wire [WIDTH-1:0] wire_d14_17;
	wire [WIDTH-1:0] wire_d14_18;
	wire [WIDTH-1:0] wire_d14_19;
	wire [WIDTH-1:0] wire_d14_20;
	wire [WIDTH-1:0] wire_d14_21;
	wire [WIDTH-1:0] wire_d14_22;
	wire [WIDTH-1:0] wire_d14_23;
	wire [WIDTH-1:0] wire_d14_24;
	wire [WIDTH-1:0] wire_d14_25;
	wire [WIDTH-1:0] wire_d14_26;
	wire [WIDTH-1:0] wire_d14_27;
	wire [WIDTH-1:0] wire_d14_28;
	wire [WIDTH-1:0] wire_d15_0;
	wire [WIDTH-1:0] wire_d15_1;
	wire [WIDTH-1:0] wire_d15_2;
	wire [WIDTH-1:0] wire_d15_3;
	wire [WIDTH-1:0] wire_d15_4;
	wire [WIDTH-1:0] wire_d15_5;
	wire [WIDTH-1:0] wire_d15_6;
	wire [WIDTH-1:0] wire_d15_7;
	wire [WIDTH-1:0] wire_d15_8;
	wire [WIDTH-1:0] wire_d15_9;
	wire [WIDTH-1:0] wire_d15_10;
	wire [WIDTH-1:0] wire_d15_11;
	wire [WIDTH-1:0] wire_d15_12;
	wire [WIDTH-1:0] wire_d15_13;
	wire [WIDTH-1:0] wire_d15_14;
	wire [WIDTH-1:0] wire_d15_15;
	wire [WIDTH-1:0] wire_d15_16;
	wire [WIDTH-1:0] wire_d15_17;
	wire [WIDTH-1:0] wire_d15_18;
	wire [WIDTH-1:0] wire_d15_19;
	wire [WIDTH-1:0] wire_d15_20;
	wire [WIDTH-1:0] wire_d15_21;
	wire [WIDTH-1:0] wire_d15_22;
	wire [WIDTH-1:0] wire_d15_23;
	wire [WIDTH-1:0] wire_d15_24;
	wire [WIDTH-1:0] wire_d15_25;
	wire [WIDTH-1:0] wire_d15_26;
	wire [WIDTH-1:0] wire_d15_27;
	wire [WIDTH-1:0] wire_d15_28;
	wire [WIDTH-1:0] wire_d16_0;
	wire [WIDTH-1:0] wire_d16_1;
	wire [WIDTH-1:0] wire_d16_2;
	wire [WIDTH-1:0] wire_d16_3;
	wire [WIDTH-1:0] wire_d16_4;
	wire [WIDTH-1:0] wire_d16_5;
	wire [WIDTH-1:0] wire_d16_6;
	wire [WIDTH-1:0] wire_d16_7;
	wire [WIDTH-1:0] wire_d16_8;
	wire [WIDTH-1:0] wire_d16_9;
	wire [WIDTH-1:0] wire_d16_10;
	wire [WIDTH-1:0] wire_d16_11;
	wire [WIDTH-1:0] wire_d16_12;
	wire [WIDTH-1:0] wire_d16_13;
	wire [WIDTH-1:0] wire_d16_14;
	wire [WIDTH-1:0] wire_d16_15;
	wire [WIDTH-1:0] wire_d16_16;
	wire [WIDTH-1:0] wire_d16_17;
	wire [WIDTH-1:0] wire_d16_18;
	wire [WIDTH-1:0] wire_d16_19;
	wire [WIDTH-1:0] wire_d16_20;
	wire [WIDTH-1:0] wire_d16_21;
	wire [WIDTH-1:0] wire_d16_22;
	wire [WIDTH-1:0] wire_d16_23;
	wire [WIDTH-1:0] wire_d16_24;
	wire [WIDTH-1:0] wire_d16_25;
	wire [WIDTH-1:0] wire_d16_26;
	wire [WIDTH-1:0] wire_d16_27;
	wire [WIDTH-1:0] wire_d16_28;
	wire [WIDTH-1:0] wire_d17_0;
	wire [WIDTH-1:0] wire_d17_1;
	wire [WIDTH-1:0] wire_d17_2;
	wire [WIDTH-1:0] wire_d17_3;
	wire [WIDTH-1:0] wire_d17_4;
	wire [WIDTH-1:0] wire_d17_5;
	wire [WIDTH-1:0] wire_d17_6;
	wire [WIDTH-1:0] wire_d17_7;
	wire [WIDTH-1:0] wire_d17_8;
	wire [WIDTH-1:0] wire_d17_9;
	wire [WIDTH-1:0] wire_d17_10;
	wire [WIDTH-1:0] wire_d17_11;
	wire [WIDTH-1:0] wire_d17_12;
	wire [WIDTH-1:0] wire_d17_13;
	wire [WIDTH-1:0] wire_d17_14;
	wire [WIDTH-1:0] wire_d17_15;
	wire [WIDTH-1:0] wire_d17_16;
	wire [WIDTH-1:0] wire_d17_17;
	wire [WIDTH-1:0] wire_d17_18;
	wire [WIDTH-1:0] wire_d17_19;
	wire [WIDTH-1:0] wire_d17_20;
	wire [WIDTH-1:0] wire_d17_21;
	wire [WIDTH-1:0] wire_d17_22;
	wire [WIDTH-1:0] wire_d17_23;
	wire [WIDTH-1:0] wire_d17_24;
	wire [WIDTH-1:0] wire_d17_25;
	wire [WIDTH-1:0] wire_d17_26;
	wire [WIDTH-1:0] wire_d17_27;
	wire [WIDTH-1:0] wire_d17_28;
	wire [WIDTH-1:0] wire_d18_0;
	wire [WIDTH-1:0] wire_d18_1;
	wire [WIDTH-1:0] wire_d18_2;
	wire [WIDTH-1:0] wire_d18_3;
	wire [WIDTH-1:0] wire_d18_4;
	wire [WIDTH-1:0] wire_d18_5;
	wire [WIDTH-1:0] wire_d18_6;
	wire [WIDTH-1:0] wire_d18_7;
	wire [WIDTH-1:0] wire_d18_8;
	wire [WIDTH-1:0] wire_d18_9;
	wire [WIDTH-1:0] wire_d18_10;
	wire [WIDTH-1:0] wire_d18_11;
	wire [WIDTH-1:0] wire_d18_12;
	wire [WIDTH-1:0] wire_d18_13;
	wire [WIDTH-1:0] wire_d18_14;
	wire [WIDTH-1:0] wire_d18_15;
	wire [WIDTH-1:0] wire_d18_16;
	wire [WIDTH-1:0] wire_d18_17;
	wire [WIDTH-1:0] wire_d18_18;
	wire [WIDTH-1:0] wire_d18_19;
	wire [WIDTH-1:0] wire_d18_20;
	wire [WIDTH-1:0] wire_d18_21;
	wire [WIDTH-1:0] wire_d18_22;
	wire [WIDTH-1:0] wire_d18_23;
	wire [WIDTH-1:0] wire_d18_24;
	wire [WIDTH-1:0] wire_d18_25;
	wire [WIDTH-1:0] wire_d18_26;
	wire [WIDTH-1:0] wire_d18_27;
	wire [WIDTH-1:0] wire_d18_28;
	wire [WIDTH-1:0] wire_d19_0;
	wire [WIDTH-1:0] wire_d19_1;
	wire [WIDTH-1:0] wire_d19_2;
	wire [WIDTH-1:0] wire_d19_3;
	wire [WIDTH-1:0] wire_d19_4;
	wire [WIDTH-1:0] wire_d19_5;
	wire [WIDTH-1:0] wire_d19_6;
	wire [WIDTH-1:0] wire_d19_7;
	wire [WIDTH-1:0] wire_d19_8;
	wire [WIDTH-1:0] wire_d19_9;
	wire [WIDTH-1:0] wire_d19_10;
	wire [WIDTH-1:0] wire_d19_11;
	wire [WIDTH-1:0] wire_d19_12;
	wire [WIDTH-1:0] wire_d19_13;
	wire [WIDTH-1:0] wire_d19_14;
	wire [WIDTH-1:0] wire_d19_15;
	wire [WIDTH-1:0] wire_d19_16;
	wire [WIDTH-1:0] wire_d19_17;
	wire [WIDTH-1:0] wire_d19_18;
	wire [WIDTH-1:0] wire_d19_19;
	wire [WIDTH-1:0] wire_d19_20;
	wire [WIDTH-1:0] wire_d19_21;
	wire [WIDTH-1:0] wire_d19_22;
	wire [WIDTH-1:0] wire_d19_23;
	wire [WIDTH-1:0] wire_d19_24;
	wire [WIDTH-1:0] wire_d19_25;
	wire [WIDTH-1:0] wire_d19_26;
	wire [WIDTH-1:0] wire_d19_27;
	wire [WIDTH-1:0] wire_d19_28;

	invertion #(.WIDTH(WIDTH)) invertion_instance100(.data_in(d_in0),.data_out(wire_d0_0),.clk(clk),.rst(rst));            //channel 1
	invertion #(.WIDTH(WIDTH)) invertion_instance101(.data_in(wire_d0_0),.data_out(wire_d0_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance102(.data_in(wire_d0_1),.data_out(wire_d0_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance103(.data_in(wire_d0_2),.data_out(wire_d0_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance104(.data_in(wire_d0_3),.data_out(wire_d0_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance105(.data_in(wire_d0_4),.data_out(wire_d0_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance106(.data_in(wire_d0_5),.data_out(wire_d0_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance107(.data_in(wire_d0_6),.data_out(wire_d0_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance108(.data_in(wire_d0_7),.data_out(wire_d0_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance109(.data_in(wire_d0_8),.data_out(wire_d0_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1010(.data_in(wire_d0_9),.data_out(wire_d0_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1011(.data_in(wire_d0_10),.data_out(wire_d0_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1012(.data_in(wire_d0_11),.data_out(wire_d0_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1013(.data_in(wire_d0_12),.data_out(wire_d0_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1014(.data_in(wire_d0_13),.data_out(wire_d0_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1015(.data_in(wire_d0_14),.data_out(wire_d0_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1016(.data_in(wire_d0_15),.data_out(wire_d0_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1017(.data_in(wire_d0_16),.data_out(wire_d0_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1018(.data_in(wire_d0_17),.data_out(wire_d0_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1019(.data_in(wire_d0_18),.data_out(wire_d0_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1020(.data_in(wire_d0_19),.data_out(wire_d0_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1021(.data_in(wire_d0_20),.data_out(wire_d0_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1022(.data_in(wire_d0_21),.data_out(wire_d0_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1023(.data_in(wire_d0_22),.data_out(wire_d0_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1024(.data_in(wire_d0_23),.data_out(wire_d0_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1025(.data_in(wire_d0_24),.data_out(wire_d0_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1026(.data_in(wire_d0_25),.data_out(wire_d0_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1027(.data_in(wire_d0_26),.data_out(wire_d0_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1028(.data_in(wire_d0_27),.data_out(wire_d0_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1029(.data_in(wire_d0_28),.data_out(d_out0),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance210(.data_in(d_in1),.data_out(wire_d1_0),.clk(clk),.rst(rst));            //channel 2
	invertion #(.WIDTH(WIDTH)) invertion_instance211(.data_in(wire_d1_0),.data_out(wire_d1_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212(.data_in(wire_d1_1),.data_out(wire_d1_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance213(.data_in(wire_d1_2),.data_out(wire_d1_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance214(.data_in(wire_d1_3),.data_out(wire_d1_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance215(.data_in(wire_d1_4),.data_out(wire_d1_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance216(.data_in(wire_d1_5),.data_out(wire_d1_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance217(.data_in(wire_d1_6),.data_out(wire_d1_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance218(.data_in(wire_d1_7),.data_out(wire_d1_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance219(.data_in(wire_d1_8),.data_out(wire_d1_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2110(.data_in(wire_d1_9),.data_out(wire_d1_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2111(.data_in(wire_d1_10),.data_out(wire_d1_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2112(.data_in(wire_d1_11),.data_out(wire_d1_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2113(.data_in(wire_d1_12),.data_out(wire_d1_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2114(.data_in(wire_d1_13),.data_out(wire_d1_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2115(.data_in(wire_d1_14),.data_out(wire_d1_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2116(.data_in(wire_d1_15),.data_out(wire_d1_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2117(.data_in(wire_d1_16),.data_out(wire_d1_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2118(.data_in(wire_d1_17),.data_out(wire_d1_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2119(.data_in(wire_d1_18),.data_out(wire_d1_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2120(.data_in(wire_d1_19),.data_out(wire_d1_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2121(.data_in(wire_d1_20),.data_out(wire_d1_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2122(.data_in(wire_d1_21),.data_out(wire_d1_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2123(.data_in(wire_d1_22),.data_out(wire_d1_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2124(.data_in(wire_d1_23),.data_out(wire_d1_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2125(.data_in(wire_d1_24),.data_out(wire_d1_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2126(.data_in(wire_d1_25),.data_out(wire_d1_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2127(.data_in(wire_d1_26),.data_out(wire_d1_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2128(.data_in(wire_d1_27),.data_out(wire_d1_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2129(.data_in(wire_d1_28),.data_out(d_out1),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance320(.data_in(d_in2),.data_out(wire_d2_0),.clk(clk),.rst(rst));            //channel 3
	large_mux #(.WIDTH(WIDTH)) large_mux_instance321(.data_in(wire_d2_0),.data_out(wire_d2_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance322(.data_in(wire_d2_1),.data_out(wire_d2_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323(.data_in(wire_d2_2),.data_out(wire_d2_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance324(.data_in(wire_d2_3),.data_out(wire_d2_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance325(.data_in(wire_d2_4),.data_out(wire_d2_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance326(.data_in(wire_d2_5),.data_out(wire_d2_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance327(.data_in(wire_d2_6),.data_out(wire_d2_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance328(.data_in(wire_d2_7),.data_out(wire_d2_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance329(.data_in(wire_d2_8),.data_out(wire_d2_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3210(.data_in(wire_d2_9),.data_out(wire_d2_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3211(.data_in(wire_d2_10),.data_out(wire_d2_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3212(.data_in(wire_d2_11),.data_out(wire_d2_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3213(.data_in(wire_d2_12),.data_out(wire_d2_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3214(.data_in(wire_d2_13),.data_out(wire_d2_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3215(.data_in(wire_d2_14),.data_out(wire_d2_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3216(.data_in(wire_d2_15),.data_out(wire_d2_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3217(.data_in(wire_d2_16),.data_out(wire_d2_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3218(.data_in(wire_d2_17),.data_out(wire_d2_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3219(.data_in(wire_d2_18),.data_out(wire_d2_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3220(.data_in(wire_d2_19),.data_out(wire_d2_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3221(.data_in(wire_d2_20),.data_out(wire_d2_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3222(.data_in(wire_d2_21),.data_out(wire_d2_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3223(.data_in(wire_d2_22),.data_out(wire_d2_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3224(.data_in(wire_d2_23),.data_out(wire_d2_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3225(.data_in(wire_d2_24),.data_out(wire_d2_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3226(.data_in(wire_d2_25),.data_out(wire_d2_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3227(.data_in(wire_d2_26),.data_out(wire_d2_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3228(.data_in(wire_d2_27),.data_out(wire_d2_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3229(.data_in(wire_d2_28),.data_out(d_out2),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance430(.data_in(d_in3),.data_out(wire_d3_0),.clk(clk),.rst(rst));            //channel 4
	register #(.WIDTH(WIDTH)) register_instance431(.data_in(wire_d3_0),.data_out(wire_d3_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance432(.data_in(wire_d3_1),.data_out(wire_d3_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance433(.data_in(wire_d3_2),.data_out(wire_d3_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434(.data_in(wire_d3_3),.data_out(wire_d3_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance435(.data_in(wire_d3_4),.data_out(wire_d3_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance436(.data_in(wire_d3_5),.data_out(wire_d3_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance437(.data_in(wire_d3_6),.data_out(wire_d3_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance438(.data_in(wire_d3_7),.data_out(wire_d3_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance439(.data_in(wire_d3_8),.data_out(wire_d3_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4310(.data_in(wire_d3_9),.data_out(wire_d3_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4311(.data_in(wire_d3_10),.data_out(wire_d3_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4312(.data_in(wire_d3_11),.data_out(wire_d3_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4313(.data_in(wire_d3_12),.data_out(wire_d3_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4314(.data_in(wire_d3_13),.data_out(wire_d3_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4315(.data_in(wire_d3_14),.data_out(wire_d3_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4316(.data_in(wire_d3_15),.data_out(wire_d3_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4317(.data_in(wire_d3_16),.data_out(wire_d3_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4318(.data_in(wire_d3_17),.data_out(wire_d3_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4319(.data_in(wire_d3_18),.data_out(wire_d3_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4320(.data_in(wire_d3_19),.data_out(wire_d3_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4321(.data_in(wire_d3_20),.data_out(wire_d3_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4322(.data_in(wire_d3_21),.data_out(wire_d3_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4323(.data_in(wire_d3_22),.data_out(wire_d3_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4324(.data_in(wire_d3_23),.data_out(wire_d3_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4325(.data_in(wire_d3_24),.data_out(wire_d3_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4326(.data_in(wire_d3_25),.data_out(wire_d3_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4327(.data_in(wire_d3_26),.data_out(wire_d3_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4328(.data_in(wire_d3_27),.data_out(wire_d3_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4329(.data_in(wire_d3_28),.data_out(d_out3),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance540(.data_in(d_in4),.data_out(wire_d4_0),.clk(clk),.rst(rst));            //channel 5
	large_mux #(.WIDTH(WIDTH)) large_mux_instance541(.data_in(wire_d4_0),.data_out(wire_d4_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance542(.data_in(wire_d4_1),.data_out(wire_d4_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance543(.data_in(wire_d4_2),.data_out(wire_d4_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance544(.data_in(wire_d4_3),.data_out(wire_d4_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance545(.data_in(wire_d4_4),.data_out(wire_d4_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance546(.data_in(wire_d4_5),.data_out(wire_d4_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance547(.data_in(wire_d4_6),.data_out(wire_d4_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance548(.data_in(wire_d4_7),.data_out(wire_d4_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance549(.data_in(wire_d4_8),.data_out(wire_d4_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5410(.data_in(wire_d4_9),.data_out(wire_d4_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5411(.data_in(wire_d4_10),.data_out(wire_d4_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5412(.data_in(wire_d4_11),.data_out(wire_d4_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5413(.data_in(wire_d4_12),.data_out(wire_d4_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5414(.data_in(wire_d4_13),.data_out(wire_d4_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5415(.data_in(wire_d4_14),.data_out(wire_d4_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5416(.data_in(wire_d4_15),.data_out(wire_d4_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5417(.data_in(wire_d4_16),.data_out(wire_d4_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5418(.data_in(wire_d4_17),.data_out(wire_d4_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5419(.data_in(wire_d4_18),.data_out(wire_d4_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5420(.data_in(wire_d4_19),.data_out(wire_d4_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5421(.data_in(wire_d4_20),.data_out(wire_d4_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5422(.data_in(wire_d4_21),.data_out(wire_d4_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5423(.data_in(wire_d4_22),.data_out(wire_d4_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5424(.data_in(wire_d4_23),.data_out(wire_d4_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5425(.data_in(wire_d4_24),.data_out(wire_d4_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5426(.data_in(wire_d4_25),.data_out(wire_d4_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5427(.data_in(wire_d4_26),.data_out(wire_d4_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5428(.data_in(wire_d4_27),.data_out(wire_d4_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5429(.data_in(wire_d4_28),.data_out(d_out4),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance650(.data_in(d_in5),.data_out(wire_d5_0),.clk(clk),.rst(rst));            //channel 6
	encoder #(.WIDTH(WIDTH)) encoder_instance651(.data_in(wire_d5_0),.data_out(wire_d5_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance652(.data_in(wire_d5_1),.data_out(wire_d5_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance653(.data_in(wire_d5_2),.data_out(wire_d5_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance654(.data_in(wire_d5_3),.data_out(wire_d5_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance655(.data_in(wire_d5_4),.data_out(wire_d5_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656(.data_in(wire_d5_5),.data_out(wire_d5_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance657(.data_in(wire_d5_6),.data_out(wire_d5_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance658(.data_in(wire_d5_7),.data_out(wire_d5_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance659(.data_in(wire_d5_8),.data_out(wire_d5_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6510(.data_in(wire_d5_9),.data_out(wire_d5_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6511(.data_in(wire_d5_10),.data_out(wire_d5_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6512(.data_in(wire_d5_11),.data_out(wire_d5_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6513(.data_in(wire_d5_12),.data_out(wire_d5_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6514(.data_in(wire_d5_13),.data_out(wire_d5_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6515(.data_in(wire_d5_14),.data_out(wire_d5_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6516(.data_in(wire_d5_15),.data_out(wire_d5_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6517(.data_in(wire_d5_16),.data_out(wire_d5_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6518(.data_in(wire_d5_17),.data_out(wire_d5_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6519(.data_in(wire_d5_18),.data_out(wire_d5_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6520(.data_in(wire_d5_19),.data_out(wire_d5_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6521(.data_in(wire_d5_20),.data_out(wire_d5_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6522(.data_in(wire_d5_21),.data_out(wire_d5_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6523(.data_in(wire_d5_22),.data_out(wire_d5_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6524(.data_in(wire_d5_23),.data_out(wire_d5_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6525(.data_in(wire_d5_24),.data_out(wire_d5_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6526(.data_in(wire_d5_25),.data_out(wire_d5_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6527(.data_in(wire_d5_26),.data_out(wire_d5_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6528(.data_in(wire_d5_27),.data_out(wire_d5_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6529(.data_in(wire_d5_28),.data_out(d_out5),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance760(.data_in(d_in6),.data_out(wire_d6_0),.clk(clk),.rst(rst));            //channel 7
	encoder #(.WIDTH(WIDTH)) encoder_instance761(.data_in(wire_d6_0),.data_out(wire_d6_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance762(.data_in(wire_d6_1),.data_out(wire_d6_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance763(.data_in(wire_d6_2),.data_out(wire_d6_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance764(.data_in(wire_d6_3),.data_out(wire_d6_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance765(.data_in(wire_d6_4),.data_out(wire_d6_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance766(.data_in(wire_d6_5),.data_out(wire_d6_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767(.data_in(wire_d6_6),.data_out(wire_d6_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance768(.data_in(wire_d6_7),.data_out(wire_d6_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance769(.data_in(wire_d6_8),.data_out(wire_d6_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7610(.data_in(wire_d6_9),.data_out(wire_d6_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7611(.data_in(wire_d6_10),.data_out(wire_d6_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7612(.data_in(wire_d6_11),.data_out(wire_d6_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7613(.data_in(wire_d6_12),.data_out(wire_d6_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7614(.data_in(wire_d6_13),.data_out(wire_d6_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7615(.data_in(wire_d6_14),.data_out(wire_d6_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7616(.data_in(wire_d6_15),.data_out(wire_d6_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7617(.data_in(wire_d6_16),.data_out(wire_d6_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7618(.data_in(wire_d6_17),.data_out(wire_d6_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7619(.data_in(wire_d6_18),.data_out(wire_d6_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7620(.data_in(wire_d6_19),.data_out(wire_d6_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7621(.data_in(wire_d6_20),.data_out(wire_d6_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7622(.data_in(wire_d6_21),.data_out(wire_d6_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7623(.data_in(wire_d6_22),.data_out(wire_d6_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7624(.data_in(wire_d6_23),.data_out(wire_d6_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7625(.data_in(wire_d6_24),.data_out(wire_d6_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7626(.data_in(wire_d6_25),.data_out(wire_d6_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7627(.data_in(wire_d6_26),.data_out(wire_d6_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7628(.data_in(wire_d6_27),.data_out(wire_d6_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7629(.data_in(wire_d6_28),.data_out(d_out6),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance870(.data_in(d_in7),.data_out(wire_d7_0),.clk(clk),.rst(rst));            //channel 8
	register #(.WIDTH(WIDTH)) register_instance871(.data_in(wire_d7_0),.data_out(wire_d7_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance872(.data_in(wire_d7_1),.data_out(wire_d7_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance873(.data_in(wire_d7_2),.data_out(wire_d7_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance874(.data_in(wire_d7_3),.data_out(wire_d7_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance875(.data_in(wire_d7_4),.data_out(wire_d7_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance876(.data_in(wire_d7_5),.data_out(wire_d7_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance877(.data_in(wire_d7_6),.data_out(wire_d7_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance878(.data_in(wire_d7_7),.data_out(wire_d7_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance879(.data_in(wire_d7_8),.data_out(wire_d7_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8710(.data_in(wire_d7_9),.data_out(wire_d7_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8711(.data_in(wire_d7_10),.data_out(wire_d7_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8712(.data_in(wire_d7_11),.data_out(wire_d7_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8713(.data_in(wire_d7_12),.data_out(wire_d7_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8714(.data_in(wire_d7_13),.data_out(wire_d7_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8715(.data_in(wire_d7_14),.data_out(wire_d7_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8716(.data_in(wire_d7_15),.data_out(wire_d7_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8717(.data_in(wire_d7_16),.data_out(wire_d7_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8718(.data_in(wire_d7_17),.data_out(wire_d7_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8719(.data_in(wire_d7_18),.data_out(wire_d7_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8720(.data_in(wire_d7_19),.data_out(wire_d7_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8721(.data_in(wire_d7_20),.data_out(wire_d7_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8722(.data_in(wire_d7_21),.data_out(wire_d7_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8723(.data_in(wire_d7_22),.data_out(wire_d7_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8724(.data_in(wire_d7_23),.data_out(wire_d7_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8725(.data_in(wire_d7_24),.data_out(wire_d7_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8726(.data_in(wire_d7_25),.data_out(wire_d7_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8727(.data_in(wire_d7_26),.data_out(wire_d7_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8728(.data_in(wire_d7_27),.data_out(wire_d7_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8729(.data_in(wire_d7_28),.data_out(d_out7),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance980(.data_in(d_in8),.data_out(wire_d8_0),.clk(clk),.rst(rst));            //channel 9
	register #(.WIDTH(WIDTH)) register_instance981(.data_in(wire_d8_0),.data_out(wire_d8_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance982(.data_in(wire_d8_1),.data_out(wire_d8_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance983(.data_in(wire_d8_2),.data_out(wire_d8_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance984(.data_in(wire_d8_3),.data_out(wire_d8_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance985(.data_in(wire_d8_4),.data_out(wire_d8_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance986(.data_in(wire_d8_5),.data_out(wire_d8_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance987(.data_in(wire_d8_6),.data_out(wire_d8_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance988(.data_in(wire_d8_7),.data_out(wire_d8_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance989(.data_in(wire_d8_8),.data_out(wire_d8_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9810(.data_in(wire_d8_9),.data_out(wire_d8_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9811(.data_in(wire_d8_10),.data_out(wire_d8_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9812(.data_in(wire_d8_11),.data_out(wire_d8_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9813(.data_in(wire_d8_12),.data_out(wire_d8_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9814(.data_in(wire_d8_13),.data_out(wire_d8_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9815(.data_in(wire_d8_14),.data_out(wire_d8_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9816(.data_in(wire_d8_15),.data_out(wire_d8_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9817(.data_in(wire_d8_16),.data_out(wire_d8_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9818(.data_in(wire_d8_17),.data_out(wire_d8_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9819(.data_in(wire_d8_18),.data_out(wire_d8_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9820(.data_in(wire_d8_19),.data_out(wire_d8_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9821(.data_in(wire_d8_20),.data_out(wire_d8_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9822(.data_in(wire_d8_21),.data_out(wire_d8_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9823(.data_in(wire_d8_22),.data_out(wire_d8_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9824(.data_in(wire_d8_23),.data_out(wire_d8_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9825(.data_in(wire_d8_24),.data_out(wire_d8_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9826(.data_in(wire_d8_25),.data_out(wire_d8_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9827(.data_in(wire_d8_26),.data_out(wire_d8_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9828(.data_in(wire_d8_27),.data_out(wire_d8_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9829(.data_in(wire_d8_28),.data_out(d_out8),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance1090(.data_in(d_in9),.data_out(wire_d9_0),.clk(clk),.rst(rst));            //channel 10
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1091(.data_in(wire_d9_0),.data_out(wire_d9_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1092(.data_in(wire_d9_1),.data_out(wire_d9_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1093(.data_in(wire_d9_2),.data_out(wire_d9_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1094(.data_in(wire_d9_3),.data_out(wire_d9_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1095(.data_in(wire_d9_4),.data_out(wire_d9_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1096(.data_in(wire_d9_5),.data_out(wire_d9_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1097(.data_in(wire_d9_6),.data_out(wire_d9_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1098(.data_in(wire_d9_7),.data_out(wire_d9_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1099(.data_in(wire_d9_8),.data_out(wire_d9_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10910(.data_in(wire_d9_9),.data_out(wire_d9_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10911(.data_in(wire_d9_10),.data_out(wire_d9_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10912(.data_in(wire_d9_11),.data_out(wire_d9_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10913(.data_in(wire_d9_12),.data_out(wire_d9_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10914(.data_in(wire_d9_13),.data_out(wire_d9_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10915(.data_in(wire_d9_14),.data_out(wire_d9_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10916(.data_in(wire_d9_15),.data_out(wire_d9_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10917(.data_in(wire_d9_16),.data_out(wire_d9_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10918(.data_in(wire_d9_17),.data_out(wire_d9_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10919(.data_in(wire_d9_18),.data_out(wire_d9_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10920(.data_in(wire_d9_19),.data_out(wire_d9_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10921(.data_in(wire_d9_20),.data_out(wire_d9_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10922(.data_in(wire_d9_21),.data_out(wire_d9_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10923(.data_in(wire_d9_22),.data_out(wire_d9_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10924(.data_in(wire_d9_23),.data_out(wire_d9_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10925(.data_in(wire_d9_24),.data_out(wire_d9_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10926(.data_in(wire_d9_25),.data_out(wire_d9_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10927(.data_in(wire_d9_26),.data_out(wire_d9_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10928(.data_in(wire_d9_27),.data_out(wire_d9_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10929(.data_in(wire_d9_28),.data_out(d_out9),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance11100(.data_in(d_in10),.data_out(wire_d10_0),.clk(clk),.rst(rst));            //channel 11
	encoder #(.WIDTH(WIDTH)) encoder_instance11101(.data_in(wire_d10_0),.data_out(wire_d10_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance11102(.data_in(wire_d10_1),.data_out(wire_d10_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance11103(.data_in(wire_d10_2),.data_out(wire_d10_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance11104(.data_in(wire_d10_3),.data_out(wire_d10_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance11105(.data_in(wire_d10_4),.data_out(wire_d10_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance11106(.data_in(wire_d10_5),.data_out(wire_d10_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance11107(.data_in(wire_d10_6),.data_out(wire_d10_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance11108(.data_in(wire_d10_7),.data_out(wire_d10_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance11109(.data_in(wire_d10_8),.data_out(wire_d10_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111010(.data_in(wire_d10_9),.data_out(wire_d10_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111011(.data_in(wire_d10_10),.data_out(wire_d10_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111012(.data_in(wire_d10_11),.data_out(wire_d10_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111013(.data_in(wire_d10_12),.data_out(wire_d10_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111014(.data_in(wire_d10_13),.data_out(wire_d10_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111015(.data_in(wire_d10_14),.data_out(wire_d10_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111016(.data_in(wire_d10_15),.data_out(wire_d10_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111017(.data_in(wire_d10_16),.data_out(wire_d10_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111018(.data_in(wire_d10_17),.data_out(wire_d10_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111019(.data_in(wire_d10_18),.data_out(wire_d10_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111020(.data_in(wire_d10_19),.data_out(wire_d10_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111021(.data_in(wire_d10_20),.data_out(wire_d10_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111022(.data_in(wire_d10_21),.data_out(wire_d10_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111023(.data_in(wire_d10_22),.data_out(wire_d10_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111024(.data_in(wire_d10_23),.data_out(wire_d10_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111025(.data_in(wire_d10_24),.data_out(wire_d10_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111026(.data_in(wire_d10_25),.data_out(wire_d10_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111027(.data_in(wire_d10_26),.data_out(wire_d10_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111028(.data_in(wire_d10_27),.data_out(wire_d10_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111029(.data_in(wire_d10_28),.data_out(d_out10),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance12110(.data_in(d_in11),.data_out(wire_d11_0),.clk(clk),.rst(rst));            //channel 12
	encoder #(.WIDTH(WIDTH)) encoder_instance12111(.data_in(wire_d11_0),.data_out(wire_d11_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance12112(.data_in(wire_d11_1),.data_out(wire_d11_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance12113(.data_in(wire_d11_2),.data_out(wire_d11_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance12114(.data_in(wire_d11_3),.data_out(wire_d11_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance12115(.data_in(wire_d11_4),.data_out(wire_d11_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance12116(.data_in(wire_d11_5),.data_out(wire_d11_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance12117(.data_in(wire_d11_6),.data_out(wire_d11_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance12118(.data_in(wire_d11_7),.data_out(wire_d11_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance12119(.data_in(wire_d11_8),.data_out(wire_d11_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121110(.data_in(wire_d11_9),.data_out(wire_d11_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121111(.data_in(wire_d11_10),.data_out(wire_d11_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121112(.data_in(wire_d11_11),.data_out(wire_d11_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121113(.data_in(wire_d11_12),.data_out(wire_d11_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121114(.data_in(wire_d11_13),.data_out(wire_d11_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121115(.data_in(wire_d11_14),.data_out(wire_d11_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121116(.data_in(wire_d11_15),.data_out(wire_d11_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121117(.data_in(wire_d11_16),.data_out(wire_d11_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121118(.data_in(wire_d11_17),.data_out(wire_d11_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121119(.data_in(wire_d11_18),.data_out(wire_d11_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121120(.data_in(wire_d11_19),.data_out(wire_d11_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121121(.data_in(wire_d11_20),.data_out(wire_d11_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121122(.data_in(wire_d11_21),.data_out(wire_d11_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121123(.data_in(wire_d11_22),.data_out(wire_d11_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121124(.data_in(wire_d11_23),.data_out(wire_d11_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121125(.data_in(wire_d11_24),.data_out(wire_d11_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121126(.data_in(wire_d11_25),.data_out(wire_d11_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121127(.data_in(wire_d11_26),.data_out(wire_d11_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121128(.data_in(wire_d11_27),.data_out(wire_d11_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121129(.data_in(wire_d11_28),.data_out(d_out11),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance13120(.data_in(d_in12),.data_out(wire_d12_0),.clk(clk),.rst(rst));            //channel 13
	invertion #(.WIDTH(WIDTH)) invertion_instance13121(.data_in(wire_d12_0),.data_out(wire_d12_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance13122(.data_in(wire_d12_1),.data_out(wire_d12_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance13123(.data_in(wire_d12_2),.data_out(wire_d12_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance13124(.data_in(wire_d12_3),.data_out(wire_d12_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance13125(.data_in(wire_d12_4),.data_out(wire_d12_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance13126(.data_in(wire_d12_5),.data_out(wire_d12_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance13127(.data_in(wire_d12_6),.data_out(wire_d12_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance13128(.data_in(wire_d12_7),.data_out(wire_d12_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance13129(.data_in(wire_d12_8),.data_out(wire_d12_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131210(.data_in(wire_d12_9),.data_out(wire_d12_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131211(.data_in(wire_d12_10),.data_out(wire_d12_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131212(.data_in(wire_d12_11),.data_out(wire_d12_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131213(.data_in(wire_d12_12),.data_out(wire_d12_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131214(.data_in(wire_d12_13),.data_out(wire_d12_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131215(.data_in(wire_d12_14),.data_out(wire_d12_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131216(.data_in(wire_d12_15),.data_out(wire_d12_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131217(.data_in(wire_d12_16),.data_out(wire_d12_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131218(.data_in(wire_d12_17),.data_out(wire_d12_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131219(.data_in(wire_d12_18),.data_out(wire_d12_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131220(.data_in(wire_d12_19),.data_out(wire_d12_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131221(.data_in(wire_d12_20),.data_out(wire_d12_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131222(.data_in(wire_d12_21),.data_out(wire_d12_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131223(.data_in(wire_d12_22),.data_out(wire_d12_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131224(.data_in(wire_d12_23),.data_out(wire_d12_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131225(.data_in(wire_d12_24),.data_out(wire_d12_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131226(.data_in(wire_d12_25),.data_out(wire_d12_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131227(.data_in(wire_d12_26),.data_out(wire_d12_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131228(.data_in(wire_d12_27),.data_out(wire_d12_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131229(.data_in(wire_d12_28),.data_out(d_out12),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance14130(.data_in(d_in13),.data_out(wire_d13_0),.clk(clk),.rst(rst));            //channel 14
	large_mux #(.WIDTH(WIDTH)) large_mux_instance14131(.data_in(wire_d13_0),.data_out(wire_d13_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance14132(.data_in(wire_d13_1),.data_out(wire_d13_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance14133(.data_in(wire_d13_2),.data_out(wire_d13_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance14134(.data_in(wire_d13_3),.data_out(wire_d13_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance14135(.data_in(wire_d13_4),.data_out(wire_d13_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance14136(.data_in(wire_d13_5),.data_out(wire_d13_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance14137(.data_in(wire_d13_6),.data_out(wire_d13_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance14138(.data_in(wire_d13_7),.data_out(wire_d13_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance14139(.data_in(wire_d13_8),.data_out(wire_d13_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141310(.data_in(wire_d13_9),.data_out(wire_d13_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141311(.data_in(wire_d13_10),.data_out(wire_d13_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141312(.data_in(wire_d13_11),.data_out(wire_d13_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141313(.data_in(wire_d13_12),.data_out(wire_d13_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141314(.data_in(wire_d13_13),.data_out(wire_d13_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141315(.data_in(wire_d13_14),.data_out(wire_d13_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141316(.data_in(wire_d13_15),.data_out(wire_d13_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141317(.data_in(wire_d13_16),.data_out(wire_d13_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141318(.data_in(wire_d13_17),.data_out(wire_d13_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141319(.data_in(wire_d13_18),.data_out(wire_d13_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141320(.data_in(wire_d13_19),.data_out(wire_d13_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141321(.data_in(wire_d13_20),.data_out(wire_d13_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141322(.data_in(wire_d13_21),.data_out(wire_d13_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141323(.data_in(wire_d13_22),.data_out(wire_d13_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141324(.data_in(wire_d13_23),.data_out(wire_d13_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141325(.data_in(wire_d13_24),.data_out(wire_d13_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141326(.data_in(wire_d13_25),.data_out(wire_d13_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141327(.data_in(wire_d13_26),.data_out(wire_d13_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141328(.data_in(wire_d13_27),.data_out(wire_d13_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141329(.data_in(wire_d13_28),.data_out(d_out13),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance15140(.data_in(d_in14),.data_out(wire_d14_0),.clk(clk),.rst(rst));            //channel 15
	invertion #(.WIDTH(WIDTH)) invertion_instance15141(.data_in(wire_d14_0),.data_out(wire_d14_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance15142(.data_in(wire_d14_1),.data_out(wire_d14_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance15143(.data_in(wire_d14_2),.data_out(wire_d14_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance15144(.data_in(wire_d14_3),.data_out(wire_d14_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance15145(.data_in(wire_d14_4),.data_out(wire_d14_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance15146(.data_in(wire_d14_5),.data_out(wire_d14_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance15147(.data_in(wire_d14_6),.data_out(wire_d14_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance15148(.data_in(wire_d14_7),.data_out(wire_d14_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance15149(.data_in(wire_d14_8),.data_out(wire_d14_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151410(.data_in(wire_d14_9),.data_out(wire_d14_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151411(.data_in(wire_d14_10),.data_out(wire_d14_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151412(.data_in(wire_d14_11),.data_out(wire_d14_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151413(.data_in(wire_d14_12),.data_out(wire_d14_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151414(.data_in(wire_d14_13),.data_out(wire_d14_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151415(.data_in(wire_d14_14),.data_out(wire_d14_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151416(.data_in(wire_d14_15),.data_out(wire_d14_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151417(.data_in(wire_d14_16),.data_out(wire_d14_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151418(.data_in(wire_d14_17),.data_out(wire_d14_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151419(.data_in(wire_d14_18),.data_out(wire_d14_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151420(.data_in(wire_d14_19),.data_out(wire_d14_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151421(.data_in(wire_d14_20),.data_out(wire_d14_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151422(.data_in(wire_d14_21),.data_out(wire_d14_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151423(.data_in(wire_d14_22),.data_out(wire_d14_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151424(.data_in(wire_d14_23),.data_out(wire_d14_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151425(.data_in(wire_d14_24),.data_out(wire_d14_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151426(.data_in(wire_d14_25),.data_out(wire_d14_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151427(.data_in(wire_d14_26),.data_out(wire_d14_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151428(.data_in(wire_d14_27),.data_out(wire_d14_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151429(.data_in(wire_d14_28),.data_out(d_out14),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance16150(.data_in(d_in15),.data_out(wire_d15_0),.clk(clk),.rst(rst));            //channel 16
	encoder #(.WIDTH(WIDTH)) encoder_instance16151(.data_in(wire_d15_0),.data_out(wire_d15_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance16152(.data_in(wire_d15_1),.data_out(wire_d15_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance16153(.data_in(wire_d15_2),.data_out(wire_d15_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance16154(.data_in(wire_d15_3),.data_out(wire_d15_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance16155(.data_in(wire_d15_4),.data_out(wire_d15_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance16156(.data_in(wire_d15_5),.data_out(wire_d15_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance16157(.data_in(wire_d15_6),.data_out(wire_d15_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance16158(.data_in(wire_d15_7),.data_out(wire_d15_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance16159(.data_in(wire_d15_8),.data_out(wire_d15_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161510(.data_in(wire_d15_9),.data_out(wire_d15_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161511(.data_in(wire_d15_10),.data_out(wire_d15_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161512(.data_in(wire_d15_11),.data_out(wire_d15_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161513(.data_in(wire_d15_12),.data_out(wire_d15_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161514(.data_in(wire_d15_13),.data_out(wire_d15_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161515(.data_in(wire_d15_14),.data_out(wire_d15_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161516(.data_in(wire_d15_15),.data_out(wire_d15_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161517(.data_in(wire_d15_16),.data_out(wire_d15_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161518(.data_in(wire_d15_17),.data_out(wire_d15_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161519(.data_in(wire_d15_18),.data_out(wire_d15_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161520(.data_in(wire_d15_19),.data_out(wire_d15_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161521(.data_in(wire_d15_20),.data_out(wire_d15_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161522(.data_in(wire_d15_21),.data_out(wire_d15_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161523(.data_in(wire_d15_22),.data_out(wire_d15_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161524(.data_in(wire_d15_23),.data_out(wire_d15_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161525(.data_in(wire_d15_24),.data_out(wire_d15_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161526(.data_in(wire_d15_25),.data_out(wire_d15_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161527(.data_in(wire_d15_26),.data_out(wire_d15_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161528(.data_in(wire_d15_27),.data_out(wire_d15_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161529(.data_in(wire_d15_28),.data_out(d_out15),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance17160(.data_in(d_in16),.data_out(wire_d16_0),.clk(clk),.rst(rst));            //channel 17
	large_mux #(.WIDTH(WIDTH)) large_mux_instance17161(.data_in(wire_d16_0),.data_out(wire_d16_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance17162(.data_in(wire_d16_1),.data_out(wire_d16_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance17163(.data_in(wire_d16_2),.data_out(wire_d16_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance17164(.data_in(wire_d16_3),.data_out(wire_d16_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance17165(.data_in(wire_d16_4),.data_out(wire_d16_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance17166(.data_in(wire_d16_5),.data_out(wire_d16_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance17167(.data_in(wire_d16_6),.data_out(wire_d16_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance17168(.data_in(wire_d16_7),.data_out(wire_d16_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance17169(.data_in(wire_d16_8),.data_out(wire_d16_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171610(.data_in(wire_d16_9),.data_out(wire_d16_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171611(.data_in(wire_d16_10),.data_out(wire_d16_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171612(.data_in(wire_d16_11),.data_out(wire_d16_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171613(.data_in(wire_d16_12),.data_out(wire_d16_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171614(.data_in(wire_d16_13),.data_out(wire_d16_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171615(.data_in(wire_d16_14),.data_out(wire_d16_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171616(.data_in(wire_d16_15),.data_out(wire_d16_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171617(.data_in(wire_d16_16),.data_out(wire_d16_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171618(.data_in(wire_d16_17),.data_out(wire_d16_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171619(.data_in(wire_d16_18),.data_out(wire_d16_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171620(.data_in(wire_d16_19),.data_out(wire_d16_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171621(.data_in(wire_d16_20),.data_out(wire_d16_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171622(.data_in(wire_d16_21),.data_out(wire_d16_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171623(.data_in(wire_d16_22),.data_out(wire_d16_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171624(.data_in(wire_d16_23),.data_out(wire_d16_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171625(.data_in(wire_d16_24),.data_out(wire_d16_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171626(.data_in(wire_d16_25),.data_out(wire_d16_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171627(.data_in(wire_d16_26),.data_out(wire_d16_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171628(.data_in(wire_d16_27),.data_out(wire_d16_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171629(.data_in(wire_d16_28),.data_out(d_out16),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance18170(.data_in(d_in17),.data_out(wire_d17_0),.clk(clk),.rst(rst));            //channel 18
	encoder #(.WIDTH(WIDTH)) encoder_instance18171(.data_in(wire_d17_0),.data_out(wire_d17_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance18172(.data_in(wire_d17_1),.data_out(wire_d17_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance18173(.data_in(wire_d17_2),.data_out(wire_d17_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance18174(.data_in(wire_d17_3),.data_out(wire_d17_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance18175(.data_in(wire_d17_4),.data_out(wire_d17_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance18176(.data_in(wire_d17_5),.data_out(wire_d17_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance18177(.data_in(wire_d17_6),.data_out(wire_d17_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance18178(.data_in(wire_d17_7),.data_out(wire_d17_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance18179(.data_in(wire_d17_8),.data_out(wire_d17_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181710(.data_in(wire_d17_9),.data_out(wire_d17_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181711(.data_in(wire_d17_10),.data_out(wire_d17_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181712(.data_in(wire_d17_11),.data_out(wire_d17_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181713(.data_in(wire_d17_12),.data_out(wire_d17_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181714(.data_in(wire_d17_13),.data_out(wire_d17_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181715(.data_in(wire_d17_14),.data_out(wire_d17_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181716(.data_in(wire_d17_15),.data_out(wire_d17_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181717(.data_in(wire_d17_16),.data_out(wire_d17_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181718(.data_in(wire_d17_17),.data_out(wire_d17_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181719(.data_in(wire_d17_18),.data_out(wire_d17_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181720(.data_in(wire_d17_19),.data_out(wire_d17_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181721(.data_in(wire_d17_20),.data_out(wire_d17_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181722(.data_in(wire_d17_21),.data_out(wire_d17_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181723(.data_in(wire_d17_22),.data_out(wire_d17_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181724(.data_in(wire_d17_23),.data_out(wire_d17_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181725(.data_in(wire_d17_24),.data_out(wire_d17_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181726(.data_in(wire_d17_25),.data_out(wire_d17_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181727(.data_in(wire_d17_26),.data_out(wire_d17_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181728(.data_in(wire_d17_27),.data_out(wire_d17_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181729(.data_in(wire_d17_28),.data_out(d_out17),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance19180(.data_in(d_in18),.data_out(wire_d18_0),.clk(clk),.rst(rst));            //channel 19
	encoder #(.WIDTH(WIDTH)) encoder_instance19181(.data_in(wire_d18_0),.data_out(wire_d18_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance19182(.data_in(wire_d18_1),.data_out(wire_d18_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance19183(.data_in(wire_d18_2),.data_out(wire_d18_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance19184(.data_in(wire_d18_3),.data_out(wire_d18_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance19185(.data_in(wire_d18_4),.data_out(wire_d18_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance19186(.data_in(wire_d18_5),.data_out(wire_d18_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance19187(.data_in(wire_d18_6),.data_out(wire_d18_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance19188(.data_in(wire_d18_7),.data_out(wire_d18_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance19189(.data_in(wire_d18_8),.data_out(wire_d18_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191810(.data_in(wire_d18_9),.data_out(wire_d18_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191811(.data_in(wire_d18_10),.data_out(wire_d18_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191812(.data_in(wire_d18_11),.data_out(wire_d18_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191813(.data_in(wire_d18_12),.data_out(wire_d18_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191814(.data_in(wire_d18_13),.data_out(wire_d18_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191815(.data_in(wire_d18_14),.data_out(wire_d18_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191816(.data_in(wire_d18_15),.data_out(wire_d18_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191817(.data_in(wire_d18_16),.data_out(wire_d18_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191818(.data_in(wire_d18_17),.data_out(wire_d18_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191819(.data_in(wire_d18_18),.data_out(wire_d18_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191820(.data_in(wire_d18_19),.data_out(wire_d18_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191821(.data_in(wire_d18_20),.data_out(wire_d18_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191822(.data_in(wire_d18_21),.data_out(wire_d18_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191823(.data_in(wire_d18_22),.data_out(wire_d18_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191824(.data_in(wire_d18_23),.data_out(wire_d18_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191825(.data_in(wire_d18_24),.data_out(wire_d18_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191826(.data_in(wire_d18_25),.data_out(wire_d18_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191827(.data_in(wire_d18_26),.data_out(wire_d18_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191828(.data_in(wire_d18_27),.data_out(wire_d18_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191829(.data_in(wire_d18_28),.data_out(d_out18),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance20190(.data_in(d_in19),.data_out(wire_d19_0),.clk(clk),.rst(rst));            //channel 20
	large_mux #(.WIDTH(WIDTH)) large_mux_instance20191(.data_in(wire_d19_0),.data_out(wire_d19_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance20192(.data_in(wire_d19_1),.data_out(wire_d19_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance20193(.data_in(wire_d19_2),.data_out(wire_d19_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance20194(.data_in(wire_d19_3),.data_out(wire_d19_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance20195(.data_in(wire_d19_4),.data_out(wire_d19_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance20196(.data_in(wire_d19_5),.data_out(wire_d19_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance20197(.data_in(wire_d19_6),.data_out(wire_d19_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance20198(.data_in(wire_d19_7),.data_out(wire_d19_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance20199(.data_in(wire_d19_8),.data_out(wire_d19_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201910(.data_in(wire_d19_9),.data_out(wire_d19_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201911(.data_in(wire_d19_10),.data_out(wire_d19_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201912(.data_in(wire_d19_11),.data_out(wire_d19_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201913(.data_in(wire_d19_12),.data_out(wire_d19_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201914(.data_in(wire_d19_13),.data_out(wire_d19_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201915(.data_in(wire_d19_14),.data_out(wire_d19_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201916(.data_in(wire_d19_15),.data_out(wire_d19_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201917(.data_in(wire_d19_16),.data_out(wire_d19_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201918(.data_in(wire_d19_17),.data_out(wire_d19_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201919(.data_in(wire_d19_18),.data_out(wire_d19_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201920(.data_in(wire_d19_19),.data_out(wire_d19_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201921(.data_in(wire_d19_20),.data_out(wire_d19_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201922(.data_in(wire_d19_21),.data_out(wire_d19_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201923(.data_in(wire_d19_22),.data_out(wire_d19_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201924(.data_in(wire_d19_23),.data_out(wire_d19_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201925(.data_in(wire_d19_24),.data_out(wire_d19_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201926(.data_in(wire_d19_25),.data_out(wire_d19_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201927(.data_in(wire_d19_26),.data_out(wire_d19_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201928(.data_in(wire_d19_27),.data_out(wire_d19_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201929(.data_in(wire_d19_28),.data_out(d_out19),.clk(clk),.rst(rst));


endmodule