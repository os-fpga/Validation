/******************** Computation *********************/

/***** package *****/
package pkg_computation;
	import globalDefinitions::*;
	
	// ---- public params ---- //		

	// ---- private params --- //	

endpackage
