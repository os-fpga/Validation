module InverseSubBytes(sub_byte,byte_out);
input [127:0] sub_byte;
output [127:0] byte_out;

function [7:0] bite;
    input [7:0] sbox_byte;

	begin  
		case(sbox_byte)
					8'h00:bite =8'h52;
					8'h01:bite =8'h09;
					8'h02:bite =8'h6a;
					8'h03:bite =8'hd5;
					8'h04:bite =8'h30;
					8'h05:bite =8'h36;
					8'h06:bite =8'ha5;
					8'h07:bite =8'h38;
					8'h08:bite =8'hbf;
					8'h09:bite =8'h40;
					8'h0a:bite =8'ha3;
					8'h0b:bite =8'h9e;
					8'h0c:bite =8'h81;
					8'h0d:bite =8'hf3;
					8'h0e:bite =8'hd7;
					8'h0f:bite =8'hfb;
					8'h10:bite =8'h7c;
					8'h11:bite =8'he3;
					8'h12:bite =8'h39;
					8'h13:bite =8'h82;
					8'h14:bite =8'h9b;
					8'h15:bite =8'h2f;
					8'h16:bite =8'hff;
					8'h17:bite =8'h87;
					8'h18:bite =8'h34;
					8'h19:bite =8'h8e;
					8'h1a:bite =8'h43;
					8'h1b:bite =8'h44;
					8'h1c:bite =8'hc4;
					8'h1d:bite =8'hde;
					8'h1e:bite =8'he9;
					8'h1f:bite =8'hcb;
					8'h20:bite =8'h54;
					8'h21:bite =8'h7b;
					8'h22:bite =8'h94;
					8'h23:bite =8'h32;
					8'h24:bite =8'ha6;
					8'h25:bite =8'hc2;
					8'h26:bite =8'h23;
					8'h27:bite =8'h3d;
					8'h28:bite =8'hee;
					8'h29:bite =8'h4c;
					8'h2a:bite =8'h95;
					8'h2b:bite =8'h0b;
					8'h2c:bite =8'h42;
					8'h2d:bite =8'hfa;
					8'h2e:bite =8'hc3;
					8'h2f:bite =8'h4e;
					8'h30:bite =8'h08;
					8'h31:bite =8'h2e;
					8'h32:bite =8'ha1;
					8'h33:bite =8'h66;
					8'h34:bite =8'h28;
					8'h35:bite =8'hd9;
					8'h36:bite =8'h24;
					8'h37:bite =8'hb2;
					8'h38:bite =8'h76;
					8'h39:bite =8'h5b;
					8'h3a:bite =8'ha2;
					8'h3b:bite =8'h49;
					8'h3c:bite =8'h6d;
					8'h3d:bite =8'h8b;
					8'h3e:bite =8'hd1;
					8'h3f:bite =8'h25;
					8'h40:bite =8'h72;
					8'h41:bite =8'hf8;
					8'h42:bite =8'hf6;
					8'h43:bite =8'h64;
					8'h44:bite =8'h86;
					8'h45:bite =8'h68;
					8'h46:bite =8'h98;
					8'h47:bite =8'h16;
					8'h48:bite =8'hd4;
					8'h49:bite =8'ha4;
					8'h4a:bite =8'h5c;
					8'h4b:bite =8'hcc;
					8'h4c:bite =8'h5d;
					8'h4d:bite =8'h65;
					8'h4e:bite =8'hb6;
					8'h4f:bite =8'h92;
					8'h50:bite =8'h6c;
					8'h51:bite =8'h70;
					8'h52:bite =8'h48;
					8'h53:bite =8'h50;
					8'h54:bite =8'hfd;
					8'h55:bite =8'hed;
					8'h56:bite =8'hb9;
					8'h57:bite =8'hda;
					8'h58:bite =8'h5e;
					8'h59:bite =8'h15;
					8'h5a:bite =8'h46;
					8'h5b:bite =8'h57;
					8'h5c:bite =8'ha7;
					8'h5d:bite =8'h8d;
					8'h5e:bite =8'h9d;
					8'h5f:bite =8'h84;
					8'h60:bite =8'h90;
					8'h61:bite =8'hd8;
					8'h62:bite =8'hab;
					8'h63:bite =8'h00;
					8'h64:bite =8'h8c;
					8'h65:bite =8'hbc;
					8'h66:bite =8'hd3;
					8'h67:bite =8'h0a;
					8'h68:bite =8'hf7;
					8'h69:bite =8'he4;
					8'h6a:bite =8'h58;
					8'h6b:bite =8'h05;
					8'h6c:bite =8'hb8;
					8'h6d:bite =8'hb3;
					8'h6e:bite =8'h45;
					8'h6f:bite =8'h06;
					8'h70:bite =8'hd0;
					8'h71:bite =8'h2c;
					8'h72:bite =8'h1e;
					8'h73:bite =8'h8f;
					8'h74:bite =8'hca;
					8'h75:bite =8'h3f;
					8'h76:bite =8'h0f;
					8'h77:bite =8'h02;
					8'h78:bite =8'hc1;
					8'h79:bite =8'haf;
					8'h7a:bite =8'hbd;
					8'h7b:bite =8'h03;
					8'h7c:bite =8'h01;
					8'h7d:bite =8'h13;
					8'h7e:bite =8'h8a;
					8'h7f:bite =8'h6b;
					8'h80:bite =8'h3a;
					8'h81:bite =8'h91;
					8'h82:bite =8'h11;
					8'h83:bite =8'h41;
					8'h84:bite =8'h4f;
					8'h85:bite =8'h67;
					8'h86:bite =8'hdc;
					8'h87:bite =8'hea;
					8'h88:bite =8'h97;
					8'h89:bite =8'hf2;
					8'h8a:bite =8'hcf;
					8'h8b:bite =8'hce;
					8'h8c:bite =8'hf0;
					8'h8d:bite =8'hb4;
					8'h8e:bite =8'he6;
					8'h8f:bite =8'h73;
					8'h90:bite =8'h96;
					8'h91:bite =8'hac;
					8'h92:bite =8'h74;
					8'h93:bite =8'h22;
					8'h94:bite =8'he7;
					8'h95:bite =8'had;
					8'h96:bite =8'h35;
					8'h97:bite =8'h85;
					8'h98:bite =8'he2;
					8'h99:bite =8'hf9;
					8'h9a:bite =8'h37;
					8'h9b:bite =8'he8;
					8'h9c:bite =8'h1c;
					8'h9d:bite =8'h75;
					8'h9e:bite =8'hdf;
					8'h9f:bite =8'h6e;
					8'ha0:bite =8'h47;
					8'ha1:bite =8'hf1;
					8'ha2:bite =8'h1a;
					8'ha3:bite =8'h71;
					8'ha4:bite =8'h1d;
					8'ha5:bite =8'h29;
					8'ha6:bite =8'hc5;
					8'ha7:bite =8'h89;
					8'ha8:bite =8'h6f;
					8'ha9:bite =8'hb7;
					8'haa:bite =8'h62;
					8'hab:bite =8'h0e;
					8'hac:bite =8'haa;
					8'had:bite =8'h18;
					8'hae:bite =8'hbe;
					8'haf:bite =8'h1b;
					8'hb0:bite =8'hfc;
					8'hb1:bite =8'h56;
					8'hb2:bite =8'h3e;
					8'hb3:bite =8'h4b;
					8'hb4:bite =8'hc6;
					8'hb5:bite =8'hd2;
					8'hb6:bite =8'h79;
					8'hb7:bite =8'h20;
					8'hb8:bite =8'h9a;
					8'hb9:bite =8'hdb;
					8'hba:bite =8'hc0;
					8'hbb:bite =8'hfe;
					8'hbc:bite =8'h78;
					8'hbd:bite =8'hcd;
					8'hbe:bite =8'h5a;
					8'hbf:bite =8'hf4;
					8'hc0:bite =8'h1f;
					8'hc1:bite =8'hdd;
					8'hc2:bite =8'ha8;
					8'hc3:bite =8'h33;
					8'hc4:bite =8'h88;
					8'hc5:bite =8'h07;
					8'hc6:bite =8'hc7;
					8'hc7:bite =8'h31;
					8'hc8:bite =8'hb1;
					8'hc9:bite =8'h12;
					8'hca:bite =8'h10;
					8'hcb:bite =8'h59;
					8'hcc:bite =8'h27;
					8'hcd:bite =8'h80;
					8'hce:bite =8'hec;
					8'hcf:bite =8'h5f;
					8'hd0:bite =8'h60;
					8'hd1:bite =8'h51;
					8'hd2:bite =8'h7f;
					8'hd3:bite =8'ha9;
					8'hd4:bite =8'h19;
					8'hd5:bite =8'hb5;
					8'hd6:bite =8'h4a;
					8'hd7:bite =8'h0d;
					8'hd8:bite =8'h2d;
					8'hd9:bite =8'he5;
					8'hda:bite =8'h7a;
					8'hdb:bite =8'h9f;
					8'hdc:bite =8'h93;
					8'hdd:bite =8'hc9;
					8'hde:bite =8'h9c;
					8'hdf:bite =8'hef;
					8'he0:bite =8'ha0;
					8'he1:bite =8'he0;
					8'he2:bite =8'h3b;
					8'he3:bite =8'h4d;
					8'he4:bite =8'hae;
					8'he5:bite =8'h2a;
					8'he6:bite =8'hf5;
					8'he7:bite =8'hb0;
					8'he8:bite =8'hc8;
					8'he9:bite =8'heb;
					8'hea:bite =8'hbb;
					8'heb:bite =8'h3c;
					8'hec:bite =8'h83;
					8'hed:bite =8'h53;
					8'hee:bite =8'h99;
					8'hef:bite =8'h61;
					8'hf0:bite =8'h17;
					8'hf1:bite =8'h2b;
					8'hf2:bite =8'h04;
					8'hf3:bite =8'h7e;
					8'hf4:bite =8'hba;
					8'hf5:bite =8'h77;
					8'hf6:bite =8'hd6;
					8'hf7:bite =8'h26;
					8'hf8:bite =8'he1;
					8'hf9:bite =8'h69;
					8'hfa:bite =8'h14;
					8'hfb:bite =8'h63;
					8'hfc:bite =8'h55;
					8'hfd:bite =8'h21;
					8'hfe:bite =8'h0c;
					8'hff:bite =8'h7d;
					endcase
	end

endfunction

genvar i;

generate
	for(i = 0; i < 128; i = i+8) 
		assign byte_out[i +:8] = bite(sub_byte[i +:8]);
endgenerate


endmodule