//`include "encoder.v"
//`include "invertion.v"
//`include "large_mux.v"
//`include "register.v"
module design32_50_70_top #(parameter WIDTH=32,CHANNEL=50) (clk, rst, in, out);

	localparam OUT_BUS=CHANNEL*WIDTH;
	input clk,rst;
	input [WIDTH-1:0] in;
	output [WIDTH-1:0] out;

	reg [WIDTH-1:0] d_in0;
	reg [WIDTH-1:0] d_in1;
	reg [WIDTH-1:0] d_in2;
	reg [WIDTH-1:0] d_in3;
	reg [WIDTH-1:0] d_in4;
	reg [WIDTH-1:0] d_in5;
	reg [WIDTH-1:0] d_in6;
	reg [WIDTH-1:0] d_in7;
	reg [WIDTH-1:0] d_in8;
	reg [WIDTH-1:0] d_in9;
	reg [WIDTH-1:0] d_in10;
	reg [WIDTH-1:0] d_in11;
	reg [WIDTH-1:0] d_in12;
	reg [WIDTH-1:0] d_in13;
	reg [WIDTH-1:0] d_in14;
	reg [WIDTH-1:0] d_in15;
	reg [WIDTH-1:0] d_in16;
	reg [WIDTH-1:0] d_in17;
	reg [WIDTH-1:0] d_in18;
	reg [WIDTH-1:0] d_in19;
	reg [WIDTH-1:0] d_in20;
	reg [WIDTH-1:0] d_in21;
	reg [WIDTH-1:0] d_in22;
	reg [WIDTH-1:0] d_in23;
	reg [WIDTH-1:0] d_in24;
	reg [WIDTH-1:0] d_in25;
	reg [WIDTH-1:0] d_in26;
	reg [WIDTH-1:0] d_in27;
	reg [WIDTH-1:0] d_in28;
	reg [WIDTH-1:0] d_in29;
	reg [WIDTH-1:0] d_in30;
	reg [WIDTH-1:0] d_in31;
	reg [WIDTH-1:0] d_in32;
	reg [WIDTH-1:0] d_in33;
	reg [WIDTH-1:0] d_in34;
	reg [WIDTH-1:0] d_in35;
	reg [WIDTH-1:0] d_in36;
	reg [WIDTH-1:0] d_in37;
	reg [WIDTH-1:0] d_in38;
	reg [WIDTH-1:0] d_in39;
	reg [WIDTH-1:0] d_in40;
	reg [WIDTH-1:0] d_in41;
	reg [WIDTH-1:0] d_in42;
	reg [WIDTH-1:0] d_in43;
	reg [WIDTH-1:0] d_in44;
	reg [WIDTH-1:0] d_in45;
	reg [WIDTH-1:0] d_in46;
	reg [WIDTH-1:0] d_in47;
	reg [WIDTH-1:0] d_in48;
	reg [WIDTH-1:0] d_in49;
	wire [WIDTH-1:0] d_out0;
	wire [WIDTH-1:0] d_out1;
	wire [WIDTH-1:0] d_out2;
	wire [WIDTH-1:0] d_out3;
	wire [WIDTH-1:0] d_out4;
	wire [WIDTH-1:0] d_out5;
	wire [WIDTH-1:0] d_out6;
	wire [WIDTH-1:0] d_out7;
	wire [WIDTH-1:0] d_out8;
	wire [WIDTH-1:0] d_out9;
	wire [WIDTH-1:0] d_out10;
	wire [WIDTH-1:0] d_out11;
	wire [WIDTH-1:0] d_out12;
	wire [WIDTH-1:0] d_out13;
	wire [WIDTH-1:0] d_out14;
	wire [WIDTH-1:0] d_out15;
	wire [WIDTH-1:0] d_out16;
	wire [WIDTH-1:0] d_out17;
	wire [WIDTH-1:0] d_out18;
	wire [WIDTH-1:0] d_out19;
	wire [WIDTH-1:0] d_out20;
	wire [WIDTH-1:0] d_out21;
	wire [WIDTH-1:0] d_out22;
	wire [WIDTH-1:0] d_out23;
	wire [WIDTH-1:0] d_out24;
	wire [WIDTH-1:0] d_out25;
	wire [WIDTH-1:0] d_out26;
	wire [WIDTH-1:0] d_out27;
	wire [WIDTH-1:0] d_out28;
	wire [WIDTH-1:0] d_out29;
	wire [WIDTH-1:0] d_out30;
	wire [WIDTH-1:0] d_out31;
	wire [WIDTH-1:0] d_out32;
	wire [WIDTH-1:0] d_out33;
	wire [WIDTH-1:0] d_out34;
	wire [WIDTH-1:0] d_out35;
	wire [WIDTH-1:0] d_out36;
	wire [WIDTH-1:0] d_out37;
	wire [WIDTH-1:0] d_out38;
	wire [WIDTH-1:0] d_out39;
	wire [WIDTH-1:0] d_out40;
	wire [WIDTH-1:0] d_out41;
	wire [WIDTH-1:0] d_out42;
	wire [WIDTH-1:0] d_out43;
	wire [WIDTH-1:0] d_out44;
	wire [WIDTH-1:0] d_out45;
	wire [WIDTH-1:0] d_out46;
	wire [WIDTH-1:0] d_out47;
	wire [WIDTH-1:0] d_out48;
	wire [WIDTH-1:0] d_out49;

	reg [OUT_BUS-1:0] tmp;

	always @ (posedge clk or posedge rst) begin
		if (rst)
			tmp <= 0;
		else
			tmp <= {tmp[OUT_BUS-(WIDTH-1):0],in};
	end

	always @ (posedge clk) begin
		d_in0 <= tmp[WIDTH-1:0];
		d_in1 <= tmp[(WIDTH*2)-1:WIDTH*1];
		d_in2 <= tmp[(WIDTH*3)-1:WIDTH*2];
		d_in3 <= tmp[(WIDTH*4)-1:WIDTH*3];
		d_in4 <= tmp[(WIDTH*5)-1:WIDTH*4];
		d_in5 <= tmp[(WIDTH*6)-1:WIDTH*5];
		d_in6 <= tmp[(WIDTH*7)-1:WIDTH*6];
		d_in7 <= tmp[(WIDTH*8)-1:WIDTH*7];
		d_in8 <= tmp[(WIDTH*9)-1:WIDTH*8];
		d_in9 <= tmp[(WIDTH*10)-1:WIDTH*9];
		d_in10 <= tmp[(WIDTH*11)-1:WIDTH*10];
		d_in11 <= tmp[(WIDTH*12)-1:WIDTH*11];
		d_in12 <= tmp[(WIDTH*13)-1:WIDTH*12];
		d_in13 <= tmp[(WIDTH*14)-1:WIDTH*13];
		d_in14 <= tmp[(WIDTH*15)-1:WIDTH*14];
		d_in15 <= tmp[(WIDTH*16)-1:WIDTH*15];
		d_in16 <= tmp[(WIDTH*17)-1:WIDTH*16];
		d_in17 <= tmp[(WIDTH*18)-1:WIDTH*17];
		d_in18 <= tmp[(WIDTH*19)-1:WIDTH*18];
		d_in19 <= tmp[(WIDTH*20)-1:WIDTH*19];
		d_in20 <= tmp[(WIDTH*21)-1:WIDTH*20];
		d_in21 <= tmp[(WIDTH*22)-1:WIDTH*21];
		d_in22 <= tmp[(WIDTH*23)-1:WIDTH*22];
		d_in23 <= tmp[(WIDTH*24)-1:WIDTH*23];
		d_in24 <= tmp[(WIDTH*25)-1:WIDTH*24];
		d_in25 <= tmp[(WIDTH*26)-1:WIDTH*25];
		d_in26 <= tmp[(WIDTH*27)-1:WIDTH*26];
		d_in27 <= tmp[(WIDTH*28)-1:WIDTH*27];
		d_in28 <= tmp[(WIDTH*29)-1:WIDTH*28];
		d_in29 <= tmp[(WIDTH*30)-1:WIDTH*29];
		d_in30 <= tmp[(WIDTH*31)-1:WIDTH*30];
		d_in31 <= tmp[(WIDTH*32)-1:WIDTH*31];
		d_in32 <= tmp[(WIDTH*33)-1:WIDTH*32];
		d_in33 <= tmp[(WIDTH*34)-1:WIDTH*33];
		d_in34 <= tmp[(WIDTH*35)-1:WIDTH*34];
		d_in35 <= tmp[(WIDTH*36)-1:WIDTH*35];
		d_in36 <= tmp[(WIDTH*37)-1:WIDTH*36];
		d_in37 <= tmp[(WIDTH*38)-1:WIDTH*37];
		d_in38 <= tmp[(WIDTH*39)-1:WIDTH*38];
		d_in39 <= tmp[(WIDTH*40)-1:WIDTH*39];
		d_in40 <= tmp[(WIDTH*41)-1:WIDTH*40];
		d_in41 <= tmp[(WIDTH*42)-1:WIDTH*41];
		d_in42 <= tmp[(WIDTH*43)-1:WIDTH*42];
		d_in43 <= tmp[(WIDTH*44)-1:WIDTH*43];
		d_in44 <= tmp[(WIDTH*45)-1:WIDTH*44];
		d_in45 <= tmp[(WIDTH*46)-1:WIDTH*45];
		d_in46 <= tmp[(WIDTH*47)-1:WIDTH*46];
		d_in47 <= tmp[(WIDTH*48)-1:WIDTH*47];
		d_in48 <= tmp[(WIDTH*49)-1:WIDTH*48];
		d_in49 <= tmp[(WIDTH*50)-1:WIDTH*49];
	end

	design32_50_70 #(.WIDTH(WIDTH)) design32_50_70_inst(.d_in0(d_in0),.d_in1(d_in1),.d_in2(d_in2),.d_in3(d_in3),.d_in4(d_in4),.d_in5(d_in5),.d_in6(d_in6),.d_in7(d_in7),.d_in8(d_in8),.d_in9(d_in9),.d_in10(d_in10),.d_in11(d_in11),.d_in12(d_in12),.d_in13(d_in13),.d_in14(d_in14),.d_in15(d_in15),.d_in16(d_in16),.d_in17(d_in17),.d_in18(d_in18),.d_in19(d_in19),.d_in20(d_in20),.d_in21(d_in21),.d_in22(d_in22),.d_in23(d_in23),.d_in24(d_in24),.d_in25(d_in25),.d_in26(d_in26),.d_in27(d_in27),.d_in28(d_in28),.d_in29(d_in29),.d_in30(d_in30),.d_in31(d_in31),.d_in32(d_in32),.d_in33(d_in33),.d_in34(d_in34),.d_in35(d_in35),.d_in36(d_in36),.d_in37(d_in37),.d_in38(d_in38),.d_in39(d_in39),.d_in40(d_in40),.d_in41(d_in41),.d_in42(d_in42),.d_in43(d_in43),.d_in44(d_in44),.d_in45(d_in45),.d_in46(d_in46),.d_in47(d_in47),.d_in48(d_in48),.d_in49(d_in49),.d_out0(d_out0),.d_out1(d_out1),.d_out2(d_out2),.d_out3(d_out3),.d_out4(d_out4),.d_out5(d_out5),.d_out6(d_out6),.d_out7(d_out7),.d_out8(d_out8),.d_out9(d_out9),.d_out10(d_out10),.d_out11(d_out11),.d_out12(d_out12),.d_out13(d_out13),.d_out14(d_out14),.d_out15(d_out15),.d_out16(d_out16),.d_out17(d_out17),.d_out18(d_out18),.d_out19(d_out19),.d_out20(d_out20),.d_out21(d_out21),.d_out22(d_out22),.d_out23(d_out23),.d_out24(d_out24),.d_out25(d_out25),.d_out26(d_out26),.d_out27(d_out27),.d_out28(d_out28),.d_out29(d_out29),.d_out30(d_out30),.d_out31(d_out31),.d_out32(d_out32),.d_out33(d_out33),.d_out34(d_out34),.d_out35(d_out35),.d_out36(d_out36),.d_out37(d_out37),.d_out38(d_out38),.d_out39(d_out39),.d_out40(d_out40),.d_out41(d_out41),.d_out42(d_out42),.d_out43(d_out43),.d_out44(d_out44),.d_out45(d_out45),.d_out46(d_out46),.d_out47(d_out47),.d_out48(d_out48),.d_out49(d_out49),.clk(clk),.rst(rst));

	assign out = d_out0^d_out1^d_out2^d_out3^d_out4^d_out5^d_out6^d_out7^d_out8^d_out9^d_out10^d_out11^d_out12^d_out13^d_out14^d_out15^d_out16^d_out17^d_out18^d_out19^d_out20^d_out21^d_out22^d_out23^d_out24^d_out25^d_out26^d_out27^d_out28^d_out29^d_out30^d_out31^d_out32^d_out33^d_out34^d_out35^d_out36^d_out37^d_out38^d_out39^d_out40^d_out41^d_out42^d_out43^d_out44^d_out45^d_out46^d_out47^d_out48^d_out49;

endmodule

module design32_50_70 #(parameter WIDTH=32) (d_in0, d_in1, d_in2, d_in3, d_in4, d_in5, d_in6, d_in7, d_in8, d_in9, d_in10, d_in11, d_in12, d_in13, d_in14, d_in15, d_in16, d_in17, d_in18, d_in19, d_in20, d_in21, d_in22, d_in23, d_in24, d_in25, d_in26, d_in27, d_in28, d_in29, d_in30, d_in31, d_in32, d_in33, d_in34, d_in35, d_in36, d_in37, d_in38, d_in39, d_in40, d_in41, d_in42, d_in43, d_in44, d_in45, d_in46, d_in47, d_in48, d_in49, d_out0, d_out1, d_out2, d_out3, d_out4, d_out5, d_out6, d_out7, d_out8, d_out9, d_out10, d_out11, d_out12, d_out13, d_out14, d_out15, d_out16, d_out17, d_out18, d_out19, d_out20, d_out21, d_out22, d_out23, d_out24, d_out25, d_out26, d_out27, d_out28, d_out29, d_out30, d_out31, d_out32, d_out33, d_out34, d_out35, d_out36, d_out37, d_out38, d_out39, d_out40, d_out41, d_out42, d_out43, d_out44, d_out45, d_out46, d_out47, d_out48, d_out49, clk, rst);
	input clk;
	input rst;
	input [WIDTH-1:0] d_in0; 
	input [WIDTH-1:0] d_in1; 
	input [WIDTH-1:0] d_in2; 
	input [WIDTH-1:0] d_in3; 
	input [WIDTH-1:0] d_in4; 
	input [WIDTH-1:0] d_in5; 
	input [WIDTH-1:0] d_in6; 
	input [WIDTH-1:0] d_in7; 
	input [WIDTH-1:0] d_in8; 
	input [WIDTH-1:0] d_in9; 
	input [WIDTH-1:0] d_in10; 
	input [WIDTH-1:0] d_in11; 
	input [WIDTH-1:0] d_in12; 
	input [WIDTH-1:0] d_in13; 
	input [WIDTH-1:0] d_in14; 
	input [WIDTH-1:0] d_in15; 
	input [WIDTH-1:0] d_in16; 
	input [WIDTH-1:0] d_in17; 
	input [WIDTH-1:0] d_in18; 
	input [WIDTH-1:0] d_in19; 
	input [WIDTH-1:0] d_in20; 
	input [WIDTH-1:0] d_in21; 
	input [WIDTH-1:0] d_in22; 
	input [WIDTH-1:0] d_in23; 
	input [WIDTH-1:0] d_in24; 
	input [WIDTH-1:0] d_in25; 
	input [WIDTH-1:0] d_in26; 
	input [WIDTH-1:0] d_in27; 
	input [WIDTH-1:0] d_in28; 
	input [WIDTH-1:0] d_in29; 
	input [WIDTH-1:0] d_in30; 
	input [WIDTH-1:0] d_in31; 
	input [WIDTH-1:0] d_in32; 
	input [WIDTH-1:0] d_in33; 
	input [WIDTH-1:0] d_in34; 
	input [WIDTH-1:0] d_in35; 
	input [WIDTH-1:0] d_in36; 
	input [WIDTH-1:0] d_in37; 
	input [WIDTH-1:0] d_in38; 
	input [WIDTH-1:0] d_in39; 
	input [WIDTH-1:0] d_in40; 
	input [WIDTH-1:0] d_in41; 
	input [WIDTH-1:0] d_in42; 
	input [WIDTH-1:0] d_in43; 
	input [WIDTH-1:0] d_in44; 
	input [WIDTH-1:0] d_in45; 
	input [WIDTH-1:0] d_in46; 
	input [WIDTH-1:0] d_in47; 
	input [WIDTH-1:0] d_in48; 
	input [WIDTH-1:0] d_in49; 
	output [WIDTH-1:0] d_out0; 
	output [WIDTH-1:0] d_out1; 
	output [WIDTH-1:0] d_out2; 
	output [WIDTH-1:0] d_out3; 
	output [WIDTH-1:0] d_out4; 
	output [WIDTH-1:0] d_out5; 
	output [WIDTH-1:0] d_out6; 
	output [WIDTH-1:0] d_out7; 
	output [WIDTH-1:0] d_out8; 
	output [WIDTH-1:0] d_out9; 
	output [WIDTH-1:0] d_out10; 
	output [WIDTH-1:0] d_out11; 
	output [WIDTH-1:0] d_out12; 
	output [WIDTH-1:0] d_out13; 
	output [WIDTH-1:0] d_out14; 
	output [WIDTH-1:0] d_out15; 
	output [WIDTH-1:0] d_out16; 
	output [WIDTH-1:0] d_out17; 
	output [WIDTH-1:0] d_out18; 
	output [WIDTH-1:0] d_out19; 
	output [WIDTH-1:0] d_out20; 
	output [WIDTH-1:0] d_out21; 
	output [WIDTH-1:0] d_out22; 
	output [WIDTH-1:0] d_out23; 
	output [WIDTH-1:0] d_out24; 
	output [WIDTH-1:0] d_out25; 
	output [WIDTH-1:0] d_out26; 
	output [WIDTH-1:0] d_out27; 
	output [WIDTH-1:0] d_out28; 
	output [WIDTH-1:0] d_out29; 
	output [WIDTH-1:0] d_out30; 
	output [WIDTH-1:0] d_out31; 
	output [WIDTH-1:0] d_out32; 
	output [WIDTH-1:0] d_out33; 
	output [WIDTH-1:0] d_out34; 
	output [WIDTH-1:0] d_out35; 
	output [WIDTH-1:0] d_out36; 
	output [WIDTH-1:0] d_out37; 
	output [WIDTH-1:0] d_out38; 
	output [WIDTH-1:0] d_out39; 
	output [WIDTH-1:0] d_out40; 
	output [WIDTH-1:0] d_out41; 
	output [WIDTH-1:0] d_out42; 
	output [WIDTH-1:0] d_out43; 
	output [WIDTH-1:0] d_out44; 
	output [WIDTH-1:0] d_out45; 
	output [WIDTH-1:0] d_out46; 
	output [WIDTH-1:0] d_out47; 
	output [WIDTH-1:0] d_out48; 
	output [WIDTH-1:0] d_out49; 

	wire [WIDTH-1:0] wire_d0_0;
	wire [WIDTH-1:0] wire_d0_1;
	wire [WIDTH-1:0] wire_d0_2;
	wire [WIDTH-1:0] wire_d0_3;
	wire [WIDTH-1:0] wire_d0_4;
	wire [WIDTH-1:0] wire_d0_5;
	wire [WIDTH-1:0] wire_d0_6;
	wire [WIDTH-1:0] wire_d0_7;
	wire [WIDTH-1:0] wire_d0_8;
	wire [WIDTH-1:0] wire_d0_9;
	wire [WIDTH-1:0] wire_d0_10;
	wire [WIDTH-1:0] wire_d0_11;
	wire [WIDTH-1:0] wire_d0_12;
	wire [WIDTH-1:0] wire_d0_13;
	wire [WIDTH-1:0] wire_d0_14;
	wire [WIDTH-1:0] wire_d0_15;
	wire [WIDTH-1:0] wire_d0_16;
	wire [WIDTH-1:0] wire_d0_17;
	wire [WIDTH-1:0] wire_d0_18;
	wire [WIDTH-1:0] wire_d0_19;
	wire [WIDTH-1:0] wire_d0_20;
	wire [WIDTH-1:0] wire_d0_21;
	wire [WIDTH-1:0] wire_d0_22;
	wire [WIDTH-1:0] wire_d0_23;
	wire [WIDTH-1:0] wire_d0_24;
	wire [WIDTH-1:0] wire_d0_25;
	wire [WIDTH-1:0] wire_d0_26;
	wire [WIDTH-1:0] wire_d0_27;
	wire [WIDTH-1:0] wire_d0_28;
	wire [WIDTH-1:0] wire_d0_29;
	wire [WIDTH-1:0] wire_d0_30;
	wire [WIDTH-1:0] wire_d0_31;
	wire [WIDTH-1:0] wire_d0_32;
	wire [WIDTH-1:0] wire_d0_33;
	wire [WIDTH-1:0] wire_d0_34;
	wire [WIDTH-1:0] wire_d0_35;
	wire [WIDTH-1:0] wire_d0_36;
	wire [WIDTH-1:0] wire_d0_37;
	wire [WIDTH-1:0] wire_d0_38;
	wire [WIDTH-1:0] wire_d0_39;
	wire [WIDTH-1:0] wire_d0_40;
	wire [WIDTH-1:0] wire_d0_41;
	wire [WIDTH-1:0] wire_d0_42;
	wire [WIDTH-1:0] wire_d0_43;
	wire [WIDTH-1:0] wire_d0_44;
	wire [WIDTH-1:0] wire_d0_45;
	wire [WIDTH-1:0] wire_d0_46;
	wire [WIDTH-1:0] wire_d0_47;
	wire [WIDTH-1:0] wire_d0_48;
	wire [WIDTH-1:0] wire_d0_49;
	wire [WIDTH-1:0] wire_d0_50;
	wire [WIDTH-1:0] wire_d0_51;
	wire [WIDTH-1:0] wire_d0_52;
	wire [WIDTH-1:0] wire_d0_53;
	wire [WIDTH-1:0] wire_d0_54;
	wire [WIDTH-1:0] wire_d0_55;
	wire [WIDTH-1:0] wire_d0_56;
	wire [WIDTH-1:0] wire_d0_57;
	wire [WIDTH-1:0] wire_d0_58;
	wire [WIDTH-1:0] wire_d0_59;
	wire [WIDTH-1:0] wire_d0_60;
	wire [WIDTH-1:0] wire_d0_61;
	wire [WIDTH-1:0] wire_d0_62;
	wire [WIDTH-1:0] wire_d0_63;
	wire [WIDTH-1:0] wire_d0_64;
	wire [WIDTH-1:0] wire_d0_65;
	wire [WIDTH-1:0] wire_d0_66;
	wire [WIDTH-1:0] wire_d0_67;
	wire [WIDTH-1:0] wire_d0_68;
	wire [WIDTH-1:0] wire_d1_0;
	wire [WIDTH-1:0] wire_d1_1;
	wire [WIDTH-1:0] wire_d1_2;
	wire [WIDTH-1:0] wire_d1_3;
	wire [WIDTH-1:0] wire_d1_4;
	wire [WIDTH-1:0] wire_d1_5;
	wire [WIDTH-1:0] wire_d1_6;
	wire [WIDTH-1:0] wire_d1_7;
	wire [WIDTH-1:0] wire_d1_8;
	wire [WIDTH-1:0] wire_d1_9;
	wire [WIDTH-1:0] wire_d1_10;
	wire [WIDTH-1:0] wire_d1_11;
	wire [WIDTH-1:0] wire_d1_12;
	wire [WIDTH-1:0] wire_d1_13;
	wire [WIDTH-1:0] wire_d1_14;
	wire [WIDTH-1:0] wire_d1_15;
	wire [WIDTH-1:0] wire_d1_16;
	wire [WIDTH-1:0] wire_d1_17;
	wire [WIDTH-1:0] wire_d1_18;
	wire [WIDTH-1:0] wire_d1_19;
	wire [WIDTH-1:0] wire_d1_20;
	wire [WIDTH-1:0] wire_d1_21;
	wire [WIDTH-1:0] wire_d1_22;
	wire [WIDTH-1:0] wire_d1_23;
	wire [WIDTH-1:0] wire_d1_24;
	wire [WIDTH-1:0] wire_d1_25;
	wire [WIDTH-1:0] wire_d1_26;
	wire [WIDTH-1:0] wire_d1_27;
	wire [WIDTH-1:0] wire_d1_28;
	wire [WIDTH-1:0] wire_d1_29;
	wire [WIDTH-1:0] wire_d1_30;
	wire [WIDTH-1:0] wire_d1_31;
	wire [WIDTH-1:0] wire_d1_32;
	wire [WIDTH-1:0] wire_d1_33;
	wire [WIDTH-1:0] wire_d1_34;
	wire [WIDTH-1:0] wire_d1_35;
	wire [WIDTH-1:0] wire_d1_36;
	wire [WIDTH-1:0] wire_d1_37;
	wire [WIDTH-1:0] wire_d1_38;
	wire [WIDTH-1:0] wire_d1_39;
	wire [WIDTH-1:0] wire_d1_40;
	wire [WIDTH-1:0] wire_d1_41;
	wire [WIDTH-1:0] wire_d1_42;
	wire [WIDTH-1:0] wire_d1_43;
	wire [WIDTH-1:0] wire_d1_44;
	wire [WIDTH-1:0] wire_d1_45;
	wire [WIDTH-1:0] wire_d1_46;
	wire [WIDTH-1:0] wire_d1_47;
	wire [WIDTH-1:0] wire_d1_48;
	wire [WIDTH-1:0] wire_d1_49;
	wire [WIDTH-1:0] wire_d1_50;
	wire [WIDTH-1:0] wire_d1_51;
	wire [WIDTH-1:0] wire_d1_52;
	wire [WIDTH-1:0] wire_d1_53;
	wire [WIDTH-1:0] wire_d1_54;
	wire [WIDTH-1:0] wire_d1_55;
	wire [WIDTH-1:0] wire_d1_56;
	wire [WIDTH-1:0] wire_d1_57;
	wire [WIDTH-1:0] wire_d1_58;
	wire [WIDTH-1:0] wire_d1_59;
	wire [WIDTH-1:0] wire_d1_60;
	wire [WIDTH-1:0] wire_d1_61;
	wire [WIDTH-1:0] wire_d1_62;
	wire [WIDTH-1:0] wire_d1_63;
	wire [WIDTH-1:0] wire_d1_64;
	wire [WIDTH-1:0] wire_d1_65;
	wire [WIDTH-1:0] wire_d1_66;
	wire [WIDTH-1:0] wire_d1_67;
	wire [WIDTH-1:0] wire_d1_68;
	wire [WIDTH-1:0] wire_d2_0;
	wire [WIDTH-1:0] wire_d2_1;
	wire [WIDTH-1:0] wire_d2_2;
	wire [WIDTH-1:0] wire_d2_3;
	wire [WIDTH-1:0] wire_d2_4;
	wire [WIDTH-1:0] wire_d2_5;
	wire [WIDTH-1:0] wire_d2_6;
	wire [WIDTH-1:0] wire_d2_7;
	wire [WIDTH-1:0] wire_d2_8;
	wire [WIDTH-1:0] wire_d2_9;
	wire [WIDTH-1:0] wire_d2_10;
	wire [WIDTH-1:0] wire_d2_11;
	wire [WIDTH-1:0] wire_d2_12;
	wire [WIDTH-1:0] wire_d2_13;
	wire [WIDTH-1:0] wire_d2_14;
	wire [WIDTH-1:0] wire_d2_15;
	wire [WIDTH-1:0] wire_d2_16;
	wire [WIDTH-1:0] wire_d2_17;
	wire [WIDTH-1:0] wire_d2_18;
	wire [WIDTH-1:0] wire_d2_19;
	wire [WIDTH-1:0] wire_d2_20;
	wire [WIDTH-1:0] wire_d2_21;
	wire [WIDTH-1:0] wire_d2_22;
	wire [WIDTH-1:0] wire_d2_23;
	wire [WIDTH-1:0] wire_d2_24;
	wire [WIDTH-1:0] wire_d2_25;
	wire [WIDTH-1:0] wire_d2_26;
	wire [WIDTH-1:0] wire_d2_27;
	wire [WIDTH-1:0] wire_d2_28;
	wire [WIDTH-1:0] wire_d2_29;
	wire [WIDTH-1:0] wire_d2_30;
	wire [WIDTH-1:0] wire_d2_31;
	wire [WIDTH-1:0] wire_d2_32;
	wire [WIDTH-1:0] wire_d2_33;
	wire [WIDTH-1:0] wire_d2_34;
	wire [WIDTH-1:0] wire_d2_35;
	wire [WIDTH-1:0] wire_d2_36;
	wire [WIDTH-1:0] wire_d2_37;
	wire [WIDTH-1:0] wire_d2_38;
	wire [WIDTH-1:0] wire_d2_39;
	wire [WIDTH-1:0] wire_d2_40;
	wire [WIDTH-1:0] wire_d2_41;
	wire [WIDTH-1:0] wire_d2_42;
	wire [WIDTH-1:0] wire_d2_43;
	wire [WIDTH-1:0] wire_d2_44;
	wire [WIDTH-1:0] wire_d2_45;
	wire [WIDTH-1:0] wire_d2_46;
	wire [WIDTH-1:0] wire_d2_47;
	wire [WIDTH-1:0] wire_d2_48;
	wire [WIDTH-1:0] wire_d2_49;
	wire [WIDTH-1:0] wire_d2_50;
	wire [WIDTH-1:0] wire_d2_51;
	wire [WIDTH-1:0] wire_d2_52;
	wire [WIDTH-1:0] wire_d2_53;
	wire [WIDTH-1:0] wire_d2_54;
	wire [WIDTH-1:0] wire_d2_55;
	wire [WIDTH-1:0] wire_d2_56;
	wire [WIDTH-1:0] wire_d2_57;
	wire [WIDTH-1:0] wire_d2_58;
	wire [WIDTH-1:0] wire_d2_59;
	wire [WIDTH-1:0] wire_d2_60;
	wire [WIDTH-1:0] wire_d2_61;
	wire [WIDTH-1:0] wire_d2_62;
	wire [WIDTH-1:0] wire_d2_63;
	wire [WIDTH-1:0] wire_d2_64;
	wire [WIDTH-1:0] wire_d2_65;
	wire [WIDTH-1:0] wire_d2_66;
	wire [WIDTH-1:0] wire_d2_67;
	wire [WIDTH-1:0] wire_d2_68;
	wire [WIDTH-1:0] wire_d3_0;
	wire [WIDTH-1:0] wire_d3_1;
	wire [WIDTH-1:0] wire_d3_2;
	wire [WIDTH-1:0] wire_d3_3;
	wire [WIDTH-1:0] wire_d3_4;
	wire [WIDTH-1:0] wire_d3_5;
	wire [WIDTH-1:0] wire_d3_6;
	wire [WIDTH-1:0] wire_d3_7;
	wire [WIDTH-1:0] wire_d3_8;
	wire [WIDTH-1:0] wire_d3_9;
	wire [WIDTH-1:0] wire_d3_10;
	wire [WIDTH-1:0] wire_d3_11;
	wire [WIDTH-1:0] wire_d3_12;
	wire [WIDTH-1:0] wire_d3_13;
	wire [WIDTH-1:0] wire_d3_14;
	wire [WIDTH-1:0] wire_d3_15;
	wire [WIDTH-1:0] wire_d3_16;
	wire [WIDTH-1:0] wire_d3_17;
	wire [WIDTH-1:0] wire_d3_18;
	wire [WIDTH-1:0] wire_d3_19;
	wire [WIDTH-1:0] wire_d3_20;
	wire [WIDTH-1:0] wire_d3_21;
	wire [WIDTH-1:0] wire_d3_22;
	wire [WIDTH-1:0] wire_d3_23;
	wire [WIDTH-1:0] wire_d3_24;
	wire [WIDTH-1:0] wire_d3_25;
	wire [WIDTH-1:0] wire_d3_26;
	wire [WIDTH-1:0] wire_d3_27;
	wire [WIDTH-1:0] wire_d3_28;
	wire [WIDTH-1:0] wire_d3_29;
	wire [WIDTH-1:0] wire_d3_30;
	wire [WIDTH-1:0] wire_d3_31;
	wire [WIDTH-1:0] wire_d3_32;
	wire [WIDTH-1:0] wire_d3_33;
	wire [WIDTH-1:0] wire_d3_34;
	wire [WIDTH-1:0] wire_d3_35;
	wire [WIDTH-1:0] wire_d3_36;
	wire [WIDTH-1:0] wire_d3_37;
	wire [WIDTH-1:0] wire_d3_38;
	wire [WIDTH-1:0] wire_d3_39;
	wire [WIDTH-1:0] wire_d3_40;
	wire [WIDTH-1:0] wire_d3_41;
	wire [WIDTH-1:0] wire_d3_42;
	wire [WIDTH-1:0] wire_d3_43;
	wire [WIDTH-1:0] wire_d3_44;
	wire [WIDTH-1:0] wire_d3_45;
	wire [WIDTH-1:0] wire_d3_46;
	wire [WIDTH-1:0] wire_d3_47;
	wire [WIDTH-1:0] wire_d3_48;
	wire [WIDTH-1:0] wire_d3_49;
	wire [WIDTH-1:0] wire_d3_50;
	wire [WIDTH-1:0] wire_d3_51;
	wire [WIDTH-1:0] wire_d3_52;
	wire [WIDTH-1:0] wire_d3_53;
	wire [WIDTH-1:0] wire_d3_54;
	wire [WIDTH-1:0] wire_d3_55;
	wire [WIDTH-1:0] wire_d3_56;
	wire [WIDTH-1:0] wire_d3_57;
	wire [WIDTH-1:0] wire_d3_58;
	wire [WIDTH-1:0] wire_d3_59;
	wire [WIDTH-1:0] wire_d3_60;
	wire [WIDTH-1:0] wire_d3_61;
	wire [WIDTH-1:0] wire_d3_62;
	wire [WIDTH-1:0] wire_d3_63;
	wire [WIDTH-1:0] wire_d3_64;
	wire [WIDTH-1:0] wire_d3_65;
	wire [WIDTH-1:0] wire_d3_66;
	wire [WIDTH-1:0] wire_d3_67;
	wire [WIDTH-1:0] wire_d3_68;
	wire [WIDTH-1:0] wire_d4_0;
	wire [WIDTH-1:0] wire_d4_1;
	wire [WIDTH-1:0] wire_d4_2;
	wire [WIDTH-1:0] wire_d4_3;
	wire [WIDTH-1:0] wire_d4_4;
	wire [WIDTH-1:0] wire_d4_5;
	wire [WIDTH-1:0] wire_d4_6;
	wire [WIDTH-1:0] wire_d4_7;
	wire [WIDTH-1:0] wire_d4_8;
	wire [WIDTH-1:0] wire_d4_9;
	wire [WIDTH-1:0] wire_d4_10;
	wire [WIDTH-1:0] wire_d4_11;
	wire [WIDTH-1:0] wire_d4_12;
	wire [WIDTH-1:0] wire_d4_13;
	wire [WIDTH-1:0] wire_d4_14;
	wire [WIDTH-1:0] wire_d4_15;
	wire [WIDTH-1:0] wire_d4_16;
	wire [WIDTH-1:0] wire_d4_17;
	wire [WIDTH-1:0] wire_d4_18;
	wire [WIDTH-1:0] wire_d4_19;
	wire [WIDTH-1:0] wire_d4_20;
	wire [WIDTH-1:0] wire_d4_21;
	wire [WIDTH-1:0] wire_d4_22;
	wire [WIDTH-1:0] wire_d4_23;
	wire [WIDTH-1:0] wire_d4_24;
	wire [WIDTH-1:0] wire_d4_25;
	wire [WIDTH-1:0] wire_d4_26;
	wire [WIDTH-1:0] wire_d4_27;
	wire [WIDTH-1:0] wire_d4_28;
	wire [WIDTH-1:0] wire_d4_29;
	wire [WIDTH-1:0] wire_d4_30;
	wire [WIDTH-1:0] wire_d4_31;
	wire [WIDTH-1:0] wire_d4_32;
	wire [WIDTH-1:0] wire_d4_33;
	wire [WIDTH-1:0] wire_d4_34;
	wire [WIDTH-1:0] wire_d4_35;
	wire [WIDTH-1:0] wire_d4_36;
	wire [WIDTH-1:0] wire_d4_37;
	wire [WIDTH-1:0] wire_d4_38;
	wire [WIDTH-1:0] wire_d4_39;
	wire [WIDTH-1:0] wire_d4_40;
	wire [WIDTH-1:0] wire_d4_41;
	wire [WIDTH-1:0] wire_d4_42;
	wire [WIDTH-1:0] wire_d4_43;
	wire [WIDTH-1:0] wire_d4_44;
	wire [WIDTH-1:0] wire_d4_45;
	wire [WIDTH-1:0] wire_d4_46;
	wire [WIDTH-1:0] wire_d4_47;
	wire [WIDTH-1:0] wire_d4_48;
	wire [WIDTH-1:0] wire_d4_49;
	wire [WIDTH-1:0] wire_d4_50;
	wire [WIDTH-1:0] wire_d4_51;
	wire [WIDTH-1:0] wire_d4_52;
	wire [WIDTH-1:0] wire_d4_53;
	wire [WIDTH-1:0] wire_d4_54;
	wire [WIDTH-1:0] wire_d4_55;
	wire [WIDTH-1:0] wire_d4_56;
	wire [WIDTH-1:0] wire_d4_57;
	wire [WIDTH-1:0] wire_d4_58;
	wire [WIDTH-1:0] wire_d4_59;
	wire [WIDTH-1:0] wire_d4_60;
	wire [WIDTH-1:0] wire_d4_61;
	wire [WIDTH-1:0] wire_d4_62;
	wire [WIDTH-1:0] wire_d4_63;
	wire [WIDTH-1:0] wire_d4_64;
	wire [WIDTH-1:0] wire_d4_65;
	wire [WIDTH-1:0] wire_d4_66;
	wire [WIDTH-1:0] wire_d4_67;
	wire [WIDTH-1:0] wire_d4_68;
	wire [WIDTH-1:0] wire_d5_0;
	wire [WIDTH-1:0] wire_d5_1;
	wire [WIDTH-1:0] wire_d5_2;
	wire [WIDTH-1:0] wire_d5_3;
	wire [WIDTH-1:0] wire_d5_4;
	wire [WIDTH-1:0] wire_d5_5;
	wire [WIDTH-1:0] wire_d5_6;
	wire [WIDTH-1:0] wire_d5_7;
	wire [WIDTH-1:0] wire_d5_8;
	wire [WIDTH-1:0] wire_d5_9;
	wire [WIDTH-1:0] wire_d5_10;
	wire [WIDTH-1:0] wire_d5_11;
	wire [WIDTH-1:0] wire_d5_12;
	wire [WIDTH-1:0] wire_d5_13;
	wire [WIDTH-1:0] wire_d5_14;
	wire [WIDTH-1:0] wire_d5_15;
	wire [WIDTH-1:0] wire_d5_16;
	wire [WIDTH-1:0] wire_d5_17;
	wire [WIDTH-1:0] wire_d5_18;
	wire [WIDTH-1:0] wire_d5_19;
	wire [WIDTH-1:0] wire_d5_20;
	wire [WIDTH-1:0] wire_d5_21;
	wire [WIDTH-1:0] wire_d5_22;
	wire [WIDTH-1:0] wire_d5_23;
	wire [WIDTH-1:0] wire_d5_24;
	wire [WIDTH-1:0] wire_d5_25;
	wire [WIDTH-1:0] wire_d5_26;
	wire [WIDTH-1:0] wire_d5_27;
	wire [WIDTH-1:0] wire_d5_28;
	wire [WIDTH-1:0] wire_d5_29;
	wire [WIDTH-1:0] wire_d5_30;
	wire [WIDTH-1:0] wire_d5_31;
	wire [WIDTH-1:0] wire_d5_32;
	wire [WIDTH-1:0] wire_d5_33;
	wire [WIDTH-1:0] wire_d5_34;
	wire [WIDTH-1:0] wire_d5_35;
	wire [WIDTH-1:0] wire_d5_36;
	wire [WIDTH-1:0] wire_d5_37;
	wire [WIDTH-1:0] wire_d5_38;
	wire [WIDTH-1:0] wire_d5_39;
	wire [WIDTH-1:0] wire_d5_40;
	wire [WIDTH-1:0] wire_d5_41;
	wire [WIDTH-1:0] wire_d5_42;
	wire [WIDTH-1:0] wire_d5_43;
	wire [WIDTH-1:0] wire_d5_44;
	wire [WIDTH-1:0] wire_d5_45;
	wire [WIDTH-1:0] wire_d5_46;
	wire [WIDTH-1:0] wire_d5_47;
	wire [WIDTH-1:0] wire_d5_48;
	wire [WIDTH-1:0] wire_d5_49;
	wire [WIDTH-1:0] wire_d5_50;
	wire [WIDTH-1:0] wire_d5_51;
	wire [WIDTH-1:0] wire_d5_52;
	wire [WIDTH-1:0] wire_d5_53;
	wire [WIDTH-1:0] wire_d5_54;
	wire [WIDTH-1:0] wire_d5_55;
	wire [WIDTH-1:0] wire_d5_56;
	wire [WIDTH-1:0] wire_d5_57;
	wire [WIDTH-1:0] wire_d5_58;
	wire [WIDTH-1:0] wire_d5_59;
	wire [WIDTH-1:0] wire_d5_60;
	wire [WIDTH-1:0] wire_d5_61;
	wire [WIDTH-1:0] wire_d5_62;
	wire [WIDTH-1:0] wire_d5_63;
	wire [WIDTH-1:0] wire_d5_64;
	wire [WIDTH-1:0] wire_d5_65;
	wire [WIDTH-1:0] wire_d5_66;
	wire [WIDTH-1:0] wire_d5_67;
	wire [WIDTH-1:0] wire_d5_68;
	wire [WIDTH-1:0] wire_d6_0;
	wire [WIDTH-1:0] wire_d6_1;
	wire [WIDTH-1:0] wire_d6_2;
	wire [WIDTH-1:0] wire_d6_3;
	wire [WIDTH-1:0] wire_d6_4;
	wire [WIDTH-1:0] wire_d6_5;
	wire [WIDTH-1:0] wire_d6_6;
	wire [WIDTH-1:0] wire_d6_7;
	wire [WIDTH-1:0] wire_d6_8;
	wire [WIDTH-1:0] wire_d6_9;
	wire [WIDTH-1:0] wire_d6_10;
	wire [WIDTH-1:0] wire_d6_11;
	wire [WIDTH-1:0] wire_d6_12;
	wire [WIDTH-1:0] wire_d6_13;
	wire [WIDTH-1:0] wire_d6_14;
	wire [WIDTH-1:0] wire_d6_15;
	wire [WIDTH-1:0] wire_d6_16;
	wire [WIDTH-1:0] wire_d6_17;
	wire [WIDTH-1:0] wire_d6_18;
	wire [WIDTH-1:0] wire_d6_19;
	wire [WIDTH-1:0] wire_d6_20;
	wire [WIDTH-1:0] wire_d6_21;
	wire [WIDTH-1:0] wire_d6_22;
	wire [WIDTH-1:0] wire_d6_23;
	wire [WIDTH-1:0] wire_d6_24;
	wire [WIDTH-1:0] wire_d6_25;
	wire [WIDTH-1:0] wire_d6_26;
	wire [WIDTH-1:0] wire_d6_27;
	wire [WIDTH-1:0] wire_d6_28;
	wire [WIDTH-1:0] wire_d6_29;
	wire [WIDTH-1:0] wire_d6_30;
	wire [WIDTH-1:0] wire_d6_31;
	wire [WIDTH-1:0] wire_d6_32;
	wire [WIDTH-1:0] wire_d6_33;
	wire [WIDTH-1:0] wire_d6_34;
	wire [WIDTH-1:0] wire_d6_35;
	wire [WIDTH-1:0] wire_d6_36;
	wire [WIDTH-1:0] wire_d6_37;
	wire [WIDTH-1:0] wire_d6_38;
	wire [WIDTH-1:0] wire_d6_39;
	wire [WIDTH-1:0] wire_d6_40;
	wire [WIDTH-1:0] wire_d6_41;
	wire [WIDTH-1:0] wire_d6_42;
	wire [WIDTH-1:0] wire_d6_43;
	wire [WIDTH-1:0] wire_d6_44;
	wire [WIDTH-1:0] wire_d6_45;
	wire [WIDTH-1:0] wire_d6_46;
	wire [WIDTH-1:0] wire_d6_47;
	wire [WIDTH-1:0] wire_d6_48;
	wire [WIDTH-1:0] wire_d6_49;
	wire [WIDTH-1:0] wire_d6_50;
	wire [WIDTH-1:0] wire_d6_51;
	wire [WIDTH-1:0] wire_d6_52;
	wire [WIDTH-1:0] wire_d6_53;
	wire [WIDTH-1:0] wire_d6_54;
	wire [WIDTH-1:0] wire_d6_55;
	wire [WIDTH-1:0] wire_d6_56;
	wire [WIDTH-1:0] wire_d6_57;
	wire [WIDTH-1:0] wire_d6_58;
	wire [WIDTH-1:0] wire_d6_59;
	wire [WIDTH-1:0] wire_d6_60;
	wire [WIDTH-1:0] wire_d6_61;
	wire [WIDTH-1:0] wire_d6_62;
	wire [WIDTH-1:0] wire_d6_63;
	wire [WIDTH-1:0] wire_d6_64;
	wire [WIDTH-1:0] wire_d6_65;
	wire [WIDTH-1:0] wire_d6_66;
	wire [WIDTH-1:0] wire_d6_67;
	wire [WIDTH-1:0] wire_d6_68;
	wire [WIDTH-1:0] wire_d7_0;
	wire [WIDTH-1:0] wire_d7_1;
	wire [WIDTH-1:0] wire_d7_2;
	wire [WIDTH-1:0] wire_d7_3;
	wire [WIDTH-1:0] wire_d7_4;
	wire [WIDTH-1:0] wire_d7_5;
	wire [WIDTH-1:0] wire_d7_6;
	wire [WIDTH-1:0] wire_d7_7;
	wire [WIDTH-1:0] wire_d7_8;
	wire [WIDTH-1:0] wire_d7_9;
	wire [WIDTH-1:0] wire_d7_10;
	wire [WIDTH-1:0] wire_d7_11;
	wire [WIDTH-1:0] wire_d7_12;
	wire [WIDTH-1:0] wire_d7_13;
	wire [WIDTH-1:0] wire_d7_14;
	wire [WIDTH-1:0] wire_d7_15;
	wire [WIDTH-1:0] wire_d7_16;
	wire [WIDTH-1:0] wire_d7_17;
	wire [WIDTH-1:0] wire_d7_18;
	wire [WIDTH-1:0] wire_d7_19;
	wire [WIDTH-1:0] wire_d7_20;
	wire [WIDTH-1:0] wire_d7_21;
	wire [WIDTH-1:0] wire_d7_22;
	wire [WIDTH-1:0] wire_d7_23;
	wire [WIDTH-1:0] wire_d7_24;
	wire [WIDTH-1:0] wire_d7_25;
	wire [WIDTH-1:0] wire_d7_26;
	wire [WIDTH-1:0] wire_d7_27;
	wire [WIDTH-1:0] wire_d7_28;
	wire [WIDTH-1:0] wire_d7_29;
	wire [WIDTH-1:0] wire_d7_30;
	wire [WIDTH-1:0] wire_d7_31;
	wire [WIDTH-1:0] wire_d7_32;
	wire [WIDTH-1:0] wire_d7_33;
	wire [WIDTH-1:0] wire_d7_34;
	wire [WIDTH-1:0] wire_d7_35;
	wire [WIDTH-1:0] wire_d7_36;
	wire [WIDTH-1:0] wire_d7_37;
	wire [WIDTH-1:0] wire_d7_38;
	wire [WIDTH-1:0] wire_d7_39;
	wire [WIDTH-1:0] wire_d7_40;
	wire [WIDTH-1:0] wire_d7_41;
	wire [WIDTH-1:0] wire_d7_42;
	wire [WIDTH-1:0] wire_d7_43;
	wire [WIDTH-1:0] wire_d7_44;
	wire [WIDTH-1:0] wire_d7_45;
	wire [WIDTH-1:0] wire_d7_46;
	wire [WIDTH-1:0] wire_d7_47;
	wire [WIDTH-1:0] wire_d7_48;
	wire [WIDTH-1:0] wire_d7_49;
	wire [WIDTH-1:0] wire_d7_50;
	wire [WIDTH-1:0] wire_d7_51;
	wire [WIDTH-1:0] wire_d7_52;
	wire [WIDTH-1:0] wire_d7_53;
	wire [WIDTH-1:0] wire_d7_54;
	wire [WIDTH-1:0] wire_d7_55;
	wire [WIDTH-1:0] wire_d7_56;
	wire [WIDTH-1:0] wire_d7_57;
	wire [WIDTH-1:0] wire_d7_58;
	wire [WIDTH-1:0] wire_d7_59;
	wire [WIDTH-1:0] wire_d7_60;
	wire [WIDTH-1:0] wire_d7_61;
	wire [WIDTH-1:0] wire_d7_62;
	wire [WIDTH-1:0] wire_d7_63;
	wire [WIDTH-1:0] wire_d7_64;
	wire [WIDTH-1:0] wire_d7_65;
	wire [WIDTH-1:0] wire_d7_66;
	wire [WIDTH-1:0] wire_d7_67;
	wire [WIDTH-1:0] wire_d7_68;
	wire [WIDTH-1:0] wire_d8_0;
	wire [WIDTH-1:0] wire_d8_1;
	wire [WIDTH-1:0] wire_d8_2;
	wire [WIDTH-1:0] wire_d8_3;
	wire [WIDTH-1:0] wire_d8_4;
	wire [WIDTH-1:0] wire_d8_5;
	wire [WIDTH-1:0] wire_d8_6;
	wire [WIDTH-1:0] wire_d8_7;
	wire [WIDTH-1:0] wire_d8_8;
	wire [WIDTH-1:0] wire_d8_9;
	wire [WIDTH-1:0] wire_d8_10;
	wire [WIDTH-1:0] wire_d8_11;
	wire [WIDTH-1:0] wire_d8_12;
	wire [WIDTH-1:0] wire_d8_13;
	wire [WIDTH-1:0] wire_d8_14;
	wire [WIDTH-1:0] wire_d8_15;
	wire [WIDTH-1:0] wire_d8_16;
	wire [WIDTH-1:0] wire_d8_17;
	wire [WIDTH-1:0] wire_d8_18;
	wire [WIDTH-1:0] wire_d8_19;
	wire [WIDTH-1:0] wire_d8_20;
	wire [WIDTH-1:0] wire_d8_21;
	wire [WIDTH-1:0] wire_d8_22;
	wire [WIDTH-1:0] wire_d8_23;
	wire [WIDTH-1:0] wire_d8_24;
	wire [WIDTH-1:0] wire_d8_25;
	wire [WIDTH-1:0] wire_d8_26;
	wire [WIDTH-1:0] wire_d8_27;
	wire [WIDTH-1:0] wire_d8_28;
	wire [WIDTH-1:0] wire_d8_29;
	wire [WIDTH-1:0] wire_d8_30;
	wire [WIDTH-1:0] wire_d8_31;
	wire [WIDTH-1:0] wire_d8_32;
	wire [WIDTH-1:0] wire_d8_33;
	wire [WIDTH-1:0] wire_d8_34;
	wire [WIDTH-1:0] wire_d8_35;
	wire [WIDTH-1:0] wire_d8_36;
	wire [WIDTH-1:0] wire_d8_37;
	wire [WIDTH-1:0] wire_d8_38;
	wire [WIDTH-1:0] wire_d8_39;
	wire [WIDTH-1:0] wire_d8_40;
	wire [WIDTH-1:0] wire_d8_41;
	wire [WIDTH-1:0] wire_d8_42;
	wire [WIDTH-1:0] wire_d8_43;
	wire [WIDTH-1:0] wire_d8_44;
	wire [WIDTH-1:0] wire_d8_45;
	wire [WIDTH-1:0] wire_d8_46;
	wire [WIDTH-1:0] wire_d8_47;
	wire [WIDTH-1:0] wire_d8_48;
	wire [WIDTH-1:0] wire_d8_49;
	wire [WIDTH-1:0] wire_d8_50;
	wire [WIDTH-1:0] wire_d8_51;
	wire [WIDTH-1:0] wire_d8_52;
	wire [WIDTH-1:0] wire_d8_53;
	wire [WIDTH-1:0] wire_d8_54;
	wire [WIDTH-1:0] wire_d8_55;
	wire [WIDTH-1:0] wire_d8_56;
	wire [WIDTH-1:0] wire_d8_57;
	wire [WIDTH-1:0] wire_d8_58;
	wire [WIDTH-1:0] wire_d8_59;
	wire [WIDTH-1:0] wire_d8_60;
	wire [WIDTH-1:0] wire_d8_61;
	wire [WIDTH-1:0] wire_d8_62;
	wire [WIDTH-1:0] wire_d8_63;
	wire [WIDTH-1:0] wire_d8_64;
	wire [WIDTH-1:0] wire_d8_65;
	wire [WIDTH-1:0] wire_d8_66;
	wire [WIDTH-1:0] wire_d8_67;
	wire [WIDTH-1:0] wire_d8_68;
	wire [WIDTH-1:0] wire_d9_0;
	wire [WIDTH-1:0] wire_d9_1;
	wire [WIDTH-1:0] wire_d9_2;
	wire [WIDTH-1:0] wire_d9_3;
	wire [WIDTH-1:0] wire_d9_4;
	wire [WIDTH-1:0] wire_d9_5;
	wire [WIDTH-1:0] wire_d9_6;
	wire [WIDTH-1:0] wire_d9_7;
	wire [WIDTH-1:0] wire_d9_8;
	wire [WIDTH-1:0] wire_d9_9;
	wire [WIDTH-1:0] wire_d9_10;
	wire [WIDTH-1:0] wire_d9_11;
	wire [WIDTH-1:0] wire_d9_12;
	wire [WIDTH-1:0] wire_d9_13;
	wire [WIDTH-1:0] wire_d9_14;
	wire [WIDTH-1:0] wire_d9_15;
	wire [WIDTH-1:0] wire_d9_16;
	wire [WIDTH-1:0] wire_d9_17;
	wire [WIDTH-1:0] wire_d9_18;
	wire [WIDTH-1:0] wire_d9_19;
	wire [WIDTH-1:0] wire_d9_20;
	wire [WIDTH-1:0] wire_d9_21;
	wire [WIDTH-1:0] wire_d9_22;
	wire [WIDTH-1:0] wire_d9_23;
	wire [WIDTH-1:0] wire_d9_24;
	wire [WIDTH-1:0] wire_d9_25;
	wire [WIDTH-1:0] wire_d9_26;
	wire [WIDTH-1:0] wire_d9_27;
	wire [WIDTH-1:0] wire_d9_28;
	wire [WIDTH-1:0] wire_d9_29;
	wire [WIDTH-1:0] wire_d9_30;
	wire [WIDTH-1:0] wire_d9_31;
	wire [WIDTH-1:0] wire_d9_32;
	wire [WIDTH-1:0] wire_d9_33;
	wire [WIDTH-1:0] wire_d9_34;
	wire [WIDTH-1:0] wire_d9_35;
	wire [WIDTH-1:0] wire_d9_36;
	wire [WIDTH-1:0] wire_d9_37;
	wire [WIDTH-1:0] wire_d9_38;
	wire [WIDTH-1:0] wire_d9_39;
	wire [WIDTH-1:0] wire_d9_40;
	wire [WIDTH-1:0] wire_d9_41;
	wire [WIDTH-1:0] wire_d9_42;
	wire [WIDTH-1:0] wire_d9_43;
	wire [WIDTH-1:0] wire_d9_44;
	wire [WIDTH-1:0] wire_d9_45;
	wire [WIDTH-1:0] wire_d9_46;
	wire [WIDTH-1:0] wire_d9_47;
	wire [WIDTH-1:0] wire_d9_48;
	wire [WIDTH-1:0] wire_d9_49;
	wire [WIDTH-1:0] wire_d9_50;
	wire [WIDTH-1:0] wire_d9_51;
	wire [WIDTH-1:0] wire_d9_52;
	wire [WIDTH-1:0] wire_d9_53;
	wire [WIDTH-1:0] wire_d9_54;
	wire [WIDTH-1:0] wire_d9_55;
	wire [WIDTH-1:0] wire_d9_56;
	wire [WIDTH-1:0] wire_d9_57;
	wire [WIDTH-1:0] wire_d9_58;
	wire [WIDTH-1:0] wire_d9_59;
	wire [WIDTH-1:0] wire_d9_60;
	wire [WIDTH-1:0] wire_d9_61;
	wire [WIDTH-1:0] wire_d9_62;
	wire [WIDTH-1:0] wire_d9_63;
	wire [WIDTH-1:0] wire_d9_64;
	wire [WIDTH-1:0] wire_d9_65;
	wire [WIDTH-1:0] wire_d9_66;
	wire [WIDTH-1:0] wire_d9_67;
	wire [WIDTH-1:0] wire_d9_68;
	wire [WIDTH-1:0] wire_d10_0;
	wire [WIDTH-1:0] wire_d10_1;
	wire [WIDTH-1:0] wire_d10_2;
	wire [WIDTH-1:0] wire_d10_3;
	wire [WIDTH-1:0] wire_d10_4;
	wire [WIDTH-1:0] wire_d10_5;
	wire [WIDTH-1:0] wire_d10_6;
	wire [WIDTH-1:0] wire_d10_7;
	wire [WIDTH-1:0] wire_d10_8;
	wire [WIDTH-1:0] wire_d10_9;
	wire [WIDTH-1:0] wire_d10_10;
	wire [WIDTH-1:0] wire_d10_11;
	wire [WIDTH-1:0] wire_d10_12;
	wire [WIDTH-1:0] wire_d10_13;
	wire [WIDTH-1:0] wire_d10_14;
	wire [WIDTH-1:0] wire_d10_15;
	wire [WIDTH-1:0] wire_d10_16;
	wire [WIDTH-1:0] wire_d10_17;
	wire [WIDTH-1:0] wire_d10_18;
	wire [WIDTH-1:0] wire_d10_19;
	wire [WIDTH-1:0] wire_d10_20;
	wire [WIDTH-1:0] wire_d10_21;
	wire [WIDTH-1:0] wire_d10_22;
	wire [WIDTH-1:0] wire_d10_23;
	wire [WIDTH-1:0] wire_d10_24;
	wire [WIDTH-1:0] wire_d10_25;
	wire [WIDTH-1:0] wire_d10_26;
	wire [WIDTH-1:0] wire_d10_27;
	wire [WIDTH-1:0] wire_d10_28;
	wire [WIDTH-1:0] wire_d10_29;
	wire [WIDTH-1:0] wire_d10_30;
	wire [WIDTH-1:0] wire_d10_31;
	wire [WIDTH-1:0] wire_d10_32;
	wire [WIDTH-1:0] wire_d10_33;
	wire [WIDTH-1:0] wire_d10_34;
	wire [WIDTH-1:0] wire_d10_35;
	wire [WIDTH-1:0] wire_d10_36;
	wire [WIDTH-1:0] wire_d10_37;
	wire [WIDTH-1:0] wire_d10_38;
	wire [WIDTH-1:0] wire_d10_39;
	wire [WIDTH-1:0] wire_d10_40;
	wire [WIDTH-1:0] wire_d10_41;
	wire [WIDTH-1:0] wire_d10_42;
	wire [WIDTH-1:0] wire_d10_43;
	wire [WIDTH-1:0] wire_d10_44;
	wire [WIDTH-1:0] wire_d10_45;
	wire [WIDTH-1:0] wire_d10_46;
	wire [WIDTH-1:0] wire_d10_47;
	wire [WIDTH-1:0] wire_d10_48;
	wire [WIDTH-1:0] wire_d10_49;
	wire [WIDTH-1:0] wire_d10_50;
	wire [WIDTH-1:0] wire_d10_51;
	wire [WIDTH-1:0] wire_d10_52;
	wire [WIDTH-1:0] wire_d10_53;
	wire [WIDTH-1:0] wire_d10_54;
	wire [WIDTH-1:0] wire_d10_55;
	wire [WIDTH-1:0] wire_d10_56;
	wire [WIDTH-1:0] wire_d10_57;
	wire [WIDTH-1:0] wire_d10_58;
	wire [WIDTH-1:0] wire_d10_59;
	wire [WIDTH-1:0] wire_d10_60;
	wire [WIDTH-1:0] wire_d10_61;
	wire [WIDTH-1:0] wire_d10_62;
	wire [WIDTH-1:0] wire_d10_63;
	wire [WIDTH-1:0] wire_d10_64;
	wire [WIDTH-1:0] wire_d10_65;
	wire [WIDTH-1:0] wire_d10_66;
	wire [WIDTH-1:0] wire_d10_67;
	wire [WIDTH-1:0] wire_d10_68;
	wire [WIDTH-1:0] wire_d11_0;
	wire [WIDTH-1:0] wire_d11_1;
	wire [WIDTH-1:0] wire_d11_2;
	wire [WIDTH-1:0] wire_d11_3;
	wire [WIDTH-1:0] wire_d11_4;
	wire [WIDTH-1:0] wire_d11_5;
	wire [WIDTH-1:0] wire_d11_6;
	wire [WIDTH-1:0] wire_d11_7;
	wire [WIDTH-1:0] wire_d11_8;
	wire [WIDTH-1:0] wire_d11_9;
	wire [WIDTH-1:0] wire_d11_10;
	wire [WIDTH-1:0] wire_d11_11;
	wire [WIDTH-1:0] wire_d11_12;
	wire [WIDTH-1:0] wire_d11_13;
	wire [WIDTH-1:0] wire_d11_14;
	wire [WIDTH-1:0] wire_d11_15;
	wire [WIDTH-1:0] wire_d11_16;
	wire [WIDTH-1:0] wire_d11_17;
	wire [WIDTH-1:0] wire_d11_18;
	wire [WIDTH-1:0] wire_d11_19;
	wire [WIDTH-1:0] wire_d11_20;
	wire [WIDTH-1:0] wire_d11_21;
	wire [WIDTH-1:0] wire_d11_22;
	wire [WIDTH-1:0] wire_d11_23;
	wire [WIDTH-1:0] wire_d11_24;
	wire [WIDTH-1:0] wire_d11_25;
	wire [WIDTH-1:0] wire_d11_26;
	wire [WIDTH-1:0] wire_d11_27;
	wire [WIDTH-1:0] wire_d11_28;
	wire [WIDTH-1:0] wire_d11_29;
	wire [WIDTH-1:0] wire_d11_30;
	wire [WIDTH-1:0] wire_d11_31;
	wire [WIDTH-1:0] wire_d11_32;
	wire [WIDTH-1:0] wire_d11_33;
	wire [WIDTH-1:0] wire_d11_34;
	wire [WIDTH-1:0] wire_d11_35;
	wire [WIDTH-1:0] wire_d11_36;
	wire [WIDTH-1:0] wire_d11_37;
	wire [WIDTH-1:0] wire_d11_38;
	wire [WIDTH-1:0] wire_d11_39;
	wire [WIDTH-1:0] wire_d11_40;
	wire [WIDTH-1:0] wire_d11_41;
	wire [WIDTH-1:0] wire_d11_42;
	wire [WIDTH-1:0] wire_d11_43;
	wire [WIDTH-1:0] wire_d11_44;
	wire [WIDTH-1:0] wire_d11_45;
	wire [WIDTH-1:0] wire_d11_46;
	wire [WIDTH-1:0] wire_d11_47;
	wire [WIDTH-1:0] wire_d11_48;
	wire [WIDTH-1:0] wire_d11_49;
	wire [WIDTH-1:0] wire_d11_50;
	wire [WIDTH-1:0] wire_d11_51;
	wire [WIDTH-1:0] wire_d11_52;
	wire [WIDTH-1:0] wire_d11_53;
	wire [WIDTH-1:0] wire_d11_54;
	wire [WIDTH-1:0] wire_d11_55;
	wire [WIDTH-1:0] wire_d11_56;
	wire [WIDTH-1:0] wire_d11_57;
	wire [WIDTH-1:0] wire_d11_58;
	wire [WIDTH-1:0] wire_d11_59;
	wire [WIDTH-1:0] wire_d11_60;
	wire [WIDTH-1:0] wire_d11_61;
	wire [WIDTH-1:0] wire_d11_62;
	wire [WIDTH-1:0] wire_d11_63;
	wire [WIDTH-1:0] wire_d11_64;
	wire [WIDTH-1:0] wire_d11_65;
	wire [WIDTH-1:0] wire_d11_66;
	wire [WIDTH-1:0] wire_d11_67;
	wire [WIDTH-1:0] wire_d11_68;
	wire [WIDTH-1:0] wire_d12_0;
	wire [WIDTH-1:0] wire_d12_1;
	wire [WIDTH-1:0] wire_d12_2;
	wire [WIDTH-1:0] wire_d12_3;
	wire [WIDTH-1:0] wire_d12_4;
	wire [WIDTH-1:0] wire_d12_5;
	wire [WIDTH-1:0] wire_d12_6;
	wire [WIDTH-1:0] wire_d12_7;
	wire [WIDTH-1:0] wire_d12_8;
	wire [WIDTH-1:0] wire_d12_9;
	wire [WIDTH-1:0] wire_d12_10;
	wire [WIDTH-1:0] wire_d12_11;
	wire [WIDTH-1:0] wire_d12_12;
	wire [WIDTH-1:0] wire_d12_13;
	wire [WIDTH-1:0] wire_d12_14;
	wire [WIDTH-1:0] wire_d12_15;
	wire [WIDTH-1:0] wire_d12_16;
	wire [WIDTH-1:0] wire_d12_17;
	wire [WIDTH-1:0] wire_d12_18;
	wire [WIDTH-1:0] wire_d12_19;
	wire [WIDTH-1:0] wire_d12_20;
	wire [WIDTH-1:0] wire_d12_21;
	wire [WIDTH-1:0] wire_d12_22;
	wire [WIDTH-1:0] wire_d12_23;
	wire [WIDTH-1:0] wire_d12_24;
	wire [WIDTH-1:0] wire_d12_25;
	wire [WIDTH-1:0] wire_d12_26;
	wire [WIDTH-1:0] wire_d12_27;
	wire [WIDTH-1:0] wire_d12_28;
	wire [WIDTH-1:0] wire_d12_29;
	wire [WIDTH-1:0] wire_d12_30;
	wire [WIDTH-1:0] wire_d12_31;
	wire [WIDTH-1:0] wire_d12_32;
	wire [WIDTH-1:0] wire_d12_33;
	wire [WIDTH-1:0] wire_d12_34;
	wire [WIDTH-1:0] wire_d12_35;
	wire [WIDTH-1:0] wire_d12_36;
	wire [WIDTH-1:0] wire_d12_37;
	wire [WIDTH-1:0] wire_d12_38;
	wire [WIDTH-1:0] wire_d12_39;
	wire [WIDTH-1:0] wire_d12_40;
	wire [WIDTH-1:0] wire_d12_41;
	wire [WIDTH-1:0] wire_d12_42;
	wire [WIDTH-1:0] wire_d12_43;
	wire [WIDTH-1:0] wire_d12_44;
	wire [WIDTH-1:0] wire_d12_45;
	wire [WIDTH-1:0] wire_d12_46;
	wire [WIDTH-1:0] wire_d12_47;
	wire [WIDTH-1:0] wire_d12_48;
	wire [WIDTH-1:0] wire_d12_49;
	wire [WIDTH-1:0] wire_d12_50;
	wire [WIDTH-1:0] wire_d12_51;
	wire [WIDTH-1:0] wire_d12_52;
	wire [WIDTH-1:0] wire_d12_53;
	wire [WIDTH-1:0] wire_d12_54;
	wire [WIDTH-1:0] wire_d12_55;
	wire [WIDTH-1:0] wire_d12_56;
	wire [WIDTH-1:0] wire_d12_57;
	wire [WIDTH-1:0] wire_d12_58;
	wire [WIDTH-1:0] wire_d12_59;
	wire [WIDTH-1:0] wire_d12_60;
	wire [WIDTH-1:0] wire_d12_61;
	wire [WIDTH-1:0] wire_d12_62;
	wire [WIDTH-1:0] wire_d12_63;
	wire [WIDTH-1:0] wire_d12_64;
	wire [WIDTH-1:0] wire_d12_65;
	wire [WIDTH-1:0] wire_d12_66;
	wire [WIDTH-1:0] wire_d12_67;
	wire [WIDTH-1:0] wire_d12_68;
	wire [WIDTH-1:0] wire_d13_0;
	wire [WIDTH-1:0] wire_d13_1;
	wire [WIDTH-1:0] wire_d13_2;
	wire [WIDTH-1:0] wire_d13_3;
	wire [WIDTH-1:0] wire_d13_4;
	wire [WIDTH-1:0] wire_d13_5;
	wire [WIDTH-1:0] wire_d13_6;
	wire [WIDTH-1:0] wire_d13_7;
	wire [WIDTH-1:0] wire_d13_8;
	wire [WIDTH-1:0] wire_d13_9;
	wire [WIDTH-1:0] wire_d13_10;
	wire [WIDTH-1:0] wire_d13_11;
	wire [WIDTH-1:0] wire_d13_12;
	wire [WIDTH-1:0] wire_d13_13;
	wire [WIDTH-1:0] wire_d13_14;
	wire [WIDTH-1:0] wire_d13_15;
	wire [WIDTH-1:0] wire_d13_16;
	wire [WIDTH-1:0] wire_d13_17;
	wire [WIDTH-1:0] wire_d13_18;
	wire [WIDTH-1:0] wire_d13_19;
	wire [WIDTH-1:0] wire_d13_20;
	wire [WIDTH-1:0] wire_d13_21;
	wire [WIDTH-1:0] wire_d13_22;
	wire [WIDTH-1:0] wire_d13_23;
	wire [WIDTH-1:0] wire_d13_24;
	wire [WIDTH-1:0] wire_d13_25;
	wire [WIDTH-1:0] wire_d13_26;
	wire [WIDTH-1:0] wire_d13_27;
	wire [WIDTH-1:0] wire_d13_28;
	wire [WIDTH-1:0] wire_d13_29;
	wire [WIDTH-1:0] wire_d13_30;
	wire [WIDTH-1:0] wire_d13_31;
	wire [WIDTH-1:0] wire_d13_32;
	wire [WIDTH-1:0] wire_d13_33;
	wire [WIDTH-1:0] wire_d13_34;
	wire [WIDTH-1:0] wire_d13_35;
	wire [WIDTH-1:0] wire_d13_36;
	wire [WIDTH-1:0] wire_d13_37;
	wire [WIDTH-1:0] wire_d13_38;
	wire [WIDTH-1:0] wire_d13_39;
	wire [WIDTH-1:0] wire_d13_40;
	wire [WIDTH-1:0] wire_d13_41;
	wire [WIDTH-1:0] wire_d13_42;
	wire [WIDTH-1:0] wire_d13_43;
	wire [WIDTH-1:0] wire_d13_44;
	wire [WIDTH-1:0] wire_d13_45;
	wire [WIDTH-1:0] wire_d13_46;
	wire [WIDTH-1:0] wire_d13_47;
	wire [WIDTH-1:0] wire_d13_48;
	wire [WIDTH-1:0] wire_d13_49;
	wire [WIDTH-1:0] wire_d13_50;
	wire [WIDTH-1:0] wire_d13_51;
	wire [WIDTH-1:0] wire_d13_52;
	wire [WIDTH-1:0] wire_d13_53;
	wire [WIDTH-1:0] wire_d13_54;
	wire [WIDTH-1:0] wire_d13_55;
	wire [WIDTH-1:0] wire_d13_56;
	wire [WIDTH-1:0] wire_d13_57;
	wire [WIDTH-1:0] wire_d13_58;
	wire [WIDTH-1:0] wire_d13_59;
	wire [WIDTH-1:0] wire_d13_60;
	wire [WIDTH-1:0] wire_d13_61;
	wire [WIDTH-1:0] wire_d13_62;
	wire [WIDTH-1:0] wire_d13_63;
	wire [WIDTH-1:0] wire_d13_64;
	wire [WIDTH-1:0] wire_d13_65;
	wire [WIDTH-1:0] wire_d13_66;
	wire [WIDTH-1:0] wire_d13_67;
	wire [WIDTH-1:0] wire_d13_68;
	wire [WIDTH-1:0] wire_d14_0;
	wire [WIDTH-1:0] wire_d14_1;
	wire [WIDTH-1:0] wire_d14_2;
	wire [WIDTH-1:0] wire_d14_3;
	wire [WIDTH-1:0] wire_d14_4;
	wire [WIDTH-1:0] wire_d14_5;
	wire [WIDTH-1:0] wire_d14_6;
	wire [WIDTH-1:0] wire_d14_7;
	wire [WIDTH-1:0] wire_d14_8;
	wire [WIDTH-1:0] wire_d14_9;
	wire [WIDTH-1:0] wire_d14_10;
	wire [WIDTH-1:0] wire_d14_11;
	wire [WIDTH-1:0] wire_d14_12;
	wire [WIDTH-1:0] wire_d14_13;
	wire [WIDTH-1:0] wire_d14_14;
	wire [WIDTH-1:0] wire_d14_15;
	wire [WIDTH-1:0] wire_d14_16;
	wire [WIDTH-1:0] wire_d14_17;
	wire [WIDTH-1:0] wire_d14_18;
	wire [WIDTH-1:0] wire_d14_19;
	wire [WIDTH-1:0] wire_d14_20;
	wire [WIDTH-1:0] wire_d14_21;
	wire [WIDTH-1:0] wire_d14_22;
	wire [WIDTH-1:0] wire_d14_23;
	wire [WIDTH-1:0] wire_d14_24;
	wire [WIDTH-1:0] wire_d14_25;
	wire [WIDTH-1:0] wire_d14_26;
	wire [WIDTH-1:0] wire_d14_27;
	wire [WIDTH-1:0] wire_d14_28;
	wire [WIDTH-1:0] wire_d14_29;
	wire [WIDTH-1:0] wire_d14_30;
	wire [WIDTH-1:0] wire_d14_31;
	wire [WIDTH-1:0] wire_d14_32;
	wire [WIDTH-1:0] wire_d14_33;
	wire [WIDTH-1:0] wire_d14_34;
	wire [WIDTH-1:0] wire_d14_35;
	wire [WIDTH-1:0] wire_d14_36;
	wire [WIDTH-1:0] wire_d14_37;
	wire [WIDTH-1:0] wire_d14_38;
	wire [WIDTH-1:0] wire_d14_39;
	wire [WIDTH-1:0] wire_d14_40;
	wire [WIDTH-1:0] wire_d14_41;
	wire [WIDTH-1:0] wire_d14_42;
	wire [WIDTH-1:0] wire_d14_43;
	wire [WIDTH-1:0] wire_d14_44;
	wire [WIDTH-1:0] wire_d14_45;
	wire [WIDTH-1:0] wire_d14_46;
	wire [WIDTH-1:0] wire_d14_47;
	wire [WIDTH-1:0] wire_d14_48;
	wire [WIDTH-1:0] wire_d14_49;
	wire [WIDTH-1:0] wire_d14_50;
	wire [WIDTH-1:0] wire_d14_51;
	wire [WIDTH-1:0] wire_d14_52;
	wire [WIDTH-1:0] wire_d14_53;
	wire [WIDTH-1:0] wire_d14_54;
	wire [WIDTH-1:0] wire_d14_55;
	wire [WIDTH-1:0] wire_d14_56;
	wire [WIDTH-1:0] wire_d14_57;
	wire [WIDTH-1:0] wire_d14_58;
	wire [WIDTH-1:0] wire_d14_59;
	wire [WIDTH-1:0] wire_d14_60;
	wire [WIDTH-1:0] wire_d14_61;
	wire [WIDTH-1:0] wire_d14_62;
	wire [WIDTH-1:0] wire_d14_63;
	wire [WIDTH-1:0] wire_d14_64;
	wire [WIDTH-1:0] wire_d14_65;
	wire [WIDTH-1:0] wire_d14_66;
	wire [WIDTH-1:0] wire_d14_67;
	wire [WIDTH-1:0] wire_d14_68;
	wire [WIDTH-1:0] wire_d15_0;
	wire [WIDTH-1:0] wire_d15_1;
	wire [WIDTH-1:0] wire_d15_2;
	wire [WIDTH-1:0] wire_d15_3;
	wire [WIDTH-1:0] wire_d15_4;
	wire [WIDTH-1:0] wire_d15_5;
	wire [WIDTH-1:0] wire_d15_6;
	wire [WIDTH-1:0] wire_d15_7;
	wire [WIDTH-1:0] wire_d15_8;
	wire [WIDTH-1:0] wire_d15_9;
	wire [WIDTH-1:0] wire_d15_10;
	wire [WIDTH-1:0] wire_d15_11;
	wire [WIDTH-1:0] wire_d15_12;
	wire [WIDTH-1:0] wire_d15_13;
	wire [WIDTH-1:0] wire_d15_14;
	wire [WIDTH-1:0] wire_d15_15;
	wire [WIDTH-1:0] wire_d15_16;
	wire [WIDTH-1:0] wire_d15_17;
	wire [WIDTH-1:0] wire_d15_18;
	wire [WIDTH-1:0] wire_d15_19;
	wire [WIDTH-1:0] wire_d15_20;
	wire [WIDTH-1:0] wire_d15_21;
	wire [WIDTH-1:0] wire_d15_22;
	wire [WIDTH-1:0] wire_d15_23;
	wire [WIDTH-1:0] wire_d15_24;
	wire [WIDTH-1:0] wire_d15_25;
	wire [WIDTH-1:0] wire_d15_26;
	wire [WIDTH-1:0] wire_d15_27;
	wire [WIDTH-1:0] wire_d15_28;
	wire [WIDTH-1:0] wire_d15_29;
	wire [WIDTH-1:0] wire_d15_30;
	wire [WIDTH-1:0] wire_d15_31;
	wire [WIDTH-1:0] wire_d15_32;
	wire [WIDTH-1:0] wire_d15_33;
	wire [WIDTH-1:0] wire_d15_34;
	wire [WIDTH-1:0] wire_d15_35;
	wire [WIDTH-1:0] wire_d15_36;
	wire [WIDTH-1:0] wire_d15_37;
	wire [WIDTH-1:0] wire_d15_38;
	wire [WIDTH-1:0] wire_d15_39;
	wire [WIDTH-1:0] wire_d15_40;
	wire [WIDTH-1:0] wire_d15_41;
	wire [WIDTH-1:0] wire_d15_42;
	wire [WIDTH-1:0] wire_d15_43;
	wire [WIDTH-1:0] wire_d15_44;
	wire [WIDTH-1:0] wire_d15_45;
	wire [WIDTH-1:0] wire_d15_46;
	wire [WIDTH-1:0] wire_d15_47;
	wire [WIDTH-1:0] wire_d15_48;
	wire [WIDTH-1:0] wire_d15_49;
	wire [WIDTH-1:0] wire_d15_50;
	wire [WIDTH-1:0] wire_d15_51;
	wire [WIDTH-1:0] wire_d15_52;
	wire [WIDTH-1:0] wire_d15_53;
	wire [WIDTH-1:0] wire_d15_54;
	wire [WIDTH-1:0] wire_d15_55;
	wire [WIDTH-1:0] wire_d15_56;
	wire [WIDTH-1:0] wire_d15_57;
	wire [WIDTH-1:0] wire_d15_58;
	wire [WIDTH-1:0] wire_d15_59;
	wire [WIDTH-1:0] wire_d15_60;
	wire [WIDTH-1:0] wire_d15_61;
	wire [WIDTH-1:0] wire_d15_62;
	wire [WIDTH-1:0] wire_d15_63;
	wire [WIDTH-1:0] wire_d15_64;
	wire [WIDTH-1:0] wire_d15_65;
	wire [WIDTH-1:0] wire_d15_66;
	wire [WIDTH-1:0] wire_d15_67;
	wire [WIDTH-1:0] wire_d15_68;
	wire [WIDTH-1:0] wire_d16_0;
	wire [WIDTH-1:0] wire_d16_1;
	wire [WIDTH-1:0] wire_d16_2;
	wire [WIDTH-1:0] wire_d16_3;
	wire [WIDTH-1:0] wire_d16_4;
	wire [WIDTH-1:0] wire_d16_5;
	wire [WIDTH-1:0] wire_d16_6;
	wire [WIDTH-1:0] wire_d16_7;
	wire [WIDTH-1:0] wire_d16_8;
	wire [WIDTH-1:0] wire_d16_9;
	wire [WIDTH-1:0] wire_d16_10;
	wire [WIDTH-1:0] wire_d16_11;
	wire [WIDTH-1:0] wire_d16_12;
	wire [WIDTH-1:0] wire_d16_13;
	wire [WIDTH-1:0] wire_d16_14;
	wire [WIDTH-1:0] wire_d16_15;
	wire [WIDTH-1:0] wire_d16_16;
	wire [WIDTH-1:0] wire_d16_17;
	wire [WIDTH-1:0] wire_d16_18;
	wire [WIDTH-1:0] wire_d16_19;
	wire [WIDTH-1:0] wire_d16_20;
	wire [WIDTH-1:0] wire_d16_21;
	wire [WIDTH-1:0] wire_d16_22;
	wire [WIDTH-1:0] wire_d16_23;
	wire [WIDTH-1:0] wire_d16_24;
	wire [WIDTH-1:0] wire_d16_25;
	wire [WIDTH-1:0] wire_d16_26;
	wire [WIDTH-1:0] wire_d16_27;
	wire [WIDTH-1:0] wire_d16_28;
	wire [WIDTH-1:0] wire_d16_29;
	wire [WIDTH-1:0] wire_d16_30;
	wire [WIDTH-1:0] wire_d16_31;
	wire [WIDTH-1:0] wire_d16_32;
	wire [WIDTH-1:0] wire_d16_33;
	wire [WIDTH-1:0] wire_d16_34;
	wire [WIDTH-1:0] wire_d16_35;
	wire [WIDTH-1:0] wire_d16_36;
	wire [WIDTH-1:0] wire_d16_37;
	wire [WIDTH-1:0] wire_d16_38;
	wire [WIDTH-1:0] wire_d16_39;
	wire [WIDTH-1:0] wire_d16_40;
	wire [WIDTH-1:0] wire_d16_41;
	wire [WIDTH-1:0] wire_d16_42;
	wire [WIDTH-1:0] wire_d16_43;
	wire [WIDTH-1:0] wire_d16_44;
	wire [WIDTH-1:0] wire_d16_45;
	wire [WIDTH-1:0] wire_d16_46;
	wire [WIDTH-1:0] wire_d16_47;
	wire [WIDTH-1:0] wire_d16_48;
	wire [WIDTH-1:0] wire_d16_49;
	wire [WIDTH-1:0] wire_d16_50;
	wire [WIDTH-1:0] wire_d16_51;
	wire [WIDTH-1:0] wire_d16_52;
	wire [WIDTH-1:0] wire_d16_53;
	wire [WIDTH-1:0] wire_d16_54;
	wire [WIDTH-1:0] wire_d16_55;
	wire [WIDTH-1:0] wire_d16_56;
	wire [WIDTH-1:0] wire_d16_57;
	wire [WIDTH-1:0] wire_d16_58;
	wire [WIDTH-1:0] wire_d16_59;
	wire [WIDTH-1:0] wire_d16_60;
	wire [WIDTH-1:0] wire_d16_61;
	wire [WIDTH-1:0] wire_d16_62;
	wire [WIDTH-1:0] wire_d16_63;
	wire [WIDTH-1:0] wire_d16_64;
	wire [WIDTH-1:0] wire_d16_65;
	wire [WIDTH-1:0] wire_d16_66;
	wire [WIDTH-1:0] wire_d16_67;
	wire [WIDTH-1:0] wire_d16_68;
	wire [WIDTH-1:0] wire_d17_0;
	wire [WIDTH-1:0] wire_d17_1;
	wire [WIDTH-1:0] wire_d17_2;
	wire [WIDTH-1:0] wire_d17_3;
	wire [WIDTH-1:0] wire_d17_4;
	wire [WIDTH-1:0] wire_d17_5;
	wire [WIDTH-1:0] wire_d17_6;
	wire [WIDTH-1:0] wire_d17_7;
	wire [WIDTH-1:0] wire_d17_8;
	wire [WIDTH-1:0] wire_d17_9;
	wire [WIDTH-1:0] wire_d17_10;
	wire [WIDTH-1:0] wire_d17_11;
	wire [WIDTH-1:0] wire_d17_12;
	wire [WIDTH-1:0] wire_d17_13;
	wire [WIDTH-1:0] wire_d17_14;
	wire [WIDTH-1:0] wire_d17_15;
	wire [WIDTH-1:0] wire_d17_16;
	wire [WIDTH-1:0] wire_d17_17;
	wire [WIDTH-1:0] wire_d17_18;
	wire [WIDTH-1:0] wire_d17_19;
	wire [WIDTH-1:0] wire_d17_20;
	wire [WIDTH-1:0] wire_d17_21;
	wire [WIDTH-1:0] wire_d17_22;
	wire [WIDTH-1:0] wire_d17_23;
	wire [WIDTH-1:0] wire_d17_24;
	wire [WIDTH-1:0] wire_d17_25;
	wire [WIDTH-1:0] wire_d17_26;
	wire [WIDTH-1:0] wire_d17_27;
	wire [WIDTH-1:0] wire_d17_28;
	wire [WIDTH-1:0] wire_d17_29;
	wire [WIDTH-1:0] wire_d17_30;
	wire [WIDTH-1:0] wire_d17_31;
	wire [WIDTH-1:0] wire_d17_32;
	wire [WIDTH-1:0] wire_d17_33;
	wire [WIDTH-1:0] wire_d17_34;
	wire [WIDTH-1:0] wire_d17_35;
	wire [WIDTH-1:0] wire_d17_36;
	wire [WIDTH-1:0] wire_d17_37;
	wire [WIDTH-1:0] wire_d17_38;
	wire [WIDTH-1:0] wire_d17_39;
	wire [WIDTH-1:0] wire_d17_40;
	wire [WIDTH-1:0] wire_d17_41;
	wire [WIDTH-1:0] wire_d17_42;
	wire [WIDTH-1:0] wire_d17_43;
	wire [WIDTH-1:0] wire_d17_44;
	wire [WIDTH-1:0] wire_d17_45;
	wire [WIDTH-1:0] wire_d17_46;
	wire [WIDTH-1:0] wire_d17_47;
	wire [WIDTH-1:0] wire_d17_48;
	wire [WIDTH-1:0] wire_d17_49;
	wire [WIDTH-1:0] wire_d17_50;
	wire [WIDTH-1:0] wire_d17_51;
	wire [WIDTH-1:0] wire_d17_52;
	wire [WIDTH-1:0] wire_d17_53;
	wire [WIDTH-1:0] wire_d17_54;
	wire [WIDTH-1:0] wire_d17_55;
	wire [WIDTH-1:0] wire_d17_56;
	wire [WIDTH-1:0] wire_d17_57;
	wire [WIDTH-1:0] wire_d17_58;
	wire [WIDTH-1:0] wire_d17_59;
	wire [WIDTH-1:0] wire_d17_60;
	wire [WIDTH-1:0] wire_d17_61;
	wire [WIDTH-1:0] wire_d17_62;
	wire [WIDTH-1:0] wire_d17_63;
	wire [WIDTH-1:0] wire_d17_64;
	wire [WIDTH-1:0] wire_d17_65;
	wire [WIDTH-1:0] wire_d17_66;
	wire [WIDTH-1:0] wire_d17_67;
	wire [WIDTH-1:0] wire_d17_68;
	wire [WIDTH-1:0] wire_d18_0;
	wire [WIDTH-1:0] wire_d18_1;
	wire [WIDTH-1:0] wire_d18_2;
	wire [WIDTH-1:0] wire_d18_3;
	wire [WIDTH-1:0] wire_d18_4;
	wire [WIDTH-1:0] wire_d18_5;
	wire [WIDTH-1:0] wire_d18_6;
	wire [WIDTH-1:0] wire_d18_7;
	wire [WIDTH-1:0] wire_d18_8;
	wire [WIDTH-1:0] wire_d18_9;
	wire [WIDTH-1:0] wire_d18_10;
	wire [WIDTH-1:0] wire_d18_11;
	wire [WIDTH-1:0] wire_d18_12;
	wire [WIDTH-1:0] wire_d18_13;
	wire [WIDTH-1:0] wire_d18_14;
	wire [WIDTH-1:0] wire_d18_15;
	wire [WIDTH-1:0] wire_d18_16;
	wire [WIDTH-1:0] wire_d18_17;
	wire [WIDTH-1:0] wire_d18_18;
	wire [WIDTH-1:0] wire_d18_19;
	wire [WIDTH-1:0] wire_d18_20;
	wire [WIDTH-1:0] wire_d18_21;
	wire [WIDTH-1:0] wire_d18_22;
	wire [WIDTH-1:0] wire_d18_23;
	wire [WIDTH-1:0] wire_d18_24;
	wire [WIDTH-1:0] wire_d18_25;
	wire [WIDTH-1:0] wire_d18_26;
	wire [WIDTH-1:0] wire_d18_27;
	wire [WIDTH-1:0] wire_d18_28;
	wire [WIDTH-1:0] wire_d18_29;
	wire [WIDTH-1:0] wire_d18_30;
	wire [WIDTH-1:0] wire_d18_31;
	wire [WIDTH-1:0] wire_d18_32;
	wire [WIDTH-1:0] wire_d18_33;
	wire [WIDTH-1:0] wire_d18_34;
	wire [WIDTH-1:0] wire_d18_35;
	wire [WIDTH-1:0] wire_d18_36;
	wire [WIDTH-1:0] wire_d18_37;
	wire [WIDTH-1:0] wire_d18_38;
	wire [WIDTH-1:0] wire_d18_39;
	wire [WIDTH-1:0] wire_d18_40;
	wire [WIDTH-1:0] wire_d18_41;
	wire [WIDTH-1:0] wire_d18_42;
	wire [WIDTH-1:0] wire_d18_43;
	wire [WIDTH-1:0] wire_d18_44;
	wire [WIDTH-1:0] wire_d18_45;
	wire [WIDTH-1:0] wire_d18_46;
	wire [WIDTH-1:0] wire_d18_47;
	wire [WIDTH-1:0] wire_d18_48;
	wire [WIDTH-1:0] wire_d18_49;
	wire [WIDTH-1:0] wire_d18_50;
	wire [WIDTH-1:0] wire_d18_51;
	wire [WIDTH-1:0] wire_d18_52;
	wire [WIDTH-1:0] wire_d18_53;
	wire [WIDTH-1:0] wire_d18_54;
	wire [WIDTH-1:0] wire_d18_55;
	wire [WIDTH-1:0] wire_d18_56;
	wire [WIDTH-1:0] wire_d18_57;
	wire [WIDTH-1:0] wire_d18_58;
	wire [WIDTH-1:0] wire_d18_59;
	wire [WIDTH-1:0] wire_d18_60;
	wire [WIDTH-1:0] wire_d18_61;
	wire [WIDTH-1:0] wire_d18_62;
	wire [WIDTH-1:0] wire_d18_63;
	wire [WIDTH-1:0] wire_d18_64;
	wire [WIDTH-1:0] wire_d18_65;
	wire [WIDTH-1:0] wire_d18_66;
	wire [WIDTH-1:0] wire_d18_67;
	wire [WIDTH-1:0] wire_d18_68;
	wire [WIDTH-1:0] wire_d19_0;
	wire [WIDTH-1:0] wire_d19_1;
	wire [WIDTH-1:0] wire_d19_2;
	wire [WIDTH-1:0] wire_d19_3;
	wire [WIDTH-1:0] wire_d19_4;
	wire [WIDTH-1:0] wire_d19_5;
	wire [WIDTH-1:0] wire_d19_6;
	wire [WIDTH-1:0] wire_d19_7;
	wire [WIDTH-1:0] wire_d19_8;
	wire [WIDTH-1:0] wire_d19_9;
	wire [WIDTH-1:0] wire_d19_10;
	wire [WIDTH-1:0] wire_d19_11;
	wire [WIDTH-1:0] wire_d19_12;
	wire [WIDTH-1:0] wire_d19_13;
	wire [WIDTH-1:0] wire_d19_14;
	wire [WIDTH-1:0] wire_d19_15;
	wire [WIDTH-1:0] wire_d19_16;
	wire [WIDTH-1:0] wire_d19_17;
	wire [WIDTH-1:0] wire_d19_18;
	wire [WIDTH-1:0] wire_d19_19;
	wire [WIDTH-1:0] wire_d19_20;
	wire [WIDTH-1:0] wire_d19_21;
	wire [WIDTH-1:0] wire_d19_22;
	wire [WIDTH-1:0] wire_d19_23;
	wire [WIDTH-1:0] wire_d19_24;
	wire [WIDTH-1:0] wire_d19_25;
	wire [WIDTH-1:0] wire_d19_26;
	wire [WIDTH-1:0] wire_d19_27;
	wire [WIDTH-1:0] wire_d19_28;
	wire [WIDTH-1:0] wire_d19_29;
	wire [WIDTH-1:0] wire_d19_30;
	wire [WIDTH-1:0] wire_d19_31;
	wire [WIDTH-1:0] wire_d19_32;
	wire [WIDTH-1:0] wire_d19_33;
	wire [WIDTH-1:0] wire_d19_34;
	wire [WIDTH-1:0] wire_d19_35;
	wire [WIDTH-1:0] wire_d19_36;
	wire [WIDTH-1:0] wire_d19_37;
	wire [WIDTH-1:0] wire_d19_38;
	wire [WIDTH-1:0] wire_d19_39;
	wire [WIDTH-1:0] wire_d19_40;
	wire [WIDTH-1:0] wire_d19_41;
	wire [WIDTH-1:0] wire_d19_42;
	wire [WIDTH-1:0] wire_d19_43;
	wire [WIDTH-1:0] wire_d19_44;
	wire [WIDTH-1:0] wire_d19_45;
	wire [WIDTH-1:0] wire_d19_46;
	wire [WIDTH-1:0] wire_d19_47;
	wire [WIDTH-1:0] wire_d19_48;
	wire [WIDTH-1:0] wire_d19_49;
	wire [WIDTH-1:0] wire_d19_50;
	wire [WIDTH-1:0] wire_d19_51;
	wire [WIDTH-1:0] wire_d19_52;
	wire [WIDTH-1:0] wire_d19_53;
	wire [WIDTH-1:0] wire_d19_54;
	wire [WIDTH-1:0] wire_d19_55;
	wire [WIDTH-1:0] wire_d19_56;
	wire [WIDTH-1:0] wire_d19_57;
	wire [WIDTH-1:0] wire_d19_58;
	wire [WIDTH-1:0] wire_d19_59;
	wire [WIDTH-1:0] wire_d19_60;
	wire [WIDTH-1:0] wire_d19_61;
	wire [WIDTH-1:0] wire_d19_62;
	wire [WIDTH-1:0] wire_d19_63;
	wire [WIDTH-1:0] wire_d19_64;
	wire [WIDTH-1:0] wire_d19_65;
	wire [WIDTH-1:0] wire_d19_66;
	wire [WIDTH-1:0] wire_d19_67;
	wire [WIDTH-1:0] wire_d19_68;
	wire [WIDTH-1:0] wire_d20_0;
	wire [WIDTH-1:0] wire_d20_1;
	wire [WIDTH-1:0] wire_d20_2;
	wire [WIDTH-1:0] wire_d20_3;
	wire [WIDTH-1:0] wire_d20_4;
	wire [WIDTH-1:0] wire_d20_5;
	wire [WIDTH-1:0] wire_d20_6;
	wire [WIDTH-1:0] wire_d20_7;
	wire [WIDTH-1:0] wire_d20_8;
	wire [WIDTH-1:0] wire_d20_9;
	wire [WIDTH-1:0] wire_d20_10;
	wire [WIDTH-1:0] wire_d20_11;
	wire [WIDTH-1:0] wire_d20_12;
	wire [WIDTH-1:0] wire_d20_13;
	wire [WIDTH-1:0] wire_d20_14;
	wire [WIDTH-1:0] wire_d20_15;
	wire [WIDTH-1:0] wire_d20_16;
	wire [WIDTH-1:0] wire_d20_17;
	wire [WIDTH-1:0] wire_d20_18;
	wire [WIDTH-1:0] wire_d20_19;
	wire [WIDTH-1:0] wire_d20_20;
	wire [WIDTH-1:0] wire_d20_21;
	wire [WIDTH-1:0] wire_d20_22;
	wire [WIDTH-1:0] wire_d20_23;
	wire [WIDTH-1:0] wire_d20_24;
	wire [WIDTH-1:0] wire_d20_25;
	wire [WIDTH-1:0] wire_d20_26;
	wire [WIDTH-1:0] wire_d20_27;
	wire [WIDTH-1:0] wire_d20_28;
	wire [WIDTH-1:0] wire_d20_29;
	wire [WIDTH-1:0] wire_d20_30;
	wire [WIDTH-1:0] wire_d20_31;
	wire [WIDTH-1:0] wire_d20_32;
	wire [WIDTH-1:0] wire_d20_33;
	wire [WIDTH-1:0] wire_d20_34;
	wire [WIDTH-1:0] wire_d20_35;
	wire [WIDTH-1:0] wire_d20_36;
	wire [WIDTH-1:0] wire_d20_37;
	wire [WIDTH-1:0] wire_d20_38;
	wire [WIDTH-1:0] wire_d20_39;
	wire [WIDTH-1:0] wire_d20_40;
	wire [WIDTH-1:0] wire_d20_41;
	wire [WIDTH-1:0] wire_d20_42;
	wire [WIDTH-1:0] wire_d20_43;
	wire [WIDTH-1:0] wire_d20_44;
	wire [WIDTH-1:0] wire_d20_45;
	wire [WIDTH-1:0] wire_d20_46;
	wire [WIDTH-1:0] wire_d20_47;
	wire [WIDTH-1:0] wire_d20_48;
	wire [WIDTH-1:0] wire_d20_49;
	wire [WIDTH-1:0] wire_d20_50;
	wire [WIDTH-1:0] wire_d20_51;
	wire [WIDTH-1:0] wire_d20_52;
	wire [WIDTH-1:0] wire_d20_53;
	wire [WIDTH-1:0] wire_d20_54;
	wire [WIDTH-1:0] wire_d20_55;
	wire [WIDTH-1:0] wire_d20_56;
	wire [WIDTH-1:0] wire_d20_57;
	wire [WIDTH-1:0] wire_d20_58;
	wire [WIDTH-1:0] wire_d20_59;
	wire [WIDTH-1:0] wire_d20_60;
	wire [WIDTH-1:0] wire_d20_61;
	wire [WIDTH-1:0] wire_d20_62;
	wire [WIDTH-1:0] wire_d20_63;
	wire [WIDTH-1:0] wire_d20_64;
	wire [WIDTH-1:0] wire_d20_65;
	wire [WIDTH-1:0] wire_d20_66;
	wire [WIDTH-1:0] wire_d20_67;
	wire [WIDTH-1:0] wire_d20_68;
	wire [WIDTH-1:0] wire_d21_0;
	wire [WIDTH-1:0] wire_d21_1;
	wire [WIDTH-1:0] wire_d21_2;
	wire [WIDTH-1:0] wire_d21_3;
	wire [WIDTH-1:0] wire_d21_4;
	wire [WIDTH-1:0] wire_d21_5;
	wire [WIDTH-1:0] wire_d21_6;
	wire [WIDTH-1:0] wire_d21_7;
	wire [WIDTH-1:0] wire_d21_8;
	wire [WIDTH-1:0] wire_d21_9;
	wire [WIDTH-1:0] wire_d21_10;
	wire [WIDTH-1:0] wire_d21_11;
	wire [WIDTH-1:0] wire_d21_12;
	wire [WIDTH-1:0] wire_d21_13;
	wire [WIDTH-1:0] wire_d21_14;
	wire [WIDTH-1:0] wire_d21_15;
	wire [WIDTH-1:0] wire_d21_16;
	wire [WIDTH-1:0] wire_d21_17;
	wire [WIDTH-1:0] wire_d21_18;
	wire [WIDTH-1:0] wire_d21_19;
	wire [WIDTH-1:0] wire_d21_20;
	wire [WIDTH-1:0] wire_d21_21;
	wire [WIDTH-1:0] wire_d21_22;
	wire [WIDTH-1:0] wire_d21_23;
	wire [WIDTH-1:0] wire_d21_24;
	wire [WIDTH-1:0] wire_d21_25;
	wire [WIDTH-1:0] wire_d21_26;
	wire [WIDTH-1:0] wire_d21_27;
	wire [WIDTH-1:0] wire_d21_28;
	wire [WIDTH-1:0] wire_d21_29;
	wire [WIDTH-1:0] wire_d21_30;
	wire [WIDTH-1:0] wire_d21_31;
	wire [WIDTH-1:0] wire_d21_32;
	wire [WIDTH-1:0] wire_d21_33;
	wire [WIDTH-1:0] wire_d21_34;
	wire [WIDTH-1:0] wire_d21_35;
	wire [WIDTH-1:0] wire_d21_36;
	wire [WIDTH-1:0] wire_d21_37;
	wire [WIDTH-1:0] wire_d21_38;
	wire [WIDTH-1:0] wire_d21_39;
	wire [WIDTH-1:0] wire_d21_40;
	wire [WIDTH-1:0] wire_d21_41;
	wire [WIDTH-1:0] wire_d21_42;
	wire [WIDTH-1:0] wire_d21_43;
	wire [WIDTH-1:0] wire_d21_44;
	wire [WIDTH-1:0] wire_d21_45;
	wire [WIDTH-1:0] wire_d21_46;
	wire [WIDTH-1:0] wire_d21_47;
	wire [WIDTH-1:0] wire_d21_48;
	wire [WIDTH-1:0] wire_d21_49;
	wire [WIDTH-1:0] wire_d21_50;
	wire [WIDTH-1:0] wire_d21_51;
	wire [WIDTH-1:0] wire_d21_52;
	wire [WIDTH-1:0] wire_d21_53;
	wire [WIDTH-1:0] wire_d21_54;
	wire [WIDTH-1:0] wire_d21_55;
	wire [WIDTH-1:0] wire_d21_56;
	wire [WIDTH-1:0] wire_d21_57;
	wire [WIDTH-1:0] wire_d21_58;
	wire [WIDTH-1:0] wire_d21_59;
	wire [WIDTH-1:0] wire_d21_60;
	wire [WIDTH-1:0] wire_d21_61;
	wire [WIDTH-1:0] wire_d21_62;
	wire [WIDTH-1:0] wire_d21_63;
	wire [WIDTH-1:0] wire_d21_64;
	wire [WIDTH-1:0] wire_d21_65;
	wire [WIDTH-1:0] wire_d21_66;
	wire [WIDTH-1:0] wire_d21_67;
	wire [WIDTH-1:0] wire_d21_68;
	wire [WIDTH-1:0] wire_d22_0;
	wire [WIDTH-1:0] wire_d22_1;
	wire [WIDTH-1:0] wire_d22_2;
	wire [WIDTH-1:0] wire_d22_3;
	wire [WIDTH-1:0] wire_d22_4;
	wire [WIDTH-1:0] wire_d22_5;
	wire [WIDTH-1:0] wire_d22_6;
	wire [WIDTH-1:0] wire_d22_7;
	wire [WIDTH-1:0] wire_d22_8;
	wire [WIDTH-1:0] wire_d22_9;
	wire [WIDTH-1:0] wire_d22_10;
	wire [WIDTH-1:0] wire_d22_11;
	wire [WIDTH-1:0] wire_d22_12;
	wire [WIDTH-1:0] wire_d22_13;
	wire [WIDTH-1:0] wire_d22_14;
	wire [WIDTH-1:0] wire_d22_15;
	wire [WIDTH-1:0] wire_d22_16;
	wire [WIDTH-1:0] wire_d22_17;
	wire [WIDTH-1:0] wire_d22_18;
	wire [WIDTH-1:0] wire_d22_19;
	wire [WIDTH-1:0] wire_d22_20;
	wire [WIDTH-1:0] wire_d22_21;
	wire [WIDTH-1:0] wire_d22_22;
	wire [WIDTH-1:0] wire_d22_23;
	wire [WIDTH-1:0] wire_d22_24;
	wire [WIDTH-1:0] wire_d22_25;
	wire [WIDTH-1:0] wire_d22_26;
	wire [WIDTH-1:0] wire_d22_27;
	wire [WIDTH-1:0] wire_d22_28;
	wire [WIDTH-1:0] wire_d22_29;
	wire [WIDTH-1:0] wire_d22_30;
	wire [WIDTH-1:0] wire_d22_31;
	wire [WIDTH-1:0] wire_d22_32;
	wire [WIDTH-1:0] wire_d22_33;
	wire [WIDTH-1:0] wire_d22_34;
	wire [WIDTH-1:0] wire_d22_35;
	wire [WIDTH-1:0] wire_d22_36;
	wire [WIDTH-1:0] wire_d22_37;
	wire [WIDTH-1:0] wire_d22_38;
	wire [WIDTH-1:0] wire_d22_39;
	wire [WIDTH-1:0] wire_d22_40;
	wire [WIDTH-1:0] wire_d22_41;
	wire [WIDTH-1:0] wire_d22_42;
	wire [WIDTH-1:0] wire_d22_43;
	wire [WIDTH-1:0] wire_d22_44;
	wire [WIDTH-1:0] wire_d22_45;
	wire [WIDTH-1:0] wire_d22_46;
	wire [WIDTH-1:0] wire_d22_47;
	wire [WIDTH-1:0] wire_d22_48;
	wire [WIDTH-1:0] wire_d22_49;
	wire [WIDTH-1:0] wire_d22_50;
	wire [WIDTH-1:0] wire_d22_51;
	wire [WIDTH-1:0] wire_d22_52;
	wire [WIDTH-1:0] wire_d22_53;
	wire [WIDTH-1:0] wire_d22_54;
	wire [WIDTH-1:0] wire_d22_55;
	wire [WIDTH-1:0] wire_d22_56;
	wire [WIDTH-1:0] wire_d22_57;
	wire [WIDTH-1:0] wire_d22_58;
	wire [WIDTH-1:0] wire_d22_59;
	wire [WIDTH-1:0] wire_d22_60;
	wire [WIDTH-1:0] wire_d22_61;
	wire [WIDTH-1:0] wire_d22_62;
	wire [WIDTH-1:0] wire_d22_63;
	wire [WIDTH-1:0] wire_d22_64;
	wire [WIDTH-1:0] wire_d22_65;
	wire [WIDTH-1:0] wire_d22_66;
	wire [WIDTH-1:0] wire_d22_67;
	wire [WIDTH-1:0] wire_d22_68;
	wire [WIDTH-1:0] wire_d23_0;
	wire [WIDTH-1:0] wire_d23_1;
	wire [WIDTH-1:0] wire_d23_2;
	wire [WIDTH-1:0] wire_d23_3;
	wire [WIDTH-1:0] wire_d23_4;
	wire [WIDTH-1:0] wire_d23_5;
	wire [WIDTH-1:0] wire_d23_6;
	wire [WIDTH-1:0] wire_d23_7;
	wire [WIDTH-1:0] wire_d23_8;
	wire [WIDTH-1:0] wire_d23_9;
	wire [WIDTH-1:0] wire_d23_10;
	wire [WIDTH-1:0] wire_d23_11;
	wire [WIDTH-1:0] wire_d23_12;
	wire [WIDTH-1:0] wire_d23_13;
	wire [WIDTH-1:0] wire_d23_14;
	wire [WIDTH-1:0] wire_d23_15;
	wire [WIDTH-1:0] wire_d23_16;
	wire [WIDTH-1:0] wire_d23_17;
	wire [WIDTH-1:0] wire_d23_18;
	wire [WIDTH-1:0] wire_d23_19;
	wire [WIDTH-1:0] wire_d23_20;
	wire [WIDTH-1:0] wire_d23_21;
	wire [WIDTH-1:0] wire_d23_22;
	wire [WIDTH-1:0] wire_d23_23;
	wire [WIDTH-1:0] wire_d23_24;
	wire [WIDTH-1:0] wire_d23_25;
	wire [WIDTH-1:0] wire_d23_26;
	wire [WIDTH-1:0] wire_d23_27;
	wire [WIDTH-1:0] wire_d23_28;
	wire [WIDTH-1:0] wire_d23_29;
	wire [WIDTH-1:0] wire_d23_30;
	wire [WIDTH-1:0] wire_d23_31;
	wire [WIDTH-1:0] wire_d23_32;
	wire [WIDTH-1:0] wire_d23_33;
	wire [WIDTH-1:0] wire_d23_34;
	wire [WIDTH-1:0] wire_d23_35;
	wire [WIDTH-1:0] wire_d23_36;
	wire [WIDTH-1:0] wire_d23_37;
	wire [WIDTH-1:0] wire_d23_38;
	wire [WIDTH-1:0] wire_d23_39;
	wire [WIDTH-1:0] wire_d23_40;
	wire [WIDTH-1:0] wire_d23_41;
	wire [WIDTH-1:0] wire_d23_42;
	wire [WIDTH-1:0] wire_d23_43;
	wire [WIDTH-1:0] wire_d23_44;
	wire [WIDTH-1:0] wire_d23_45;
	wire [WIDTH-1:0] wire_d23_46;
	wire [WIDTH-1:0] wire_d23_47;
	wire [WIDTH-1:0] wire_d23_48;
	wire [WIDTH-1:0] wire_d23_49;
	wire [WIDTH-1:0] wire_d23_50;
	wire [WIDTH-1:0] wire_d23_51;
	wire [WIDTH-1:0] wire_d23_52;
	wire [WIDTH-1:0] wire_d23_53;
	wire [WIDTH-1:0] wire_d23_54;
	wire [WIDTH-1:0] wire_d23_55;
	wire [WIDTH-1:0] wire_d23_56;
	wire [WIDTH-1:0] wire_d23_57;
	wire [WIDTH-1:0] wire_d23_58;
	wire [WIDTH-1:0] wire_d23_59;
	wire [WIDTH-1:0] wire_d23_60;
	wire [WIDTH-1:0] wire_d23_61;
	wire [WIDTH-1:0] wire_d23_62;
	wire [WIDTH-1:0] wire_d23_63;
	wire [WIDTH-1:0] wire_d23_64;
	wire [WIDTH-1:0] wire_d23_65;
	wire [WIDTH-1:0] wire_d23_66;
	wire [WIDTH-1:0] wire_d23_67;
	wire [WIDTH-1:0] wire_d23_68;
	wire [WIDTH-1:0] wire_d24_0;
	wire [WIDTH-1:0] wire_d24_1;
	wire [WIDTH-1:0] wire_d24_2;
	wire [WIDTH-1:0] wire_d24_3;
	wire [WIDTH-1:0] wire_d24_4;
	wire [WIDTH-1:0] wire_d24_5;
	wire [WIDTH-1:0] wire_d24_6;
	wire [WIDTH-1:0] wire_d24_7;
	wire [WIDTH-1:0] wire_d24_8;
	wire [WIDTH-1:0] wire_d24_9;
	wire [WIDTH-1:0] wire_d24_10;
	wire [WIDTH-1:0] wire_d24_11;
	wire [WIDTH-1:0] wire_d24_12;
	wire [WIDTH-1:0] wire_d24_13;
	wire [WIDTH-1:0] wire_d24_14;
	wire [WIDTH-1:0] wire_d24_15;
	wire [WIDTH-1:0] wire_d24_16;
	wire [WIDTH-1:0] wire_d24_17;
	wire [WIDTH-1:0] wire_d24_18;
	wire [WIDTH-1:0] wire_d24_19;
	wire [WIDTH-1:0] wire_d24_20;
	wire [WIDTH-1:0] wire_d24_21;
	wire [WIDTH-1:0] wire_d24_22;
	wire [WIDTH-1:0] wire_d24_23;
	wire [WIDTH-1:0] wire_d24_24;
	wire [WIDTH-1:0] wire_d24_25;
	wire [WIDTH-1:0] wire_d24_26;
	wire [WIDTH-1:0] wire_d24_27;
	wire [WIDTH-1:0] wire_d24_28;
	wire [WIDTH-1:0] wire_d24_29;
	wire [WIDTH-1:0] wire_d24_30;
	wire [WIDTH-1:0] wire_d24_31;
	wire [WIDTH-1:0] wire_d24_32;
	wire [WIDTH-1:0] wire_d24_33;
	wire [WIDTH-1:0] wire_d24_34;
	wire [WIDTH-1:0] wire_d24_35;
	wire [WIDTH-1:0] wire_d24_36;
	wire [WIDTH-1:0] wire_d24_37;
	wire [WIDTH-1:0] wire_d24_38;
	wire [WIDTH-1:0] wire_d24_39;
	wire [WIDTH-1:0] wire_d24_40;
	wire [WIDTH-1:0] wire_d24_41;
	wire [WIDTH-1:0] wire_d24_42;
	wire [WIDTH-1:0] wire_d24_43;
	wire [WIDTH-1:0] wire_d24_44;
	wire [WIDTH-1:0] wire_d24_45;
	wire [WIDTH-1:0] wire_d24_46;
	wire [WIDTH-1:0] wire_d24_47;
	wire [WIDTH-1:0] wire_d24_48;
	wire [WIDTH-1:0] wire_d24_49;
	wire [WIDTH-1:0] wire_d24_50;
	wire [WIDTH-1:0] wire_d24_51;
	wire [WIDTH-1:0] wire_d24_52;
	wire [WIDTH-1:0] wire_d24_53;
	wire [WIDTH-1:0] wire_d24_54;
	wire [WIDTH-1:0] wire_d24_55;
	wire [WIDTH-1:0] wire_d24_56;
	wire [WIDTH-1:0] wire_d24_57;
	wire [WIDTH-1:0] wire_d24_58;
	wire [WIDTH-1:0] wire_d24_59;
	wire [WIDTH-1:0] wire_d24_60;
	wire [WIDTH-1:0] wire_d24_61;
	wire [WIDTH-1:0] wire_d24_62;
	wire [WIDTH-1:0] wire_d24_63;
	wire [WIDTH-1:0] wire_d24_64;
	wire [WIDTH-1:0] wire_d24_65;
	wire [WIDTH-1:0] wire_d24_66;
	wire [WIDTH-1:0] wire_d24_67;
	wire [WIDTH-1:0] wire_d24_68;
	wire [WIDTH-1:0] wire_d25_0;
	wire [WIDTH-1:0] wire_d25_1;
	wire [WIDTH-1:0] wire_d25_2;
	wire [WIDTH-1:0] wire_d25_3;
	wire [WIDTH-1:0] wire_d25_4;
	wire [WIDTH-1:0] wire_d25_5;
	wire [WIDTH-1:0] wire_d25_6;
	wire [WIDTH-1:0] wire_d25_7;
	wire [WIDTH-1:0] wire_d25_8;
	wire [WIDTH-1:0] wire_d25_9;
	wire [WIDTH-1:0] wire_d25_10;
	wire [WIDTH-1:0] wire_d25_11;
	wire [WIDTH-1:0] wire_d25_12;
	wire [WIDTH-1:0] wire_d25_13;
	wire [WIDTH-1:0] wire_d25_14;
	wire [WIDTH-1:0] wire_d25_15;
	wire [WIDTH-1:0] wire_d25_16;
	wire [WIDTH-1:0] wire_d25_17;
	wire [WIDTH-1:0] wire_d25_18;
	wire [WIDTH-1:0] wire_d25_19;
	wire [WIDTH-1:0] wire_d25_20;
	wire [WIDTH-1:0] wire_d25_21;
	wire [WIDTH-1:0] wire_d25_22;
	wire [WIDTH-1:0] wire_d25_23;
	wire [WIDTH-1:0] wire_d25_24;
	wire [WIDTH-1:0] wire_d25_25;
	wire [WIDTH-1:0] wire_d25_26;
	wire [WIDTH-1:0] wire_d25_27;
	wire [WIDTH-1:0] wire_d25_28;
	wire [WIDTH-1:0] wire_d25_29;
	wire [WIDTH-1:0] wire_d25_30;
	wire [WIDTH-1:0] wire_d25_31;
	wire [WIDTH-1:0] wire_d25_32;
	wire [WIDTH-1:0] wire_d25_33;
	wire [WIDTH-1:0] wire_d25_34;
	wire [WIDTH-1:0] wire_d25_35;
	wire [WIDTH-1:0] wire_d25_36;
	wire [WIDTH-1:0] wire_d25_37;
	wire [WIDTH-1:0] wire_d25_38;
	wire [WIDTH-1:0] wire_d25_39;
	wire [WIDTH-1:0] wire_d25_40;
	wire [WIDTH-1:0] wire_d25_41;
	wire [WIDTH-1:0] wire_d25_42;
	wire [WIDTH-1:0] wire_d25_43;
	wire [WIDTH-1:0] wire_d25_44;
	wire [WIDTH-1:0] wire_d25_45;
	wire [WIDTH-1:0] wire_d25_46;
	wire [WIDTH-1:0] wire_d25_47;
	wire [WIDTH-1:0] wire_d25_48;
	wire [WIDTH-1:0] wire_d25_49;
	wire [WIDTH-1:0] wire_d25_50;
	wire [WIDTH-1:0] wire_d25_51;
	wire [WIDTH-1:0] wire_d25_52;
	wire [WIDTH-1:0] wire_d25_53;
	wire [WIDTH-1:0] wire_d25_54;
	wire [WIDTH-1:0] wire_d25_55;
	wire [WIDTH-1:0] wire_d25_56;
	wire [WIDTH-1:0] wire_d25_57;
	wire [WIDTH-1:0] wire_d25_58;
	wire [WIDTH-1:0] wire_d25_59;
	wire [WIDTH-1:0] wire_d25_60;
	wire [WIDTH-1:0] wire_d25_61;
	wire [WIDTH-1:0] wire_d25_62;
	wire [WIDTH-1:0] wire_d25_63;
	wire [WIDTH-1:0] wire_d25_64;
	wire [WIDTH-1:0] wire_d25_65;
	wire [WIDTH-1:0] wire_d25_66;
	wire [WIDTH-1:0] wire_d25_67;
	wire [WIDTH-1:0] wire_d25_68;
	wire [WIDTH-1:0] wire_d26_0;
	wire [WIDTH-1:0] wire_d26_1;
	wire [WIDTH-1:0] wire_d26_2;
	wire [WIDTH-1:0] wire_d26_3;
	wire [WIDTH-1:0] wire_d26_4;
	wire [WIDTH-1:0] wire_d26_5;
	wire [WIDTH-1:0] wire_d26_6;
	wire [WIDTH-1:0] wire_d26_7;
	wire [WIDTH-1:0] wire_d26_8;
	wire [WIDTH-1:0] wire_d26_9;
	wire [WIDTH-1:0] wire_d26_10;
	wire [WIDTH-1:0] wire_d26_11;
	wire [WIDTH-1:0] wire_d26_12;
	wire [WIDTH-1:0] wire_d26_13;
	wire [WIDTH-1:0] wire_d26_14;
	wire [WIDTH-1:0] wire_d26_15;
	wire [WIDTH-1:0] wire_d26_16;
	wire [WIDTH-1:0] wire_d26_17;
	wire [WIDTH-1:0] wire_d26_18;
	wire [WIDTH-1:0] wire_d26_19;
	wire [WIDTH-1:0] wire_d26_20;
	wire [WIDTH-1:0] wire_d26_21;
	wire [WIDTH-1:0] wire_d26_22;
	wire [WIDTH-1:0] wire_d26_23;
	wire [WIDTH-1:0] wire_d26_24;
	wire [WIDTH-1:0] wire_d26_25;
	wire [WIDTH-1:0] wire_d26_26;
	wire [WIDTH-1:0] wire_d26_27;
	wire [WIDTH-1:0] wire_d26_28;
	wire [WIDTH-1:0] wire_d26_29;
	wire [WIDTH-1:0] wire_d26_30;
	wire [WIDTH-1:0] wire_d26_31;
	wire [WIDTH-1:0] wire_d26_32;
	wire [WIDTH-1:0] wire_d26_33;
	wire [WIDTH-1:0] wire_d26_34;
	wire [WIDTH-1:0] wire_d26_35;
	wire [WIDTH-1:0] wire_d26_36;
	wire [WIDTH-1:0] wire_d26_37;
	wire [WIDTH-1:0] wire_d26_38;
	wire [WIDTH-1:0] wire_d26_39;
	wire [WIDTH-1:0] wire_d26_40;
	wire [WIDTH-1:0] wire_d26_41;
	wire [WIDTH-1:0] wire_d26_42;
	wire [WIDTH-1:0] wire_d26_43;
	wire [WIDTH-1:0] wire_d26_44;
	wire [WIDTH-1:0] wire_d26_45;
	wire [WIDTH-1:0] wire_d26_46;
	wire [WIDTH-1:0] wire_d26_47;
	wire [WIDTH-1:0] wire_d26_48;
	wire [WIDTH-1:0] wire_d26_49;
	wire [WIDTH-1:0] wire_d26_50;
	wire [WIDTH-1:0] wire_d26_51;
	wire [WIDTH-1:0] wire_d26_52;
	wire [WIDTH-1:0] wire_d26_53;
	wire [WIDTH-1:0] wire_d26_54;
	wire [WIDTH-1:0] wire_d26_55;
	wire [WIDTH-1:0] wire_d26_56;
	wire [WIDTH-1:0] wire_d26_57;
	wire [WIDTH-1:0] wire_d26_58;
	wire [WIDTH-1:0] wire_d26_59;
	wire [WIDTH-1:0] wire_d26_60;
	wire [WIDTH-1:0] wire_d26_61;
	wire [WIDTH-1:0] wire_d26_62;
	wire [WIDTH-1:0] wire_d26_63;
	wire [WIDTH-1:0] wire_d26_64;
	wire [WIDTH-1:0] wire_d26_65;
	wire [WIDTH-1:0] wire_d26_66;
	wire [WIDTH-1:0] wire_d26_67;
	wire [WIDTH-1:0] wire_d26_68;
	wire [WIDTH-1:0] wire_d27_0;
	wire [WIDTH-1:0] wire_d27_1;
	wire [WIDTH-1:0] wire_d27_2;
	wire [WIDTH-1:0] wire_d27_3;
	wire [WIDTH-1:0] wire_d27_4;
	wire [WIDTH-1:0] wire_d27_5;
	wire [WIDTH-1:0] wire_d27_6;
	wire [WIDTH-1:0] wire_d27_7;
	wire [WIDTH-1:0] wire_d27_8;
	wire [WIDTH-1:0] wire_d27_9;
	wire [WIDTH-1:0] wire_d27_10;
	wire [WIDTH-1:0] wire_d27_11;
	wire [WIDTH-1:0] wire_d27_12;
	wire [WIDTH-1:0] wire_d27_13;
	wire [WIDTH-1:0] wire_d27_14;
	wire [WIDTH-1:0] wire_d27_15;
	wire [WIDTH-1:0] wire_d27_16;
	wire [WIDTH-1:0] wire_d27_17;
	wire [WIDTH-1:0] wire_d27_18;
	wire [WIDTH-1:0] wire_d27_19;
	wire [WIDTH-1:0] wire_d27_20;
	wire [WIDTH-1:0] wire_d27_21;
	wire [WIDTH-1:0] wire_d27_22;
	wire [WIDTH-1:0] wire_d27_23;
	wire [WIDTH-1:0] wire_d27_24;
	wire [WIDTH-1:0] wire_d27_25;
	wire [WIDTH-1:0] wire_d27_26;
	wire [WIDTH-1:0] wire_d27_27;
	wire [WIDTH-1:0] wire_d27_28;
	wire [WIDTH-1:0] wire_d27_29;
	wire [WIDTH-1:0] wire_d27_30;
	wire [WIDTH-1:0] wire_d27_31;
	wire [WIDTH-1:0] wire_d27_32;
	wire [WIDTH-1:0] wire_d27_33;
	wire [WIDTH-1:0] wire_d27_34;
	wire [WIDTH-1:0] wire_d27_35;
	wire [WIDTH-1:0] wire_d27_36;
	wire [WIDTH-1:0] wire_d27_37;
	wire [WIDTH-1:0] wire_d27_38;
	wire [WIDTH-1:0] wire_d27_39;
	wire [WIDTH-1:0] wire_d27_40;
	wire [WIDTH-1:0] wire_d27_41;
	wire [WIDTH-1:0] wire_d27_42;
	wire [WIDTH-1:0] wire_d27_43;
	wire [WIDTH-1:0] wire_d27_44;
	wire [WIDTH-1:0] wire_d27_45;
	wire [WIDTH-1:0] wire_d27_46;
	wire [WIDTH-1:0] wire_d27_47;
	wire [WIDTH-1:0] wire_d27_48;
	wire [WIDTH-1:0] wire_d27_49;
	wire [WIDTH-1:0] wire_d27_50;
	wire [WIDTH-1:0] wire_d27_51;
	wire [WIDTH-1:0] wire_d27_52;
	wire [WIDTH-1:0] wire_d27_53;
	wire [WIDTH-1:0] wire_d27_54;
	wire [WIDTH-1:0] wire_d27_55;
	wire [WIDTH-1:0] wire_d27_56;
	wire [WIDTH-1:0] wire_d27_57;
	wire [WIDTH-1:0] wire_d27_58;
	wire [WIDTH-1:0] wire_d27_59;
	wire [WIDTH-1:0] wire_d27_60;
	wire [WIDTH-1:0] wire_d27_61;
	wire [WIDTH-1:0] wire_d27_62;
	wire [WIDTH-1:0] wire_d27_63;
	wire [WIDTH-1:0] wire_d27_64;
	wire [WIDTH-1:0] wire_d27_65;
	wire [WIDTH-1:0] wire_d27_66;
	wire [WIDTH-1:0] wire_d27_67;
	wire [WIDTH-1:0] wire_d27_68;
	wire [WIDTH-1:0] wire_d28_0;
	wire [WIDTH-1:0] wire_d28_1;
	wire [WIDTH-1:0] wire_d28_2;
	wire [WIDTH-1:0] wire_d28_3;
	wire [WIDTH-1:0] wire_d28_4;
	wire [WIDTH-1:0] wire_d28_5;
	wire [WIDTH-1:0] wire_d28_6;
	wire [WIDTH-1:0] wire_d28_7;
	wire [WIDTH-1:0] wire_d28_8;
	wire [WIDTH-1:0] wire_d28_9;
	wire [WIDTH-1:0] wire_d28_10;
	wire [WIDTH-1:0] wire_d28_11;
	wire [WIDTH-1:0] wire_d28_12;
	wire [WIDTH-1:0] wire_d28_13;
	wire [WIDTH-1:0] wire_d28_14;
	wire [WIDTH-1:0] wire_d28_15;
	wire [WIDTH-1:0] wire_d28_16;
	wire [WIDTH-1:0] wire_d28_17;
	wire [WIDTH-1:0] wire_d28_18;
	wire [WIDTH-1:0] wire_d28_19;
	wire [WIDTH-1:0] wire_d28_20;
	wire [WIDTH-1:0] wire_d28_21;
	wire [WIDTH-1:0] wire_d28_22;
	wire [WIDTH-1:0] wire_d28_23;
	wire [WIDTH-1:0] wire_d28_24;
	wire [WIDTH-1:0] wire_d28_25;
	wire [WIDTH-1:0] wire_d28_26;
	wire [WIDTH-1:0] wire_d28_27;
	wire [WIDTH-1:0] wire_d28_28;
	wire [WIDTH-1:0] wire_d28_29;
	wire [WIDTH-1:0] wire_d28_30;
	wire [WIDTH-1:0] wire_d28_31;
	wire [WIDTH-1:0] wire_d28_32;
	wire [WIDTH-1:0] wire_d28_33;
	wire [WIDTH-1:0] wire_d28_34;
	wire [WIDTH-1:0] wire_d28_35;
	wire [WIDTH-1:0] wire_d28_36;
	wire [WIDTH-1:0] wire_d28_37;
	wire [WIDTH-1:0] wire_d28_38;
	wire [WIDTH-1:0] wire_d28_39;
	wire [WIDTH-1:0] wire_d28_40;
	wire [WIDTH-1:0] wire_d28_41;
	wire [WIDTH-1:0] wire_d28_42;
	wire [WIDTH-1:0] wire_d28_43;
	wire [WIDTH-1:0] wire_d28_44;
	wire [WIDTH-1:0] wire_d28_45;
	wire [WIDTH-1:0] wire_d28_46;
	wire [WIDTH-1:0] wire_d28_47;
	wire [WIDTH-1:0] wire_d28_48;
	wire [WIDTH-1:0] wire_d28_49;
	wire [WIDTH-1:0] wire_d28_50;
	wire [WIDTH-1:0] wire_d28_51;
	wire [WIDTH-1:0] wire_d28_52;
	wire [WIDTH-1:0] wire_d28_53;
	wire [WIDTH-1:0] wire_d28_54;
	wire [WIDTH-1:0] wire_d28_55;
	wire [WIDTH-1:0] wire_d28_56;
	wire [WIDTH-1:0] wire_d28_57;
	wire [WIDTH-1:0] wire_d28_58;
	wire [WIDTH-1:0] wire_d28_59;
	wire [WIDTH-1:0] wire_d28_60;
	wire [WIDTH-1:0] wire_d28_61;
	wire [WIDTH-1:0] wire_d28_62;
	wire [WIDTH-1:0] wire_d28_63;
	wire [WIDTH-1:0] wire_d28_64;
	wire [WIDTH-1:0] wire_d28_65;
	wire [WIDTH-1:0] wire_d28_66;
	wire [WIDTH-1:0] wire_d28_67;
	wire [WIDTH-1:0] wire_d28_68;
	wire [WIDTH-1:0] wire_d29_0;
	wire [WIDTH-1:0] wire_d29_1;
	wire [WIDTH-1:0] wire_d29_2;
	wire [WIDTH-1:0] wire_d29_3;
	wire [WIDTH-1:0] wire_d29_4;
	wire [WIDTH-1:0] wire_d29_5;
	wire [WIDTH-1:0] wire_d29_6;
	wire [WIDTH-1:0] wire_d29_7;
	wire [WIDTH-1:0] wire_d29_8;
	wire [WIDTH-1:0] wire_d29_9;
	wire [WIDTH-1:0] wire_d29_10;
	wire [WIDTH-1:0] wire_d29_11;
	wire [WIDTH-1:0] wire_d29_12;
	wire [WIDTH-1:0] wire_d29_13;
	wire [WIDTH-1:0] wire_d29_14;
	wire [WIDTH-1:0] wire_d29_15;
	wire [WIDTH-1:0] wire_d29_16;
	wire [WIDTH-1:0] wire_d29_17;
	wire [WIDTH-1:0] wire_d29_18;
	wire [WIDTH-1:0] wire_d29_19;
	wire [WIDTH-1:0] wire_d29_20;
	wire [WIDTH-1:0] wire_d29_21;
	wire [WIDTH-1:0] wire_d29_22;
	wire [WIDTH-1:0] wire_d29_23;
	wire [WIDTH-1:0] wire_d29_24;
	wire [WIDTH-1:0] wire_d29_25;
	wire [WIDTH-1:0] wire_d29_26;
	wire [WIDTH-1:0] wire_d29_27;
	wire [WIDTH-1:0] wire_d29_28;
	wire [WIDTH-1:0] wire_d29_29;
	wire [WIDTH-1:0] wire_d29_30;
	wire [WIDTH-1:0] wire_d29_31;
	wire [WIDTH-1:0] wire_d29_32;
	wire [WIDTH-1:0] wire_d29_33;
	wire [WIDTH-1:0] wire_d29_34;
	wire [WIDTH-1:0] wire_d29_35;
	wire [WIDTH-1:0] wire_d29_36;
	wire [WIDTH-1:0] wire_d29_37;
	wire [WIDTH-1:0] wire_d29_38;
	wire [WIDTH-1:0] wire_d29_39;
	wire [WIDTH-1:0] wire_d29_40;
	wire [WIDTH-1:0] wire_d29_41;
	wire [WIDTH-1:0] wire_d29_42;
	wire [WIDTH-1:0] wire_d29_43;
	wire [WIDTH-1:0] wire_d29_44;
	wire [WIDTH-1:0] wire_d29_45;
	wire [WIDTH-1:0] wire_d29_46;
	wire [WIDTH-1:0] wire_d29_47;
	wire [WIDTH-1:0] wire_d29_48;
	wire [WIDTH-1:0] wire_d29_49;
	wire [WIDTH-1:0] wire_d29_50;
	wire [WIDTH-1:0] wire_d29_51;
	wire [WIDTH-1:0] wire_d29_52;
	wire [WIDTH-1:0] wire_d29_53;
	wire [WIDTH-1:0] wire_d29_54;
	wire [WIDTH-1:0] wire_d29_55;
	wire [WIDTH-1:0] wire_d29_56;
	wire [WIDTH-1:0] wire_d29_57;
	wire [WIDTH-1:0] wire_d29_58;
	wire [WIDTH-1:0] wire_d29_59;
	wire [WIDTH-1:0] wire_d29_60;
	wire [WIDTH-1:0] wire_d29_61;
	wire [WIDTH-1:0] wire_d29_62;
	wire [WIDTH-1:0] wire_d29_63;
	wire [WIDTH-1:0] wire_d29_64;
	wire [WIDTH-1:0] wire_d29_65;
	wire [WIDTH-1:0] wire_d29_66;
	wire [WIDTH-1:0] wire_d29_67;
	wire [WIDTH-1:0] wire_d29_68;
	wire [WIDTH-1:0] wire_d30_0;
	wire [WIDTH-1:0] wire_d30_1;
	wire [WIDTH-1:0] wire_d30_2;
	wire [WIDTH-1:0] wire_d30_3;
	wire [WIDTH-1:0] wire_d30_4;
	wire [WIDTH-1:0] wire_d30_5;
	wire [WIDTH-1:0] wire_d30_6;
	wire [WIDTH-1:0] wire_d30_7;
	wire [WIDTH-1:0] wire_d30_8;
	wire [WIDTH-1:0] wire_d30_9;
	wire [WIDTH-1:0] wire_d30_10;
	wire [WIDTH-1:0] wire_d30_11;
	wire [WIDTH-1:0] wire_d30_12;
	wire [WIDTH-1:0] wire_d30_13;
	wire [WIDTH-1:0] wire_d30_14;
	wire [WIDTH-1:0] wire_d30_15;
	wire [WIDTH-1:0] wire_d30_16;
	wire [WIDTH-1:0] wire_d30_17;
	wire [WIDTH-1:0] wire_d30_18;
	wire [WIDTH-1:0] wire_d30_19;
	wire [WIDTH-1:0] wire_d30_20;
	wire [WIDTH-1:0] wire_d30_21;
	wire [WIDTH-1:0] wire_d30_22;
	wire [WIDTH-1:0] wire_d30_23;
	wire [WIDTH-1:0] wire_d30_24;
	wire [WIDTH-1:0] wire_d30_25;
	wire [WIDTH-1:0] wire_d30_26;
	wire [WIDTH-1:0] wire_d30_27;
	wire [WIDTH-1:0] wire_d30_28;
	wire [WIDTH-1:0] wire_d30_29;
	wire [WIDTH-1:0] wire_d30_30;
	wire [WIDTH-1:0] wire_d30_31;
	wire [WIDTH-1:0] wire_d30_32;
	wire [WIDTH-1:0] wire_d30_33;
	wire [WIDTH-1:0] wire_d30_34;
	wire [WIDTH-1:0] wire_d30_35;
	wire [WIDTH-1:0] wire_d30_36;
	wire [WIDTH-1:0] wire_d30_37;
	wire [WIDTH-1:0] wire_d30_38;
	wire [WIDTH-1:0] wire_d30_39;
	wire [WIDTH-1:0] wire_d30_40;
	wire [WIDTH-1:0] wire_d30_41;
	wire [WIDTH-1:0] wire_d30_42;
	wire [WIDTH-1:0] wire_d30_43;
	wire [WIDTH-1:0] wire_d30_44;
	wire [WIDTH-1:0] wire_d30_45;
	wire [WIDTH-1:0] wire_d30_46;
	wire [WIDTH-1:0] wire_d30_47;
	wire [WIDTH-1:0] wire_d30_48;
	wire [WIDTH-1:0] wire_d30_49;
	wire [WIDTH-1:0] wire_d30_50;
	wire [WIDTH-1:0] wire_d30_51;
	wire [WIDTH-1:0] wire_d30_52;
	wire [WIDTH-1:0] wire_d30_53;
	wire [WIDTH-1:0] wire_d30_54;
	wire [WIDTH-1:0] wire_d30_55;
	wire [WIDTH-1:0] wire_d30_56;
	wire [WIDTH-1:0] wire_d30_57;
	wire [WIDTH-1:0] wire_d30_58;
	wire [WIDTH-1:0] wire_d30_59;
	wire [WIDTH-1:0] wire_d30_60;
	wire [WIDTH-1:0] wire_d30_61;
	wire [WIDTH-1:0] wire_d30_62;
	wire [WIDTH-1:0] wire_d30_63;
	wire [WIDTH-1:0] wire_d30_64;
	wire [WIDTH-1:0] wire_d30_65;
	wire [WIDTH-1:0] wire_d30_66;
	wire [WIDTH-1:0] wire_d30_67;
	wire [WIDTH-1:0] wire_d30_68;
	wire [WIDTH-1:0] wire_d31_0;
	wire [WIDTH-1:0] wire_d31_1;
	wire [WIDTH-1:0] wire_d31_2;
	wire [WIDTH-1:0] wire_d31_3;
	wire [WIDTH-1:0] wire_d31_4;
	wire [WIDTH-1:0] wire_d31_5;
	wire [WIDTH-1:0] wire_d31_6;
	wire [WIDTH-1:0] wire_d31_7;
	wire [WIDTH-1:0] wire_d31_8;
	wire [WIDTH-1:0] wire_d31_9;
	wire [WIDTH-1:0] wire_d31_10;
	wire [WIDTH-1:0] wire_d31_11;
	wire [WIDTH-1:0] wire_d31_12;
	wire [WIDTH-1:0] wire_d31_13;
	wire [WIDTH-1:0] wire_d31_14;
	wire [WIDTH-1:0] wire_d31_15;
	wire [WIDTH-1:0] wire_d31_16;
	wire [WIDTH-1:0] wire_d31_17;
	wire [WIDTH-1:0] wire_d31_18;
	wire [WIDTH-1:0] wire_d31_19;
	wire [WIDTH-1:0] wire_d31_20;
	wire [WIDTH-1:0] wire_d31_21;
	wire [WIDTH-1:0] wire_d31_22;
	wire [WIDTH-1:0] wire_d31_23;
	wire [WIDTH-1:0] wire_d31_24;
	wire [WIDTH-1:0] wire_d31_25;
	wire [WIDTH-1:0] wire_d31_26;
	wire [WIDTH-1:0] wire_d31_27;
	wire [WIDTH-1:0] wire_d31_28;
	wire [WIDTH-1:0] wire_d31_29;
	wire [WIDTH-1:0] wire_d31_30;
	wire [WIDTH-1:0] wire_d31_31;
	wire [WIDTH-1:0] wire_d31_32;
	wire [WIDTH-1:0] wire_d31_33;
	wire [WIDTH-1:0] wire_d31_34;
	wire [WIDTH-1:0] wire_d31_35;
	wire [WIDTH-1:0] wire_d31_36;
	wire [WIDTH-1:0] wire_d31_37;
	wire [WIDTH-1:0] wire_d31_38;
	wire [WIDTH-1:0] wire_d31_39;
	wire [WIDTH-1:0] wire_d31_40;
	wire [WIDTH-1:0] wire_d31_41;
	wire [WIDTH-1:0] wire_d31_42;
	wire [WIDTH-1:0] wire_d31_43;
	wire [WIDTH-1:0] wire_d31_44;
	wire [WIDTH-1:0] wire_d31_45;
	wire [WIDTH-1:0] wire_d31_46;
	wire [WIDTH-1:0] wire_d31_47;
	wire [WIDTH-1:0] wire_d31_48;
	wire [WIDTH-1:0] wire_d31_49;
	wire [WIDTH-1:0] wire_d31_50;
	wire [WIDTH-1:0] wire_d31_51;
	wire [WIDTH-1:0] wire_d31_52;
	wire [WIDTH-1:0] wire_d31_53;
	wire [WIDTH-1:0] wire_d31_54;
	wire [WIDTH-1:0] wire_d31_55;
	wire [WIDTH-1:0] wire_d31_56;
	wire [WIDTH-1:0] wire_d31_57;
	wire [WIDTH-1:0] wire_d31_58;
	wire [WIDTH-1:0] wire_d31_59;
	wire [WIDTH-1:0] wire_d31_60;
	wire [WIDTH-1:0] wire_d31_61;
	wire [WIDTH-1:0] wire_d31_62;
	wire [WIDTH-1:0] wire_d31_63;
	wire [WIDTH-1:0] wire_d31_64;
	wire [WIDTH-1:0] wire_d31_65;
	wire [WIDTH-1:0] wire_d31_66;
	wire [WIDTH-1:0] wire_d31_67;
	wire [WIDTH-1:0] wire_d31_68;
	wire [WIDTH-1:0] wire_d32_0;
	wire [WIDTH-1:0] wire_d32_1;
	wire [WIDTH-1:0] wire_d32_2;
	wire [WIDTH-1:0] wire_d32_3;
	wire [WIDTH-1:0] wire_d32_4;
	wire [WIDTH-1:0] wire_d32_5;
	wire [WIDTH-1:0] wire_d32_6;
	wire [WIDTH-1:0] wire_d32_7;
	wire [WIDTH-1:0] wire_d32_8;
	wire [WIDTH-1:0] wire_d32_9;
	wire [WIDTH-1:0] wire_d32_10;
	wire [WIDTH-1:0] wire_d32_11;
	wire [WIDTH-1:0] wire_d32_12;
	wire [WIDTH-1:0] wire_d32_13;
	wire [WIDTH-1:0] wire_d32_14;
	wire [WIDTH-1:0] wire_d32_15;
	wire [WIDTH-1:0] wire_d32_16;
	wire [WIDTH-1:0] wire_d32_17;
	wire [WIDTH-1:0] wire_d32_18;
	wire [WIDTH-1:0] wire_d32_19;
	wire [WIDTH-1:0] wire_d32_20;
	wire [WIDTH-1:0] wire_d32_21;
	wire [WIDTH-1:0] wire_d32_22;
	wire [WIDTH-1:0] wire_d32_23;
	wire [WIDTH-1:0] wire_d32_24;
	wire [WIDTH-1:0] wire_d32_25;
	wire [WIDTH-1:0] wire_d32_26;
	wire [WIDTH-1:0] wire_d32_27;
	wire [WIDTH-1:0] wire_d32_28;
	wire [WIDTH-1:0] wire_d32_29;
	wire [WIDTH-1:0] wire_d32_30;
	wire [WIDTH-1:0] wire_d32_31;
	wire [WIDTH-1:0] wire_d32_32;
	wire [WIDTH-1:0] wire_d32_33;
	wire [WIDTH-1:0] wire_d32_34;
	wire [WIDTH-1:0] wire_d32_35;
	wire [WIDTH-1:0] wire_d32_36;
	wire [WIDTH-1:0] wire_d32_37;
	wire [WIDTH-1:0] wire_d32_38;
	wire [WIDTH-1:0] wire_d32_39;
	wire [WIDTH-1:0] wire_d32_40;
	wire [WIDTH-1:0] wire_d32_41;
	wire [WIDTH-1:0] wire_d32_42;
	wire [WIDTH-1:0] wire_d32_43;
	wire [WIDTH-1:0] wire_d32_44;
	wire [WIDTH-1:0] wire_d32_45;
	wire [WIDTH-1:0] wire_d32_46;
	wire [WIDTH-1:0] wire_d32_47;
	wire [WIDTH-1:0] wire_d32_48;
	wire [WIDTH-1:0] wire_d32_49;
	wire [WIDTH-1:0] wire_d32_50;
	wire [WIDTH-1:0] wire_d32_51;
	wire [WIDTH-1:0] wire_d32_52;
	wire [WIDTH-1:0] wire_d32_53;
	wire [WIDTH-1:0] wire_d32_54;
	wire [WIDTH-1:0] wire_d32_55;
	wire [WIDTH-1:0] wire_d32_56;
	wire [WIDTH-1:0] wire_d32_57;
	wire [WIDTH-1:0] wire_d32_58;
	wire [WIDTH-1:0] wire_d32_59;
	wire [WIDTH-1:0] wire_d32_60;
	wire [WIDTH-1:0] wire_d32_61;
	wire [WIDTH-1:0] wire_d32_62;
	wire [WIDTH-1:0] wire_d32_63;
	wire [WIDTH-1:0] wire_d32_64;
	wire [WIDTH-1:0] wire_d32_65;
	wire [WIDTH-1:0] wire_d32_66;
	wire [WIDTH-1:0] wire_d32_67;
	wire [WIDTH-1:0] wire_d32_68;
	wire [WIDTH-1:0] wire_d33_0;
	wire [WIDTH-1:0] wire_d33_1;
	wire [WIDTH-1:0] wire_d33_2;
	wire [WIDTH-1:0] wire_d33_3;
	wire [WIDTH-1:0] wire_d33_4;
	wire [WIDTH-1:0] wire_d33_5;
	wire [WIDTH-1:0] wire_d33_6;
	wire [WIDTH-1:0] wire_d33_7;
	wire [WIDTH-1:0] wire_d33_8;
	wire [WIDTH-1:0] wire_d33_9;
	wire [WIDTH-1:0] wire_d33_10;
	wire [WIDTH-1:0] wire_d33_11;
	wire [WIDTH-1:0] wire_d33_12;
	wire [WIDTH-1:0] wire_d33_13;
	wire [WIDTH-1:0] wire_d33_14;
	wire [WIDTH-1:0] wire_d33_15;
	wire [WIDTH-1:0] wire_d33_16;
	wire [WIDTH-1:0] wire_d33_17;
	wire [WIDTH-1:0] wire_d33_18;
	wire [WIDTH-1:0] wire_d33_19;
	wire [WIDTH-1:0] wire_d33_20;
	wire [WIDTH-1:0] wire_d33_21;
	wire [WIDTH-1:0] wire_d33_22;
	wire [WIDTH-1:0] wire_d33_23;
	wire [WIDTH-1:0] wire_d33_24;
	wire [WIDTH-1:0] wire_d33_25;
	wire [WIDTH-1:0] wire_d33_26;
	wire [WIDTH-1:0] wire_d33_27;
	wire [WIDTH-1:0] wire_d33_28;
	wire [WIDTH-1:0] wire_d33_29;
	wire [WIDTH-1:0] wire_d33_30;
	wire [WIDTH-1:0] wire_d33_31;
	wire [WIDTH-1:0] wire_d33_32;
	wire [WIDTH-1:0] wire_d33_33;
	wire [WIDTH-1:0] wire_d33_34;
	wire [WIDTH-1:0] wire_d33_35;
	wire [WIDTH-1:0] wire_d33_36;
	wire [WIDTH-1:0] wire_d33_37;
	wire [WIDTH-1:0] wire_d33_38;
	wire [WIDTH-1:0] wire_d33_39;
	wire [WIDTH-1:0] wire_d33_40;
	wire [WIDTH-1:0] wire_d33_41;
	wire [WIDTH-1:0] wire_d33_42;
	wire [WIDTH-1:0] wire_d33_43;
	wire [WIDTH-1:0] wire_d33_44;
	wire [WIDTH-1:0] wire_d33_45;
	wire [WIDTH-1:0] wire_d33_46;
	wire [WIDTH-1:0] wire_d33_47;
	wire [WIDTH-1:0] wire_d33_48;
	wire [WIDTH-1:0] wire_d33_49;
	wire [WIDTH-1:0] wire_d33_50;
	wire [WIDTH-1:0] wire_d33_51;
	wire [WIDTH-1:0] wire_d33_52;
	wire [WIDTH-1:0] wire_d33_53;
	wire [WIDTH-1:0] wire_d33_54;
	wire [WIDTH-1:0] wire_d33_55;
	wire [WIDTH-1:0] wire_d33_56;
	wire [WIDTH-1:0] wire_d33_57;
	wire [WIDTH-1:0] wire_d33_58;
	wire [WIDTH-1:0] wire_d33_59;
	wire [WIDTH-1:0] wire_d33_60;
	wire [WIDTH-1:0] wire_d33_61;
	wire [WIDTH-1:0] wire_d33_62;
	wire [WIDTH-1:0] wire_d33_63;
	wire [WIDTH-1:0] wire_d33_64;
	wire [WIDTH-1:0] wire_d33_65;
	wire [WIDTH-1:0] wire_d33_66;
	wire [WIDTH-1:0] wire_d33_67;
	wire [WIDTH-1:0] wire_d33_68;
	wire [WIDTH-1:0] wire_d34_0;
	wire [WIDTH-1:0] wire_d34_1;
	wire [WIDTH-1:0] wire_d34_2;
	wire [WIDTH-1:0] wire_d34_3;
	wire [WIDTH-1:0] wire_d34_4;
	wire [WIDTH-1:0] wire_d34_5;
	wire [WIDTH-1:0] wire_d34_6;
	wire [WIDTH-1:0] wire_d34_7;
	wire [WIDTH-1:0] wire_d34_8;
	wire [WIDTH-1:0] wire_d34_9;
	wire [WIDTH-1:0] wire_d34_10;
	wire [WIDTH-1:0] wire_d34_11;
	wire [WIDTH-1:0] wire_d34_12;
	wire [WIDTH-1:0] wire_d34_13;
	wire [WIDTH-1:0] wire_d34_14;
	wire [WIDTH-1:0] wire_d34_15;
	wire [WIDTH-1:0] wire_d34_16;
	wire [WIDTH-1:0] wire_d34_17;
	wire [WIDTH-1:0] wire_d34_18;
	wire [WIDTH-1:0] wire_d34_19;
	wire [WIDTH-1:0] wire_d34_20;
	wire [WIDTH-1:0] wire_d34_21;
	wire [WIDTH-1:0] wire_d34_22;
	wire [WIDTH-1:0] wire_d34_23;
	wire [WIDTH-1:0] wire_d34_24;
	wire [WIDTH-1:0] wire_d34_25;
	wire [WIDTH-1:0] wire_d34_26;
	wire [WIDTH-1:0] wire_d34_27;
	wire [WIDTH-1:0] wire_d34_28;
	wire [WIDTH-1:0] wire_d34_29;
	wire [WIDTH-1:0] wire_d34_30;
	wire [WIDTH-1:0] wire_d34_31;
	wire [WIDTH-1:0] wire_d34_32;
	wire [WIDTH-1:0] wire_d34_33;
	wire [WIDTH-1:0] wire_d34_34;
	wire [WIDTH-1:0] wire_d34_35;
	wire [WIDTH-1:0] wire_d34_36;
	wire [WIDTH-1:0] wire_d34_37;
	wire [WIDTH-1:0] wire_d34_38;
	wire [WIDTH-1:0] wire_d34_39;
	wire [WIDTH-1:0] wire_d34_40;
	wire [WIDTH-1:0] wire_d34_41;
	wire [WIDTH-1:0] wire_d34_42;
	wire [WIDTH-1:0] wire_d34_43;
	wire [WIDTH-1:0] wire_d34_44;
	wire [WIDTH-1:0] wire_d34_45;
	wire [WIDTH-1:0] wire_d34_46;
	wire [WIDTH-1:0] wire_d34_47;
	wire [WIDTH-1:0] wire_d34_48;
	wire [WIDTH-1:0] wire_d34_49;
	wire [WIDTH-1:0] wire_d34_50;
	wire [WIDTH-1:0] wire_d34_51;
	wire [WIDTH-1:0] wire_d34_52;
	wire [WIDTH-1:0] wire_d34_53;
	wire [WIDTH-1:0] wire_d34_54;
	wire [WIDTH-1:0] wire_d34_55;
	wire [WIDTH-1:0] wire_d34_56;
	wire [WIDTH-1:0] wire_d34_57;
	wire [WIDTH-1:0] wire_d34_58;
	wire [WIDTH-1:0] wire_d34_59;
	wire [WIDTH-1:0] wire_d34_60;
	wire [WIDTH-1:0] wire_d34_61;
	wire [WIDTH-1:0] wire_d34_62;
	wire [WIDTH-1:0] wire_d34_63;
	wire [WIDTH-1:0] wire_d34_64;
	wire [WIDTH-1:0] wire_d34_65;
	wire [WIDTH-1:0] wire_d34_66;
	wire [WIDTH-1:0] wire_d34_67;
	wire [WIDTH-1:0] wire_d34_68;
	wire [WIDTH-1:0] wire_d35_0;
	wire [WIDTH-1:0] wire_d35_1;
	wire [WIDTH-1:0] wire_d35_2;
	wire [WIDTH-1:0] wire_d35_3;
	wire [WIDTH-1:0] wire_d35_4;
	wire [WIDTH-1:0] wire_d35_5;
	wire [WIDTH-1:0] wire_d35_6;
	wire [WIDTH-1:0] wire_d35_7;
	wire [WIDTH-1:0] wire_d35_8;
	wire [WIDTH-1:0] wire_d35_9;
	wire [WIDTH-1:0] wire_d35_10;
	wire [WIDTH-1:0] wire_d35_11;
	wire [WIDTH-1:0] wire_d35_12;
	wire [WIDTH-1:0] wire_d35_13;
	wire [WIDTH-1:0] wire_d35_14;
	wire [WIDTH-1:0] wire_d35_15;
	wire [WIDTH-1:0] wire_d35_16;
	wire [WIDTH-1:0] wire_d35_17;
	wire [WIDTH-1:0] wire_d35_18;
	wire [WIDTH-1:0] wire_d35_19;
	wire [WIDTH-1:0] wire_d35_20;
	wire [WIDTH-1:0] wire_d35_21;
	wire [WIDTH-1:0] wire_d35_22;
	wire [WIDTH-1:0] wire_d35_23;
	wire [WIDTH-1:0] wire_d35_24;
	wire [WIDTH-1:0] wire_d35_25;
	wire [WIDTH-1:0] wire_d35_26;
	wire [WIDTH-1:0] wire_d35_27;
	wire [WIDTH-1:0] wire_d35_28;
	wire [WIDTH-1:0] wire_d35_29;
	wire [WIDTH-1:0] wire_d35_30;
	wire [WIDTH-1:0] wire_d35_31;
	wire [WIDTH-1:0] wire_d35_32;
	wire [WIDTH-1:0] wire_d35_33;
	wire [WIDTH-1:0] wire_d35_34;
	wire [WIDTH-1:0] wire_d35_35;
	wire [WIDTH-1:0] wire_d35_36;
	wire [WIDTH-1:0] wire_d35_37;
	wire [WIDTH-1:0] wire_d35_38;
	wire [WIDTH-1:0] wire_d35_39;
	wire [WIDTH-1:0] wire_d35_40;
	wire [WIDTH-1:0] wire_d35_41;
	wire [WIDTH-1:0] wire_d35_42;
	wire [WIDTH-1:0] wire_d35_43;
	wire [WIDTH-1:0] wire_d35_44;
	wire [WIDTH-1:0] wire_d35_45;
	wire [WIDTH-1:0] wire_d35_46;
	wire [WIDTH-1:0] wire_d35_47;
	wire [WIDTH-1:0] wire_d35_48;
	wire [WIDTH-1:0] wire_d35_49;
	wire [WIDTH-1:0] wire_d35_50;
	wire [WIDTH-1:0] wire_d35_51;
	wire [WIDTH-1:0] wire_d35_52;
	wire [WIDTH-1:0] wire_d35_53;
	wire [WIDTH-1:0] wire_d35_54;
	wire [WIDTH-1:0] wire_d35_55;
	wire [WIDTH-1:0] wire_d35_56;
	wire [WIDTH-1:0] wire_d35_57;
	wire [WIDTH-1:0] wire_d35_58;
	wire [WIDTH-1:0] wire_d35_59;
	wire [WIDTH-1:0] wire_d35_60;
	wire [WIDTH-1:0] wire_d35_61;
	wire [WIDTH-1:0] wire_d35_62;
	wire [WIDTH-1:0] wire_d35_63;
	wire [WIDTH-1:0] wire_d35_64;
	wire [WIDTH-1:0] wire_d35_65;
	wire [WIDTH-1:0] wire_d35_66;
	wire [WIDTH-1:0] wire_d35_67;
	wire [WIDTH-1:0] wire_d35_68;
	wire [WIDTH-1:0] wire_d36_0;
	wire [WIDTH-1:0] wire_d36_1;
	wire [WIDTH-1:0] wire_d36_2;
	wire [WIDTH-1:0] wire_d36_3;
	wire [WIDTH-1:0] wire_d36_4;
	wire [WIDTH-1:0] wire_d36_5;
	wire [WIDTH-1:0] wire_d36_6;
	wire [WIDTH-1:0] wire_d36_7;
	wire [WIDTH-1:0] wire_d36_8;
	wire [WIDTH-1:0] wire_d36_9;
	wire [WIDTH-1:0] wire_d36_10;
	wire [WIDTH-1:0] wire_d36_11;
	wire [WIDTH-1:0] wire_d36_12;
	wire [WIDTH-1:0] wire_d36_13;
	wire [WIDTH-1:0] wire_d36_14;
	wire [WIDTH-1:0] wire_d36_15;
	wire [WIDTH-1:0] wire_d36_16;
	wire [WIDTH-1:0] wire_d36_17;
	wire [WIDTH-1:0] wire_d36_18;
	wire [WIDTH-1:0] wire_d36_19;
	wire [WIDTH-1:0] wire_d36_20;
	wire [WIDTH-1:0] wire_d36_21;
	wire [WIDTH-1:0] wire_d36_22;
	wire [WIDTH-1:0] wire_d36_23;
	wire [WIDTH-1:0] wire_d36_24;
	wire [WIDTH-1:0] wire_d36_25;
	wire [WIDTH-1:0] wire_d36_26;
	wire [WIDTH-1:0] wire_d36_27;
	wire [WIDTH-1:0] wire_d36_28;
	wire [WIDTH-1:0] wire_d36_29;
	wire [WIDTH-1:0] wire_d36_30;
	wire [WIDTH-1:0] wire_d36_31;
	wire [WIDTH-1:0] wire_d36_32;
	wire [WIDTH-1:0] wire_d36_33;
	wire [WIDTH-1:0] wire_d36_34;
	wire [WIDTH-1:0] wire_d36_35;
	wire [WIDTH-1:0] wire_d36_36;
	wire [WIDTH-1:0] wire_d36_37;
	wire [WIDTH-1:0] wire_d36_38;
	wire [WIDTH-1:0] wire_d36_39;
	wire [WIDTH-1:0] wire_d36_40;
	wire [WIDTH-1:0] wire_d36_41;
	wire [WIDTH-1:0] wire_d36_42;
	wire [WIDTH-1:0] wire_d36_43;
	wire [WIDTH-1:0] wire_d36_44;
	wire [WIDTH-1:0] wire_d36_45;
	wire [WIDTH-1:0] wire_d36_46;
	wire [WIDTH-1:0] wire_d36_47;
	wire [WIDTH-1:0] wire_d36_48;
	wire [WIDTH-1:0] wire_d36_49;
	wire [WIDTH-1:0] wire_d36_50;
	wire [WIDTH-1:0] wire_d36_51;
	wire [WIDTH-1:0] wire_d36_52;
	wire [WIDTH-1:0] wire_d36_53;
	wire [WIDTH-1:0] wire_d36_54;
	wire [WIDTH-1:0] wire_d36_55;
	wire [WIDTH-1:0] wire_d36_56;
	wire [WIDTH-1:0] wire_d36_57;
	wire [WIDTH-1:0] wire_d36_58;
	wire [WIDTH-1:0] wire_d36_59;
	wire [WIDTH-1:0] wire_d36_60;
	wire [WIDTH-1:0] wire_d36_61;
	wire [WIDTH-1:0] wire_d36_62;
	wire [WIDTH-1:0] wire_d36_63;
	wire [WIDTH-1:0] wire_d36_64;
	wire [WIDTH-1:0] wire_d36_65;
	wire [WIDTH-1:0] wire_d36_66;
	wire [WIDTH-1:0] wire_d36_67;
	wire [WIDTH-1:0] wire_d36_68;
	wire [WIDTH-1:0] wire_d37_0;
	wire [WIDTH-1:0] wire_d37_1;
	wire [WIDTH-1:0] wire_d37_2;
	wire [WIDTH-1:0] wire_d37_3;
	wire [WIDTH-1:0] wire_d37_4;
	wire [WIDTH-1:0] wire_d37_5;
	wire [WIDTH-1:0] wire_d37_6;
	wire [WIDTH-1:0] wire_d37_7;
	wire [WIDTH-1:0] wire_d37_8;
	wire [WIDTH-1:0] wire_d37_9;
	wire [WIDTH-1:0] wire_d37_10;
	wire [WIDTH-1:0] wire_d37_11;
	wire [WIDTH-1:0] wire_d37_12;
	wire [WIDTH-1:0] wire_d37_13;
	wire [WIDTH-1:0] wire_d37_14;
	wire [WIDTH-1:0] wire_d37_15;
	wire [WIDTH-1:0] wire_d37_16;
	wire [WIDTH-1:0] wire_d37_17;
	wire [WIDTH-1:0] wire_d37_18;
	wire [WIDTH-1:0] wire_d37_19;
	wire [WIDTH-1:0] wire_d37_20;
	wire [WIDTH-1:0] wire_d37_21;
	wire [WIDTH-1:0] wire_d37_22;
	wire [WIDTH-1:0] wire_d37_23;
	wire [WIDTH-1:0] wire_d37_24;
	wire [WIDTH-1:0] wire_d37_25;
	wire [WIDTH-1:0] wire_d37_26;
	wire [WIDTH-1:0] wire_d37_27;
	wire [WIDTH-1:0] wire_d37_28;
	wire [WIDTH-1:0] wire_d37_29;
	wire [WIDTH-1:0] wire_d37_30;
	wire [WIDTH-1:0] wire_d37_31;
	wire [WIDTH-1:0] wire_d37_32;
	wire [WIDTH-1:0] wire_d37_33;
	wire [WIDTH-1:0] wire_d37_34;
	wire [WIDTH-1:0] wire_d37_35;
	wire [WIDTH-1:0] wire_d37_36;
	wire [WIDTH-1:0] wire_d37_37;
	wire [WIDTH-1:0] wire_d37_38;
	wire [WIDTH-1:0] wire_d37_39;
	wire [WIDTH-1:0] wire_d37_40;
	wire [WIDTH-1:0] wire_d37_41;
	wire [WIDTH-1:0] wire_d37_42;
	wire [WIDTH-1:0] wire_d37_43;
	wire [WIDTH-1:0] wire_d37_44;
	wire [WIDTH-1:0] wire_d37_45;
	wire [WIDTH-1:0] wire_d37_46;
	wire [WIDTH-1:0] wire_d37_47;
	wire [WIDTH-1:0] wire_d37_48;
	wire [WIDTH-1:0] wire_d37_49;
	wire [WIDTH-1:0] wire_d37_50;
	wire [WIDTH-1:0] wire_d37_51;
	wire [WIDTH-1:0] wire_d37_52;
	wire [WIDTH-1:0] wire_d37_53;
	wire [WIDTH-1:0] wire_d37_54;
	wire [WIDTH-1:0] wire_d37_55;
	wire [WIDTH-1:0] wire_d37_56;
	wire [WIDTH-1:0] wire_d37_57;
	wire [WIDTH-1:0] wire_d37_58;
	wire [WIDTH-1:0] wire_d37_59;
	wire [WIDTH-1:0] wire_d37_60;
	wire [WIDTH-1:0] wire_d37_61;
	wire [WIDTH-1:0] wire_d37_62;
	wire [WIDTH-1:0] wire_d37_63;
	wire [WIDTH-1:0] wire_d37_64;
	wire [WIDTH-1:0] wire_d37_65;
	wire [WIDTH-1:0] wire_d37_66;
	wire [WIDTH-1:0] wire_d37_67;
	wire [WIDTH-1:0] wire_d37_68;
	wire [WIDTH-1:0] wire_d38_0;
	wire [WIDTH-1:0] wire_d38_1;
	wire [WIDTH-1:0] wire_d38_2;
	wire [WIDTH-1:0] wire_d38_3;
	wire [WIDTH-1:0] wire_d38_4;
	wire [WIDTH-1:0] wire_d38_5;
	wire [WIDTH-1:0] wire_d38_6;
	wire [WIDTH-1:0] wire_d38_7;
	wire [WIDTH-1:0] wire_d38_8;
	wire [WIDTH-1:0] wire_d38_9;
	wire [WIDTH-1:0] wire_d38_10;
	wire [WIDTH-1:0] wire_d38_11;
	wire [WIDTH-1:0] wire_d38_12;
	wire [WIDTH-1:0] wire_d38_13;
	wire [WIDTH-1:0] wire_d38_14;
	wire [WIDTH-1:0] wire_d38_15;
	wire [WIDTH-1:0] wire_d38_16;
	wire [WIDTH-1:0] wire_d38_17;
	wire [WIDTH-1:0] wire_d38_18;
	wire [WIDTH-1:0] wire_d38_19;
	wire [WIDTH-1:0] wire_d38_20;
	wire [WIDTH-1:0] wire_d38_21;
	wire [WIDTH-1:0] wire_d38_22;
	wire [WIDTH-1:0] wire_d38_23;
	wire [WIDTH-1:0] wire_d38_24;
	wire [WIDTH-1:0] wire_d38_25;
	wire [WIDTH-1:0] wire_d38_26;
	wire [WIDTH-1:0] wire_d38_27;
	wire [WIDTH-1:0] wire_d38_28;
	wire [WIDTH-1:0] wire_d38_29;
	wire [WIDTH-1:0] wire_d38_30;
	wire [WIDTH-1:0] wire_d38_31;
	wire [WIDTH-1:0] wire_d38_32;
	wire [WIDTH-1:0] wire_d38_33;
	wire [WIDTH-1:0] wire_d38_34;
	wire [WIDTH-1:0] wire_d38_35;
	wire [WIDTH-1:0] wire_d38_36;
	wire [WIDTH-1:0] wire_d38_37;
	wire [WIDTH-1:0] wire_d38_38;
	wire [WIDTH-1:0] wire_d38_39;
	wire [WIDTH-1:0] wire_d38_40;
	wire [WIDTH-1:0] wire_d38_41;
	wire [WIDTH-1:0] wire_d38_42;
	wire [WIDTH-1:0] wire_d38_43;
	wire [WIDTH-1:0] wire_d38_44;
	wire [WIDTH-1:0] wire_d38_45;
	wire [WIDTH-1:0] wire_d38_46;
	wire [WIDTH-1:0] wire_d38_47;
	wire [WIDTH-1:0] wire_d38_48;
	wire [WIDTH-1:0] wire_d38_49;
	wire [WIDTH-1:0] wire_d38_50;
	wire [WIDTH-1:0] wire_d38_51;
	wire [WIDTH-1:0] wire_d38_52;
	wire [WIDTH-1:0] wire_d38_53;
	wire [WIDTH-1:0] wire_d38_54;
	wire [WIDTH-1:0] wire_d38_55;
	wire [WIDTH-1:0] wire_d38_56;
	wire [WIDTH-1:0] wire_d38_57;
	wire [WIDTH-1:0] wire_d38_58;
	wire [WIDTH-1:0] wire_d38_59;
	wire [WIDTH-1:0] wire_d38_60;
	wire [WIDTH-1:0] wire_d38_61;
	wire [WIDTH-1:0] wire_d38_62;
	wire [WIDTH-1:0] wire_d38_63;
	wire [WIDTH-1:0] wire_d38_64;
	wire [WIDTH-1:0] wire_d38_65;
	wire [WIDTH-1:0] wire_d38_66;
	wire [WIDTH-1:0] wire_d38_67;
	wire [WIDTH-1:0] wire_d38_68;
	wire [WIDTH-1:0] wire_d39_0;
	wire [WIDTH-1:0] wire_d39_1;
	wire [WIDTH-1:0] wire_d39_2;
	wire [WIDTH-1:0] wire_d39_3;
	wire [WIDTH-1:0] wire_d39_4;
	wire [WIDTH-1:0] wire_d39_5;
	wire [WIDTH-1:0] wire_d39_6;
	wire [WIDTH-1:0] wire_d39_7;
	wire [WIDTH-1:0] wire_d39_8;
	wire [WIDTH-1:0] wire_d39_9;
	wire [WIDTH-1:0] wire_d39_10;
	wire [WIDTH-1:0] wire_d39_11;
	wire [WIDTH-1:0] wire_d39_12;
	wire [WIDTH-1:0] wire_d39_13;
	wire [WIDTH-1:0] wire_d39_14;
	wire [WIDTH-1:0] wire_d39_15;
	wire [WIDTH-1:0] wire_d39_16;
	wire [WIDTH-1:0] wire_d39_17;
	wire [WIDTH-1:0] wire_d39_18;
	wire [WIDTH-1:0] wire_d39_19;
	wire [WIDTH-1:0] wire_d39_20;
	wire [WIDTH-1:0] wire_d39_21;
	wire [WIDTH-1:0] wire_d39_22;
	wire [WIDTH-1:0] wire_d39_23;
	wire [WIDTH-1:0] wire_d39_24;
	wire [WIDTH-1:0] wire_d39_25;
	wire [WIDTH-1:0] wire_d39_26;
	wire [WIDTH-1:0] wire_d39_27;
	wire [WIDTH-1:0] wire_d39_28;
	wire [WIDTH-1:0] wire_d39_29;
	wire [WIDTH-1:0] wire_d39_30;
	wire [WIDTH-1:0] wire_d39_31;
	wire [WIDTH-1:0] wire_d39_32;
	wire [WIDTH-1:0] wire_d39_33;
	wire [WIDTH-1:0] wire_d39_34;
	wire [WIDTH-1:0] wire_d39_35;
	wire [WIDTH-1:0] wire_d39_36;
	wire [WIDTH-1:0] wire_d39_37;
	wire [WIDTH-1:0] wire_d39_38;
	wire [WIDTH-1:0] wire_d39_39;
	wire [WIDTH-1:0] wire_d39_40;
	wire [WIDTH-1:0] wire_d39_41;
	wire [WIDTH-1:0] wire_d39_42;
	wire [WIDTH-1:0] wire_d39_43;
	wire [WIDTH-1:0] wire_d39_44;
	wire [WIDTH-1:0] wire_d39_45;
	wire [WIDTH-1:0] wire_d39_46;
	wire [WIDTH-1:0] wire_d39_47;
	wire [WIDTH-1:0] wire_d39_48;
	wire [WIDTH-1:0] wire_d39_49;
	wire [WIDTH-1:0] wire_d39_50;
	wire [WIDTH-1:0] wire_d39_51;
	wire [WIDTH-1:0] wire_d39_52;
	wire [WIDTH-1:0] wire_d39_53;
	wire [WIDTH-1:0] wire_d39_54;
	wire [WIDTH-1:0] wire_d39_55;
	wire [WIDTH-1:0] wire_d39_56;
	wire [WIDTH-1:0] wire_d39_57;
	wire [WIDTH-1:0] wire_d39_58;
	wire [WIDTH-1:0] wire_d39_59;
	wire [WIDTH-1:0] wire_d39_60;
	wire [WIDTH-1:0] wire_d39_61;
	wire [WIDTH-1:0] wire_d39_62;
	wire [WIDTH-1:0] wire_d39_63;
	wire [WIDTH-1:0] wire_d39_64;
	wire [WIDTH-1:0] wire_d39_65;
	wire [WIDTH-1:0] wire_d39_66;
	wire [WIDTH-1:0] wire_d39_67;
	wire [WIDTH-1:0] wire_d39_68;
	wire [WIDTH-1:0] wire_d40_0;
	wire [WIDTH-1:0] wire_d40_1;
	wire [WIDTH-1:0] wire_d40_2;
	wire [WIDTH-1:0] wire_d40_3;
	wire [WIDTH-1:0] wire_d40_4;
	wire [WIDTH-1:0] wire_d40_5;
	wire [WIDTH-1:0] wire_d40_6;
	wire [WIDTH-1:0] wire_d40_7;
	wire [WIDTH-1:0] wire_d40_8;
	wire [WIDTH-1:0] wire_d40_9;
	wire [WIDTH-1:0] wire_d40_10;
	wire [WIDTH-1:0] wire_d40_11;
	wire [WIDTH-1:0] wire_d40_12;
	wire [WIDTH-1:0] wire_d40_13;
	wire [WIDTH-1:0] wire_d40_14;
	wire [WIDTH-1:0] wire_d40_15;
	wire [WIDTH-1:0] wire_d40_16;
	wire [WIDTH-1:0] wire_d40_17;
	wire [WIDTH-1:0] wire_d40_18;
	wire [WIDTH-1:0] wire_d40_19;
	wire [WIDTH-1:0] wire_d40_20;
	wire [WIDTH-1:0] wire_d40_21;
	wire [WIDTH-1:0] wire_d40_22;
	wire [WIDTH-1:0] wire_d40_23;
	wire [WIDTH-1:0] wire_d40_24;
	wire [WIDTH-1:0] wire_d40_25;
	wire [WIDTH-1:0] wire_d40_26;
	wire [WIDTH-1:0] wire_d40_27;
	wire [WIDTH-1:0] wire_d40_28;
	wire [WIDTH-1:0] wire_d40_29;
	wire [WIDTH-1:0] wire_d40_30;
	wire [WIDTH-1:0] wire_d40_31;
	wire [WIDTH-1:0] wire_d40_32;
	wire [WIDTH-1:0] wire_d40_33;
	wire [WIDTH-1:0] wire_d40_34;
	wire [WIDTH-1:0] wire_d40_35;
	wire [WIDTH-1:0] wire_d40_36;
	wire [WIDTH-1:0] wire_d40_37;
	wire [WIDTH-1:0] wire_d40_38;
	wire [WIDTH-1:0] wire_d40_39;
	wire [WIDTH-1:0] wire_d40_40;
	wire [WIDTH-1:0] wire_d40_41;
	wire [WIDTH-1:0] wire_d40_42;
	wire [WIDTH-1:0] wire_d40_43;
	wire [WIDTH-1:0] wire_d40_44;
	wire [WIDTH-1:0] wire_d40_45;
	wire [WIDTH-1:0] wire_d40_46;
	wire [WIDTH-1:0] wire_d40_47;
	wire [WIDTH-1:0] wire_d40_48;
	wire [WIDTH-1:0] wire_d40_49;
	wire [WIDTH-1:0] wire_d40_50;
	wire [WIDTH-1:0] wire_d40_51;
	wire [WIDTH-1:0] wire_d40_52;
	wire [WIDTH-1:0] wire_d40_53;
	wire [WIDTH-1:0] wire_d40_54;
	wire [WIDTH-1:0] wire_d40_55;
	wire [WIDTH-1:0] wire_d40_56;
	wire [WIDTH-1:0] wire_d40_57;
	wire [WIDTH-1:0] wire_d40_58;
	wire [WIDTH-1:0] wire_d40_59;
	wire [WIDTH-1:0] wire_d40_60;
	wire [WIDTH-1:0] wire_d40_61;
	wire [WIDTH-1:0] wire_d40_62;
	wire [WIDTH-1:0] wire_d40_63;
	wire [WIDTH-1:0] wire_d40_64;
	wire [WIDTH-1:0] wire_d40_65;
	wire [WIDTH-1:0] wire_d40_66;
	wire [WIDTH-1:0] wire_d40_67;
	wire [WIDTH-1:0] wire_d40_68;
	wire [WIDTH-1:0] wire_d41_0;
	wire [WIDTH-1:0] wire_d41_1;
	wire [WIDTH-1:0] wire_d41_2;
	wire [WIDTH-1:0] wire_d41_3;
	wire [WIDTH-1:0] wire_d41_4;
	wire [WIDTH-1:0] wire_d41_5;
	wire [WIDTH-1:0] wire_d41_6;
	wire [WIDTH-1:0] wire_d41_7;
	wire [WIDTH-1:0] wire_d41_8;
	wire [WIDTH-1:0] wire_d41_9;
	wire [WIDTH-1:0] wire_d41_10;
	wire [WIDTH-1:0] wire_d41_11;
	wire [WIDTH-1:0] wire_d41_12;
	wire [WIDTH-1:0] wire_d41_13;
	wire [WIDTH-1:0] wire_d41_14;
	wire [WIDTH-1:0] wire_d41_15;
	wire [WIDTH-1:0] wire_d41_16;
	wire [WIDTH-1:0] wire_d41_17;
	wire [WIDTH-1:0] wire_d41_18;
	wire [WIDTH-1:0] wire_d41_19;
	wire [WIDTH-1:0] wire_d41_20;
	wire [WIDTH-1:0] wire_d41_21;
	wire [WIDTH-1:0] wire_d41_22;
	wire [WIDTH-1:0] wire_d41_23;
	wire [WIDTH-1:0] wire_d41_24;
	wire [WIDTH-1:0] wire_d41_25;
	wire [WIDTH-1:0] wire_d41_26;
	wire [WIDTH-1:0] wire_d41_27;
	wire [WIDTH-1:0] wire_d41_28;
	wire [WIDTH-1:0] wire_d41_29;
	wire [WIDTH-1:0] wire_d41_30;
	wire [WIDTH-1:0] wire_d41_31;
	wire [WIDTH-1:0] wire_d41_32;
	wire [WIDTH-1:0] wire_d41_33;
	wire [WIDTH-1:0] wire_d41_34;
	wire [WIDTH-1:0] wire_d41_35;
	wire [WIDTH-1:0] wire_d41_36;
	wire [WIDTH-1:0] wire_d41_37;
	wire [WIDTH-1:0] wire_d41_38;
	wire [WIDTH-1:0] wire_d41_39;
	wire [WIDTH-1:0] wire_d41_40;
	wire [WIDTH-1:0] wire_d41_41;
	wire [WIDTH-1:0] wire_d41_42;
	wire [WIDTH-1:0] wire_d41_43;
	wire [WIDTH-1:0] wire_d41_44;
	wire [WIDTH-1:0] wire_d41_45;
	wire [WIDTH-1:0] wire_d41_46;
	wire [WIDTH-1:0] wire_d41_47;
	wire [WIDTH-1:0] wire_d41_48;
	wire [WIDTH-1:0] wire_d41_49;
	wire [WIDTH-1:0] wire_d41_50;
	wire [WIDTH-1:0] wire_d41_51;
	wire [WIDTH-1:0] wire_d41_52;
	wire [WIDTH-1:0] wire_d41_53;
	wire [WIDTH-1:0] wire_d41_54;
	wire [WIDTH-1:0] wire_d41_55;
	wire [WIDTH-1:0] wire_d41_56;
	wire [WIDTH-1:0] wire_d41_57;
	wire [WIDTH-1:0] wire_d41_58;
	wire [WIDTH-1:0] wire_d41_59;
	wire [WIDTH-1:0] wire_d41_60;
	wire [WIDTH-1:0] wire_d41_61;
	wire [WIDTH-1:0] wire_d41_62;
	wire [WIDTH-1:0] wire_d41_63;
	wire [WIDTH-1:0] wire_d41_64;
	wire [WIDTH-1:0] wire_d41_65;
	wire [WIDTH-1:0] wire_d41_66;
	wire [WIDTH-1:0] wire_d41_67;
	wire [WIDTH-1:0] wire_d41_68;
	wire [WIDTH-1:0] wire_d42_0;
	wire [WIDTH-1:0] wire_d42_1;
	wire [WIDTH-1:0] wire_d42_2;
	wire [WIDTH-1:0] wire_d42_3;
	wire [WIDTH-1:0] wire_d42_4;
	wire [WIDTH-1:0] wire_d42_5;
	wire [WIDTH-1:0] wire_d42_6;
	wire [WIDTH-1:0] wire_d42_7;
	wire [WIDTH-1:0] wire_d42_8;
	wire [WIDTH-1:0] wire_d42_9;
	wire [WIDTH-1:0] wire_d42_10;
	wire [WIDTH-1:0] wire_d42_11;
	wire [WIDTH-1:0] wire_d42_12;
	wire [WIDTH-1:0] wire_d42_13;
	wire [WIDTH-1:0] wire_d42_14;
	wire [WIDTH-1:0] wire_d42_15;
	wire [WIDTH-1:0] wire_d42_16;
	wire [WIDTH-1:0] wire_d42_17;
	wire [WIDTH-1:0] wire_d42_18;
	wire [WIDTH-1:0] wire_d42_19;
	wire [WIDTH-1:0] wire_d42_20;
	wire [WIDTH-1:0] wire_d42_21;
	wire [WIDTH-1:0] wire_d42_22;
	wire [WIDTH-1:0] wire_d42_23;
	wire [WIDTH-1:0] wire_d42_24;
	wire [WIDTH-1:0] wire_d42_25;
	wire [WIDTH-1:0] wire_d42_26;
	wire [WIDTH-1:0] wire_d42_27;
	wire [WIDTH-1:0] wire_d42_28;
	wire [WIDTH-1:0] wire_d42_29;
	wire [WIDTH-1:0] wire_d42_30;
	wire [WIDTH-1:0] wire_d42_31;
	wire [WIDTH-1:0] wire_d42_32;
	wire [WIDTH-1:0] wire_d42_33;
	wire [WIDTH-1:0] wire_d42_34;
	wire [WIDTH-1:0] wire_d42_35;
	wire [WIDTH-1:0] wire_d42_36;
	wire [WIDTH-1:0] wire_d42_37;
	wire [WIDTH-1:0] wire_d42_38;
	wire [WIDTH-1:0] wire_d42_39;
	wire [WIDTH-1:0] wire_d42_40;
	wire [WIDTH-1:0] wire_d42_41;
	wire [WIDTH-1:0] wire_d42_42;
	wire [WIDTH-1:0] wire_d42_43;
	wire [WIDTH-1:0] wire_d42_44;
	wire [WIDTH-1:0] wire_d42_45;
	wire [WIDTH-1:0] wire_d42_46;
	wire [WIDTH-1:0] wire_d42_47;
	wire [WIDTH-1:0] wire_d42_48;
	wire [WIDTH-1:0] wire_d42_49;
	wire [WIDTH-1:0] wire_d42_50;
	wire [WIDTH-1:0] wire_d42_51;
	wire [WIDTH-1:0] wire_d42_52;
	wire [WIDTH-1:0] wire_d42_53;
	wire [WIDTH-1:0] wire_d42_54;
	wire [WIDTH-1:0] wire_d42_55;
	wire [WIDTH-1:0] wire_d42_56;
	wire [WIDTH-1:0] wire_d42_57;
	wire [WIDTH-1:0] wire_d42_58;
	wire [WIDTH-1:0] wire_d42_59;
	wire [WIDTH-1:0] wire_d42_60;
	wire [WIDTH-1:0] wire_d42_61;
	wire [WIDTH-1:0] wire_d42_62;
	wire [WIDTH-1:0] wire_d42_63;
	wire [WIDTH-1:0] wire_d42_64;
	wire [WIDTH-1:0] wire_d42_65;
	wire [WIDTH-1:0] wire_d42_66;
	wire [WIDTH-1:0] wire_d42_67;
	wire [WIDTH-1:0] wire_d42_68;
	wire [WIDTH-1:0] wire_d43_0;
	wire [WIDTH-1:0] wire_d43_1;
	wire [WIDTH-1:0] wire_d43_2;
	wire [WIDTH-1:0] wire_d43_3;
	wire [WIDTH-1:0] wire_d43_4;
	wire [WIDTH-1:0] wire_d43_5;
	wire [WIDTH-1:0] wire_d43_6;
	wire [WIDTH-1:0] wire_d43_7;
	wire [WIDTH-1:0] wire_d43_8;
	wire [WIDTH-1:0] wire_d43_9;
	wire [WIDTH-1:0] wire_d43_10;
	wire [WIDTH-1:0] wire_d43_11;
	wire [WIDTH-1:0] wire_d43_12;
	wire [WIDTH-1:0] wire_d43_13;
	wire [WIDTH-1:0] wire_d43_14;
	wire [WIDTH-1:0] wire_d43_15;
	wire [WIDTH-1:0] wire_d43_16;
	wire [WIDTH-1:0] wire_d43_17;
	wire [WIDTH-1:0] wire_d43_18;
	wire [WIDTH-1:0] wire_d43_19;
	wire [WIDTH-1:0] wire_d43_20;
	wire [WIDTH-1:0] wire_d43_21;
	wire [WIDTH-1:0] wire_d43_22;
	wire [WIDTH-1:0] wire_d43_23;
	wire [WIDTH-1:0] wire_d43_24;
	wire [WIDTH-1:0] wire_d43_25;
	wire [WIDTH-1:0] wire_d43_26;
	wire [WIDTH-1:0] wire_d43_27;
	wire [WIDTH-1:0] wire_d43_28;
	wire [WIDTH-1:0] wire_d43_29;
	wire [WIDTH-1:0] wire_d43_30;
	wire [WIDTH-1:0] wire_d43_31;
	wire [WIDTH-1:0] wire_d43_32;
	wire [WIDTH-1:0] wire_d43_33;
	wire [WIDTH-1:0] wire_d43_34;
	wire [WIDTH-1:0] wire_d43_35;
	wire [WIDTH-1:0] wire_d43_36;
	wire [WIDTH-1:0] wire_d43_37;
	wire [WIDTH-1:0] wire_d43_38;
	wire [WIDTH-1:0] wire_d43_39;
	wire [WIDTH-1:0] wire_d43_40;
	wire [WIDTH-1:0] wire_d43_41;
	wire [WIDTH-1:0] wire_d43_42;
	wire [WIDTH-1:0] wire_d43_43;
	wire [WIDTH-1:0] wire_d43_44;
	wire [WIDTH-1:0] wire_d43_45;
	wire [WIDTH-1:0] wire_d43_46;
	wire [WIDTH-1:0] wire_d43_47;
	wire [WIDTH-1:0] wire_d43_48;
	wire [WIDTH-1:0] wire_d43_49;
	wire [WIDTH-1:0] wire_d43_50;
	wire [WIDTH-1:0] wire_d43_51;
	wire [WIDTH-1:0] wire_d43_52;
	wire [WIDTH-1:0] wire_d43_53;
	wire [WIDTH-1:0] wire_d43_54;
	wire [WIDTH-1:0] wire_d43_55;
	wire [WIDTH-1:0] wire_d43_56;
	wire [WIDTH-1:0] wire_d43_57;
	wire [WIDTH-1:0] wire_d43_58;
	wire [WIDTH-1:0] wire_d43_59;
	wire [WIDTH-1:0] wire_d43_60;
	wire [WIDTH-1:0] wire_d43_61;
	wire [WIDTH-1:0] wire_d43_62;
	wire [WIDTH-1:0] wire_d43_63;
	wire [WIDTH-1:0] wire_d43_64;
	wire [WIDTH-1:0] wire_d43_65;
	wire [WIDTH-1:0] wire_d43_66;
	wire [WIDTH-1:0] wire_d43_67;
	wire [WIDTH-1:0] wire_d43_68;
	wire [WIDTH-1:0] wire_d44_0;
	wire [WIDTH-1:0] wire_d44_1;
	wire [WIDTH-1:0] wire_d44_2;
	wire [WIDTH-1:0] wire_d44_3;
	wire [WIDTH-1:0] wire_d44_4;
	wire [WIDTH-1:0] wire_d44_5;
	wire [WIDTH-1:0] wire_d44_6;
	wire [WIDTH-1:0] wire_d44_7;
	wire [WIDTH-1:0] wire_d44_8;
	wire [WIDTH-1:0] wire_d44_9;
	wire [WIDTH-1:0] wire_d44_10;
	wire [WIDTH-1:0] wire_d44_11;
	wire [WIDTH-1:0] wire_d44_12;
	wire [WIDTH-1:0] wire_d44_13;
	wire [WIDTH-1:0] wire_d44_14;
	wire [WIDTH-1:0] wire_d44_15;
	wire [WIDTH-1:0] wire_d44_16;
	wire [WIDTH-1:0] wire_d44_17;
	wire [WIDTH-1:0] wire_d44_18;
	wire [WIDTH-1:0] wire_d44_19;
	wire [WIDTH-1:0] wire_d44_20;
	wire [WIDTH-1:0] wire_d44_21;
	wire [WIDTH-1:0] wire_d44_22;
	wire [WIDTH-1:0] wire_d44_23;
	wire [WIDTH-1:0] wire_d44_24;
	wire [WIDTH-1:0] wire_d44_25;
	wire [WIDTH-1:0] wire_d44_26;
	wire [WIDTH-1:0] wire_d44_27;
	wire [WIDTH-1:0] wire_d44_28;
	wire [WIDTH-1:0] wire_d44_29;
	wire [WIDTH-1:0] wire_d44_30;
	wire [WIDTH-1:0] wire_d44_31;
	wire [WIDTH-1:0] wire_d44_32;
	wire [WIDTH-1:0] wire_d44_33;
	wire [WIDTH-1:0] wire_d44_34;
	wire [WIDTH-1:0] wire_d44_35;
	wire [WIDTH-1:0] wire_d44_36;
	wire [WIDTH-1:0] wire_d44_37;
	wire [WIDTH-1:0] wire_d44_38;
	wire [WIDTH-1:0] wire_d44_39;
	wire [WIDTH-1:0] wire_d44_40;
	wire [WIDTH-1:0] wire_d44_41;
	wire [WIDTH-1:0] wire_d44_42;
	wire [WIDTH-1:0] wire_d44_43;
	wire [WIDTH-1:0] wire_d44_44;
	wire [WIDTH-1:0] wire_d44_45;
	wire [WIDTH-1:0] wire_d44_46;
	wire [WIDTH-1:0] wire_d44_47;
	wire [WIDTH-1:0] wire_d44_48;
	wire [WIDTH-1:0] wire_d44_49;
	wire [WIDTH-1:0] wire_d44_50;
	wire [WIDTH-1:0] wire_d44_51;
	wire [WIDTH-1:0] wire_d44_52;
	wire [WIDTH-1:0] wire_d44_53;
	wire [WIDTH-1:0] wire_d44_54;
	wire [WIDTH-1:0] wire_d44_55;
	wire [WIDTH-1:0] wire_d44_56;
	wire [WIDTH-1:0] wire_d44_57;
	wire [WIDTH-1:0] wire_d44_58;
	wire [WIDTH-1:0] wire_d44_59;
	wire [WIDTH-1:0] wire_d44_60;
	wire [WIDTH-1:0] wire_d44_61;
	wire [WIDTH-1:0] wire_d44_62;
	wire [WIDTH-1:0] wire_d44_63;
	wire [WIDTH-1:0] wire_d44_64;
	wire [WIDTH-1:0] wire_d44_65;
	wire [WIDTH-1:0] wire_d44_66;
	wire [WIDTH-1:0] wire_d44_67;
	wire [WIDTH-1:0] wire_d44_68;
	wire [WIDTH-1:0] wire_d45_0;
	wire [WIDTH-1:0] wire_d45_1;
	wire [WIDTH-1:0] wire_d45_2;
	wire [WIDTH-1:0] wire_d45_3;
	wire [WIDTH-1:0] wire_d45_4;
	wire [WIDTH-1:0] wire_d45_5;
	wire [WIDTH-1:0] wire_d45_6;
	wire [WIDTH-1:0] wire_d45_7;
	wire [WIDTH-1:0] wire_d45_8;
	wire [WIDTH-1:0] wire_d45_9;
	wire [WIDTH-1:0] wire_d45_10;
	wire [WIDTH-1:0] wire_d45_11;
	wire [WIDTH-1:0] wire_d45_12;
	wire [WIDTH-1:0] wire_d45_13;
	wire [WIDTH-1:0] wire_d45_14;
	wire [WIDTH-1:0] wire_d45_15;
	wire [WIDTH-1:0] wire_d45_16;
	wire [WIDTH-1:0] wire_d45_17;
	wire [WIDTH-1:0] wire_d45_18;
	wire [WIDTH-1:0] wire_d45_19;
	wire [WIDTH-1:0] wire_d45_20;
	wire [WIDTH-1:0] wire_d45_21;
	wire [WIDTH-1:0] wire_d45_22;
	wire [WIDTH-1:0] wire_d45_23;
	wire [WIDTH-1:0] wire_d45_24;
	wire [WIDTH-1:0] wire_d45_25;
	wire [WIDTH-1:0] wire_d45_26;
	wire [WIDTH-1:0] wire_d45_27;
	wire [WIDTH-1:0] wire_d45_28;
	wire [WIDTH-1:0] wire_d45_29;
	wire [WIDTH-1:0] wire_d45_30;
	wire [WIDTH-1:0] wire_d45_31;
	wire [WIDTH-1:0] wire_d45_32;
	wire [WIDTH-1:0] wire_d45_33;
	wire [WIDTH-1:0] wire_d45_34;
	wire [WIDTH-1:0] wire_d45_35;
	wire [WIDTH-1:0] wire_d45_36;
	wire [WIDTH-1:0] wire_d45_37;
	wire [WIDTH-1:0] wire_d45_38;
	wire [WIDTH-1:0] wire_d45_39;
	wire [WIDTH-1:0] wire_d45_40;
	wire [WIDTH-1:0] wire_d45_41;
	wire [WIDTH-1:0] wire_d45_42;
	wire [WIDTH-1:0] wire_d45_43;
	wire [WIDTH-1:0] wire_d45_44;
	wire [WIDTH-1:0] wire_d45_45;
	wire [WIDTH-1:0] wire_d45_46;
	wire [WIDTH-1:0] wire_d45_47;
	wire [WIDTH-1:0] wire_d45_48;
	wire [WIDTH-1:0] wire_d45_49;
	wire [WIDTH-1:0] wire_d45_50;
	wire [WIDTH-1:0] wire_d45_51;
	wire [WIDTH-1:0] wire_d45_52;
	wire [WIDTH-1:0] wire_d45_53;
	wire [WIDTH-1:0] wire_d45_54;
	wire [WIDTH-1:0] wire_d45_55;
	wire [WIDTH-1:0] wire_d45_56;
	wire [WIDTH-1:0] wire_d45_57;
	wire [WIDTH-1:0] wire_d45_58;
	wire [WIDTH-1:0] wire_d45_59;
	wire [WIDTH-1:0] wire_d45_60;
	wire [WIDTH-1:0] wire_d45_61;
	wire [WIDTH-1:0] wire_d45_62;
	wire [WIDTH-1:0] wire_d45_63;
	wire [WIDTH-1:0] wire_d45_64;
	wire [WIDTH-1:0] wire_d45_65;
	wire [WIDTH-1:0] wire_d45_66;
	wire [WIDTH-1:0] wire_d45_67;
	wire [WIDTH-1:0] wire_d45_68;
	wire [WIDTH-1:0] wire_d46_0;
	wire [WIDTH-1:0] wire_d46_1;
	wire [WIDTH-1:0] wire_d46_2;
	wire [WIDTH-1:0] wire_d46_3;
	wire [WIDTH-1:0] wire_d46_4;
	wire [WIDTH-1:0] wire_d46_5;
	wire [WIDTH-1:0] wire_d46_6;
	wire [WIDTH-1:0] wire_d46_7;
	wire [WIDTH-1:0] wire_d46_8;
	wire [WIDTH-1:0] wire_d46_9;
	wire [WIDTH-1:0] wire_d46_10;
	wire [WIDTH-1:0] wire_d46_11;
	wire [WIDTH-1:0] wire_d46_12;
	wire [WIDTH-1:0] wire_d46_13;
	wire [WIDTH-1:0] wire_d46_14;
	wire [WIDTH-1:0] wire_d46_15;
	wire [WIDTH-1:0] wire_d46_16;
	wire [WIDTH-1:0] wire_d46_17;
	wire [WIDTH-1:0] wire_d46_18;
	wire [WIDTH-1:0] wire_d46_19;
	wire [WIDTH-1:0] wire_d46_20;
	wire [WIDTH-1:0] wire_d46_21;
	wire [WIDTH-1:0] wire_d46_22;
	wire [WIDTH-1:0] wire_d46_23;
	wire [WIDTH-1:0] wire_d46_24;
	wire [WIDTH-1:0] wire_d46_25;
	wire [WIDTH-1:0] wire_d46_26;
	wire [WIDTH-1:0] wire_d46_27;
	wire [WIDTH-1:0] wire_d46_28;
	wire [WIDTH-1:0] wire_d46_29;
	wire [WIDTH-1:0] wire_d46_30;
	wire [WIDTH-1:0] wire_d46_31;
	wire [WIDTH-1:0] wire_d46_32;
	wire [WIDTH-1:0] wire_d46_33;
	wire [WIDTH-1:0] wire_d46_34;
	wire [WIDTH-1:0] wire_d46_35;
	wire [WIDTH-1:0] wire_d46_36;
	wire [WIDTH-1:0] wire_d46_37;
	wire [WIDTH-1:0] wire_d46_38;
	wire [WIDTH-1:0] wire_d46_39;
	wire [WIDTH-1:0] wire_d46_40;
	wire [WIDTH-1:0] wire_d46_41;
	wire [WIDTH-1:0] wire_d46_42;
	wire [WIDTH-1:0] wire_d46_43;
	wire [WIDTH-1:0] wire_d46_44;
	wire [WIDTH-1:0] wire_d46_45;
	wire [WIDTH-1:0] wire_d46_46;
	wire [WIDTH-1:0] wire_d46_47;
	wire [WIDTH-1:0] wire_d46_48;
	wire [WIDTH-1:0] wire_d46_49;
	wire [WIDTH-1:0] wire_d46_50;
	wire [WIDTH-1:0] wire_d46_51;
	wire [WIDTH-1:0] wire_d46_52;
	wire [WIDTH-1:0] wire_d46_53;
	wire [WIDTH-1:0] wire_d46_54;
	wire [WIDTH-1:0] wire_d46_55;
	wire [WIDTH-1:0] wire_d46_56;
	wire [WIDTH-1:0] wire_d46_57;
	wire [WIDTH-1:0] wire_d46_58;
	wire [WIDTH-1:0] wire_d46_59;
	wire [WIDTH-1:0] wire_d46_60;
	wire [WIDTH-1:0] wire_d46_61;
	wire [WIDTH-1:0] wire_d46_62;
	wire [WIDTH-1:0] wire_d46_63;
	wire [WIDTH-1:0] wire_d46_64;
	wire [WIDTH-1:0] wire_d46_65;
	wire [WIDTH-1:0] wire_d46_66;
	wire [WIDTH-1:0] wire_d46_67;
	wire [WIDTH-1:0] wire_d46_68;
	wire [WIDTH-1:0] wire_d47_0;
	wire [WIDTH-1:0] wire_d47_1;
	wire [WIDTH-1:0] wire_d47_2;
	wire [WIDTH-1:0] wire_d47_3;
	wire [WIDTH-1:0] wire_d47_4;
	wire [WIDTH-1:0] wire_d47_5;
	wire [WIDTH-1:0] wire_d47_6;
	wire [WIDTH-1:0] wire_d47_7;
	wire [WIDTH-1:0] wire_d47_8;
	wire [WIDTH-1:0] wire_d47_9;
	wire [WIDTH-1:0] wire_d47_10;
	wire [WIDTH-1:0] wire_d47_11;
	wire [WIDTH-1:0] wire_d47_12;
	wire [WIDTH-1:0] wire_d47_13;
	wire [WIDTH-1:0] wire_d47_14;
	wire [WIDTH-1:0] wire_d47_15;
	wire [WIDTH-1:0] wire_d47_16;
	wire [WIDTH-1:0] wire_d47_17;
	wire [WIDTH-1:0] wire_d47_18;
	wire [WIDTH-1:0] wire_d47_19;
	wire [WIDTH-1:0] wire_d47_20;
	wire [WIDTH-1:0] wire_d47_21;
	wire [WIDTH-1:0] wire_d47_22;
	wire [WIDTH-1:0] wire_d47_23;
	wire [WIDTH-1:0] wire_d47_24;
	wire [WIDTH-1:0] wire_d47_25;
	wire [WIDTH-1:0] wire_d47_26;
	wire [WIDTH-1:0] wire_d47_27;
	wire [WIDTH-1:0] wire_d47_28;
	wire [WIDTH-1:0] wire_d47_29;
	wire [WIDTH-1:0] wire_d47_30;
	wire [WIDTH-1:0] wire_d47_31;
	wire [WIDTH-1:0] wire_d47_32;
	wire [WIDTH-1:0] wire_d47_33;
	wire [WIDTH-1:0] wire_d47_34;
	wire [WIDTH-1:0] wire_d47_35;
	wire [WIDTH-1:0] wire_d47_36;
	wire [WIDTH-1:0] wire_d47_37;
	wire [WIDTH-1:0] wire_d47_38;
	wire [WIDTH-1:0] wire_d47_39;
	wire [WIDTH-1:0] wire_d47_40;
	wire [WIDTH-1:0] wire_d47_41;
	wire [WIDTH-1:0] wire_d47_42;
	wire [WIDTH-1:0] wire_d47_43;
	wire [WIDTH-1:0] wire_d47_44;
	wire [WIDTH-1:0] wire_d47_45;
	wire [WIDTH-1:0] wire_d47_46;
	wire [WIDTH-1:0] wire_d47_47;
	wire [WIDTH-1:0] wire_d47_48;
	wire [WIDTH-1:0] wire_d47_49;
	wire [WIDTH-1:0] wire_d47_50;
	wire [WIDTH-1:0] wire_d47_51;
	wire [WIDTH-1:0] wire_d47_52;
	wire [WIDTH-1:0] wire_d47_53;
	wire [WIDTH-1:0] wire_d47_54;
	wire [WIDTH-1:0] wire_d47_55;
	wire [WIDTH-1:0] wire_d47_56;
	wire [WIDTH-1:0] wire_d47_57;
	wire [WIDTH-1:0] wire_d47_58;
	wire [WIDTH-1:0] wire_d47_59;
	wire [WIDTH-1:0] wire_d47_60;
	wire [WIDTH-1:0] wire_d47_61;
	wire [WIDTH-1:0] wire_d47_62;
	wire [WIDTH-1:0] wire_d47_63;
	wire [WIDTH-1:0] wire_d47_64;
	wire [WIDTH-1:0] wire_d47_65;
	wire [WIDTH-1:0] wire_d47_66;
	wire [WIDTH-1:0] wire_d47_67;
	wire [WIDTH-1:0] wire_d47_68;
	wire [WIDTH-1:0] wire_d48_0;
	wire [WIDTH-1:0] wire_d48_1;
	wire [WIDTH-1:0] wire_d48_2;
	wire [WIDTH-1:0] wire_d48_3;
	wire [WIDTH-1:0] wire_d48_4;
	wire [WIDTH-1:0] wire_d48_5;
	wire [WIDTH-1:0] wire_d48_6;
	wire [WIDTH-1:0] wire_d48_7;
	wire [WIDTH-1:0] wire_d48_8;
	wire [WIDTH-1:0] wire_d48_9;
	wire [WIDTH-1:0] wire_d48_10;
	wire [WIDTH-1:0] wire_d48_11;
	wire [WIDTH-1:0] wire_d48_12;
	wire [WIDTH-1:0] wire_d48_13;
	wire [WIDTH-1:0] wire_d48_14;
	wire [WIDTH-1:0] wire_d48_15;
	wire [WIDTH-1:0] wire_d48_16;
	wire [WIDTH-1:0] wire_d48_17;
	wire [WIDTH-1:0] wire_d48_18;
	wire [WIDTH-1:0] wire_d48_19;
	wire [WIDTH-1:0] wire_d48_20;
	wire [WIDTH-1:0] wire_d48_21;
	wire [WIDTH-1:0] wire_d48_22;
	wire [WIDTH-1:0] wire_d48_23;
	wire [WIDTH-1:0] wire_d48_24;
	wire [WIDTH-1:0] wire_d48_25;
	wire [WIDTH-1:0] wire_d48_26;
	wire [WIDTH-1:0] wire_d48_27;
	wire [WIDTH-1:0] wire_d48_28;
	wire [WIDTH-1:0] wire_d48_29;
	wire [WIDTH-1:0] wire_d48_30;
	wire [WIDTH-1:0] wire_d48_31;
	wire [WIDTH-1:0] wire_d48_32;
	wire [WIDTH-1:0] wire_d48_33;
	wire [WIDTH-1:0] wire_d48_34;
	wire [WIDTH-1:0] wire_d48_35;
	wire [WIDTH-1:0] wire_d48_36;
	wire [WIDTH-1:0] wire_d48_37;
	wire [WIDTH-1:0] wire_d48_38;
	wire [WIDTH-1:0] wire_d48_39;
	wire [WIDTH-1:0] wire_d48_40;
	wire [WIDTH-1:0] wire_d48_41;
	wire [WIDTH-1:0] wire_d48_42;
	wire [WIDTH-1:0] wire_d48_43;
	wire [WIDTH-1:0] wire_d48_44;
	wire [WIDTH-1:0] wire_d48_45;
	wire [WIDTH-1:0] wire_d48_46;
	wire [WIDTH-1:0] wire_d48_47;
	wire [WIDTH-1:0] wire_d48_48;
	wire [WIDTH-1:0] wire_d48_49;
	wire [WIDTH-1:0] wire_d48_50;
	wire [WIDTH-1:0] wire_d48_51;
	wire [WIDTH-1:0] wire_d48_52;
	wire [WIDTH-1:0] wire_d48_53;
	wire [WIDTH-1:0] wire_d48_54;
	wire [WIDTH-1:0] wire_d48_55;
	wire [WIDTH-1:0] wire_d48_56;
	wire [WIDTH-1:0] wire_d48_57;
	wire [WIDTH-1:0] wire_d48_58;
	wire [WIDTH-1:0] wire_d48_59;
	wire [WIDTH-1:0] wire_d48_60;
	wire [WIDTH-1:0] wire_d48_61;
	wire [WIDTH-1:0] wire_d48_62;
	wire [WIDTH-1:0] wire_d48_63;
	wire [WIDTH-1:0] wire_d48_64;
	wire [WIDTH-1:0] wire_d48_65;
	wire [WIDTH-1:0] wire_d48_66;
	wire [WIDTH-1:0] wire_d48_67;
	wire [WIDTH-1:0] wire_d48_68;
	wire [WIDTH-1:0] wire_d49_0;
	wire [WIDTH-1:0] wire_d49_1;
	wire [WIDTH-1:0] wire_d49_2;
	wire [WIDTH-1:0] wire_d49_3;
	wire [WIDTH-1:0] wire_d49_4;
	wire [WIDTH-1:0] wire_d49_5;
	wire [WIDTH-1:0] wire_d49_6;
	wire [WIDTH-1:0] wire_d49_7;
	wire [WIDTH-1:0] wire_d49_8;
	wire [WIDTH-1:0] wire_d49_9;
	wire [WIDTH-1:0] wire_d49_10;
	wire [WIDTH-1:0] wire_d49_11;
	wire [WIDTH-1:0] wire_d49_12;
	wire [WIDTH-1:0] wire_d49_13;
	wire [WIDTH-1:0] wire_d49_14;
	wire [WIDTH-1:0] wire_d49_15;
	wire [WIDTH-1:0] wire_d49_16;
	wire [WIDTH-1:0] wire_d49_17;
	wire [WIDTH-1:0] wire_d49_18;
	wire [WIDTH-1:0] wire_d49_19;
	wire [WIDTH-1:0] wire_d49_20;
	wire [WIDTH-1:0] wire_d49_21;
	wire [WIDTH-1:0] wire_d49_22;
	wire [WIDTH-1:0] wire_d49_23;
	wire [WIDTH-1:0] wire_d49_24;
	wire [WIDTH-1:0] wire_d49_25;
	wire [WIDTH-1:0] wire_d49_26;
	wire [WIDTH-1:0] wire_d49_27;
	wire [WIDTH-1:0] wire_d49_28;
	wire [WIDTH-1:0] wire_d49_29;
	wire [WIDTH-1:0] wire_d49_30;
	wire [WIDTH-1:0] wire_d49_31;
	wire [WIDTH-1:0] wire_d49_32;
	wire [WIDTH-1:0] wire_d49_33;
	wire [WIDTH-1:0] wire_d49_34;
	wire [WIDTH-1:0] wire_d49_35;
	wire [WIDTH-1:0] wire_d49_36;
	wire [WIDTH-1:0] wire_d49_37;
	wire [WIDTH-1:0] wire_d49_38;
	wire [WIDTH-1:0] wire_d49_39;
	wire [WIDTH-1:0] wire_d49_40;
	wire [WIDTH-1:0] wire_d49_41;
	wire [WIDTH-1:0] wire_d49_42;
	wire [WIDTH-1:0] wire_d49_43;
	wire [WIDTH-1:0] wire_d49_44;
	wire [WIDTH-1:0] wire_d49_45;
	wire [WIDTH-1:0] wire_d49_46;
	wire [WIDTH-1:0] wire_d49_47;
	wire [WIDTH-1:0] wire_d49_48;
	wire [WIDTH-1:0] wire_d49_49;
	wire [WIDTH-1:0] wire_d49_50;
	wire [WIDTH-1:0] wire_d49_51;
	wire [WIDTH-1:0] wire_d49_52;
	wire [WIDTH-1:0] wire_d49_53;
	wire [WIDTH-1:0] wire_d49_54;
	wire [WIDTH-1:0] wire_d49_55;
	wire [WIDTH-1:0] wire_d49_56;
	wire [WIDTH-1:0] wire_d49_57;
	wire [WIDTH-1:0] wire_d49_58;
	wire [WIDTH-1:0] wire_d49_59;
	wire [WIDTH-1:0] wire_d49_60;
	wire [WIDTH-1:0] wire_d49_61;
	wire [WIDTH-1:0] wire_d49_62;
	wire [WIDTH-1:0] wire_d49_63;
	wire [WIDTH-1:0] wire_d49_64;
	wire [WIDTH-1:0] wire_d49_65;
	wire [WIDTH-1:0] wire_d49_66;
	wire [WIDTH-1:0] wire_d49_67;
	wire [WIDTH-1:0] wire_d49_68;

	register #(.WIDTH(WIDTH)) register_instance100(.data_in(d_in0),.data_out(wire_d0_0),.clk(clk),.rst(rst));            //channel 1
	invertion #(.WIDTH(WIDTH)) invertion_instance101(.data_in(wire_d0_0),.data_out(wire_d0_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance102(.data_in(wire_d0_1),.data_out(wire_d0_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance103(.data_in(wire_d0_2),.data_out(wire_d0_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance104(.data_in(wire_d0_3),.data_out(wire_d0_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance105(.data_in(wire_d0_4),.data_out(wire_d0_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance106(.data_in(wire_d0_5),.data_out(wire_d0_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance107(.data_in(wire_d0_6),.data_out(wire_d0_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance108(.data_in(wire_d0_7),.data_out(wire_d0_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance109(.data_in(wire_d0_8),.data_out(wire_d0_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1010(.data_in(wire_d0_9),.data_out(wire_d0_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1011(.data_in(wire_d0_10),.data_out(wire_d0_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1012(.data_in(wire_d0_11),.data_out(wire_d0_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1013(.data_in(wire_d0_12),.data_out(wire_d0_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1014(.data_in(wire_d0_13),.data_out(wire_d0_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1015(.data_in(wire_d0_14),.data_out(wire_d0_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1016(.data_in(wire_d0_15),.data_out(wire_d0_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1017(.data_in(wire_d0_16),.data_out(wire_d0_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1018(.data_in(wire_d0_17),.data_out(wire_d0_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1019(.data_in(wire_d0_18),.data_out(wire_d0_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1020(.data_in(wire_d0_19),.data_out(wire_d0_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1021(.data_in(wire_d0_20),.data_out(wire_d0_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1022(.data_in(wire_d0_21),.data_out(wire_d0_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1023(.data_in(wire_d0_22),.data_out(wire_d0_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1024(.data_in(wire_d0_23),.data_out(wire_d0_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1025(.data_in(wire_d0_24),.data_out(wire_d0_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1026(.data_in(wire_d0_25),.data_out(wire_d0_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1027(.data_in(wire_d0_26),.data_out(wire_d0_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1028(.data_in(wire_d0_27),.data_out(wire_d0_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1029(.data_in(wire_d0_28),.data_out(wire_d0_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1030(.data_in(wire_d0_29),.data_out(wire_d0_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1031(.data_in(wire_d0_30),.data_out(wire_d0_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1032(.data_in(wire_d0_31),.data_out(wire_d0_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1033(.data_in(wire_d0_32),.data_out(wire_d0_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1034(.data_in(wire_d0_33),.data_out(wire_d0_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1035(.data_in(wire_d0_34),.data_out(wire_d0_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1036(.data_in(wire_d0_35),.data_out(wire_d0_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1037(.data_in(wire_d0_36),.data_out(wire_d0_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1038(.data_in(wire_d0_37),.data_out(wire_d0_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1039(.data_in(wire_d0_38),.data_out(wire_d0_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1040(.data_in(wire_d0_39),.data_out(wire_d0_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1041(.data_in(wire_d0_40),.data_out(wire_d0_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1042(.data_in(wire_d0_41),.data_out(wire_d0_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1043(.data_in(wire_d0_42),.data_out(wire_d0_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1044(.data_in(wire_d0_43),.data_out(wire_d0_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1045(.data_in(wire_d0_44),.data_out(wire_d0_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1046(.data_in(wire_d0_45),.data_out(wire_d0_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1047(.data_in(wire_d0_46),.data_out(wire_d0_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1048(.data_in(wire_d0_47),.data_out(wire_d0_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1049(.data_in(wire_d0_48),.data_out(wire_d0_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1050(.data_in(wire_d0_49),.data_out(wire_d0_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1051(.data_in(wire_d0_50),.data_out(wire_d0_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1052(.data_in(wire_d0_51),.data_out(wire_d0_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1053(.data_in(wire_d0_52),.data_out(wire_d0_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1054(.data_in(wire_d0_53),.data_out(wire_d0_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1055(.data_in(wire_d0_54),.data_out(wire_d0_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1056(.data_in(wire_d0_55),.data_out(wire_d0_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1057(.data_in(wire_d0_56),.data_out(wire_d0_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1058(.data_in(wire_d0_57),.data_out(wire_d0_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1059(.data_in(wire_d0_58),.data_out(wire_d0_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1060(.data_in(wire_d0_59),.data_out(wire_d0_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1061(.data_in(wire_d0_60),.data_out(wire_d0_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1062(.data_in(wire_d0_61),.data_out(wire_d0_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1063(.data_in(wire_d0_62),.data_out(wire_d0_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1064(.data_in(wire_d0_63),.data_out(wire_d0_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1065(.data_in(wire_d0_64),.data_out(wire_d0_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1066(.data_in(wire_d0_65),.data_out(wire_d0_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1067(.data_in(wire_d0_66),.data_out(wire_d0_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1068(.data_in(wire_d0_67),.data_out(wire_d0_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1069(.data_in(wire_d0_68),.data_out(d_out0),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance210(.data_in(d_in1),.data_out(wire_d1_0),.clk(clk),.rst(rst));            //channel 2
	register #(.WIDTH(WIDTH)) register_instance211(.data_in(wire_d1_0),.data_out(wire_d1_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212(.data_in(wire_d1_1),.data_out(wire_d1_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance213(.data_in(wire_d1_2),.data_out(wire_d1_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance214(.data_in(wire_d1_3),.data_out(wire_d1_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance215(.data_in(wire_d1_4),.data_out(wire_d1_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance216(.data_in(wire_d1_5),.data_out(wire_d1_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance217(.data_in(wire_d1_6),.data_out(wire_d1_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance218(.data_in(wire_d1_7),.data_out(wire_d1_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance219(.data_in(wire_d1_8),.data_out(wire_d1_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2110(.data_in(wire_d1_9),.data_out(wire_d1_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2111(.data_in(wire_d1_10),.data_out(wire_d1_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2112(.data_in(wire_d1_11),.data_out(wire_d1_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2113(.data_in(wire_d1_12),.data_out(wire_d1_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2114(.data_in(wire_d1_13),.data_out(wire_d1_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2115(.data_in(wire_d1_14),.data_out(wire_d1_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2116(.data_in(wire_d1_15),.data_out(wire_d1_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2117(.data_in(wire_d1_16),.data_out(wire_d1_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2118(.data_in(wire_d1_17),.data_out(wire_d1_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2119(.data_in(wire_d1_18),.data_out(wire_d1_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2120(.data_in(wire_d1_19),.data_out(wire_d1_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2121(.data_in(wire_d1_20),.data_out(wire_d1_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2122(.data_in(wire_d1_21),.data_out(wire_d1_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2123(.data_in(wire_d1_22),.data_out(wire_d1_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2124(.data_in(wire_d1_23),.data_out(wire_d1_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2125(.data_in(wire_d1_24),.data_out(wire_d1_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2126(.data_in(wire_d1_25),.data_out(wire_d1_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2127(.data_in(wire_d1_26),.data_out(wire_d1_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2128(.data_in(wire_d1_27),.data_out(wire_d1_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2129(.data_in(wire_d1_28),.data_out(wire_d1_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2130(.data_in(wire_d1_29),.data_out(wire_d1_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2131(.data_in(wire_d1_30),.data_out(wire_d1_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2132(.data_in(wire_d1_31),.data_out(wire_d1_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2133(.data_in(wire_d1_32),.data_out(wire_d1_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2134(.data_in(wire_d1_33),.data_out(wire_d1_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2135(.data_in(wire_d1_34),.data_out(wire_d1_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2136(.data_in(wire_d1_35),.data_out(wire_d1_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2137(.data_in(wire_d1_36),.data_out(wire_d1_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2138(.data_in(wire_d1_37),.data_out(wire_d1_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2139(.data_in(wire_d1_38),.data_out(wire_d1_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2140(.data_in(wire_d1_39),.data_out(wire_d1_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2141(.data_in(wire_d1_40),.data_out(wire_d1_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2142(.data_in(wire_d1_41),.data_out(wire_d1_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2143(.data_in(wire_d1_42),.data_out(wire_d1_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2144(.data_in(wire_d1_43),.data_out(wire_d1_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2145(.data_in(wire_d1_44),.data_out(wire_d1_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2146(.data_in(wire_d1_45),.data_out(wire_d1_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2147(.data_in(wire_d1_46),.data_out(wire_d1_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2148(.data_in(wire_d1_47),.data_out(wire_d1_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2149(.data_in(wire_d1_48),.data_out(wire_d1_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2150(.data_in(wire_d1_49),.data_out(wire_d1_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2151(.data_in(wire_d1_50),.data_out(wire_d1_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2152(.data_in(wire_d1_51),.data_out(wire_d1_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2153(.data_in(wire_d1_52),.data_out(wire_d1_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2154(.data_in(wire_d1_53),.data_out(wire_d1_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2155(.data_in(wire_d1_54),.data_out(wire_d1_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2156(.data_in(wire_d1_55),.data_out(wire_d1_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2157(.data_in(wire_d1_56),.data_out(wire_d1_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2158(.data_in(wire_d1_57),.data_out(wire_d1_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2159(.data_in(wire_d1_58),.data_out(wire_d1_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2160(.data_in(wire_d1_59),.data_out(wire_d1_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2161(.data_in(wire_d1_60),.data_out(wire_d1_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2162(.data_in(wire_d1_61),.data_out(wire_d1_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2163(.data_in(wire_d1_62),.data_out(wire_d1_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2164(.data_in(wire_d1_63),.data_out(wire_d1_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2165(.data_in(wire_d1_64),.data_out(wire_d1_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2166(.data_in(wire_d1_65),.data_out(wire_d1_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2167(.data_in(wire_d1_66),.data_out(wire_d1_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2168(.data_in(wire_d1_67),.data_out(wire_d1_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2169(.data_in(wire_d1_68),.data_out(d_out1),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance320(.data_in(d_in2),.data_out(wire_d2_0),.clk(clk),.rst(rst));            //channel 3
	invertion #(.WIDTH(WIDTH)) invertion_instance321(.data_in(wire_d2_0),.data_out(wire_d2_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance322(.data_in(wire_d2_1),.data_out(wire_d2_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323(.data_in(wire_d2_2),.data_out(wire_d2_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance324(.data_in(wire_d2_3),.data_out(wire_d2_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance325(.data_in(wire_d2_4),.data_out(wire_d2_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance326(.data_in(wire_d2_5),.data_out(wire_d2_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance327(.data_in(wire_d2_6),.data_out(wire_d2_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance328(.data_in(wire_d2_7),.data_out(wire_d2_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance329(.data_in(wire_d2_8),.data_out(wire_d2_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3210(.data_in(wire_d2_9),.data_out(wire_d2_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3211(.data_in(wire_d2_10),.data_out(wire_d2_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3212(.data_in(wire_d2_11),.data_out(wire_d2_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3213(.data_in(wire_d2_12),.data_out(wire_d2_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3214(.data_in(wire_d2_13),.data_out(wire_d2_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3215(.data_in(wire_d2_14),.data_out(wire_d2_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3216(.data_in(wire_d2_15),.data_out(wire_d2_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3217(.data_in(wire_d2_16),.data_out(wire_d2_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3218(.data_in(wire_d2_17),.data_out(wire_d2_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3219(.data_in(wire_d2_18),.data_out(wire_d2_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3220(.data_in(wire_d2_19),.data_out(wire_d2_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3221(.data_in(wire_d2_20),.data_out(wire_d2_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3222(.data_in(wire_d2_21),.data_out(wire_d2_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3223(.data_in(wire_d2_22),.data_out(wire_d2_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3224(.data_in(wire_d2_23),.data_out(wire_d2_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3225(.data_in(wire_d2_24),.data_out(wire_d2_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3226(.data_in(wire_d2_25),.data_out(wire_d2_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3227(.data_in(wire_d2_26),.data_out(wire_d2_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3228(.data_in(wire_d2_27),.data_out(wire_d2_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3229(.data_in(wire_d2_28),.data_out(wire_d2_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3230(.data_in(wire_d2_29),.data_out(wire_d2_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3231(.data_in(wire_d2_30),.data_out(wire_d2_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3232(.data_in(wire_d2_31),.data_out(wire_d2_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3233(.data_in(wire_d2_32),.data_out(wire_d2_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3234(.data_in(wire_d2_33),.data_out(wire_d2_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3235(.data_in(wire_d2_34),.data_out(wire_d2_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3236(.data_in(wire_d2_35),.data_out(wire_d2_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3237(.data_in(wire_d2_36),.data_out(wire_d2_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3238(.data_in(wire_d2_37),.data_out(wire_d2_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3239(.data_in(wire_d2_38),.data_out(wire_d2_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3240(.data_in(wire_d2_39),.data_out(wire_d2_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3241(.data_in(wire_d2_40),.data_out(wire_d2_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3242(.data_in(wire_d2_41),.data_out(wire_d2_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3243(.data_in(wire_d2_42),.data_out(wire_d2_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3244(.data_in(wire_d2_43),.data_out(wire_d2_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3245(.data_in(wire_d2_44),.data_out(wire_d2_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3246(.data_in(wire_d2_45),.data_out(wire_d2_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3247(.data_in(wire_d2_46),.data_out(wire_d2_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3248(.data_in(wire_d2_47),.data_out(wire_d2_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3249(.data_in(wire_d2_48),.data_out(wire_d2_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3250(.data_in(wire_d2_49),.data_out(wire_d2_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3251(.data_in(wire_d2_50),.data_out(wire_d2_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3252(.data_in(wire_d2_51),.data_out(wire_d2_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3253(.data_in(wire_d2_52),.data_out(wire_d2_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3254(.data_in(wire_d2_53),.data_out(wire_d2_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3255(.data_in(wire_d2_54),.data_out(wire_d2_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3256(.data_in(wire_d2_55),.data_out(wire_d2_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3257(.data_in(wire_d2_56),.data_out(wire_d2_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3258(.data_in(wire_d2_57),.data_out(wire_d2_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3259(.data_in(wire_d2_58),.data_out(wire_d2_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3260(.data_in(wire_d2_59),.data_out(wire_d2_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3261(.data_in(wire_d2_60),.data_out(wire_d2_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3262(.data_in(wire_d2_61),.data_out(wire_d2_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3263(.data_in(wire_d2_62),.data_out(wire_d2_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3264(.data_in(wire_d2_63),.data_out(wire_d2_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3265(.data_in(wire_d2_64),.data_out(wire_d2_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3266(.data_in(wire_d2_65),.data_out(wire_d2_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3267(.data_in(wire_d2_66),.data_out(wire_d2_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3268(.data_in(wire_d2_67),.data_out(wire_d2_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3269(.data_in(wire_d2_68),.data_out(d_out2),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance430(.data_in(d_in3),.data_out(wire_d3_0),.clk(clk),.rst(rst));            //channel 4
	encoder #(.WIDTH(WIDTH)) encoder_instance431(.data_in(wire_d3_0),.data_out(wire_d3_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance432(.data_in(wire_d3_1),.data_out(wire_d3_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance433(.data_in(wire_d3_2),.data_out(wire_d3_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434(.data_in(wire_d3_3),.data_out(wire_d3_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance435(.data_in(wire_d3_4),.data_out(wire_d3_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance436(.data_in(wire_d3_5),.data_out(wire_d3_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance437(.data_in(wire_d3_6),.data_out(wire_d3_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance438(.data_in(wire_d3_7),.data_out(wire_d3_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance439(.data_in(wire_d3_8),.data_out(wire_d3_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4310(.data_in(wire_d3_9),.data_out(wire_d3_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4311(.data_in(wire_d3_10),.data_out(wire_d3_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4312(.data_in(wire_d3_11),.data_out(wire_d3_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4313(.data_in(wire_d3_12),.data_out(wire_d3_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4314(.data_in(wire_d3_13),.data_out(wire_d3_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4315(.data_in(wire_d3_14),.data_out(wire_d3_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4316(.data_in(wire_d3_15),.data_out(wire_d3_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4317(.data_in(wire_d3_16),.data_out(wire_d3_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4318(.data_in(wire_d3_17),.data_out(wire_d3_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4319(.data_in(wire_d3_18),.data_out(wire_d3_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4320(.data_in(wire_d3_19),.data_out(wire_d3_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4321(.data_in(wire_d3_20),.data_out(wire_d3_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4322(.data_in(wire_d3_21),.data_out(wire_d3_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4323(.data_in(wire_d3_22),.data_out(wire_d3_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4324(.data_in(wire_d3_23),.data_out(wire_d3_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4325(.data_in(wire_d3_24),.data_out(wire_d3_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4326(.data_in(wire_d3_25),.data_out(wire_d3_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4327(.data_in(wire_d3_26),.data_out(wire_d3_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4328(.data_in(wire_d3_27),.data_out(wire_d3_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4329(.data_in(wire_d3_28),.data_out(wire_d3_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4330(.data_in(wire_d3_29),.data_out(wire_d3_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4331(.data_in(wire_d3_30),.data_out(wire_d3_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4332(.data_in(wire_d3_31),.data_out(wire_d3_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4333(.data_in(wire_d3_32),.data_out(wire_d3_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4334(.data_in(wire_d3_33),.data_out(wire_d3_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4335(.data_in(wire_d3_34),.data_out(wire_d3_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4336(.data_in(wire_d3_35),.data_out(wire_d3_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4337(.data_in(wire_d3_36),.data_out(wire_d3_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4338(.data_in(wire_d3_37),.data_out(wire_d3_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4339(.data_in(wire_d3_38),.data_out(wire_d3_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4340(.data_in(wire_d3_39),.data_out(wire_d3_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4341(.data_in(wire_d3_40),.data_out(wire_d3_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4342(.data_in(wire_d3_41),.data_out(wire_d3_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4343(.data_in(wire_d3_42),.data_out(wire_d3_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4344(.data_in(wire_d3_43),.data_out(wire_d3_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4345(.data_in(wire_d3_44),.data_out(wire_d3_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4346(.data_in(wire_d3_45),.data_out(wire_d3_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4347(.data_in(wire_d3_46),.data_out(wire_d3_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4348(.data_in(wire_d3_47),.data_out(wire_d3_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4349(.data_in(wire_d3_48),.data_out(wire_d3_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4350(.data_in(wire_d3_49),.data_out(wire_d3_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4351(.data_in(wire_d3_50),.data_out(wire_d3_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4352(.data_in(wire_d3_51),.data_out(wire_d3_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4353(.data_in(wire_d3_52),.data_out(wire_d3_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4354(.data_in(wire_d3_53),.data_out(wire_d3_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4355(.data_in(wire_d3_54),.data_out(wire_d3_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4356(.data_in(wire_d3_55),.data_out(wire_d3_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4357(.data_in(wire_d3_56),.data_out(wire_d3_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4358(.data_in(wire_d3_57),.data_out(wire_d3_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4359(.data_in(wire_d3_58),.data_out(wire_d3_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4360(.data_in(wire_d3_59),.data_out(wire_d3_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4361(.data_in(wire_d3_60),.data_out(wire_d3_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4362(.data_in(wire_d3_61),.data_out(wire_d3_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4363(.data_in(wire_d3_62),.data_out(wire_d3_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4364(.data_in(wire_d3_63),.data_out(wire_d3_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4365(.data_in(wire_d3_64),.data_out(wire_d3_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4366(.data_in(wire_d3_65),.data_out(wire_d3_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4367(.data_in(wire_d3_66),.data_out(wire_d3_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4368(.data_in(wire_d3_67),.data_out(wire_d3_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4369(.data_in(wire_d3_68),.data_out(d_out3),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance540(.data_in(d_in4),.data_out(wire_d4_0),.clk(clk),.rst(rst));            //channel 5
	register #(.WIDTH(WIDTH)) register_instance541(.data_in(wire_d4_0),.data_out(wire_d4_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance542(.data_in(wire_d4_1),.data_out(wire_d4_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance543(.data_in(wire_d4_2),.data_out(wire_d4_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance544(.data_in(wire_d4_3),.data_out(wire_d4_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545(.data_in(wire_d4_4),.data_out(wire_d4_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance546(.data_in(wire_d4_5),.data_out(wire_d4_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance547(.data_in(wire_d4_6),.data_out(wire_d4_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance548(.data_in(wire_d4_7),.data_out(wire_d4_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance549(.data_in(wire_d4_8),.data_out(wire_d4_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5410(.data_in(wire_d4_9),.data_out(wire_d4_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5411(.data_in(wire_d4_10),.data_out(wire_d4_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5412(.data_in(wire_d4_11),.data_out(wire_d4_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5413(.data_in(wire_d4_12),.data_out(wire_d4_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5414(.data_in(wire_d4_13),.data_out(wire_d4_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5415(.data_in(wire_d4_14),.data_out(wire_d4_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5416(.data_in(wire_d4_15),.data_out(wire_d4_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5417(.data_in(wire_d4_16),.data_out(wire_d4_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5418(.data_in(wire_d4_17),.data_out(wire_d4_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5419(.data_in(wire_d4_18),.data_out(wire_d4_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5420(.data_in(wire_d4_19),.data_out(wire_d4_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5421(.data_in(wire_d4_20),.data_out(wire_d4_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5422(.data_in(wire_d4_21),.data_out(wire_d4_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5423(.data_in(wire_d4_22),.data_out(wire_d4_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5424(.data_in(wire_d4_23),.data_out(wire_d4_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5425(.data_in(wire_d4_24),.data_out(wire_d4_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5426(.data_in(wire_d4_25),.data_out(wire_d4_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5427(.data_in(wire_d4_26),.data_out(wire_d4_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5428(.data_in(wire_d4_27),.data_out(wire_d4_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5429(.data_in(wire_d4_28),.data_out(wire_d4_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5430(.data_in(wire_d4_29),.data_out(wire_d4_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5431(.data_in(wire_d4_30),.data_out(wire_d4_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5432(.data_in(wire_d4_31),.data_out(wire_d4_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5433(.data_in(wire_d4_32),.data_out(wire_d4_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5434(.data_in(wire_d4_33),.data_out(wire_d4_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5435(.data_in(wire_d4_34),.data_out(wire_d4_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5436(.data_in(wire_d4_35),.data_out(wire_d4_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5437(.data_in(wire_d4_36),.data_out(wire_d4_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5438(.data_in(wire_d4_37),.data_out(wire_d4_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5439(.data_in(wire_d4_38),.data_out(wire_d4_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5440(.data_in(wire_d4_39),.data_out(wire_d4_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5441(.data_in(wire_d4_40),.data_out(wire_d4_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5442(.data_in(wire_d4_41),.data_out(wire_d4_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5443(.data_in(wire_d4_42),.data_out(wire_d4_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5444(.data_in(wire_d4_43),.data_out(wire_d4_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5445(.data_in(wire_d4_44),.data_out(wire_d4_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5446(.data_in(wire_d4_45),.data_out(wire_d4_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5447(.data_in(wire_d4_46),.data_out(wire_d4_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5448(.data_in(wire_d4_47),.data_out(wire_d4_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5449(.data_in(wire_d4_48),.data_out(wire_d4_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5450(.data_in(wire_d4_49),.data_out(wire_d4_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5451(.data_in(wire_d4_50),.data_out(wire_d4_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5452(.data_in(wire_d4_51),.data_out(wire_d4_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5453(.data_in(wire_d4_52),.data_out(wire_d4_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5454(.data_in(wire_d4_53),.data_out(wire_d4_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5455(.data_in(wire_d4_54),.data_out(wire_d4_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5456(.data_in(wire_d4_55),.data_out(wire_d4_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5457(.data_in(wire_d4_56),.data_out(wire_d4_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5458(.data_in(wire_d4_57),.data_out(wire_d4_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5459(.data_in(wire_d4_58),.data_out(wire_d4_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5460(.data_in(wire_d4_59),.data_out(wire_d4_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5461(.data_in(wire_d4_60),.data_out(wire_d4_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5462(.data_in(wire_d4_61),.data_out(wire_d4_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5463(.data_in(wire_d4_62),.data_out(wire_d4_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5464(.data_in(wire_d4_63),.data_out(wire_d4_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5465(.data_in(wire_d4_64),.data_out(wire_d4_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5466(.data_in(wire_d4_65),.data_out(wire_d4_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5467(.data_in(wire_d4_66),.data_out(wire_d4_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5468(.data_in(wire_d4_67),.data_out(wire_d4_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5469(.data_in(wire_d4_68),.data_out(d_out4),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance650(.data_in(d_in5),.data_out(wire_d5_0),.clk(clk),.rst(rst));            //channel 6
	encoder #(.WIDTH(WIDTH)) encoder_instance651(.data_in(wire_d5_0),.data_out(wire_d5_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance652(.data_in(wire_d5_1),.data_out(wire_d5_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance653(.data_in(wire_d5_2),.data_out(wire_d5_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance654(.data_in(wire_d5_3),.data_out(wire_d5_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance655(.data_in(wire_d5_4),.data_out(wire_d5_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance656(.data_in(wire_d5_5),.data_out(wire_d5_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance657(.data_in(wire_d5_6),.data_out(wire_d5_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance658(.data_in(wire_d5_7),.data_out(wire_d5_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance659(.data_in(wire_d5_8),.data_out(wire_d5_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6510(.data_in(wire_d5_9),.data_out(wire_d5_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6511(.data_in(wire_d5_10),.data_out(wire_d5_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6512(.data_in(wire_d5_11),.data_out(wire_d5_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6513(.data_in(wire_d5_12),.data_out(wire_d5_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6514(.data_in(wire_d5_13),.data_out(wire_d5_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6515(.data_in(wire_d5_14),.data_out(wire_d5_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6516(.data_in(wire_d5_15),.data_out(wire_d5_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6517(.data_in(wire_d5_16),.data_out(wire_d5_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6518(.data_in(wire_d5_17),.data_out(wire_d5_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6519(.data_in(wire_d5_18),.data_out(wire_d5_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6520(.data_in(wire_d5_19),.data_out(wire_d5_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6521(.data_in(wire_d5_20),.data_out(wire_d5_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6522(.data_in(wire_d5_21),.data_out(wire_d5_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6523(.data_in(wire_d5_22),.data_out(wire_d5_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6524(.data_in(wire_d5_23),.data_out(wire_d5_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6525(.data_in(wire_d5_24),.data_out(wire_d5_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6526(.data_in(wire_d5_25),.data_out(wire_d5_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6527(.data_in(wire_d5_26),.data_out(wire_d5_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6528(.data_in(wire_d5_27),.data_out(wire_d5_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6529(.data_in(wire_d5_28),.data_out(wire_d5_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6530(.data_in(wire_d5_29),.data_out(wire_d5_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6531(.data_in(wire_d5_30),.data_out(wire_d5_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6532(.data_in(wire_d5_31),.data_out(wire_d5_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6533(.data_in(wire_d5_32),.data_out(wire_d5_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6534(.data_in(wire_d5_33),.data_out(wire_d5_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6535(.data_in(wire_d5_34),.data_out(wire_d5_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6536(.data_in(wire_d5_35),.data_out(wire_d5_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6537(.data_in(wire_d5_36),.data_out(wire_d5_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6538(.data_in(wire_d5_37),.data_out(wire_d5_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6539(.data_in(wire_d5_38),.data_out(wire_d5_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6540(.data_in(wire_d5_39),.data_out(wire_d5_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6541(.data_in(wire_d5_40),.data_out(wire_d5_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6542(.data_in(wire_d5_41),.data_out(wire_d5_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6543(.data_in(wire_d5_42),.data_out(wire_d5_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6544(.data_in(wire_d5_43),.data_out(wire_d5_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6545(.data_in(wire_d5_44),.data_out(wire_d5_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6546(.data_in(wire_d5_45),.data_out(wire_d5_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6547(.data_in(wire_d5_46),.data_out(wire_d5_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6548(.data_in(wire_d5_47),.data_out(wire_d5_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6549(.data_in(wire_d5_48),.data_out(wire_d5_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6550(.data_in(wire_d5_49),.data_out(wire_d5_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6551(.data_in(wire_d5_50),.data_out(wire_d5_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6552(.data_in(wire_d5_51),.data_out(wire_d5_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6553(.data_in(wire_d5_52),.data_out(wire_d5_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6554(.data_in(wire_d5_53),.data_out(wire_d5_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6555(.data_in(wire_d5_54),.data_out(wire_d5_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6556(.data_in(wire_d5_55),.data_out(wire_d5_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6557(.data_in(wire_d5_56),.data_out(wire_d5_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6558(.data_in(wire_d5_57),.data_out(wire_d5_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6559(.data_in(wire_d5_58),.data_out(wire_d5_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6560(.data_in(wire_d5_59),.data_out(wire_d5_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6561(.data_in(wire_d5_60),.data_out(wire_d5_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6562(.data_in(wire_d5_61),.data_out(wire_d5_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6563(.data_in(wire_d5_62),.data_out(wire_d5_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6564(.data_in(wire_d5_63),.data_out(wire_d5_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6565(.data_in(wire_d5_64),.data_out(wire_d5_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6566(.data_in(wire_d5_65),.data_out(wire_d5_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6567(.data_in(wire_d5_66),.data_out(wire_d5_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6568(.data_in(wire_d5_67),.data_out(wire_d5_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6569(.data_in(wire_d5_68),.data_out(d_out5),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance760(.data_in(d_in6),.data_out(wire_d6_0),.clk(clk),.rst(rst));            //channel 7
	encoder #(.WIDTH(WIDTH)) encoder_instance761(.data_in(wire_d6_0),.data_out(wire_d6_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance762(.data_in(wire_d6_1),.data_out(wire_d6_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance763(.data_in(wire_d6_2),.data_out(wire_d6_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance764(.data_in(wire_d6_3),.data_out(wire_d6_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance765(.data_in(wire_d6_4),.data_out(wire_d6_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance766(.data_in(wire_d6_5),.data_out(wire_d6_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767(.data_in(wire_d6_6),.data_out(wire_d6_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance768(.data_in(wire_d6_7),.data_out(wire_d6_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance769(.data_in(wire_d6_8),.data_out(wire_d6_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7610(.data_in(wire_d6_9),.data_out(wire_d6_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7611(.data_in(wire_d6_10),.data_out(wire_d6_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7612(.data_in(wire_d6_11),.data_out(wire_d6_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7613(.data_in(wire_d6_12),.data_out(wire_d6_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7614(.data_in(wire_d6_13),.data_out(wire_d6_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7615(.data_in(wire_d6_14),.data_out(wire_d6_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7616(.data_in(wire_d6_15),.data_out(wire_d6_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7617(.data_in(wire_d6_16),.data_out(wire_d6_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7618(.data_in(wire_d6_17),.data_out(wire_d6_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7619(.data_in(wire_d6_18),.data_out(wire_d6_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7620(.data_in(wire_d6_19),.data_out(wire_d6_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7621(.data_in(wire_d6_20),.data_out(wire_d6_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7622(.data_in(wire_d6_21),.data_out(wire_d6_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7623(.data_in(wire_d6_22),.data_out(wire_d6_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7624(.data_in(wire_d6_23),.data_out(wire_d6_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7625(.data_in(wire_d6_24),.data_out(wire_d6_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7626(.data_in(wire_d6_25),.data_out(wire_d6_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7627(.data_in(wire_d6_26),.data_out(wire_d6_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7628(.data_in(wire_d6_27),.data_out(wire_d6_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7629(.data_in(wire_d6_28),.data_out(wire_d6_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7630(.data_in(wire_d6_29),.data_out(wire_d6_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7631(.data_in(wire_d6_30),.data_out(wire_d6_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7632(.data_in(wire_d6_31),.data_out(wire_d6_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7633(.data_in(wire_d6_32),.data_out(wire_d6_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7634(.data_in(wire_d6_33),.data_out(wire_d6_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7635(.data_in(wire_d6_34),.data_out(wire_d6_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7636(.data_in(wire_d6_35),.data_out(wire_d6_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7637(.data_in(wire_d6_36),.data_out(wire_d6_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7638(.data_in(wire_d6_37),.data_out(wire_d6_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7639(.data_in(wire_d6_38),.data_out(wire_d6_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7640(.data_in(wire_d6_39),.data_out(wire_d6_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7641(.data_in(wire_d6_40),.data_out(wire_d6_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7642(.data_in(wire_d6_41),.data_out(wire_d6_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7643(.data_in(wire_d6_42),.data_out(wire_d6_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7644(.data_in(wire_d6_43),.data_out(wire_d6_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7645(.data_in(wire_d6_44),.data_out(wire_d6_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7646(.data_in(wire_d6_45),.data_out(wire_d6_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7647(.data_in(wire_d6_46),.data_out(wire_d6_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7648(.data_in(wire_d6_47),.data_out(wire_d6_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7649(.data_in(wire_d6_48),.data_out(wire_d6_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7650(.data_in(wire_d6_49),.data_out(wire_d6_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7651(.data_in(wire_d6_50),.data_out(wire_d6_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7652(.data_in(wire_d6_51),.data_out(wire_d6_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7653(.data_in(wire_d6_52),.data_out(wire_d6_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7654(.data_in(wire_d6_53),.data_out(wire_d6_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7655(.data_in(wire_d6_54),.data_out(wire_d6_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7656(.data_in(wire_d6_55),.data_out(wire_d6_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7657(.data_in(wire_d6_56),.data_out(wire_d6_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7658(.data_in(wire_d6_57),.data_out(wire_d6_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7659(.data_in(wire_d6_58),.data_out(wire_d6_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7660(.data_in(wire_d6_59),.data_out(wire_d6_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7661(.data_in(wire_d6_60),.data_out(wire_d6_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7662(.data_in(wire_d6_61),.data_out(wire_d6_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7663(.data_in(wire_d6_62),.data_out(wire_d6_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7664(.data_in(wire_d6_63),.data_out(wire_d6_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7665(.data_in(wire_d6_64),.data_out(wire_d6_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7666(.data_in(wire_d6_65),.data_out(wire_d6_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7667(.data_in(wire_d6_66),.data_out(wire_d6_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7668(.data_in(wire_d6_67),.data_out(wire_d6_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7669(.data_in(wire_d6_68),.data_out(d_out6),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance870(.data_in(d_in7),.data_out(wire_d7_0),.clk(clk),.rst(rst));            //channel 8
	encoder #(.WIDTH(WIDTH)) encoder_instance871(.data_in(wire_d7_0),.data_out(wire_d7_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance872(.data_in(wire_d7_1),.data_out(wire_d7_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance873(.data_in(wire_d7_2),.data_out(wire_d7_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance874(.data_in(wire_d7_3),.data_out(wire_d7_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance875(.data_in(wire_d7_4),.data_out(wire_d7_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance876(.data_in(wire_d7_5),.data_out(wire_d7_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance877(.data_in(wire_d7_6),.data_out(wire_d7_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878(.data_in(wire_d7_7),.data_out(wire_d7_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance879(.data_in(wire_d7_8),.data_out(wire_d7_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8710(.data_in(wire_d7_9),.data_out(wire_d7_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8711(.data_in(wire_d7_10),.data_out(wire_d7_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8712(.data_in(wire_d7_11),.data_out(wire_d7_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8713(.data_in(wire_d7_12),.data_out(wire_d7_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8714(.data_in(wire_d7_13),.data_out(wire_d7_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8715(.data_in(wire_d7_14),.data_out(wire_d7_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8716(.data_in(wire_d7_15),.data_out(wire_d7_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8717(.data_in(wire_d7_16),.data_out(wire_d7_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8718(.data_in(wire_d7_17),.data_out(wire_d7_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8719(.data_in(wire_d7_18),.data_out(wire_d7_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8720(.data_in(wire_d7_19),.data_out(wire_d7_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8721(.data_in(wire_d7_20),.data_out(wire_d7_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8722(.data_in(wire_d7_21),.data_out(wire_d7_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8723(.data_in(wire_d7_22),.data_out(wire_d7_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8724(.data_in(wire_d7_23),.data_out(wire_d7_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8725(.data_in(wire_d7_24),.data_out(wire_d7_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8726(.data_in(wire_d7_25),.data_out(wire_d7_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8727(.data_in(wire_d7_26),.data_out(wire_d7_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8728(.data_in(wire_d7_27),.data_out(wire_d7_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8729(.data_in(wire_d7_28),.data_out(wire_d7_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8730(.data_in(wire_d7_29),.data_out(wire_d7_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8731(.data_in(wire_d7_30),.data_out(wire_d7_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8732(.data_in(wire_d7_31),.data_out(wire_d7_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8733(.data_in(wire_d7_32),.data_out(wire_d7_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8734(.data_in(wire_d7_33),.data_out(wire_d7_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8735(.data_in(wire_d7_34),.data_out(wire_d7_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8736(.data_in(wire_d7_35),.data_out(wire_d7_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8737(.data_in(wire_d7_36),.data_out(wire_d7_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8738(.data_in(wire_d7_37),.data_out(wire_d7_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8739(.data_in(wire_d7_38),.data_out(wire_d7_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8740(.data_in(wire_d7_39),.data_out(wire_d7_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8741(.data_in(wire_d7_40),.data_out(wire_d7_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8742(.data_in(wire_d7_41),.data_out(wire_d7_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8743(.data_in(wire_d7_42),.data_out(wire_d7_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8744(.data_in(wire_d7_43),.data_out(wire_d7_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8745(.data_in(wire_d7_44),.data_out(wire_d7_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8746(.data_in(wire_d7_45),.data_out(wire_d7_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8747(.data_in(wire_d7_46),.data_out(wire_d7_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8748(.data_in(wire_d7_47),.data_out(wire_d7_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8749(.data_in(wire_d7_48),.data_out(wire_d7_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8750(.data_in(wire_d7_49),.data_out(wire_d7_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8751(.data_in(wire_d7_50),.data_out(wire_d7_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8752(.data_in(wire_d7_51),.data_out(wire_d7_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8753(.data_in(wire_d7_52),.data_out(wire_d7_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8754(.data_in(wire_d7_53),.data_out(wire_d7_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8755(.data_in(wire_d7_54),.data_out(wire_d7_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8756(.data_in(wire_d7_55),.data_out(wire_d7_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8757(.data_in(wire_d7_56),.data_out(wire_d7_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8758(.data_in(wire_d7_57),.data_out(wire_d7_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8759(.data_in(wire_d7_58),.data_out(wire_d7_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8760(.data_in(wire_d7_59),.data_out(wire_d7_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8761(.data_in(wire_d7_60),.data_out(wire_d7_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8762(.data_in(wire_d7_61),.data_out(wire_d7_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8763(.data_in(wire_d7_62),.data_out(wire_d7_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8764(.data_in(wire_d7_63),.data_out(wire_d7_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8765(.data_in(wire_d7_64),.data_out(wire_d7_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8766(.data_in(wire_d7_65),.data_out(wire_d7_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8767(.data_in(wire_d7_66),.data_out(wire_d7_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8768(.data_in(wire_d7_67),.data_out(wire_d7_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8769(.data_in(wire_d7_68),.data_out(d_out7),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance980(.data_in(d_in8),.data_out(wire_d8_0),.clk(clk),.rst(rst));            //channel 9
	register #(.WIDTH(WIDTH)) register_instance981(.data_in(wire_d8_0),.data_out(wire_d8_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance982(.data_in(wire_d8_1),.data_out(wire_d8_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance983(.data_in(wire_d8_2),.data_out(wire_d8_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance984(.data_in(wire_d8_3),.data_out(wire_d8_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance985(.data_in(wire_d8_4),.data_out(wire_d8_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance986(.data_in(wire_d8_5),.data_out(wire_d8_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance987(.data_in(wire_d8_6),.data_out(wire_d8_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance988(.data_in(wire_d8_7),.data_out(wire_d8_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance989(.data_in(wire_d8_8),.data_out(wire_d8_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9810(.data_in(wire_d8_9),.data_out(wire_d8_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9811(.data_in(wire_d8_10),.data_out(wire_d8_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9812(.data_in(wire_d8_11),.data_out(wire_d8_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9813(.data_in(wire_d8_12),.data_out(wire_d8_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9814(.data_in(wire_d8_13),.data_out(wire_d8_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9815(.data_in(wire_d8_14),.data_out(wire_d8_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9816(.data_in(wire_d8_15),.data_out(wire_d8_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9817(.data_in(wire_d8_16),.data_out(wire_d8_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9818(.data_in(wire_d8_17),.data_out(wire_d8_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9819(.data_in(wire_d8_18),.data_out(wire_d8_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9820(.data_in(wire_d8_19),.data_out(wire_d8_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9821(.data_in(wire_d8_20),.data_out(wire_d8_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9822(.data_in(wire_d8_21),.data_out(wire_d8_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9823(.data_in(wire_d8_22),.data_out(wire_d8_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9824(.data_in(wire_d8_23),.data_out(wire_d8_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9825(.data_in(wire_d8_24),.data_out(wire_d8_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9826(.data_in(wire_d8_25),.data_out(wire_d8_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9827(.data_in(wire_d8_26),.data_out(wire_d8_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9828(.data_in(wire_d8_27),.data_out(wire_d8_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9829(.data_in(wire_d8_28),.data_out(wire_d8_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9830(.data_in(wire_d8_29),.data_out(wire_d8_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9831(.data_in(wire_d8_30),.data_out(wire_d8_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9832(.data_in(wire_d8_31),.data_out(wire_d8_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9833(.data_in(wire_d8_32),.data_out(wire_d8_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9834(.data_in(wire_d8_33),.data_out(wire_d8_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9835(.data_in(wire_d8_34),.data_out(wire_d8_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9836(.data_in(wire_d8_35),.data_out(wire_d8_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9837(.data_in(wire_d8_36),.data_out(wire_d8_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9838(.data_in(wire_d8_37),.data_out(wire_d8_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9839(.data_in(wire_d8_38),.data_out(wire_d8_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9840(.data_in(wire_d8_39),.data_out(wire_d8_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9841(.data_in(wire_d8_40),.data_out(wire_d8_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9842(.data_in(wire_d8_41),.data_out(wire_d8_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9843(.data_in(wire_d8_42),.data_out(wire_d8_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9844(.data_in(wire_d8_43),.data_out(wire_d8_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9845(.data_in(wire_d8_44),.data_out(wire_d8_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9846(.data_in(wire_d8_45),.data_out(wire_d8_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9847(.data_in(wire_d8_46),.data_out(wire_d8_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9848(.data_in(wire_d8_47),.data_out(wire_d8_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9849(.data_in(wire_d8_48),.data_out(wire_d8_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9850(.data_in(wire_d8_49),.data_out(wire_d8_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9851(.data_in(wire_d8_50),.data_out(wire_d8_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9852(.data_in(wire_d8_51),.data_out(wire_d8_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9853(.data_in(wire_d8_52),.data_out(wire_d8_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9854(.data_in(wire_d8_53),.data_out(wire_d8_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9855(.data_in(wire_d8_54),.data_out(wire_d8_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9856(.data_in(wire_d8_55),.data_out(wire_d8_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9857(.data_in(wire_d8_56),.data_out(wire_d8_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9858(.data_in(wire_d8_57),.data_out(wire_d8_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9859(.data_in(wire_d8_58),.data_out(wire_d8_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9860(.data_in(wire_d8_59),.data_out(wire_d8_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9861(.data_in(wire_d8_60),.data_out(wire_d8_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9862(.data_in(wire_d8_61),.data_out(wire_d8_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9863(.data_in(wire_d8_62),.data_out(wire_d8_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9864(.data_in(wire_d8_63),.data_out(wire_d8_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9865(.data_in(wire_d8_64),.data_out(wire_d8_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9866(.data_in(wire_d8_65),.data_out(wire_d8_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9867(.data_in(wire_d8_66),.data_out(wire_d8_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9868(.data_in(wire_d8_67),.data_out(wire_d8_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9869(.data_in(wire_d8_68),.data_out(d_out8),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance1090(.data_in(d_in9),.data_out(wire_d9_0),.clk(clk),.rst(rst));            //channel 10
	invertion #(.WIDTH(WIDTH)) invertion_instance1091(.data_in(wire_d9_0),.data_out(wire_d9_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1092(.data_in(wire_d9_1),.data_out(wire_d9_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1093(.data_in(wire_d9_2),.data_out(wire_d9_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1094(.data_in(wire_d9_3),.data_out(wire_d9_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1095(.data_in(wire_d9_4),.data_out(wire_d9_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1096(.data_in(wire_d9_5),.data_out(wire_d9_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1097(.data_in(wire_d9_6),.data_out(wire_d9_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1098(.data_in(wire_d9_7),.data_out(wire_d9_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1099(.data_in(wire_d9_8),.data_out(wire_d9_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10910(.data_in(wire_d9_9),.data_out(wire_d9_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10911(.data_in(wire_d9_10),.data_out(wire_d9_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10912(.data_in(wire_d9_11),.data_out(wire_d9_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10913(.data_in(wire_d9_12),.data_out(wire_d9_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10914(.data_in(wire_d9_13),.data_out(wire_d9_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10915(.data_in(wire_d9_14),.data_out(wire_d9_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10916(.data_in(wire_d9_15),.data_out(wire_d9_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10917(.data_in(wire_d9_16),.data_out(wire_d9_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10918(.data_in(wire_d9_17),.data_out(wire_d9_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10919(.data_in(wire_d9_18),.data_out(wire_d9_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10920(.data_in(wire_d9_19),.data_out(wire_d9_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10921(.data_in(wire_d9_20),.data_out(wire_d9_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10922(.data_in(wire_d9_21),.data_out(wire_d9_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10923(.data_in(wire_d9_22),.data_out(wire_d9_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10924(.data_in(wire_d9_23),.data_out(wire_d9_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10925(.data_in(wire_d9_24),.data_out(wire_d9_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10926(.data_in(wire_d9_25),.data_out(wire_d9_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10927(.data_in(wire_d9_26),.data_out(wire_d9_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10928(.data_in(wire_d9_27),.data_out(wire_d9_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10929(.data_in(wire_d9_28),.data_out(wire_d9_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10930(.data_in(wire_d9_29),.data_out(wire_d9_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10931(.data_in(wire_d9_30),.data_out(wire_d9_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10932(.data_in(wire_d9_31),.data_out(wire_d9_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10933(.data_in(wire_d9_32),.data_out(wire_d9_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10934(.data_in(wire_d9_33),.data_out(wire_d9_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10935(.data_in(wire_d9_34),.data_out(wire_d9_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10936(.data_in(wire_d9_35),.data_out(wire_d9_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10937(.data_in(wire_d9_36),.data_out(wire_d9_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10938(.data_in(wire_d9_37),.data_out(wire_d9_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10939(.data_in(wire_d9_38),.data_out(wire_d9_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10940(.data_in(wire_d9_39),.data_out(wire_d9_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10941(.data_in(wire_d9_40),.data_out(wire_d9_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10942(.data_in(wire_d9_41),.data_out(wire_d9_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10943(.data_in(wire_d9_42),.data_out(wire_d9_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10944(.data_in(wire_d9_43),.data_out(wire_d9_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10945(.data_in(wire_d9_44),.data_out(wire_d9_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10946(.data_in(wire_d9_45),.data_out(wire_d9_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10947(.data_in(wire_d9_46),.data_out(wire_d9_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10948(.data_in(wire_d9_47),.data_out(wire_d9_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10949(.data_in(wire_d9_48),.data_out(wire_d9_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10950(.data_in(wire_d9_49),.data_out(wire_d9_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10951(.data_in(wire_d9_50),.data_out(wire_d9_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10952(.data_in(wire_d9_51),.data_out(wire_d9_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10953(.data_in(wire_d9_52),.data_out(wire_d9_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10954(.data_in(wire_d9_53),.data_out(wire_d9_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10955(.data_in(wire_d9_54),.data_out(wire_d9_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10956(.data_in(wire_d9_55),.data_out(wire_d9_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10957(.data_in(wire_d9_56),.data_out(wire_d9_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10958(.data_in(wire_d9_57),.data_out(wire_d9_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10959(.data_in(wire_d9_58),.data_out(wire_d9_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10960(.data_in(wire_d9_59),.data_out(wire_d9_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10961(.data_in(wire_d9_60),.data_out(wire_d9_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10962(.data_in(wire_d9_61),.data_out(wire_d9_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10963(.data_in(wire_d9_62),.data_out(wire_d9_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10964(.data_in(wire_d9_63),.data_out(wire_d9_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10965(.data_in(wire_d9_64),.data_out(wire_d9_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10966(.data_in(wire_d9_65),.data_out(wire_d9_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10967(.data_in(wire_d9_66),.data_out(wire_d9_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10968(.data_in(wire_d9_67),.data_out(wire_d9_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10969(.data_in(wire_d9_68),.data_out(d_out9),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance11100(.data_in(d_in10),.data_out(wire_d10_0),.clk(clk),.rst(rst));            //channel 11
	encoder #(.WIDTH(WIDTH)) encoder_instance11101(.data_in(wire_d10_0),.data_out(wire_d10_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance11102(.data_in(wire_d10_1),.data_out(wire_d10_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance11103(.data_in(wire_d10_2),.data_out(wire_d10_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance11104(.data_in(wire_d10_3),.data_out(wire_d10_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance11105(.data_in(wire_d10_4),.data_out(wire_d10_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance11106(.data_in(wire_d10_5),.data_out(wire_d10_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance11107(.data_in(wire_d10_6),.data_out(wire_d10_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance11108(.data_in(wire_d10_7),.data_out(wire_d10_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance11109(.data_in(wire_d10_8),.data_out(wire_d10_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111010(.data_in(wire_d10_9),.data_out(wire_d10_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111011(.data_in(wire_d10_10),.data_out(wire_d10_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111012(.data_in(wire_d10_11),.data_out(wire_d10_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111013(.data_in(wire_d10_12),.data_out(wire_d10_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111014(.data_in(wire_d10_13),.data_out(wire_d10_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111015(.data_in(wire_d10_14),.data_out(wire_d10_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111016(.data_in(wire_d10_15),.data_out(wire_d10_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111017(.data_in(wire_d10_16),.data_out(wire_d10_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111018(.data_in(wire_d10_17),.data_out(wire_d10_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111019(.data_in(wire_d10_18),.data_out(wire_d10_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111020(.data_in(wire_d10_19),.data_out(wire_d10_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111021(.data_in(wire_d10_20),.data_out(wire_d10_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111022(.data_in(wire_d10_21),.data_out(wire_d10_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111023(.data_in(wire_d10_22),.data_out(wire_d10_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111024(.data_in(wire_d10_23),.data_out(wire_d10_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111025(.data_in(wire_d10_24),.data_out(wire_d10_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111026(.data_in(wire_d10_25),.data_out(wire_d10_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111027(.data_in(wire_d10_26),.data_out(wire_d10_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111028(.data_in(wire_d10_27),.data_out(wire_d10_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111029(.data_in(wire_d10_28),.data_out(wire_d10_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111030(.data_in(wire_d10_29),.data_out(wire_d10_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111031(.data_in(wire_d10_30),.data_out(wire_d10_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111032(.data_in(wire_d10_31),.data_out(wire_d10_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111033(.data_in(wire_d10_32),.data_out(wire_d10_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111034(.data_in(wire_d10_33),.data_out(wire_d10_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111035(.data_in(wire_d10_34),.data_out(wire_d10_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111036(.data_in(wire_d10_35),.data_out(wire_d10_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111037(.data_in(wire_d10_36),.data_out(wire_d10_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111038(.data_in(wire_d10_37),.data_out(wire_d10_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111039(.data_in(wire_d10_38),.data_out(wire_d10_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111040(.data_in(wire_d10_39),.data_out(wire_d10_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111041(.data_in(wire_d10_40),.data_out(wire_d10_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111042(.data_in(wire_d10_41),.data_out(wire_d10_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111043(.data_in(wire_d10_42),.data_out(wire_d10_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111044(.data_in(wire_d10_43),.data_out(wire_d10_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111045(.data_in(wire_d10_44),.data_out(wire_d10_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111046(.data_in(wire_d10_45),.data_out(wire_d10_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111047(.data_in(wire_d10_46),.data_out(wire_d10_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111048(.data_in(wire_d10_47),.data_out(wire_d10_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111049(.data_in(wire_d10_48),.data_out(wire_d10_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111050(.data_in(wire_d10_49),.data_out(wire_d10_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111051(.data_in(wire_d10_50),.data_out(wire_d10_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111052(.data_in(wire_d10_51),.data_out(wire_d10_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111053(.data_in(wire_d10_52),.data_out(wire_d10_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111054(.data_in(wire_d10_53),.data_out(wire_d10_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111055(.data_in(wire_d10_54),.data_out(wire_d10_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111056(.data_in(wire_d10_55),.data_out(wire_d10_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111057(.data_in(wire_d10_56),.data_out(wire_d10_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111058(.data_in(wire_d10_57),.data_out(wire_d10_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111059(.data_in(wire_d10_58),.data_out(wire_d10_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111060(.data_in(wire_d10_59),.data_out(wire_d10_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111061(.data_in(wire_d10_60),.data_out(wire_d10_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111062(.data_in(wire_d10_61),.data_out(wire_d10_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111063(.data_in(wire_d10_62),.data_out(wire_d10_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111064(.data_in(wire_d10_63),.data_out(wire_d10_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111065(.data_in(wire_d10_64),.data_out(wire_d10_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111066(.data_in(wire_d10_65),.data_out(wire_d10_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111067(.data_in(wire_d10_66),.data_out(wire_d10_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111068(.data_in(wire_d10_67),.data_out(wire_d10_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111069(.data_in(wire_d10_68),.data_out(d_out10),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance12110(.data_in(d_in11),.data_out(wire_d11_0),.clk(clk),.rst(rst));            //channel 12
	invertion #(.WIDTH(WIDTH)) invertion_instance12111(.data_in(wire_d11_0),.data_out(wire_d11_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance12112(.data_in(wire_d11_1),.data_out(wire_d11_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance12113(.data_in(wire_d11_2),.data_out(wire_d11_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance12114(.data_in(wire_d11_3),.data_out(wire_d11_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance12115(.data_in(wire_d11_4),.data_out(wire_d11_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance12116(.data_in(wire_d11_5),.data_out(wire_d11_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance12117(.data_in(wire_d11_6),.data_out(wire_d11_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance12118(.data_in(wire_d11_7),.data_out(wire_d11_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance12119(.data_in(wire_d11_8),.data_out(wire_d11_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121110(.data_in(wire_d11_9),.data_out(wire_d11_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121111(.data_in(wire_d11_10),.data_out(wire_d11_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121112(.data_in(wire_d11_11),.data_out(wire_d11_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121113(.data_in(wire_d11_12),.data_out(wire_d11_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121114(.data_in(wire_d11_13),.data_out(wire_d11_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121115(.data_in(wire_d11_14),.data_out(wire_d11_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121116(.data_in(wire_d11_15),.data_out(wire_d11_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121117(.data_in(wire_d11_16),.data_out(wire_d11_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121118(.data_in(wire_d11_17),.data_out(wire_d11_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121119(.data_in(wire_d11_18),.data_out(wire_d11_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121120(.data_in(wire_d11_19),.data_out(wire_d11_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121121(.data_in(wire_d11_20),.data_out(wire_d11_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121122(.data_in(wire_d11_21),.data_out(wire_d11_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121123(.data_in(wire_d11_22),.data_out(wire_d11_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121124(.data_in(wire_d11_23),.data_out(wire_d11_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121125(.data_in(wire_d11_24),.data_out(wire_d11_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121126(.data_in(wire_d11_25),.data_out(wire_d11_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121127(.data_in(wire_d11_26),.data_out(wire_d11_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121128(.data_in(wire_d11_27),.data_out(wire_d11_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121129(.data_in(wire_d11_28),.data_out(wire_d11_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121130(.data_in(wire_d11_29),.data_out(wire_d11_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121131(.data_in(wire_d11_30),.data_out(wire_d11_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121132(.data_in(wire_d11_31),.data_out(wire_d11_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121133(.data_in(wire_d11_32),.data_out(wire_d11_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121134(.data_in(wire_d11_33),.data_out(wire_d11_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121135(.data_in(wire_d11_34),.data_out(wire_d11_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121136(.data_in(wire_d11_35),.data_out(wire_d11_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121137(.data_in(wire_d11_36),.data_out(wire_d11_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121138(.data_in(wire_d11_37),.data_out(wire_d11_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121139(.data_in(wire_d11_38),.data_out(wire_d11_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121140(.data_in(wire_d11_39),.data_out(wire_d11_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121141(.data_in(wire_d11_40),.data_out(wire_d11_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121142(.data_in(wire_d11_41),.data_out(wire_d11_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121143(.data_in(wire_d11_42),.data_out(wire_d11_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121144(.data_in(wire_d11_43),.data_out(wire_d11_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121145(.data_in(wire_d11_44),.data_out(wire_d11_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121146(.data_in(wire_d11_45),.data_out(wire_d11_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121147(.data_in(wire_d11_46),.data_out(wire_d11_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121148(.data_in(wire_d11_47),.data_out(wire_d11_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121149(.data_in(wire_d11_48),.data_out(wire_d11_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121150(.data_in(wire_d11_49),.data_out(wire_d11_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121151(.data_in(wire_d11_50),.data_out(wire_d11_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121152(.data_in(wire_d11_51),.data_out(wire_d11_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121153(.data_in(wire_d11_52),.data_out(wire_d11_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121154(.data_in(wire_d11_53),.data_out(wire_d11_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121155(.data_in(wire_d11_54),.data_out(wire_d11_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121156(.data_in(wire_d11_55),.data_out(wire_d11_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121157(.data_in(wire_d11_56),.data_out(wire_d11_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121158(.data_in(wire_d11_57),.data_out(wire_d11_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121159(.data_in(wire_d11_58),.data_out(wire_d11_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121160(.data_in(wire_d11_59),.data_out(wire_d11_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121161(.data_in(wire_d11_60),.data_out(wire_d11_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121162(.data_in(wire_d11_61),.data_out(wire_d11_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121163(.data_in(wire_d11_62),.data_out(wire_d11_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121164(.data_in(wire_d11_63),.data_out(wire_d11_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121165(.data_in(wire_d11_64),.data_out(wire_d11_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121166(.data_in(wire_d11_65),.data_out(wire_d11_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121167(.data_in(wire_d11_66),.data_out(wire_d11_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121168(.data_in(wire_d11_67),.data_out(wire_d11_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121169(.data_in(wire_d11_68),.data_out(d_out11),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance13120(.data_in(d_in12),.data_out(wire_d12_0),.clk(clk),.rst(rst));            //channel 13
	invertion #(.WIDTH(WIDTH)) invertion_instance13121(.data_in(wire_d12_0),.data_out(wire_d12_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance13122(.data_in(wire_d12_1),.data_out(wire_d12_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance13123(.data_in(wire_d12_2),.data_out(wire_d12_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance13124(.data_in(wire_d12_3),.data_out(wire_d12_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance13125(.data_in(wire_d12_4),.data_out(wire_d12_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance13126(.data_in(wire_d12_5),.data_out(wire_d12_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance13127(.data_in(wire_d12_6),.data_out(wire_d12_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance13128(.data_in(wire_d12_7),.data_out(wire_d12_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance13129(.data_in(wire_d12_8),.data_out(wire_d12_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131210(.data_in(wire_d12_9),.data_out(wire_d12_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131211(.data_in(wire_d12_10),.data_out(wire_d12_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131212(.data_in(wire_d12_11),.data_out(wire_d12_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131213(.data_in(wire_d12_12),.data_out(wire_d12_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131214(.data_in(wire_d12_13),.data_out(wire_d12_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131215(.data_in(wire_d12_14),.data_out(wire_d12_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131216(.data_in(wire_d12_15),.data_out(wire_d12_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131217(.data_in(wire_d12_16),.data_out(wire_d12_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131218(.data_in(wire_d12_17),.data_out(wire_d12_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131219(.data_in(wire_d12_18),.data_out(wire_d12_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131220(.data_in(wire_d12_19),.data_out(wire_d12_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131221(.data_in(wire_d12_20),.data_out(wire_d12_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131222(.data_in(wire_d12_21),.data_out(wire_d12_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131223(.data_in(wire_d12_22),.data_out(wire_d12_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131224(.data_in(wire_d12_23),.data_out(wire_d12_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131225(.data_in(wire_d12_24),.data_out(wire_d12_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131226(.data_in(wire_d12_25),.data_out(wire_d12_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131227(.data_in(wire_d12_26),.data_out(wire_d12_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131228(.data_in(wire_d12_27),.data_out(wire_d12_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131229(.data_in(wire_d12_28),.data_out(wire_d12_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131230(.data_in(wire_d12_29),.data_out(wire_d12_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131231(.data_in(wire_d12_30),.data_out(wire_d12_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131232(.data_in(wire_d12_31),.data_out(wire_d12_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131233(.data_in(wire_d12_32),.data_out(wire_d12_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131234(.data_in(wire_d12_33),.data_out(wire_d12_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131235(.data_in(wire_d12_34),.data_out(wire_d12_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131236(.data_in(wire_d12_35),.data_out(wire_d12_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131237(.data_in(wire_d12_36),.data_out(wire_d12_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131238(.data_in(wire_d12_37),.data_out(wire_d12_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131239(.data_in(wire_d12_38),.data_out(wire_d12_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131240(.data_in(wire_d12_39),.data_out(wire_d12_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131241(.data_in(wire_d12_40),.data_out(wire_d12_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131242(.data_in(wire_d12_41),.data_out(wire_d12_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131243(.data_in(wire_d12_42),.data_out(wire_d12_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131244(.data_in(wire_d12_43),.data_out(wire_d12_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131245(.data_in(wire_d12_44),.data_out(wire_d12_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131246(.data_in(wire_d12_45),.data_out(wire_d12_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131247(.data_in(wire_d12_46),.data_out(wire_d12_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131248(.data_in(wire_d12_47),.data_out(wire_d12_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131249(.data_in(wire_d12_48),.data_out(wire_d12_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131250(.data_in(wire_d12_49),.data_out(wire_d12_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131251(.data_in(wire_d12_50),.data_out(wire_d12_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131252(.data_in(wire_d12_51),.data_out(wire_d12_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131253(.data_in(wire_d12_52),.data_out(wire_d12_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131254(.data_in(wire_d12_53),.data_out(wire_d12_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131255(.data_in(wire_d12_54),.data_out(wire_d12_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131256(.data_in(wire_d12_55),.data_out(wire_d12_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131257(.data_in(wire_d12_56),.data_out(wire_d12_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131258(.data_in(wire_d12_57),.data_out(wire_d12_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131259(.data_in(wire_d12_58),.data_out(wire_d12_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131260(.data_in(wire_d12_59),.data_out(wire_d12_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131261(.data_in(wire_d12_60),.data_out(wire_d12_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131262(.data_in(wire_d12_61),.data_out(wire_d12_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131263(.data_in(wire_d12_62),.data_out(wire_d12_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131264(.data_in(wire_d12_63),.data_out(wire_d12_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131265(.data_in(wire_d12_64),.data_out(wire_d12_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131266(.data_in(wire_d12_65),.data_out(wire_d12_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131267(.data_in(wire_d12_66),.data_out(wire_d12_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131268(.data_in(wire_d12_67),.data_out(wire_d12_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131269(.data_in(wire_d12_68),.data_out(d_out12),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance14130(.data_in(d_in13),.data_out(wire_d13_0),.clk(clk),.rst(rst));            //channel 14
	invertion #(.WIDTH(WIDTH)) invertion_instance14131(.data_in(wire_d13_0),.data_out(wire_d13_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance14132(.data_in(wire_d13_1),.data_out(wire_d13_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance14133(.data_in(wire_d13_2),.data_out(wire_d13_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance14134(.data_in(wire_d13_3),.data_out(wire_d13_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance14135(.data_in(wire_d13_4),.data_out(wire_d13_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance14136(.data_in(wire_d13_5),.data_out(wire_d13_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance14137(.data_in(wire_d13_6),.data_out(wire_d13_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance14138(.data_in(wire_d13_7),.data_out(wire_d13_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance14139(.data_in(wire_d13_8),.data_out(wire_d13_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141310(.data_in(wire_d13_9),.data_out(wire_d13_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141311(.data_in(wire_d13_10),.data_out(wire_d13_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141312(.data_in(wire_d13_11),.data_out(wire_d13_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141313(.data_in(wire_d13_12),.data_out(wire_d13_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141314(.data_in(wire_d13_13),.data_out(wire_d13_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141315(.data_in(wire_d13_14),.data_out(wire_d13_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141316(.data_in(wire_d13_15),.data_out(wire_d13_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141317(.data_in(wire_d13_16),.data_out(wire_d13_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141318(.data_in(wire_d13_17),.data_out(wire_d13_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141319(.data_in(wire_d13_18),.data_out(wire_d13_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141320(.data_in(wire_d13_19),.data_out(wire_d13_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141321(.data_in(wire_d13_20),.data_out(wire_d13_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141322(.data_in(wire_d13_21),.data_out(wire_d13_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141323(.data_in(wire_d13_22),.data_out(wire_d13_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141324(.data_in(wire_d13_23),.data_out(wire_d13_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141325(.data_in(wire_d13_24),.data_out(wire_d13_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141326(.data_in(wire_d13_25),.data_out(wire_d13_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141327(.data_in(wire_d13_26),.data_out(wire_d13_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141328(.data_in(wire_d13_27),.data_out(wire_d13_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141329(.data_in(wire_d13_28),.data_out(wire_d13_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141330(.data_in(wire_d13_29),.data_out(wire_d13_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141331(.data_in(wire_d13_30),.data_out(wire_d13_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141332(.data_in(wire_d13_31),.data_out(wire_d13_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141333(.data_in(wire_d13_32),.data_out(wire_d13_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141334(.data_in(wire_d13_33),.data_out(wire_d13_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141335(.data_in(wire_d13_34),.data_out(wire_d13_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141336(.data_in(wire_d13_35),.data_out(wire_d13_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141337(.data_in(wire_d13_36),.data_out(wire_d13_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141338(.data_in(wire_d13_37),.data_out(wire_d13_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141339(.data_in(wire_d13_38),.data_out(wire_d13_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141340(.data_in(wire_d13_39),.data_out(wire_d13_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141341(.data_in(wire_d13_40),.data_out(wire_d13_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141342(.data_in(wire_d13_41),.data_out(wire_d13_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141343(.data_in(wire_d13_42),.data_out(wire_d13_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141344(.data_in(wire_d13_43),.data_out(wire_d13_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141345(.data_in(wire_d13_44),.data_out(wire_d13_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141346(.data_in(wire_d13_45),.data_out(wire_d13_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141347(.data_in(wire_d13_46),.data_out(wire_d13_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141348(.data_in(wire_d13_47),.data_out(wire_d13_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141349(.data_in(wire_d13_48),.data_out(wire_d13_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141350(.data_in(wire_d13_49),.data_out(wire_d13_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141351(.data_in(wire_d13_50),.data_out(wire_d13_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141352(.data_in(wire_d13_51),.data_out(wire_d13_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141353(.data_in(wire_d13_52),.data_out(wire_d13_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141354(.data_in(wire_d13_53),.data_out(wire_d13_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141355(.data_in(wire_d13_54),.data_out(wire_d13_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141356(.data_in(wire_d13_55),.data_out(wire_d13_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141357(.data_in(wire_d13_56),.data_out(wire_d13_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141358(.data_in(wire_d13_57),.data_out(wire_d13_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141359(.data_in(wire_d13_58),.data_out(wire_d13_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141360(.data_in(wire_d13_59),.data_out(wire_d13_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141361(.data_in(wire_d13_60),.data_out(wire_d13_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141362(.data_in(wire_d13_61),.data_out(wire_d13_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141363(.data_in(wire_d13_62),.data_out(wire_d13_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141364(.data_in(wire_d13_63),.data_out(wire_d13_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141365(.data_in(wire_d13_64),.data_out(wire_d13_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141366(.data_in(wire_d13_65),.data_out(wire_d13_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141367(.data_in(wire_d13_66),.data_out(wire_d13_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141368(.data_in(wire_d13_67),.data_out(wire_d13_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141369(.data_in(wire_d13_68),.data_out(d_out13),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance15140(.data_in(d_in14),.data_out(wire_d14_0),.clk(clk),.rst(rst));            //channel 15
	encoder #(.WIDTH(WIDTH)) encoder_instance15141(.data_in(wire_d14_0),.data_out(wire_d14_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance15142(.data_in(wire_d14_1),.data_out(wire_d14_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance15143(.data_in(wire_d14_2),.data_out(wire_d14_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance15144(.data_in(wire_d14_3),.data_out(wire_d14_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance15145(.data_in(wire_d14_4),.data_out(wire_d14_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance15146(.data_in(wire_d14_5),.data_out(wire_d14_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance15147(.data_in(wire_d14_6),.data_out(wire_d14_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance15148(.data_in(wire_d14_7),.data_out(wire_d14_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance15149(.data_in(wire_d14_8),.data_out(wire_d14_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151410(.data_in(wire_d14_9),.data_out(wire_d14_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151411(.data_in(wire_d14_10),.data_out(wire_d14_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151412(.data_in(wire_d14_11),.data_out(wire_d14_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151413(.data_in(wire_d14_12),.data_out(wire_d14_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151414(.data_in(wire_d14_13),.data_out(wire_d14_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151415(.data_in(wire_d14_14),.data_out(wire_d14_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151416(.data_in(wire_d14_15),.data_out(wire_d14_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151417(.data_in(wire_d14_16),.data_out(wire_d14_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151418(.data_in(wire_d14_17),.data_out(wire_d14_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151419(.data_in(wire_d14_18),.data_out(wire_d14_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151420(.data_in(wire_d14_19),.data_out(wire_d14_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151421(.data_in(wire_d14_20),.data_out(wire_d14_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151422(.data_in(wire_d14_21),.data_out(wire_d14_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151423(.data_in(wire_d14_22),.data_out(wire_d14_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151424(.data_in(wire_d14_23),.data_out(wire_d14_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151425(.data_in(wire_d14_24),.data_out(wire_d14_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151426(.data_in(wire_d14_25),.data_out(wire_d14_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151427(.data_in(wire_d14_26),.data_out(wire_d14_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151428(.data_in(wire_d14_27),.data_out(wire_d14_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151429(.data_in(wire_d14_28),.data_out(wire_d14_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151430(.data_in(wire_d14_29),.data_out(wire_d14_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151431(.data_in(wire_d14_30),.data_out(wire_d14_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151432(.data_in(wire_d14_31),.data_out(wire_d14_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151433(.data_in(wire_d14_32),.data_out(wire_d14_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151434(.data_in(wire_d14_33),.data_out(wire_d14_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151435(.data_in(wire_d14_34),.data_out(wire_d14_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151436(.data_in(wire_d14_35),.data_out(wire_d14_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151437(.data_in(wire_d14_36),.data_out(wire_d14_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151438(.data_in(wire_d14_37),.data_out(wire_d14_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151439(.data_in(wire_d14_38),.data_out(wire_d14_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151440(.data_in(wire_d14_39),.data_out(wire_d14_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151441(.data_in(wire_d14_40),.data_out(wire_d14_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151442(.data_in(wire_d14_41),.data_out(wire_d14_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151443(.data_in(wire_d14_42),.data_out(wire_d14_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151444(.data_in(wire_d14_43),.data_out(wire_d14_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151445(.data_in(wire_d14_44),.data_out(wire_d14_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151446(.data_in(wire_d14_45),.data_out(wire_d14_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151447(.data_in(wire_d14_46),.data_out(wire_d14_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151448(.data_in(wire_d14_47),.data_out(wire_d14_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151449(.data_in(wire_d14_48),.data_out(wire_d14_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151450(.data_in(wire_d14_49),.data_out(wire_d14_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151451(.data_in(wire_d14_50),.data_out(wire_d14_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151452(.data_in(wire_d14_51),.data_out(wire_d14_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151453(.data_in(wire_d14_52),.data_out(wire_d14_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151454(.data_in(wire_d14_53),.data_out(wire_d14_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151455(.data_in(wire_d14_54),.data_out(wire_d14_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151456(.data_in(wire_d14_55),.data_out(wire_d14_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151457(.data_in(wire_d14_56),.data_out(wire_d14_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151458(.data_in(wire_d14_57),.data_out(wire_d14_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151459(.data_in(wire_d14_58),.data_out(wire_d14_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151460(.data_in(wire_d14_59),.data_out(wire_d14_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151461(.data_in(wire_d14_60),.data_out(wire_d14_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151462(.data_in(wire_d14_61),.data_out(wire_d14_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151463(.data_in(wire_d14_62),.data_out(wire_d14_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151464(.data_in(wire_d14_63),.data_out(wire_d14_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151465(.data_in(wire_d14_64),.data_out(wire_d14_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151466(.data_in(wire_d14_65),.data_out(wire_d14_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151467(.data_in(wire_d14_66),.data_out(wire_d14_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151468(.data_in(wire_d14_67),.data_out(wire_d14_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151469(.data_in(wire_d14_68),.data_out(d_out14),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance16150(.data_in(d_in15),.data_out(wire_d15_0),.clk(clk),.rst(rst));            //channel 16
	large_mux #(.WIDTH(WIDTH)) large_mux_instance16151(.data_in(wire_d15_0),.data_out(wire_d15_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance16152(.data_in(wire_d15_1),.data_out(wire_d15_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance16153(.data_in(wire_d15_2),.data_out(wire_d15_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance16154(.data_in(wire_d15_3),.data_out(wire_d15_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance16155(.data_in(wire_d15_4),.data_out(wire_d15_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance16156(.data_in(wire_d15_5),.data_out(wire_d15_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance16157(.data_in(wire_d15_6),.data_out(wire_d15_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance16158(.data_in(wire_d15_7),.data_out(wire_d15_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance16159(.data_in(wire_d15_8),.data_out(wire_d15_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161510(.data_in(wire_d15_9),.data_out(wire_d15_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161511(.data_in(wire_d15_10),.data_out(wire_d15_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161512(.data_in(wire_d15_11),.data_out(wire_d15_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161513(.data_in(wire_d15_12),.data_out(wire_d15_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161514(.data_in(wire_d15_13),.data_out(wire_d15_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161515(.data_in(wire_d15_14),.data_out(wire_d15_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161516(.data_in(wire_d15_15),.data_out(wire_d15_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161517(.data_in(wire_d15_16),.data_out(wire_d15_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161518(.data_in(wire_d15_17),.data_out(wire_d15_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161519(.data_in(wire_d15_18),.data_out(wire_d15_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161520(.data_in(wire_d15_19),.data_out(wire_d15_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161521(.data_in(wire_d15_20),.data_out(wire_d15_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161522(.data_in(wire_d15_21),.data_out(wire_d15_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161523(.data_in(wire_d15_22),.data_out(wire_d15_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161524(.data_in(wire_d15_23),.data_out(wire_d15_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161525(.data_in(wire_d15_24),.data_out(wire_d15_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161526(.data_in(wire_d15_25),.data_out(wire_d15_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161527(.data_in(wire_d15_26),.data_out(wire_d15_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161528(.data_in(wire_d15_27),.data_out(wire_d15_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161529(.data_in(wire_d15_28),.data_out(wire_d15_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161530(.data_in(wire_d15_29),.data_out(wire_d15_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161531(.data_in(wire_d15_30),.data_out(wire_d15_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161532(.data_in(wire_d15_31),.data_out(wire_d15_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161533(.data_in(wire_d15_32),.data_out(wire_d15_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161534(.data_in(wire_d15_33),.data_out(wire_d15_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161535(.data_in(wire_d15_34),.data_out(wire_d15_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161536(.data_in(wire_d15_35),.data_out(wire_d15_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161537(.data_in(wire_d15_36),.data_out(wire_d15_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161538(.data_in(wire_d15_37),.data_out(wire_d15_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161539(.data_in(wire_d15_38),.data_out(wire_d15_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161540(.data_in(wire_d15_39),.data_out(wire_d15_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161541(.data_in(wire_d15_40),.data_out(wire_d15_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161542(.data_in(wire_d15_41),.data_out(wire_d15_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161543(.data_in(wire_d15_42),.data_out(wire_d15_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161544(.data_in(wire_d15_43),.data_out(wire_d15_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161545(.data_in(wire_d15_44),.data_out(wire_d15_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161546(.data_in(wire_d15_45),.data_out(wire_d15_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161547(.data_in(wire_d15_46),.data_out(wire_d15_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161548(.data_in(wire_d15_47),.data_out(wire_d15_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161549(.data_in(wire_d15_48),.data_out(wire_d15_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161550(.data_in(wire_d15_49),.data_out(wire_d15_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161551(.data_in(wire_d15_50),.data_out(wire_d15_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161552(.data_in(wire_d15_51),.data_out(wire_d15_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161553(.data_in(wire_d15_52),.data_out(wire_d15_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161554(.data_in(wire_d15_53),.data_out(wire_d15_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161555(.data_in(wire_d15_54),.data_out(wire_d15_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161556(.data_in(wire_d15_55),.data_out(wire_d15_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161557(.data_in(wire_d15_56),.data_out(wire_d15_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161558(.data_in(wire_d15_57),.data_out(wire_d15_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161559(.data_in(wire_d15_58),.data_out(wire_d15_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161560(.data_in(wire_d15_59),.data_out(wire_d15_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161561(.data_in(wire_d15_60),.data_out(wire_d15_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161562(.data_in(wire_d15_61),.data_out(wire_d15_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161563(.data_in(wire_d15_62),.data_out(wire_d15_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161564(.data_in(wire_d15_63),.data_out(wire_d15_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161565(.data_in(wire_d15_64),.data_out(wire_d15_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161566(.data_in(wire_d15_65),.data_out(wire_d15_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161567(.data_in(wire_d15_66),.data_out(wire_d15_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161568(.data_in(wire_d15_67),.data_out(wire_d15_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161569(.data_in(wire_d15_68),.data_out(d_out15),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance17160(.data_in(d_in16),.data_out(wire_d16_0),.clk(clk),.rst(rst));            //channel 17
	encoder #(.WIDTH(WIDTH)) encoder_instance17161(.data_in(wire_d16_0),.data_out(wire_d16_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance17162(.data_in(wire_d16_1),.data_out(wire_d16_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance17163(.data_in(wire_d16_2),.data_out(wire_d16_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance17164(.data_in(wire_d16_3),.data_out(wire_d16_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance17165(.data_in(wire_d16_4),.data_out(wire_d16_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance17166(.data_in(wire_d16_5),.data_out(wire_d16_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance17167(.data_in(wire_d16_6),.data_out(wire_d16_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance17168(.data_in(wire_d16_7),.data_out(wire_d16_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance17169(.data_in(wire_d16_8),.data_out(wire_d16_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171610(.data_in(wire_d16_9),.data_out(wire_d16_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171611(.data_in(wire_d16_10),.data_out(wire_d16_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171612(.data_in(wire_d16_11),.data_out(wire_d16_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171613(.data_in(wire_d16_12),.data_out(wire_d16_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171614(.data_in(wire_d16_13),.data_out(wire_d16_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171615(.data_in(wire_d16_14),.data_out(wire_d16_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171616(.data_in(wire_d16_15),.data_out(wire_d16_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171617(.data_in(wire_d16_16),.data_out(wire_d16_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171618(.data_in(wire_d16_17),.data_out(wire_d16_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171619(.data_in(wire_d16_18),.data_out(wire_d16_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171620(.data_in(wire_d16_19),.data_out(wire_d16_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171621(.data_in(wire_d16_20),.data_out(wire_d16_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171622(.data_in(wire_d16_21),.data_out(wire_d16_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171623(.data_in(wire_d16_22),.data_out(wire_d16_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171624(.data_in(wire_d16_23),.data_out(wire_d16_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171625(.data_in(wire_d16_24),.data_out(wire_d16_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171626(.data_in(wire_d16_25),.data_out(wire_d16_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171627(.data_in(wire_d16_26),.data_out(wire_d16_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171628(.data_in(wire_d16_27),.data_out(wire_d16_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171629(.data_in(wire_d16_28),.data_out(wire_d16_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171630(.data_in(wire_d16_29),.data_out(wire_d16_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171631(.data_in(wire_d16_30),.data_out(wire_d16_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171632(.data_in(wire_d16_31),.data_out(wire_d16_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171633(.data_in(wire_d16_32),.data_out(wire_d16_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171634(.data_in(wire_d16_33),.data_out(wire_d16_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171635(.data_in(wire_d16_34),.data_out(wire_d16_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171636(.data_in(wire_d16_35),.data_out(wire_d16_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171637(.data_in(wire_d16_36),.data_out(wire_d16_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171638(.data_in(wire_d16_37),.data_out(wire_d16_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171639(.data_in(wire_d16_38),.data_out(wire_d16_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171640(.data_in(wire_d16_39),.data_out(wire_d16_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171641(.data_in(wire_d16_40),.data_out(wire_d16_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171642(.data_in(wire_d16_41),.data_out(wire_d16_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171643(.data_in(wire_d16_42),.data_out(wire_d16_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171644(.data_in(wire_d16_43),.data_out(wire_d16_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171645(.data_in(wire_d16_44),.data_out(wire_d16_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171646(.data_in(wire_d16_45),.data_out(wire_d16_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171647(.data_in(wire_d16_46),.data_out(wire_d16_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171648(.data_in(wire_d16_47),.data_out(wire_d16_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171649(.data_in(wire_d16_48),.data_out(wire_d16_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171650(.data_in(wire_d16_49),.data_out(wire_d16_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171651(.data_in(wire_d16_50),.data_out(wire_d16_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171652(.data_in(wire_d16_51),.data_out(wire_d16_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171653(.data_in(wire_d16_52),.data_out(wire_d16_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171654(.data_in(wire_d16_53),.data_out(wire_d16_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171655(.data_in(wire_d16_54),.data_out(wire_d16_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171656(.data_in(wire_d16_55),.data_out(wire_d16_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171657(.data_in(wire_d16_56),.data_out(wire_d16_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171658(.data_in(wire_d16_57),.data_out(wire_d16_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171659(.data_in(wire_d16_58),.data_out(wire_d16_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171660(.data_in(wire_d16_59),.data_out(wire_d16_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171661(.data_in(wire_d16_60),.data_out(wire_d16_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171662(.data_in(wire_d16_61),.data_out(wire_d16_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171663(.data_in(wire_d16_62),.data_out(wire_d16_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171664(.data_in(wire_d16_63),.data_out(wire_d16_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171665(.data_in(wire_d16_64),.data_out(wire_d16_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171666(.data_in(wire_d16_65),.data_out(wire_d16_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171667(.data_in(wire_d16_66),.data_out(wire_d16_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171668(.data_in(wire_d16_67),.data_out(wire_d16_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171669(.data_in(wire_d16_68),.data_out(d_out16),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance18170(.data_in(d_in17),.data_out(wire_d17_0),.clk(clk),.rst(rst));            //channel 18
	register #(.WIDTH(WIDTH)) register_instance18171(.data_in(wire_d17_0),.data_out(wire_d17_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance18172(.data_in(wire_d17_1),.data_out(wire_d17_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance18173(.data_in(wire_d17_2),.data_out(wire_d17_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance18174(.data_in(wire_d17_3),.data_out(wire_d17_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance18175(.data_in(wire_d17_4),.data_out(wire_d17_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance18176(.data_in(wire_d17_5),.data_out(wire_d17_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance18177(.data_in(wire_d17_6),.data_out(wire_d17_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance18178(.data_in(wire_d17_7),.data_out(wire_d17_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance18179(.data_in(wire_d17_8),.data_out(wire_d17_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181710(.data_in(wire_d17_9),.data_out(wire_d17_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181711(.data_in(wire_d17_10),.data_out(wire_d17_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181712(.data_in(wire_d17_11),.data_out(wire_d17_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181713(.data_in(wire_d17_12),.data_out(wire_d17_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181714(.data_in(wire_d17_13),.data_out(wire_d17_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181715(.data_in(wire_d17_14),.data_out(wire_d17_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181716(.data_in(wire_d17_15),.data_out(wire_d17_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181717(.data_in(wire_d17_16),.data_out(wire_d17_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181718(.data_in(wire_d17_17),.data_out(wire_d17_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181719(.data_in(wire_d17_18),.data_out(wire_d17_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181720(.data_in(wire_d17_19),.data_out(wire_d17_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181721(.data_in(wire_d17_20),.data_out(wire_d17_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181722(.data_in(wire_d17_21),.data_out(wire_d17_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181723(.data_in(wire_d17_22),.data_out(wire_d17_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181724(.data_in(wire_d17_23),.data_out(wire_d17_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181725(.data_in(wire_d17_24),.data_out(wire_d17_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181726(.data_in(wire_d17_25),.data_out(wire_d17_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181727(.data_in(wire_d17_26),.data_out(wire_d17_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181728(.data_in(wire_d17_27),.data_out(wire_d17_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181729(.data_in(wire_d17_28),.data_out(wire_d17_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181730(.data_in(wire_d17_29),.data_out(wire_d17_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181731(.data_in(wire_d17_30),.data_out(wire_d17_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181732(.data_in(wire_d17_31),.data_out(wire_d17_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181733(.data_in(wire_d17_32),.data_out(wire_d17_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181734(.data_in(wire_d17_33),.data_out(wire_d17_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181735(.data_in(wire_d17_34),.data_out(wire_d17_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181736(.data_in(wire_d17_35),.data_out(wire_d17_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181737(.data_in(wire_d17_36),.data_out(wire_d17_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181738(.data_in(wire_d17_37),.data_out(wire_d17_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181739(.data_in(wire_d17_38),.data_out(wire_d17_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181740(.data_in(wire_d17_39),.data_out(wire_d17_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181741(.data_in(wire_d17_40),.data_out(wire_d17_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181742(.data_in(wire_d17_41),.data_out(wire_d17_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181743(.data_in(wire_d17_42),.data_out(wire_d17_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181744(.data_in(wire_d17_43),.data_out(wire_d17_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181745(.data_in(wire_d17_44),.data_out(wire_d17_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181746(.data_in(wire_d17_45),.data_out(wire_d17_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181747(.data_in(wire_d17_46),.data_out(wire_d17_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181748(.data_in(wire_d17_47),.data_out(wire_d17_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181749(.data_in(wire_d17_48),.data_out(wire_d17_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181750(.data_in(wire_d17_49),.data_out(wire_d17_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181751(.data_in(wire_d17_50),.data_out(wire_d17_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181752(.data_in(wire_d17_51),.data_out(wire_d17_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181753(.data_in(wire_d17_52),.data_out(wire_d17_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181754(.data_in(wire_d17_53),.data_out(wire_d17_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181755(.data_in(wire_d17_54),.data_out(wire_d17_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181756(.data_in(wire_d17_55),.data_out(wire_d17_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181757(.data_in(wire_d17_56),.data_out(wire_d17_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181758(.data_in(wire_d17_57),.data_out(wire_d17_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181759(.data_in(wire_d17_58),.data_out(wire_d17_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181760(.data_in(wire_d17_59),.data_out(wire_d17_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181761(.data_in(wire_d17_60),.data_out(wire_d17_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181762(.data_in(wire_d17_61),.data_out(wire_d17_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181763(.data_in(wire_d17_62),.data_out(wire_d17_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181764(.data_in(wire_d17_63),.data_out(wire_d17_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181765(.data_in(wire_d17_64),.data_out(wire_d17_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181766(.data_in(wire_d17_65),.data_out(wire_d17_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181767(.data_in(wire_d17_66),.data_out(wire_d17_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181768(.data_in(wire_d17_67),.data_out(wire_d17_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181769(.data_in(wire_d17_68),.data_out(d_out17),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance19180(.data_in(d_in18),.data_out(wire_d18_0),.clk(clk),.rst(rst));            //channel 19
	encoder #(.WIDTH(WIDTH)) encoder_instance19181(.data_in(wire_d18_0),.data_out(wire_d18_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance19182(.data_in(wire_d18_1),.data_out(wire_d18_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance19183(.data_in(wire_d18_2),.data_out(wire_d18_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance19184(.data_in(wire_d18_3),.data_out(wire_d18_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance19185(.data_in(wire_d18_4),.data_out(wire_d18_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance19186(.data_in(wire_d18_5),.data_out(wire_d18_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance19187(.data_in(wire_d18_6),.data_out(wire_d18_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance19188(.data_in(wire_d18_7),.data_out(wire_d18_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance19189(.data_in(wire_d18_8),.data_out(wire_d18_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191810(.data_in(wire_d18_9),.data_out(wire_d18_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191811(.data_in(wire_d18_10),.data_out(wire_d18_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191812(.data_in(wire_d18_11),.data_out(wire_d18_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191813(.data_in(wire_d18_12),.data_out(wire_d18_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191814(.data_in(wire_d18_13),.data_out(wire_d18_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191815(.data_in(wire_d18_14),.data_out(wire_d18_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191816(.data_in(wire_d18_15),.data_out(wire_d18_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191817(.data_in(wire_d18_16),.data_out(wire_d18_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191818(.data_in(wire_d18_17),.data_out(wire_d18_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191819(.data_in(wire_d18_18),.data_out(wire_d18_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191820(.data_in(wire_d18_19),.data_out(wire_d18_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191821(.data_in(wire_d18_20),.data_out(wire_d18_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191822(.data_in(wire_d18_21),.data_out(wire_d18_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191823(.data_in(wire_d18_22),.data_out(wire_d18_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191824(.data_in(wire_d18_23),.data_out(wire_d18_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191825(.data_in(wire_d18_24),.data_out(wire_d18_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191826(.data_in(wire_d18_25),.data_out(wire_d18_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191827(.data_in(wire_d18_26),.data_out(wire_d18_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191828(.data_in(wire_d18_27),.data_out(wire_d18_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191829(.data_in(wire_d18_28),.data_out(wire_d18_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191830(.data_in(wire_d18_29),.data_out(wire_d18_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191831(.data_in(wire_d18_30),.data_out(wire_d18_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191832(.data_in(wire_d18_31),.data_out(wire_d18_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191833(.data_in(wire_d18_32),.data_out(wire_d18_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191834(.data_in(wire_d18_33),.data_out(wire_d18_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191835(.data_in(wire_d18_34),.data_out(wire_d18_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191836(.data_in(wire_d18_35),.data_out(wire_d18_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191837(.data_in(wire_d18_36),.data_out(wire_d18_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191838(.data_in(wire_d18_37),.data_out(wire_d18_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191839(.data_in(wire_d18_38),.data_out(wire_d18_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191840(.data_in(wire_d18_39),.data_out(wire_d18_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191841(.data_in(wire_d18_40),.data_out(wire_d18_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191842(.data_in(wire_d18_41),.data_out(wire_d18_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191843(.data_in(wire_d18_42),.data_out(wire_d18_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191844(.data_in(wire_d18_43),.data_out(wire_d18_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191845(.data_in(wire_d18_44),.data_out(wire_d18_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191846(.data_in(wire_d18_45),.data_out(wire_d18_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191847(.data_in(wire_d18_46),.data_out(wire_d18_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191848(.data_in(wire_d18_47),.data_out(wire_d18_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191849(.data_in(wire_d18_48),.data_out(wire_d18_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191850(.data_in(wire_d18_49),.data_out(wire_d18_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191851(.data_in(wire_d18_50),.data_out(wire_d18_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191852(.data_in(wire_d18_51),.data_out(wire_d18_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191853(.data_in(wire_d18_52),.data_out(wire_d18_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191854(.data_in(wire_d18_53),.data_out(wire_d18_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191855(.data_in(wire_d18_54),.data_out(wire_d18_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191856(.data_in(wire_d18_55),.data_out(wire_d18_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191857(.data_in(wire_d18_56),.data_out(wire_d18_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191858(.data_in(wire_d18_57),.data_out(wire_d18_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191859(.data_in(wire_d18_58),.data_out(wire_d18_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191860(.data_in(wire_d18_59),.data_out(wire_d18_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191861(.data_in(wire_d18_60),.data_out(wire_d18_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191862(.data_in(wire_d18_61),.data_out(wire_d18_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191863(.data_in(wire_d18_62),.data_out(wire_d18_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191864(.data_in(wire_d18_63),.data_out(wire_d18_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191865(.data_in(wire_d18_64),.data_out(wire_d18_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191866(.data_in(wire_d18_65),.data_out(wire_d18_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191867(.data_in(wire_d18_66),.data_out(wire_d18_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191868(.data_in(wire_d18_67),.data_out(wire_d18_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191869(.data_in(wire_d18_68),.data_out(d_out18),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance20190(.data_in(d_in19),.data_out(wire_d19_0),.clk(clk),.rst(rst));            //channel 20
	large_mux #(.WIDTH(WIDTH)) large_mux_instance20191(.data_in(wire_d19_0),.data_out(wire_d19_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance20192(.data_in(wire_d19_1),.data_out(wire_d19_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance20193(.data_in(wire_d19_2),.data_out(wire_d19_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance20194(.data_in(wire_d19_3),.data_out(wire_d19_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance20195(.data_in(wire_d19_4),.data_out(wire_d19_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance20196(.data_in(wire_d19_5),.data_out(wire_d19_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance20197(.data_in(wire_d19_6),.data_out(wire_d19_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance20198(.data_in(wire_d19_7),.data_out(wire_d19_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance20199(.data_in(wire_d19_8),.data_out(wire_d19_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201910(.data_in(wire_d19_9),.data_out(wire_d19_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201911(.data_in(wire_d19_10),.data_out(wire_d19_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201912(.data_in(wire_d19_11),.data_out(wire_d19_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201913(.data_in(wire_d19_12),.data_out(wire_d19_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201914(.data_in(wire_d19_13),.data_out(wire_d19_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201915(.data_in(wire_d19_14),.data_out(wire_d19_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201916(.data_in(wire_d19_15),.data_out(wire_d19_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201917(.data_in(wire_d19_16),.data_out(wire_d19_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201918(.data_in(wire_d19_17),.data_out(wire_d19_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201919(.data_in(wire_d19_18),.data_out(wire_d19_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201920(.data_in(wire_d19_19),.data_out(wire_d19_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201921(.data_in(wire_d19_20),.data_out(wire_d19_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201922(.data_in(wire_d19_21),.data_out(wire_d19_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201923(.data_in(wire_d19_22),.data_out(wire_d19_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201924(.data_in(wire_d19_23),.data_out(wire_d19_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201925(.data_in(wire_d19_24),.data_out(wire_d19_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201926(.data_in(wire_d19_25),.data_out(wire_d19_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201927(.data_in(wire_d19_26),.data_out(wire_d19_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201928(.data_in(wire_d19_27),.data_out(wire_d19_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201929(.data_in(wire_d19_28),.data_out(wire_d19_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201930(.data_in(wire_d19_29),.data_out(wire_d19_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201931(.data_in(wire_d19_30),.data_out(wire_d19_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201932(.data_in(wire_d19_31),.data_out(wire_d19_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201933(.data_in(wire_d19_32),.data_out(wire_d19_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201934(.data_in(wire_d19_33),.data_out(wire_d19_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201935(.data_in(wire_d19_34),.data_out(wire_d19_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201936(.data_in(wire_d19_35),.data_out(wire_d19_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201937(.data_in(wire_d19_36),.data_out(wire_d19_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201938(.data_in(wire_d19_37),.data_out(wire_d19_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201939(.data_in(wire_d19_38),.data_out(wire_d19_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201940(.data_in(wire_d19_39),.data_out(wire_d19_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201941(.data_in(wire_d19_40),.data_out(wire_d19_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201942(.data_in(wire_d19_41),.data_out(wire_d19_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201943(.data_in(wire_d19_42),.data_out(wire_d19_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201944(.data_in(wire_d19_43),.data_out(wire_d19_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201945(.data_in(wire_d19_44),.data_out(wire_d19_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201946(.data_in(wire_d19_45),.data_out(wire_d19_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201947(.data_in(wire_d19_46),.data_out(wire_d19_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201948(.data_in(wire_d19_47),.data_out(wire_d19_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201949(.data_in(wire_d19_48),.data_out(wire_d19_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201950(.data_in(wire_d19_49),.data_out(wire_d19_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201951(.data_in(wire_d19_50),.data_out(wire_d19_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201952(.data_in(wire_d19_51),.data_out(wire_d19_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201953(.data_in(wire_d19_52),.data_out(wire_d19_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201954(.data_in(wire_d19_53),.data_out(wire_d19_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201955(.data_in(wire_d19_54),.data_out(wire_d19_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201956(.data_in(wire_d19_55),.data_out(wire_d19_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201957(.data_in(wire_d19_56),.data_out(wire_d19_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201958(.data_in(wire_d19_57),.data_out(wire_d19_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201959(.data_in(wire_d19_58),.data_out(wire_d19_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201960(.data_in(wire_d19_59),.data_out(wire_d19_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201961(.data_in(wire_d19_60),.data_out(wire_d19_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201962(.data_in(wire_d19_61),.data_out(wire_d19_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201963(.data_in(wire_d19_62),.data_out(wire_d19_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201964(.data_in(wire_d19_63),.data_out(wire_d19_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201965(.data_in(wire_d19_64),.data_out(wire_d19_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201966(.data_in(wire_d19_65),.data_out(wire_d19_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201967(.data_in(wire_d19_66),.data_out(wire_d19_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201968(.data_in(wire_d19_67),.data_out(wire_d19_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201969(.data_in(wire_d19_68),.data_out(d_out19),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance21200(.data_in(d_in20),.data_out(wire_d20_0),.clk(clk),.rst(rst));            //channel 21
	register #(.WIDTH(WIDTH)) register_instance21201(.data_in(wire_d20_0),.data_out(wire_d20_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance21202(.data_in(wire_d20_1),.data_out(wire_d20_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance21203(.data_in(wire_d20_2),.data_out(wire_d20_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21204(.data_in(wire_d20_3),.data_out(wire_d20_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance21205(.data_in(wire_d20_4),.data_out(wire_d20_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21206(.data_in(wire_d20_5),.data_out(wire_d20_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance21207(.data_in(wire_d20_6),.data_out(wire_d20_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance21208(.data_in(wire_d20_7),.data_out(wire_d20_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21209(.data_in(wire_d20_8),.data_out(wire_d20_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212010(.data_in(wire_d20_9),.data_out(wire_d20_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212011(.data_in(wire_d20_10),.data_out(wire_d20_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212012(.data_in(wire_d20_11),.data_out(wire_d20_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212013(.data_in(wire_d20_12),.data_out(wire_d20_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212014(.data_in(wire_d20_13),.data_out(wire_d20_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212015(.data_in(wire_d20_14),.data_out(wire_d20_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212016(.data_in(wire_d20_15),.data_out(wire_d20_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212017(.data_in(wire_d20_16),.data_out(wire_d20_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212018(.data_in(wire_d20_17),.data_out(wire_d20_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212019(.data_in(wire_d20_18),.data_out(wire_d20_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212020(.data_in(wire_d20_19),.data_out(wire_d20_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212021(.data_in(wire_d20_20),.data_out(wire_d20_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212022(.data_in(wire_d20_21),.data_out(wire_d20_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212023(.data_in(wire_d20_22),.data_out(wire_d20_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212024(.data_in(wire_d20_23),.data_out(wire_d20_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212025(.data_in(wire_d20_24),.data_out(wire_d20_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212026(.data_in(wire_d20_25),.data_out(wire_d20_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212027(.data_in(wire_d20_26),.data_out(wire_d20_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212028(.data_in(wire_d20_27),.data_out(wire_d20_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212029(.data_in(wire_d20_28),.data_out(wire_d20_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212030(.data_in(wire_d20_29),.data_out(wire_d20_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212031(.data_in(wire_d20_30),.data_out(wire_d20_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212032(.data_in(wire_d20_31),.data_out(wire_d20_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212033(.data_in(wire_d20_32),.data_out(wire_d20_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212034(.data_in(wire_d20_33),.data_out(wire_d20_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212035(.data_in(wire_d20_34),.data_out(wire_d20_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212036(.data_in(wire_d20_35),.data_out(wire_d20_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212037(.data_in(wire_d20_36),.data_out(wire_d20_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212038(.data_in(wire_d20_37),.data_out(wire_d20_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212039(.data_in(wire_d20_38),.data_out(wire_d20_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212040(.data_in(wire_d20_39),.data_out(wire_d20_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212041(.data_in(wire_d20_40),.data_out(wire_d20_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212042(.data_in(wire_d20_41),.data_out(wire_d20_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212043(.data_in(wire_d20_42),.data_out(wire_d20_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212044(.data_in(wire_d20_43),.data_out(wire_d20_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212045(.data_in(wire_d20_44),.data_out(wire_d20_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212046(.data_in(wire_d20_45),.data_out(wire_d20_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212047(.data_in(wire_d20_46),.data_out(wire_d20_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212048(.data_in(wire_d20_47),.data_out(wire_d20_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212049(.data_in(wire_d20_48),.data_out(wire_d20_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212050(.data_in(wire_d20_49),.data_out(wire_d20_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212051(.data_in(wire_d20_50),.data_out(wire_d20_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212052(.data_in(wire_d20_51),.data_out(wire_d20_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212053(.data_in(wire_d20_52),.data_out(wire_d20_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212054(.data_in(wire_d20_53),.data_out(wire_d20_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212055(.data_in(wire_d20_54),.data_out(wire_d20_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212056(.data_in(wire_d20_55),.data_out(wire_d20_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212057(.data_in(wire_d20_56),.data_out(wire_d20_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212058(.data_in(wire_d20_57),.data_out(wire_d20_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212059(.data_in(wire_d20_58),.data_out(wire_d20_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212060(.data_in(wire_d20_59),.data_out(wire_d20_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212061(.data_in(wire_d20_60),.data_out(wire_d20_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212062(.data_in(wire_d20_61),.data_out(wire_d20_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212063(.data_in(wire_d20_62),.data_out(wire_d20_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212064(.data_in(wire_d20_63),.data_out(wire_d20_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212065(.data_in(wire_d20_64),.data_out(wire_d20_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212066(.data_in(wire_d20_65),.data_out(wire_d20_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212067(.data_in(wire_d20_66),.data_out(wire_d20_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212068(.data_in(wire_d20_67),.data_out(wire_d20_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212069(.data_in(wire_d20_68),.data_out(d_out20),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance22210(.data_in(d_in21),.data_out(wire_d21_0),.clk(clk),.rst(rst));            //channel 22
	encoder #(.WIDTH(WIDTH)) encoder_instance22211(.data_in(wire_d21_0),.data_out(wire_d21_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance22212(.data_in(wire_d21_1),.data_out(wire_d21_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance22213(.data_in(wire_d21_2),.data_out(wire_d21_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance22214(.data_in(wire_d21_3),.data_out(wire_d21_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance22215(.data_in(wire_d21_4),.data_out(wire_d21_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance22216(.data_in(wire_d21_5),.data_out(wire_d21_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance22217(.data_in(wire_d21_6),.data_out(wire_d21_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance22218(.data_in(wire_d21_7),.data_out(wire_d21_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance22219(.data_in(wire_d21_8),.data_out(wire_d21_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222110(.data_in(wire_d21_9),.data_out(wire_d21_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222111(.data_in(wire_d21_10),.data_out(wire_d21_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222112(.data_in(wire_d21_11),.data_out(wire_d21_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222113(.data_in(wire_d21_12),.data_out(wire_d21_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222114(.data_in(wire_d21_13),.data_out(wire_d21_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222115(.data_in(wire_d21_14),.data_out(wire_d21_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222116(.data_in(wire_d21_15),.data_out(wire_d21_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222117(.data_in(wire_d21_16),.data_out(wire_d21_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222118(.data_in(wire_d21_17),.data_out(wire_d21_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222119(.data_in(wire_d21_18),.data_out(wire_d21_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222120(.data_in(wire_d21_19),.data_out(wire_d21_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222121(.data_in(wire_d21_20),.data_out(wire_d21_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222122(.data_in(wire_d21_21),.data_out(wire_d21_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222123(.data_in(wire_d21_22),.data_out(wire_d21_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222124(.data_in(wire_d21_23),.data_out(wire_d21_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222125(.data_in(wire_d21_24),.data_out(wire_d21_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222126(.data_in(wire_d21_25),.data_out(wire_d21_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222127(.data_in(wire_d21_26),.data_out(wire_d21_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222128(.data_in(wire_d21_27),.data_out(wire_d21_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222129(.data_in(wire_d21_28),.data_out(wire_d21_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222130(.data_in(wire_d21_29),.data_out(wire_d21_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222131(.data_in(wire_d21_30),.data_out(wire_d21_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222132(.data_in(wire_d21_31),.data_out(wire_d21_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222133(.data_in(wire_d21_32),.data_out(wire_d21_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222134(.data_in(wire_d21_33),.data_out(wire_d21_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222135(.data_in(wire_d21_34),.data_out(wire_d21_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222136(.data_in(wire_d21_35),.data_out(wire_d21_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222137(.data_in(wire_d21_36),.data_out(wire_d21_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222138(.data_in(wire_d21_37),.data_out(wire_d21_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222139(.data_in(wire_d21_38),.data_out(wire_d21_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222140(.data_in(wire_d21_39),.data_out(wire_d21_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222141(.data_in(wire_d21_40),.data_out(wire_d21_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222142(.data_in(wire_d21_41),.data_out(wire_d21_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222143(.data_in(wire_d21_42),.data_out(wire_d21_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222144(.data_in(wire_d21_43),.data_out(wire_d21_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222145(.data_in(wire_d21_44),.data_out(wire_d21_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222146(.data_in(wire_d21_45),.data_out(wire_d21_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222147(.data_in(wire_d21_46),.data_out(wire_d21_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222148(.data_in(wire_d21_47),.data_out(wire_d21_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222149(.data_in(wire_d21_48),.data_out(wire_d21_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222150(.data_in(wire_d21_49),.data_out(wire_d21_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222151(.data_in(wire_d21_50),.data_out(wire_d21_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222152(.data_in(wire_d21_51),.data_out(wire_d21_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222153(.data_in(wire_d21_52),.data_out(wire_d21_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222154(.data_in(wire_d21_53),.data_out(wire_d21_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222155(.data_in(wire_d21_54),.data_out(wire_d21_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222156(.data_in(wire_d21_55),.data_out(wire_d21_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222157(.data_in(wire_d21_56),.data_out(wire_d21_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222158(.data_in(wire_d21_57),.data_out(wire_d21_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222159(.data_in(wire_d21_58),.data_out(wire_d21_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222160(.data_in(wire_d21_59),.data_out(wire_d21_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222161(.data_in(wire_d21_60),.data_out(wire_d21_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222162(.data_in(wire_d21_61),.data_out(wire_d21_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222163(.data_in(wire_d21_62),.data_out(wire_d21_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222164(.data_in(wire_d21_63),.data_out(wire_d21_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222165(.data_in(wire_d21_64),.data_out(wire_d21_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222166(.data_in(wire_d21_65),.data_out(wire_d21_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222167(.data_in(wire_d21_66),.data_out(wire_d21_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222168(.data_in(wire_d21_67),.data_out(wire_d21_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222169(.data_in(wire_d21_68),.data_out(d_out21),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance23220(.data_in(d_in22),.data_out(wire_d22_0),.clk(clk),.rst(rst));            //channel 23
	large_mux #(.WIDTH(WIDTH)) large_mux_instance23221(.data_in(wire_d22_0),.data_out(wire_d22_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance23222(.data_in(wire_d22_1),.data_out(wire_d22_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance23223(.data_in(wire_d22_2),.data_out(wire_d22_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance23224(.data_in(wire_d22_3),.data_out(wire_d22_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance23225(.data_in(wire_d22_4),.data_out(wire_d22_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance23226(.data_in(wire_d22_5),.data_out(wire_d22_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance23227(.data_in(wire_d22_6),.data_out(wire_d22_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance23228(.data_in(wire_d22_7),.data_out(wire_d22_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance23229(.data_in(wire_d22_8),.data_out(wire_d22_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232210(.data_in(wire_d22_9),.data_out(wire_d22_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232211(.data_in(wire_d22_10),.data_out(wire_d22_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232212(.data_in(wire_d22_11),.data_out(wire_d22_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232213(.data_in(wire_d22_12),.data_out(wire_d22_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232214(.data_in(wire_d22_13),.data_out(wire_d22_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232215(.data_in(wire_d22_14),.data_out(wire_d22_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232216(.data_in(wire_d22_15),.data_out(wire_d22_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232217(.data_in(wire_d22_16),.data_out(wire_d22_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232218(.data_in(wire_d22_17),.data_out(wire_d22_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232219(.data_in(wire_d22_18),.data_out(wire_d22_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232220(.data_in(wire_d22_19),.data_out(wire_d22_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232221(.data_in(wire_d22_20),.data_out(wire_d22_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232222(.data_in(wire_d22_21),.data_out(wire_d22_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232223(.data_in(wire_d22_22),.data_out(wire_d22_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232224(.data_in(wire_d22_23),.data_out(wire_d22_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232225(.data_in(wire_d22_24),.data_out(wire_d22_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232226(.data_in(wire_d22_25),.data_out(wire_d22_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232227(.data_in(wire_d22_26),.data_out(wire_d22_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232228(.data_in(wire_d22_27),.data_out(wire_d22_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232229(.data_in(wire_d22_28),.data_out(wire_d22_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232230(.data_in(wire_d22_29),.data_out(wire_d22_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232231(.data_in(wire_d22_30),.data_out(wire_d22_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232232(.data_in(wire_d22_31),.data_out(wire_d22_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232233(.data_in(wire_d22_32),.data_out(wire_d22_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232234(.data_in(wire_d22_33),.data_out(wire_d22_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232235(.data_in(wire_d22_34),.data_out(wire_d22_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232236(.data_in(wire_d22_35),.data_out(wire_d22_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232237(.data_in(wire_d22_36),.data_out(wire_d22_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232238(.data_in(wire_d22_37),.data_out(wire_d22_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232239(.data_in(wire_d22_38),.data_out(wire_d22_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232240(.data_in(wire_d22_39),.data_out(wire_d22_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232241(.data_in(wire_d22_40),.data_out(wire_d22_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232242(.data_in(wire_d22_41),.data_out(wire_d22_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232243(.data_in(wire_d22_42),.data_out(wire_d22_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232244(.data_in(wire_d22_43),.data_out(wire_d22_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232245(.data_in(wire_d22_44),.data_out(wire_d22_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232246(.data_in(wire_d22_45),.data_out(wire_d22_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232247(.data_in(wire_d22_46),.data_out(wire_d22_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232248(.data_in(wire_d22_47),.data_out(wire_d22_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232249(.data_in(wire_d22_48),.data_out(wire_d22_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232250(.data_in(wire_d22_49),.data_out(wire_d22_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232251(.data_in(wire_d22_50),.data_out(wire_d22_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232252(.data_in(wire_d22_51),.data_out(wire_d22_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232253(.data_in(wire_d22_52),.data_out(wire_d22_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232254(.data_in(wire_d22_53),.data_out(wire_d22_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232255(.data_in(wire_d22_54),.data_out(wire_d22_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232256(.data_in(wire_d22_55),.data_out(wire_d22_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232257(.data_in(wire_d22_56),.data_out(wire_d22_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232258(.data_in(wire_d22_57),.data_out(wire_d22_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232259(.data_in(wire_d22_58),.data_out(wire_d22_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232260(.data_in(wire_d22_59),.data_out(wire_d22_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232261(.data_in(wire_d22_60),.data_out(wire_d22_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232262(.data_in(wire_d22_61),.data_out(wire_d22_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232263(.data_in(wire_d22_62),.data_out(wire_d22_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232264(.data_in(wire_d22_63),.data_out(wire_d22_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232265(.data_in(wire_d22_64),.data_out(wire_d22_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232266(.data_in(wire_d22_65),.data_out(wire_d22_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232267(.data_in(wire_d22_66),.data_out(wire_d22_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232268(.data_in(wire_d22_67),.data_out(wire_d22_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232269(.data_in(wire_d22_68),.data_out(d_out22),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance24230(.data_in(d_in23),.data_out(wire_d23_0),.clk(clk),.rst(rst));            //channel 24
	large_mux #(.WIDTH(WIDTH)) large_mux_instance24231(.data_in(wire_d23_0),.data_out(wire_d23_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance24232(.data_in(wire_d23_1),.data_out(wire_d23_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance24233(.data_in(wire_d23_2),.data_out(wire_d23_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance24234(.data_in(wire_d23_3),.data_out(wire_d23_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance24235(.data_in(wire_d23_4),.data_out(wire_d23_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance24236(.data_in(wire_d23_5),.data_out(wire_d23_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance24237(.data_in(wire_d23_6),.data_out(wire_d23_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance24238(.data_in(wire_d23_7),.data_out(wire_d23_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance24239(.data_in(wire_d23_8),.data_out(wire_d23_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242310(.data_in(wire_d23_9),.data_out(wire_d23_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242311(.data_in(wire_d23_10),.data_out(wire_d23_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242312(.data_in(wire_d23_11),.data_out(wire_d23_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242313(.data_in(wire_d23_12),.data_out(wire_d23_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242314(.data_in(wire_d23_13),.data_out(wire_d23_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242315(.data_in(wire_d23_14),.data_out(wire_d23_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242316(.data_in(wire_d23_15),.data_out(wire_d23_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242317(.data_in(wire_d23_16),.data_out(wire_d23_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242318(.data_in(wire_d23_17),.data_out(wire_d23_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242319(.data_in(wire_d23_18),.data_out(wire_d23_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242320(.data_in(wire_d23_19),.data_out(wire_d23_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242321(.data_in(wire_d23_20),.data_out(wire_d23_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242322(.data_in(wire_d23_21),.data_out(wire_d23_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242323(.data_in(wire_d23_22),.data_out(wire_d23_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242324(.data_in(wire_d23_23),.data_out(wire_d23_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242325(.data_in(wire_d23_24),.data_out(wire_d23_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242326(.data_in(wire_d23_25),.data_out(wire_d23_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242327(.data_in(wire_d23_26),.data_out(wire_d23_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242328(.data_in(wire_d23_27),.data_out(wire_d23_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242329(.data_in(wire_d23_28),.data_out(wire_d23_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242330(.data_in(wire_d23_29),.data_out(wire_d23_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242331(.data_in(wire_d23_30),.data_out(wire_d23_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242332(.data_in(wire_d23_31),.data_out(wire_d23_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242333(.data_in(wire_d23_32),.data_out(wire_d23_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242334(.data_in(wire_d23_33),.data_out(wire_d23_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242335(.data_in(wire_d23_34),.data_out(wire_d23_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242336(.data_in(wire_d23_35),.data_out(wire_d23_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242337(.data_in(wire_d23_36),.data_out(wire_d23_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242338(.data_in(wire_d23_37),.data_out(wire_d23_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242339(.data_in(wire_d23_38),.data_out(wire_d23_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242340(.data_in(wire_d23_39),.data_out(wire_d23_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242341(.data_in(wire_d23_40),.data_out(wire_d23_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242342(.data_in(wire_d23_41),.data_out(wire_d23_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242343(.data_in(wire_d23_42),.data_out(wire_d23_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242344(.data_in(wire_d23_43),.data_out(wire_d23_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242345(.data_in(wire_d23_44),.data_out(wire_d23_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242346(.data_in(wire_d23_45),.data_out(wire_d23_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242347(.data_in(wire_d23_46),.data_out(wire_d23_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242348(.data_in(wire_d23_47),.data_out(wire_d23_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242349(.data_in(wire_d23_48),.data_out(wire_d23_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242350(.data_in(wire_d23_49),.data_out(wire_d23_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242351(.data_in(wire_d23_50),.data_out(wire_d23_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242352(.data_in(wire_d23_51),.data_out(wire_d23_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242353(.data_in(wire_d23_52),.data_out(wire_d23_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242354(.data_in(wire_d23_53),.data_out(wire_d23_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242355(.data_in(wire_d23_54),.data_out(wire_d23_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242356(.data_in(wire_d23_55),.data_out(wire_d23_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242357(.data_in(wire_d23_56),.data_out(wire_d23_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242358(.data_in(wire_d23_57),.data_out(wire_d23_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242359(.data_in(wire_d23_58),.data_out(wire_d23_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242360(.data_in(wire_d23_59),.data_out(wire_d23_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242361(.data_in(wire_d23_60),.data_out(wire_d23_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242362(.data_in(wire_d23_61),.data_out(wire_d23_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242363(.data_in(wire_d23_62),.data_out(wire_d23_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242364(.data_in(wire_d23_63),.data_out(wire_d23_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242365(.data_in(wire_d23_64),.data_out(wire_d23_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242366(.data_in(wire_d23_65),.data_out(wire_d23_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242367(.data_in(wire_d23_66),.data_out(wire_d23_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242368(.data_in(wire_d23_67),.data_out(wire_d23_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242369(.data_in(wire_d23_68),.data_out(d_out23),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance25240(.data_in(d_in24),.data_out(wire_d24_0),.clk(clk),.rst(rst));            //channel 25
	encoder #(.WIDTH(WIDTH)) encoder_instance25241(.data_in(wire_d24_0),.data_out(wire_d24_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance25242(.data_in(wire_d24_1),.data_out(wire_d24_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance25243(.data_in(wire_d24_2),.data_out(wire_d24_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance25244(.data_in(wire_d24_3),.data_out(wire_d24_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance25245(.data_in(wire_d24_4),.data_out(wire_d24_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance25246(.data_in(wire_d24_5),.data_out(wire_d24_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance25247(.data_in(wire_d24_6),.data_out(wire_d24_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance25248(.data_in(wire_d24_7),.data_out(wire_d24_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance25249(.data_in(wire_d24_8),.data_out(wire_d24_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252410(.data_in(wire_d24_9),.data_out(wire_d24_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252411(.data_in(wire_d24_10),.data_out(wire_d24_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252412(.data_in(wire_d24_11),.data_out(wire_d24_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252413(.data_in(wire_d24_12),.data_out(wire_d24_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252414(.data_in(wire_d24_13),.data_out(wire_d24_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252415(.data_in(wire_d24_14),.data_out(wire_d24_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252416(.data_in(wire_d24_15),.data_out(wire_d24_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252417(.data_in(wire_d24_16),.data_out(wire_d24_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252418(.data_in(wire_d24_17),.data_out(wire_d24_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252419(.data_in(wire_d24_18),.data_out(wire_d24_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252420(.data_in(wire_d24_19),.data_out(wire_d24_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252421(.data_in(wire_d24_20),.data_out(wire_d24_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252422(.data_in(wire_d24_21),.data_out(wire_d24_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252423(.data_in(wire_d24_22),.data_out(wire_d24_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252424(.data_in(wire_d24_23),.data_out(wire_d24_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252425(.data_in(wire_d24_24),.data_out(wire_d24_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252426(.data_in(wire_d24_25),.data_out(wire_d24_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252427(.data_in(wire_d24_26),.data_out(wire_d24_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252428(.data_in(wire_d24_27),.data_out(wire_d24_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252429(.data_in(wire_d24_28),.data_out(wire_d24_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252430(.data_in(wire_d24_29),.data_out(wire_d24_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252431(.data_in(wire_d24_30),.data_out(wire_d24_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252432(.data_in(wire_d24_31),.data_out(wire_d24_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252433(.data_in(wire_d24_32),.data_out(wire_d24_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252434(.data_in(wire_d24_33),.data_out(wire_d24_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252435(.data_in(wire_d24_34),.data_out(wire_d24_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252436(.data_in(wire_d24_35),.data_out(wire_d24_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252437(.data_in(wire_d24_36),.data_out(wire_d24_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252438(.data_in(wire_d24_37),.data_out(wire_d24_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252439(.data_in(wire_d24_38),.data_out(wire_d24_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252440(.data_in(wire_d24_39),.data_out(wire_d24_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252441(.data_in(wire_d24_40),.data_out(wire_d24_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252442(.data_in(wire_d24_41),.data_out(wire_d24_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252443(.data_in(wire_d24_42),.data_out(wire_d24_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252444(.data_in(wire_d24_43),.data_out(wire_d24_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252445(.data_in(wire_d24_44),.data_out(wire_d24_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252446(.data_in(wire_d24_45),.data_out(wire_d24_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252447(.data_in(wire_d24_46),.data_out(wire_d24_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252448(.data_in(wire_d24_47),.data_out(wire_d24_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252449(.data_in(wire_d24_48),.data_out(wire_d24_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252450(.data_in(wire_d24_49),.data_out(wire_d24_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252451(.data_in(wire_d24_50),.data_out(wire_d24_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252452(.data_in(wire_d24_51),.data_out(wire_d24_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252453(.data_in(wire_d24_52),.data_out(wire_d24_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252454(.data_in(wire_d24_53),.data_out(wire_d24_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252455(.data_in(wire_d24_54),.data_out(wire_d24_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252456(.data_in(wire_d24_55),.data_out(wire_d24_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252457(.data_in(wire_d24_56),.data_out(wire_d24_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252458(.data_in(wire_d24_57),.data_out(wire_d24_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252459(.data_in(wire_d24_58),.data_out(wire_d24_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252460(.data_in(wire_d24_59),.data_out(wire_d24_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252461(.data_in(wire_d24_60),.data_out(wire_d24_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252462(.data_in(wire_d24_61),.data_out(wire_d24_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252463(.data_in(wire_d24_62),.data_out(wire_d24_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252464(.data_in(wire_d24_63),.data_out(wire_d24_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252465(.data_in(wire_d24_64),.data_out(wire_d24_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252466(.data_in(wire_d24_65),.data_out(wire_d24_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252467(.data_in(wire_d24_66),.data_out(wire_d24_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252468(.data_in(wire_d24_67),.data_out(wire_d24_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252469(.data_in(wire_d24_68),.data_out(d_out24),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance26250(.data_in(d_in25),.data_out(wire_d25_0),.clk(clk),.rst(rst));            //channel 26
	large_mux #(.WIDTH(WIDTH)) large_mux_instance26251(.data_in(wire_d25_0),.data_out(wire_d25_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance26252(.data_in(wire_d25_1),.data_out(wire_d25_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance26253(.data_in(wire_d25_2),.data_out(wire_d25_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance26254(.data_in(wire_d25_3),.data_out(wire_d25_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance26255(.data_in(wire_d25_4),.data_out(wire_d25_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance26256(.data_in(wire_d25_5),.data_out(wire_d25_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance26257(.data_in(wire_d25_6),.data_out(wire_d25_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance26258(.data_in(wire_d25_7),.data_out(wire_d25_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance26259(.data_in(wire_d25_8),.data_out(wire_d25_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262510(.data_in(wire_d25_9),.data_out(wire_d25_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262511(.data_in(wire_d25_10),.data_out(wire_d25_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262512(.data_in(wire_d25_11),.data_out(wire_d25_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262513(.data_in(wire_d25_12),.data_out(wire_d25_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262514(.data_in(wire_d25_13),.data_out(wire_d25_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262515(.data_in(wire_d25_14),.data_out(wire_d25_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262516(.data_in(wire_d25_15),.data_out(wire_d25_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262517(.data_in(wire_d25_16),.data_out(wire_d25_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262518(.data_in(wire_d25_17),.data_out(wire_d25_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262519(.data_in(wire_d25_18),.data_out(wire_d25_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262520(.data_in(wire_d25_19),.data_out(wire_d25_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262521(.data_in(wire_d25_20),.data_out(wire_d25_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262522(.data_in(wire_d25_21),.data_out(wire_d25_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262523(.data_in(wire_d25_22),.data_out(wire_d25_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262524(.data_in(wire_d25_23),.data_out(wire_d25_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262525(.data_in(wire_d25_24),.data_out(wire_d25_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262526(.data_in(wire_d25_25),.data_out(wire_d25_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262527(.data_in(wire_d25_26),.data_out(wire_d25_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262528(.data_in(wire_d25_27),.data_out(wire_d25_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262529(.data_in(wire_d25_28),.data_out(wire_d25_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262530(.data_in(wire_d25_29),.data_out(wire_d25_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262531(.data_in(wire_d25_30),.data_out(wire_d25_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262532(.data_in(wire_d25_31),.data_out(wire_d25_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262533(.data_in(wire_d25_32),.data_out(wire_d25_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262534(.data_in(wire_d25_33),.data_out(wire_d25_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262535(.data_in(wire_d25_34),.data_out(wire_d25_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262536(.data_in(wire_d25_35),.data_out(wire_d25_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262537(.data_in(wire_d25_36),.data_out(wire_d25_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262538(.data_in(wire_d25_37),.data_out(wire_d25_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262539(.data_in(wire_d25_38),.data_out(wire_d25_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262540(.data_in(wire_d25_39),.data_out(wire_d25_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262541(.data_in(wire_d25_40),.data_out(wire_d25_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262542(.data_in(wire_d25_41),.data_out(wire_d25_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262543(.data_in(wire_d25_42),.data_out(wire_d25_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262544(.data_in(wire_d25_43),.data_out(wire_d25_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262545(.data_in(wire_d25_44),.data_out(wire_d25_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262546(.data_in(wire_d25_45),.data_out(wire_d25_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262547(.data_in(wire_d25_46),.data_out(wire_d25_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262548(.data_in(wire_d25_47),.data_out(wire_d25_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262549(.data_in(wire_d25_48),.data_out(wire_d25_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262550(.data_in(wire_d25_49),.data_out(wire_d25_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262551(.data_in(wire_d25_50),.data_out(wire_d25_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262552(.data_in(wire_d25_51),.data_out(wire_d25_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262553(.data_in(wire_d25_52),.data_out(wire_d25_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262554(.data_in(wire_d25_53),.data_out(wire_d25_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262555(.data_in(wire_d25_54),.data_out(wire_d25_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262556(.data_in(wire_d25_55),.data_out(wire_d25_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262557(.data_in(wire_d25_56),.data_out(wire_d25_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262558(.data_in(wire_d25_57),.data_out(wire_d25_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262559(.data_in(wire_d25_58),.data_out(wire_d25_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262560(.data_in(wire_d25_59),.data_out(wire_d25_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262561(.data_in(wire_d25_60),.data_out(wire_d25_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262562(.data_in(wire_d25_61),.data_out(wire_d25_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262563(.data_in(wire_d25_62),.data_out(wire_d25_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262564(.data_in(wire_d25_63),.data_out(wire_d25_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262565(.data_in(wire_d25_64),.data_out(wire_d25_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262566(.data_in(wire_d25_65),.data_out(wire_d25_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262567(.data_in(wire_d25_66),.data_out(wire_d25_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262568(.data_in(wire_d25_67),.data_out(wire_d25_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262569(.data_in(wire_d25_68),.data_out(d_out25),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance27260(.data_in(d_in26),.data_out(wire_d26_0),.clk(clk),.rst(rst));            //channel 27
	encoder #(.WIDTH(WIDTH)) encoder_instance27261(.data_in(wire_d26_0),.data_out(wire_d26_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance27262(.data_in(wire_d26_1),.data_out(wire_d26_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance27263(.data_in(wire_d26_2),.data_out(wire_d26_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance27264(.data_in(wire_d26_3),.data_out(wire_d26_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance27265(.data_in(wire_d26_4),.data_out(wire_d26_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance27266(.data_in(wire_d26_5),.data_out(wire_d26_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance27267(.data_in(wire_d26_6),.data_out(wire_d26_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance27268(.data_in(wire_d26_7),.data_out(wire_d26_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance27269(.data_in(wire_d26_8),.data_out(wire_d26_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272610(.data_in(wire_d26_9),.data_out(wire_d26_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272611(.data_in(wire_d26_10),.data_out(wire_d26_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272612(.data_in(wire_d26_11),.data_out(wire_d26_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272613(.data_in(wire_d26_12),.data_out(wire_d26_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272614(.data_in(wire_d26_13),.data_out(wire_d26_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272615(.data_in(wire_d26_14),.data_out(wire_d26_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272616(.data_in(wire_d26_15),.data_out(wire_d26_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272617(.data_in(wire_d26_16),.data_out(wire_d26_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272618(.data_in(wire_d26_17),.data_out(wire_d26_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272619(.data_in(wire_d26_18),.data_out(wire_d26_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272620(.data_in(wire_d26_19),.data_out(wire_d26_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272621(.data_in(wire_d26_20),.data_out(wire_d26_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272622(.data_in(wire_d26_21),.data_out(wire_d26_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272623(.data_in(wire_d26_22),.data_out(wire_d26_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272624(.data_in(wire_d26_23),.data_out(wire_d26_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272625(.data_in(wire_d26_24),.data_out(wire_d26_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272626(.data_in(wire_d26_25),.data_out(wire_d26_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272627(.data_in(wire_d26_26),.data_out(wire_d26_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272628(.data_in(wire_d26_27),.data_out(wire_d26_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272629(.data_in(wire_d26_28),.data_out(wire_d26_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272630(.data_in(wire_d26_29),.data_out(wire_d26_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272631(.data_in(wire_d26_30),.data_out(wire_d26_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272632(.data_in(wire_d26_31),.data_out(wire_d26_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272633(.data_in(wire_d26_32),.data_out(wire_d26_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272634(.data_in(wire_d26_33),.data_out(wire_d26_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272635(.data_in(wire_d26_34),.data_out(wire_d26_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272636(.data_in(wire_d26_35),.data_out(wire_d26_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272637(.data_in(wire_d26_36),.data_out(wire_d26_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272638(.data_in(wire_d26_37),.data_out(wire_d26_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272639(.data_in(wire_d26_38),.data_out(wire_d26_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272640(.data_in(wire_d26_39),.data_out(wire_d26_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272641(.data_in(wire_d26_40),.data_out(wire_d26_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272642(.data_in(wire_d26_41),.data_out(wire_d26_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272643(.data_in(wire_d26_42),.data_out(wire_d26_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272644(.data_in(wire_d26_43),.data_out(wire_d26_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272645(.data_in(wire_d26_44),.data_out(wire_d26_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272646(.data_in(wire_d26_45),.data_out(wire_d26_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272647(.data_in(wire_d26_46),.data_out(wire_d26_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272648(.data_in(wire_d26_47),.data_out(wire_d26_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272649(.data_in(wire_d26_48),.data_out(wire_d26_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272650(.data_in(wire_d26_49),.data_out(wire_d26_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272651(.data_in(wire_d26_50),.data_out(wire_d26_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272652(.data_in(wire_d26_51),.data_out(wire_d26_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272653(.data_in(wire_d26_52),.data_out(wire_d26_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272654(.data_in(wire_d26_53),.data_out(wire_d26_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272655(.data_in(wire_d26_54),.data_out(wire_d26_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272656(.data_in(wire_d26_55),.data_out(wire_d26_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272657(.data_in(wire_d26_56),.data_out(wire_d26_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272658(.data_in(wire_d26_57),.data_out(wire_d26_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272659(.data_in(wire_d26_58),.data_out(wire_d26_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272660(.data_in(wire_d26_59),.data_out(wire_d26_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272661(.data_in(wire_d26_60),.data_out(wire_d26_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272662(.data_in(wire_d26_61),.data_out(wire_d26_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272663(.data_in(wire_d26_62),.data_out(wire_d26_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272664(.data_in(wire_d26_63),.data_out(wire_d26_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272665(.data_in(wire_d26_64),.data_out(wire_d26_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272666(.data_in(wire_d26_65),.data_out(wire_d26_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272667(.data_in(wire_d26_66),.data_out(wire_d26_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272668(.data_in(wire_d26_67),.data_out(wire_d26_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272669(.data_in(wire_d26_68),.data_out(d_out26),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance28270(.data_in(d_in27),.data_out(wire_d27_0),.clk(clk),.rst(rst));            //channel 28
	register #(.WIDTH(WIDTH)) register_instance28271(.data_in(wire_d27_0),.data_out(wire_d27_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance28272(.data_in(wire_d27_1),.data_out(wire_d27_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance28273(.data_in(wire_d27_2),.data_out(wire_d27_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance28274(.data_in(wire_d27_3),.data_out(wire_d27_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance28275(.data_in(wire_d27_4),.data_out(wire_d27_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance28276(.data_in(wire_d27_5),.data_out(wire_d27_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance28277(.data_in(wire_d27_6),.data_out(wire_d27_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance28278(.data_in(wire_d27_7),.data_out(wire_d27_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance28279(.data_in(wire_d27_8),.data_out(wire_d27_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282710(.data_in(wire_d27_9),.data_out(wire_d27_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282711(.data_in(wire_d27_10),.data_out(wire_d27_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282712(.data_in(wire_d27_11),.data_out(wire_d27_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282713(.data_in(wire_d27_12),.data_out(wire_d27_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282714(.data_in(wire_d27_13),.data_out(wire_d27_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282715(.data_in(wire_d27_14),.data_out(wire_d27_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282716(.data_in(wire_d27_15),.data_out(wire_d27_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282717(.data_in(wire_d27_16),.data_out(wire_d27_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282718(.data_in(wire_d27_17),.data_out(wire_d27_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282719(.data_in(wire_d27_18),.data_out(wire_d27_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282720(.data_in(wire_d27_19),.data_out(wire_d27_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282721(.data_in(wire_d27_20),.data_out(wire_d27_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282722(.data_in(wire_d27_21),.data_out(wire_d27_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282723(.data_in(wire_d27_22),.data_out(wire_d27_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282724(.data_in(wire_d27_23),.data_out(wire_d27_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282725(.data_in(wire_d27_24),.data_out(wire_d27_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282726(.data_in(wire_d27_25),.data_out(wire_d27_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282727(.data_in(wire_d27_26),.data_out(wire_d27_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282728(.data_in(wire_d27_27),.data_out(wire_d27_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282729(.data_in(wire_d27_28),.data_out(wire_d27_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282730(.data_in(wire_d27_29),.data_out(wire_d27_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282731(.data_in(wire_d27_30),.data_out(wire_d27_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282732(.data_in(wire_d27_31),.data_out(wire_d27_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282733(.data_in(wire_d27_32),.data_out(wire_d27_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282734(.data_in(wire_d27_33),.data_out(wire_d27_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282735(.data_in(wire_d27_34),.data_out(wire_d27_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282736(.data_in(wire_d27_35),.data_out(wire_d27_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282737(.data_in(wire_d27_36),.data_out(wire_d27_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282738(.data_in(wire_d27_37),.data_out(wire_d27_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282739(.data_in(wire_d27_38),.data_out(wire_d27_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282740(.data_in(wire_d27_39),.data_out(wire_d27_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282741(.data_in(wire_d27_40),.data_out(wire_d27_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282742(.data_in(wire_d27_41),.data_out(wire_d27_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282743(.data_in(wire_d27_42),.data_out(wire_d27_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282744(.data_in(wire_d27_43),.data_out(wire_d27_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282745(.data_in(wire_d27_44),.data_out(wire_d27_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282746(.data_in(wire_d27_45),.data_out(wire_d27_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282747(.data_in(wire_d27_46),.data_out(wire_d27_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282748(.data_in(wire_d27_47),.data_out(wire_d27_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282749(.data_in(wire_d27_48),.data_out(wire_d27_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282750(.data_in(wire_d27_49),.data_out(wire_d27_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282751(.data_in(wire_d27_50),.data_out(wire_d27_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282752(.data_in(wire_d27_51),.data_out(wire_d27_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282753(.data_in(wire_d27_52),.data_out(wire_d27_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282754(.data_in(wire_d27_53),.data_out(wire_d27_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282755(.data_in(wire_d27_54),.data_out(wire_d27_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282756(.data_in(wire_d27_55),.data_out(wire_d27_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282757(.data_in(wire_d27_56),.data_out(wire_d27_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282758(.data_in(wire_d27_57),.data_out(wire_d27_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282759(.data_in(wire_d27_58),.data_out(wire_d27_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282760(.data_in(wire_d27_59),.data_out(wire_d27_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282761(.data_in(wire_d27_60),.data_out(wire_d27_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282762(.data_in(wire_d27_61),.data_out(wire_d27_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282763(.data_in(wire_d27_62),.data_out(wire_d27_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282764(.data_in(wire_d27_63),.data_out(wire_d27_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282765(.data_in(wire_d27_64),.data_out(wire_d27_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282766(.data_in(wire_d27_65),.data_out(wire_d27_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282767(.data_in(wire_d27_66),.data_out(wire_d27_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282768(.data_in(wire_d27_67),.data_out(wire_d27_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282769(.data_in(wire_d27_68),.data_out(d_out27),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance29280(.data_in(d_in28),.data_out(wire_d28_0),.clk(clk),.rst(rst));            //channel 29
	large_mux #(.WIDTH(WIDTH)) large_mux_instance29281(.data_in(wire_d28_0),.data_out(wire_d28_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance29282(.data_in(wire_d28_1),.data_out(wire_d28_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance29283(.data_in(wire_d28_2),.data_out(wire_d28_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance29284(.data_in(wire_d28_3),.data_out(wire_d28_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance29285(.data_in(wire_d28_4),.data_out(wire_d28_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance29286(.data_in(wire_d28_5),.data_out(wire_d28_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance29287(.data_in(wire_d28_6),.data_out(wire_d28_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance29288(.data_in(wire_d28_7),.data_out(wire_d28_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance29289(.data_in(wire_d28_8),.data_out(wire_d28_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292810(.data_in(wire_d28_9),.data_out(wire_d28_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292811(.data_in(wire_d28_10),.data_out(wire_d28_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292812(.data_in(wire_d28_11),.data_out(wire_d28_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292813(.data_in(wire_d28_12),.data_out(wire_d28_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292814(.data_in(wire_d28_13),.data_out(wire_d28_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292815(.data_in(wire_d28_14),.data_out(wire_d28_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292816(.data_in(wire_d28_15),.data_out(wire_d28_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292817(.data_in(wire_d28_16),.data_out(wire_d28_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292818(.data_in(wire_d28_17),.data_out(wire_d28_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292819(.data_in(wire_d28_18),.data_out(wire_d28_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292820(.data_in(wire_d28_19),.data_out(wire_d28_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292821(.data_in(wire_d28_20),.data_out(wire_d28_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292822(.data_in(wire_d28_21),.data_out(wire_d28_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292823(.data_in(wire_d28_22),.data_out(wire_d28_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292824(.data_in(wire_d28_23),.data_out(wire_d28_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292825(.data_in(wire_d28_24),.data_out(wire_d28_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292826(.data_in(wire_d28_25),.data_out(wire_d28_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292827(.data_in(wire_d28_26),.data_out(wire_d28_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292828(.data_in(wire_d28_27),.data_out(wire_d28_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292829(.data_in(wire_d28_28),.data_out(wire_d28_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292830(.data_in(wire_d28_29),.data_out(wire_d28_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292831(.data_in(wire_d28_30),.data_out(wire_d28_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292832(.data_in(wire_d28_31),.data_out(wire_d28_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292833(.data_in(wire_d28_32),.data_out(wire_d28_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292834(.data_in(wire_d28_33),.data_out(wire_d28_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292835(.data_in(wire_d28_34),.data_out(wire_d28_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292836(.data_in(wire_d28_35),.data_out(wire_d28_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292837(.data_in(wire_d28_36),.data_out(wire_d28_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292838(.data_in(wire_d28_37),.data_out(wire_d28_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292839(.data_in(wire_d28_38),.data_out(wire_d28_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292840(.data_in(wire_d28_39),.data_out(wire_d28_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292841(.data_in(wire_d28_40),.data_out(wire_d28_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292842(.data_in(wire_d28_41),.data_out(wire_d28_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292843(.data_in(wire_d28_42),.data_out(wire_d28_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292844(.data_in(wire_d28_43),.data_out(wire_d28_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292845(.data_in(wire_d28_44),.data_out(wire_d28_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292846(.data_in(wire_d28_45),.data_out(wire_d28_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292847(.data_in(wire_d28_46),.data_out(wire_d28_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292848(.data_in(wire_d28_47),.data_out(wire_d28_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292849(.data_in(wire_d28_48),.data_out(wire_d28_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292850(.data_in(wire_d28_49),.data_out(wire_d28_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292851(.data_in(wire_d28_50),.data_out(wire_d28_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292852(.data_in(wire_d28_51),.data_out(wire_d28_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292853(.data_in(wire_d28_52),.data_out(wire_d28_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292854(.data_in(wire_d28_53),.data_out(wire_d28_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292855(.data_in(wire_d28_54),.data_out(wire_d28_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292856(.data_in(wire_d28_55),.data_out(wire_d28_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292857(.data_in(wire_d28_56),.data_out(wire_d28_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292858(.data_in(wire_d28_57),.data_out(wire_d28_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292859(.data_in(wire_d28_58),.data_out(wire_d28_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292860(.data_in(wire_d28_59),.data_out(wire_d28_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292861(.data_in(wire_d28_60),.data_out(wire_d28_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292862(.data_in(wire_d28_61),.data_out(wire_d28_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292863(.data_in(wire_d28_62),.data_out(wire_d28_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292864(.data_in(wire_d28_63),.data_out(wire_d28_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292865(.data_in(wire_d28_64),.data_out(wire_d28_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292866(.data_in(wire_d28_65),.data_out(wire_d28_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292867(.data_in(wire_d28_66),.data_out(wire_d28_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292868(.data_in(wire_d28_67),.data_out(wire_d28_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292869(.data_in(wire_d28_68),.data_out(d_out28),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance30290(.data_in(d_in29),.data_out(wire_d29_0),.clk(clk),.rst(rst));            //channel 30
	register #(.WIDTH(WIDTH)) register_instance30291(.data_in(wire_d29_0),.data_out(wire_d29_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance30292(.data_in(wire_d29_1),.data_out(wire_d29_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance30293(.data_in(wire_d29_2),.data_out(wire_d29_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance30294(.data_in(wire_d29_3),.data_out(wire_d29_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance30295(.data_in(wire_d29_4),.data_out(wire_d29_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance30296(.data_in(wire_d29_5),.data_out(wire_d29_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance30297(.data_in(wire_d29_6),.data_out(wire_d29_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance30298(.data_in(wire_d29_7),.data_out(wire_d29_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance30299(.data_in(wire_d29_8),.data_out(wire_d29_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302910(.data_in(wire_d29_9),.data_out(wire_d29_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302911(.data_in(wire_d29_10),.data_out(wire_d29_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302912(.data_in(wire_d29_11),.data_out(wire_d29_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302913(.data_in(wire_d29_12),.data_out(wire_d29_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302914(.data_in(wire_d29_13),.data_out(wire_d29_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302915(.data_in(wire_d29_14),.data_out(wire_d29_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302916(.data_in(wire_d29_15),.data_out(wire_d29_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302917(.data_in(wire_d29_16),.data_out(wire_d29_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302918(.data_in(wire_d29_17),.data_out(wire_d29_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302919(.data_in(wire_d29_18),.data_out(wire_d29_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302920(.data_in(wire_d29_19),.data_out(wire_d29_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302921(.data_in(wire_d29_20),.data_out(wire_d29_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302922(.data_in(wire_d29_21),.data_out(wire_d29_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302923(.data_in(wire_d29_22),.data_out(wire_d29_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302924(.data_in(wire_d29_23),.data_out(wire_d29_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302925(.data_in(wire_d29_24),.data_out(wire_d29_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302926(.data_in(wire_d29_25),.data_out(wire_d29_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302927(.data_in(wire_d29_26),.data_out(wire_d29_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302928(.data_in(wire_d29_27),.data_out(wire_d29_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302929(.data_in(wire_d29_28),.data_out(wire_d29_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302930(.data_in(wire_d29_29),.data_out(wire_d29_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302931(.data_in(wire_d29_30),.data_out(wire_d29_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302932(.data_in(wire_d29_31),.data_out(wire_d29_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302933(.data_in(wire_d29_32),.data_out(wire_d29_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302934(.data_in(wire_d29_33),.data_out(wire_d29_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302935(.data_in(wire_d29_34),.data_out(wire_d29_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302936(.data_in(wire_d29_35),.data_out(wire_d29_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302937(.data_in(wire_d29_36),.data_out(wire_d29_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302938(.data_in(wire_d29_37),.data_out(wire_d29_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302939(.data_in(wire_d29_38),.data_out(wire_d29_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302940(.data_in(wire_d29_39),.data_out(wire_d29_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302941(.data_in(wire_d29_40),.data_out(wire_d29_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302942(.data_in(wire_d29_41),.data_out(wire_d29_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302943(.data_in(wire_d29_42),.data_out(wire_d29_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302944(.data_in(wire_d29_43),.data_out(wire_d29_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302945(.data_in(wire_d29_44),.data_out(wire_d29_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302946(.data_in(wire_d29_45),.data_out(wire_d29_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302947(.data_in(wire_d29_46),.data_out(wire_d29_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302948(.data_in(wire_d29_47),.data_out(wire_d29_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302949(.data_in(wire_d29_48),.data_out(wire_d29_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302950(.data_in(wire_d29_49),.data_out(wire_d29_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302951(.data_in(wire_d29_50),.data_out(wire_d29_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302952(.data_in(wire_d29_51),.data_out(wire_d29_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302953(.data_in(wire_d29_52),.data_out(wire_d29_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302954(.data_in(wire_d29_53),.data_out(wire_d29_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302955(.data_in(wire_d29_54),.data_out(wire_d29_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302956(.data_in(wire_d29_55),.data_out(wire_d29_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302957(.data_in(wire_d29_56),.data_out(wire_d29_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302958(.data_in(wire_d29_57),.data_out(wire_d29_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302959(.data_in(wire_d29_58),.data_out(wire_d29_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302960(.data_in(wire_d29_59),.data_out(wire_d29_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302961(.data_in(wire_d29_60),.data_out(wire_d29_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302962(.data_in(wire_d29_61),.data_out(wire_d29_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302963(.data_in(wire_d29_62),.data_out(wire_d29_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302964(.data_in(wire_d29_63),.data_out(wire_d29_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302965(.data_in(wire_d29_64),.data_out(wire_d29_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302966(.data_in(wire_d29_65),.data_out(wire_d29_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302967(.data_in(wire_d29_66),.data_out(wire_d29_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302968(.data_in(wire_d29_67),.data_out(wire_d29_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302969(.data_in(wire_d29_68),.data_out(d_out29),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance31300(.data_in(d_in30),.data_out(wire_d30_0),.clk(clk),.rst(rst));            //channel 31
	large_mux #(.WIDTH(WIDTH)) large_mux_instance31301(.data_in(wire_d30_0),.data_out(wire_d30_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance31302(.data_in(wire_d30_1),.data_out(wire_d30_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance31303(.data_in(wire_d30_2),.data_out(wire_d30_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance31304(.data_in(wire_d30_3),.data_out(wire_d30_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance31305(.data_in(wire_d30_4),.data_out(wire_d30_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance31306(.data_in(wire_d30_5),.data_out(wire_d30_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance31307(.data_in(wire_d30_6),.data_out(wire_d30_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance31308(.data_in(wire_d30_7),.data_out(wire_d30_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance31309(.data_in(wire_d30_8),.data_out(wire_d30_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313010(.data_in(wire_d30_9),.data_out(wire_d30_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313011(.data_in(wire_d30_10),.data_out(wire_d30_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313012(.data_in(wire_d30_11),.data_out(wire_d30_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313013(.data_in(wire_d30_12),.data_out(wire_d30_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313014(.data_in(wire_d30_13),.data_out(wire_d30_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313015(.data_in(wire_d30_14),.data_out(wire_d30_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313016(.data_in(wire_d30_15),.data_out(wire_d30_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313017(.data_in(wire_d30_16),.data_out(wire_d30_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313018(.data_in(wire_d30_17),.data_out(wire_d30_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313019(.data_in(wire_d30_18),.data_out(wire_d30_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313020(.data_in(wire_d30_19),.data_out(wire_d30_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313021(.data_in(wire_d30_20),.data_out(wire_d30_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313022(.data_in(wire_d30_21),.data_out(wire_d30_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313023(.data_in(wire_d30_22),.data_out(wire_d30_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313024(.data_in(wire_d30_23),.data_out(wire_d30_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313025(.data_in(wire_d30_24),.data_out(wire_d30_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313026(.data_in(wire_d30_25),.data_out(wire_d30_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313027(.data_in(wire_d30_26),.data_out(wire_d30_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313028(.data_in(wire_d30_27),.data_out(wire_d30_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313029(.data_in(wire_d30_28),.data_out(wire_d30_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313030(.data_in(wire_d30_29),.data_out(wire_d30_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313031(.data_in(wire_d30_30),.data_out(wire_d30_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313032(.data_in(wire_d30_31),.data_out(wire_d30_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313033(.data_in(wire_d30_32),.data_out(wire_d30_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313034(.data_in(wire_d30_33),.data_out(wire_d30_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313035(.data_in(wire_d30_34),.data_out(wire_d30_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313036(.data_in(wire_d30_35),.data_out(wire_d30_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313037(.data_in(wire_d30_36),.data_out(wire_d30_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313038(.data_in(wire_d30_37),.data_out(wire_d30_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313039(.data_in(wire_d30_38),.data_out(wire_d30_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313040(.data_in(wire_d30_39),.data_out(wire_d30_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313041(.data_in(wire_d30_40),.data_out(wire_d30_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313042(.data_in(wire_d30_41),.data_out(wire_d30_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313043(.data_in(wire_d30_42),.data_out(wire_d30_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313044(.data_in(wire_d30_43),.data_out(wire_d30_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313045(.data_in(wire_d30_44),.data_out(wire_d30_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313046(.data_in(wire_d30_45),.data_out(wire_d30_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313047(.data_in(wire_d30_46),.data_out(wire_d30_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313048(.data_in(wire_d30_47),.data_out(wire_d30_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313049(.data_in(wire_d30_48),.data_out(wire_d30_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313050(.data_in(wire_d30_49),.data_out(wire_d30_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313051(.data_in(wire_d30_50),.data_out(wire_d30_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313052(.data_in(wire_d30_51),.data_out(wire_d30_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313053(.data_in(wire_d30_52),.data_out(wire_d30_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313054(.data_in(wire_d30_53),.data_out(wire_d30_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313055(.data_in(wire_d30_54),.data_out(wire_d30_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313056(.data_in(wire_d30_55),.data_out(wire_d30_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313057(.data_in(wire_d30_56),.data_out(wire_d30_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313058(.data_in(wire_d30_57),.data_out(wire_d30_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313059(.data_in(wire_d30_58),.data_out(wire_d30_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313060(.data_in(wire_d30_59),.data_out(wire_d30_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313061(.data_in(wire_d30_60),.data_out(wire_d30_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313062(.data_in(wire_d30_61),.data_out(wire_d30_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313063(.data_in(wire_d30_62),.data_out(wire_d30_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance313064(.data_in(wire_d30_63),.data_out(wire_d30_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313065(.data_in(wire_d30_64),.data_out(wire_d30_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313066(.data_in(wire_d30_65),.data_out(wire_d30_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance313067(.data_in(wire_d30_66),.data_out(wire_d30_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance313068(.data_in(wire_d30_67),.data_out(wire_d30_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance313069(.data_in(wire_d30_68),.data_out(d_out30),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance32310(.data_in(d_in31),.data_out(wire_d31_0),.clk(clk),.rst(rst));            //channel 32
	encoder #(.WIDTH(WIDTH)) encoder_instance32311(.data_in(wire_d31_0),.data_out(wire_d31_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance32312(.data_in(wire_d31_1),.data_out(wire_d31_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance32313(.data_in(wire_d31_2),.data_out(wire_d31_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance32314(.data_in(wire_d31_3),.data_out(wire_d31_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance32315(.data_in(wire_d31_4),.data_out(wire_d31_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance32316(.data_in(wire_d31_5),.data_out(wire_d31_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance32317(.data_in(wire_d31_6),.data_out(wire_d31_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance32318(.data_in(wire_d31_7),.data_out(wire_d31_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32319(.data_in(wire_d31_8),.data_out(wire_d31_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323110(.data_in(wire_d31_9),.data_out(wire_d31_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323111(.data_in(wire_d31_10),.data_out(wire_d31_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323112(.data_in(wire_d31_11),.data_out(wire_d31_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323113(.data_in(wire_d31_12),.data_out(wire_d31_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323114(.data_in(wire_d31_13),.data_out(wire_d31_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323115(.data_in(wire_d31_14),.data_out(wire_d31_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323116(.data_in(wire_d31_15),.data_out(wire_d31_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323117(.data_in(wire_d31_16),.data_out(wire_d31_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323118(.data_in(wire_d31_17),.data_out(wire_d31_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323119(.data_in(wire_d31_18),.data_out(wire_d31_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323120(.data_in(wire_d31_19),.data_out(wire_d31_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323121(.data_in(wire_d31_20),.data_out(wire_d31_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323122(.data_in(wire_d31_21),.data_out(wire_d31_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323123(.data_in(wire_d31_22),.data_out(wire_d31_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323124(.data_in(wire_d31_23),.data_out(wire_d31_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323125(.data_in(wire_d31_24),.data_out(wire_d31_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323126(.data_in(wire_d31_25),.data_out(wire_d31_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323127(.data_in(wire_d31_26),.data_out(wire_d31_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323128(.data_in(wire_d31_27),.data_out(wire_d31_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323129(.data_in(wire_d31_28),.data_out(wire_d31_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323130(.data_in(wire_d31_29),.data_out(wire_d31_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323131(.data_in(wire_d31_30),.data_out(wire_d31_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323132(.data_in(wire_d31_31),.data_out(wire_d31_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323133(.data_in(wire_d31_32),.data_out(wire_d31_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323134(.data_in(wire_d31_33),.data_out(wire_d31_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323135(.data_in(wire_d31_34),.data_out(wire_d31_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323136(.data_in(wire_d31_35),.data_out(wire_d31_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323137(.data_in(wire_d31_36),.data_out(wire_d31_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323138(.data_in(wire_d31_37),.data_out(wire_d31_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323139(.data_in(wire_d31_38),.data_out(wire_d31_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323140(.data_in(wire_d31_39),.data_out(wire_d31_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323141(.data_in(wire_d31_40),.data_out(wire_d31_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323142(.data_in(wire_d31_41),.data_out(wire_d31_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323143(.data_in(wire_d31_42),.data_out(wire_d31_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323144(.data_in(wire_d31_43),.data_out(wire_d31_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323145(.data_in(wire_d31_44),.data_out(wire_d31_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323146(.data_in(wire_d31_45),.data_out(wire_d31_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323147(.data_in(wire_d31_46),.data_out(wire_d31_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323148(.data_in(wire_d31_47),.data_out(wire_d31_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323149(.data_in(wire_d31_48),.data_out(wire_d31_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323150(.data_in(wire_d31_49),.data_out(wire_d31_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323151(.data_in(wire_d31_50),.data_out(wire_d31_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323152(.data_in(wire_d31_51),.data_out(wire_d31_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323153(.data_in(wire_d31_52),.data_out(wire_d31_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323154(.data_in(wire_d31_53),.data_out(wire_d31_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323155(.data_in(wire_d31_54),.data_out(wire_d31_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323156(.data_in(wire_d31_55),.data_out(wire_d31_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323157(.data_in(wire_d31_56),.data_out(wire_d31_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323158(.data_in(wire_d31_57),.data_out(wire_d31_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323159(.data_in(wire_d31_58),.data_out(wire_d31_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323160(.data_in(wire_d31_59),.data_out(wire_d31_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance323161(.data_in(wire_d31_60),.data_out(wire_d31_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323162(.data_in(wire_d31_61),.data_out(wire_d31_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323163(.data_in(wire_d31_62),.data_out(wire_d31_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323164(.data_in(wire_d31_63),.data_out(wire_d31_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323165(.data_in(wire_d31_64),.data_out(wire_d31_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323166(.data_in(wire_d31_65),.data_out(wire_d31_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323167(.data_in(wire_d31_66),.data_out(wire_d31_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance323168(.data_in(wire_d31_67),.data_out(wire_d31_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323169(.data_in(wire_d31_68),.data_out(d_out31),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance33320(.data_in(d_in32),.data_out(wire_d32_0),.clk(clk),.rst(rst));            //channel 33
	invertion #(.WIDTH(WIDTH)) invertion_instance33321(.data_in(wire_d32_0),.data_out(wire_d32_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance33322(.data_in(wire_d32_1),.data_out(wire_d32_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance33323(.data_in(wire_d32_2),.data_out(wire_d32_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance33324(.data_in(wire_d32_3),.data_out(wire_d32_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance33325(.data_in(wire_d32_4),.data_out(wire_d32_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance33326(.data_in(wire_d32_5),.data_out(wire_d32_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance33327(.data_in(wire_d32_6),.data_out(wire_d32_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance33328(.data_in(wire_d32_7),.data_out(wire_d32_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance33329(.data_in(wire_d32_8),.data_out(wire_d32_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333210(.data_in(wire_d32_9),.data_out(wire_d32_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333211(.data_in(wire_d32_10),.data_out(wire_d32_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333212(.data_in(wire_d32_11),.data_out(wire_d32_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333213(.data_in(wire_d32_12),.data_out(wire_d32_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333214(.data_in(wire_d32_13),.data_out(wire_d32_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333215(.data_in(wire_d32_14),.data_out(wire_d32_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333216(.data_in(wire_d32_15),.data_out(wire_d32_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333217(.data_in(wire_d32_16),.data_out(wire_d32_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333218(.data_in(wire_d32_17),.data_out(wire_d32_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333219(.data_in(wire_d32_18),.data_out(wire_d32_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333220(.data_in(wire_d32_19),.data_out(wire_d32_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333221(.data_in(wire_d32_20),.data_out(wire_d32_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333222(.data_in(wire_d32_21),.data_out(wire_d32_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333223(.data_in(wire_d32_22),.data_out(wire_d32_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333224(.data_in(wire_d32_23),.data_out(wire_d32_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333225(.data_in(wire_d32_24),.data_out(wire_d32_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333226(.data_in(wire_d32_25),.data_out(wire_d32_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333227(.data_in(wire_d32_26),.data_out(wire_d32_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333228(.data_in(wire_d32_27),.data_out(wire_d32_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333229(.data_in(wire_d32_28),.data_out(wire_d32_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333230(.data_in(wire_d32_29),.data_out(wire_d32_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333231(.data_in(wire_d32_30),.data_out(wire_d32_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333232(.data_in(wire_d32_31),.data_out(wire_d32_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333233(.data_in(wire_d32_32),.data_out(wire_d32_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333234(.data_in(wire_d32_33),.data_out(wire_d32_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333235(.data_in(wire_d32_34),.data_out(wire_d32_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333236(.data_in(wire_d32_35),.data_out(wire_d32_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333237(.data_in(wire_d32_36),.data_out(wire_d32_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333238(.data_in(wire_d32_37),.data_out(wire_d32_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333239(.data_in(wire_d32_38),.data_out(wire_d32_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333240(.data_in(wire_d32_39),.data_out(wire_d32_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333241(.data_in(wire_d32_40),.data_out(wire_d32_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333242(.data_in(wire_d32_41),.data_out(wire_d32_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333243(.data_in(wire_d32_42),.data_out(wire_d32_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333244(.data_in(wire_d32_43),.data_out(wire_d32_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333245(.data_in(wire_d32_44),.data_out(wire_d32_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333246(.data_in(wire_d32_45),.data_out(wire_d32_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333247(.data_in(wire_d32_46),.data_out(wire_d32_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333248(.data_in(wire_d32_47),.data_out(wire_d32_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333249(.data_in(wire_d32_48),.data_out(wire_d32_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333250(.data_in(wire_d32_49),.data_out(wire_d32_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333251(.data_in(wire_d32_50),.data_out(wire_d32_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333252(.data_in(wire_d32_51),.data_out(wire_d32_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333253(.data_in(wire_d32_52),.data_out(wire_d32_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333254(.data_in(wire_d32_53),.data_out(wire_d32_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333255(.data_in(wire_d32_54),.data_out(wire_d32_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333256(.data_in(wire_d32_55),.data_out(wire_d32_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333257(.data_in(wire_d32_56),.data_out(wire_d32_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333258(.data_in(wire_d32_57),.data_out(wire_d32_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333259(.data_in(wire_d32_58),.data_out(wire_d32_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333260(.data_in(wire_d32_59),.data_out(wire_d32_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333261(.data_in(wire_d32_60),.data_out(wire_d32_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333262(.data_in(wire_d32_61),.data_out(wire_d32_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333263(.data_in(wire_d32_62),.data_out(wire_d32_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance333264(.data_in(wire_d32_63),.data_out(wire_d32_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333265(.data_in(wire_d32_64),.data_out(wire_d32_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance333266(.data_in(wire_d32_65),.data_out(wire_d32_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333267(.data_in(wire_d32_66),.data_out(wire_d32_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance333268(.data_in(wire_d32_67),.data_out(wire_d32_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance333269(.data_in(wire_d32_68),.data_out(d_out32),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance34330(.data_in(d_in33),.data_out(wire_d33_0),.clk(clk),.rst(rst));            //channel 34
	encoder #(.WIDTH(WIDTH)) encoder_instance34331(.data_in(wire_d33_0),.data_out(wire_d33_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance34332(.data_in(wire_d33_1),.data_out(wire_d33_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance34333(.data_in(wire_d33_2),.data_out(wire_d33_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance34334(.data_in(wire_d33_3),.data_out(wire_d33_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance34335(.data_in(wire_d33_4),.data_out(wire_d33_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance34336(.data_in(wire_d33_5),.data_out(wire_d33_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance34337(.data_in(wire_d33_6),.data_out(wire_d33_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance34338(.data_in(wire_d33_7),.data_out(wire_d33_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance34339(.data_in(wire_d33_8),.data_out(wire_d33_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343310(.data_in(wire_d33_9),.data_out(wire_d33_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343311(.data_in(wire_d33_10),.data_out(wire_d33_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343312(.data_in(wire_d33_11),.data_out(wire_d33_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343313(.data_in(wire_d33_12),.data_out(wire_d33_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343314(.data_in(wire_d33_13),.data_out(wire_d33_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343315(.data_in(wire_d33_14),.data_out(wire_d33_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343316(.data_in(wire_d33_15),.data_out(wire_d33_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343317(.data_in(wire_d33_16),.data_out(wire_d33_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343318(.data_in(wire_d33_17),.data_out(wire_d33_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343319(.data_in(wire_d33_18),.data_out(wire_d33_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343320(.data_in(wire_d33_19),.data_out(wire_d33_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343321(.data_in(wire_d33_20),.data_out(wire_d33_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343322(.data_in(wire_d33_21),.data_out(wire_d33_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343323(.data_in(wire_d33_22),.data_out(wire_d33_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343324(.data_in(wire_d33_23),.data_out(wire_d33_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343325(.data_in(wire_d33_24),.data_out(wire_d33_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343326(.data_in(wire_d33_25),.data_out(wire_d33_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343327(.data_in(wire_d33_26),.data_out(wire_d33_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343328(.data_in(wire_d33_27),.data_out(wire_d33_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343329(.data_in(wire_d33_28),.data_out(wire_d33_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343330(.data_in(wire_d33_29),.data_out(wire_d33_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343331(.data_in(wire_d33_30),.data_out(wire_d33_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343332(.data_in(wire_d33_31),.data_out(wire_d33_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343333(.data_in(wire_d33_32),.data_out(wire_d33_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343334(.data_in(wire_d33_33),.data_out(wire_d33_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343335(.data_in(wire_d33_34),.data_out(wire_d33_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343336(.data_in(wire_d33_35),.data_out(wire_d33_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343337(.data_in(wire_d33_36),.data_out(wire_d33_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343338(.data_in(wire_d33_37),.data_out(wire_d33_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343339(.data_in(wire_d33_38),.data_out(wire_d33_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343340(.data_in(wire_d33_39),.data_out(wire_d33_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343341(.data_in(wire_d33_40),.data_out(wire_d33_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343342(.data_in(wire_d33_41),.data_out(wire_d33_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343343(.data_in(wire_d33_42),.data_out(wire_d33_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343344(.data_in(wire_d33_43),.data_out(wire_d33_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343345(.data_in(wire_d33_44),.data_out(wire_d33_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343346(.data_in(wire_d33_45),.data_out(wire_d33_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343347(.data_in(wire_d33_46),.data_out(wire_d33_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343348(.data_in(wire_d33_47),.data_out(wire_d33_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343349(.data_in(wire_d33_48),.data_out(wire_d33_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343350(.data_in(wire_d33_49),.data_out(wire_d33_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343351(.data_in(wire_d33_50),.data_out(wire_d33_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343352(.data_in(wire_d33_51),.data_out(wire_d33_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343353(.data_in(wire_d33_52),.data_out(wire_d33_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343354(.data_in(wire_d33_53),.data_out(wire_d33_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343355(.data_in(wire_d33_54),.data_out(wire_d33_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343356(.data_in(wire_d33_55),.data_out(wire_d33_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343357(.data_in(wire_d33_56),.data_out(wire_d33_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343358(.data_in(wire_d33_57),.data_out(wire_d33_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343359(.data_in(wire_d33_58),.data_out(wire_d33_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343360(.data_in(wire_d33_59),.data_out(wire_d33_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance343361(.data_in(wire_d33_60),.data_out(wire_d33_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343362(.data_in(wire_d33_61),.data_out(wire_d33_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343363(.data_in(wire_d33_62),.data_out(wire_d33_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343364(.data_in(wire_d33_63),.data_out(wire_d33_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance343365(.data_in(wire_d33_64),.data_out(wire_d33_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance343366(.data_in(wire_d33_65),.data_out(wire_d33_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343367(.data_in(wire_d33_66),.data_out(wire_d33_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343368(.data_in(wire_d33_67),.data_out(wire_d33_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance343369(.data_in(wire_d33_68),.data_out(d_out33),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance35340(.data_in(d_in34),.data_out(wire_d34_0),.clk(clk),.rst(rst));            //channel 35
	register #(.WIDTH(WIDTH)) register_instance35341(.data_in(wire_d34_0),.data_out(wire_d34_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance35342(.data_in(wire_d34_1),.data_out(wire_d34_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance35343(.data_in(wire_d34_2),.data_out(wire_d34_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance35344(.data_in(wire_d34_3),.data_out(wire_d34_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance35345(.data_in(wire_d34_4),.data_out(wire_d34_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance35346(.data_in(wire_d34_5),.data_out(wire_d34_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance35347(.data_in(wire_d34_6),.data_out(wire_d34_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance35348(.data_in(wire_d34_7),.data_out(wire_d34_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance35349(.data_in(wire_d34_8),.data_out(wire_d34_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353410(.data_in(wire_d34_9),.data_out(wire_d34_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353411(.data_in(wire_d34_10),.data_out(wire_d34_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353412(.data_in(wire_d34_11),.data_out(wire_d34_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353413(.data_in(wire_d34_12),.data_out(wire_d34_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353414(.data_in(wire_d34_13),.data_out(wire_d34_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353415(.data_in(wire_d34_14),.data_out(wire_d34_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353416(.data_in(wire_d34_15),.data_out(wire_d34_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353417(.data_in(wire_d34_16),.data_out(wire_d34_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353418(.data_in(wire_d34_17),.data_out(wire_d34_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353419(.data_in(wire_d34_18),.data_out(wire_d34_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353420(.data_in(wire_d34_19),.data_out(wire_d34_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353421(.data_in(wire_d34_20),.data_out(wire_d34_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353422(.data_in(wire_d34_21),.data_out(wire_d34_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353423(.data_in(wire_d34_22),.data_out(wire_d34_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353424(.data_in(wire_d34_23),.data_out(wire_d34_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353425(.data_in(wire_d34_24),.data_out(wire_d34_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353426(.data_in(wire_d34_25),.data_out(wire_d34_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353427(.data_in(wire_d34_26),.data_out(wire_d34_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353428(.data_in(wire_d34_27),.data_out(wire_d34_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353429(.data_in(wire_d34_28),.data_out(wire_d34_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353430(.data_in(wire_d34_29),.data_out(wire_d34_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353431(.data_in(wire_d34_30),.data_out(wire_d34_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353432(.data_in(wire_d34_31),.data_out(wire_d34_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353433(.data_in(wire_d34_32),.data_out(wire_d34_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353434(.data_in(wire_d34_33),.data_out(wire_d34_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353435(.data_in(wire_d34_34),.data_out(wire_d34_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353436(.data_in(wire_d34_35),.data_out(wire_d34_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353437(.data_in(wire_d34_36),.data_out(wire_d34_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353438(.data_in(wire_d34_37),.data_out(wire_d34_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353439(.data_in(wire_d34_38),.data_out(wire_d34_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353440(.data_in(wire_d34_39),.data_out(wire_d34_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353441(.data_in(wire_d34_40),.data_out(wire_d34_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353442(.data_in(wire_d34_41),.data_out(wire_d34_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353443(.data_in(wire_d34_42),.data_out(wire_d34_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353444(.data_in(wire_d34_43),.data_out(wire_d34_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353445(.data_in(wire_d34_44),.data_out(wire_d34_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353446(.data_in(wire_d34_45),.data_out(wire_d34_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353447(.data_in(wire_d34_46),.data_out(wire_d34_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353448(.data_in(wire_d34_47),.data_out(wire_d34_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353449(.data_in(wire_d34_48),.data_out(wire_d34_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353450(.data_in(wire_d34_49),.data_out(wire_d34_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353451(.data_in(wire_d34_50),.data_out(wire_d34_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353452(.data_in(wire_d34_51),.data_out(wire_d34_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353453(.data_in(wire_d34_52),.data_out(wire_d34_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353454(.data_in(wire_d34_53),.data_out(wire_d34_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353455(.data_in(wire_d34_54),.data_out(wire_d34_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353456(.data_in(wire_d34_55),.data_out(wire_d34_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353457(.data_in(wire_d34_56),.data_out(wire_d34_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353458(.data_in(wire_d34_57),.data_out(wire_d34_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353459(.data_in(wire_d34_58),.data_out(wire_d34_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353460(.data_in(wire_d34_59),.data_out(wire_d34_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353461(.data_in(wire_d34_60),.data_out(wire_d34_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353462(.data_in(wire_d34_61),.data_out(wire_d34_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance353463(.data_in(wire_d34_62),.data_out(wire_d34_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353464(.data_in(wire_d34_63),.data_out(wire_d34_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance353465(.data_in(wire_d34_64),.data_out(wire_d34_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance353466(.data_in(wire_d34_65),.data_out(wire_d34_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353467(.data_in(wire_d34_66),.data_out(wire_d34_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353468(.data_in(wire_d34_67),.data_out(wire_d34_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance353469(.data_in(wire_d34_68),.data_out(d_out34),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance36350(.data_in(d_in35),.data_out(wire_d35_0),.clk(clk),.rst(rst));            //channel 36
	encoder #(.WIDTH(WIDTH)) encoder_instance36351(.data_in(wire_d35_0),.data_out(wire_d35_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance36352(.data_in(wire_d35_1),.data_out(wire_d35_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance36353(.data_in(wire_d35_2),.data_out(wire_d35_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance36354(.data_in(wire_d35_3),.data_out(wire_d35_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance36355(.data_in(wire_d35_4),.data_out(wire_d35_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance36356(.data_in(wire_d35_5),.data_out(wire_d35_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance36357(.data_in(wire_d35_6),.data_out(wire_d35_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance36358(.data_in(wire_d35_7),.data_out(wire_d35_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance36359(.data_in(wire_d35_8),.data_out(wire_d35_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363510(.data_in(wire_d35_9),.data_out(wire_d35_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363511(.data_in(wire_d35_10),.data_out(wire_d35_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363512(.data_in(wire_d35_11),.data_out(wire_d35_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363513(.data_in(wire_d35_12),.data_out(wire_d35_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363514(.data_in(wire_d35_13),.data_out(wire_d35_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363515(.data_in(wire_d35_14),.data_out(wire_d35_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363516(.data_in(wire_d35_15),.data_out(wire_d35_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363517(.data_in(wire_d35_16),.data_out(wire_d35_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363518(.data_in(wire_d35_17),.data_out(wire_d35_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363519(.data_in(wire_d35_18),.data_out(wire_d35_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363520(.data_in(wire_d35_19),.data_out(wire_d35_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363521(.data_in(wire_d35_20),.data_out(wire_d35_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363522(.data_in(wire_d35_21),.data_out(wire_d35_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363523(.data_in(wire_d35_22),.data_out(wire_d35_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363524(.data_in(wire_d35_23),.data_out(wire_d35_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363525(.data_in(wire_d35_24),.data_out(wire_d35_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363526(.data_in(wire_d35_25),.data_out(wire_d35_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363527(.data_in(wire_d35_26),.data_out(wire_d35_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363528(.data_in(wire_d35_27),.data_out(wire_d35_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363529(.data_in(wire_d35_28),.data_out(wire_d35_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363530(.data_in(wire_d35_29),.data_out(wire_d35_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363531(.data_in(wire_d35_30),.data_out(wire_d35_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363532(.data_in(wire_d35_31),.data_out(wire_d35_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363533(.data_in(wire_d35_32),.data_out(wire_d35_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363534(.data_in(wire_d35_33),.data_out(wire_d35_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363535(.data_in(wire_d35_34),.data_out(wire_d35_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363536(.data_in(wire_d35_35),.data_out(wire_d35_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363537(.data_in(wire_d35_36),.data_out(wire_d35_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363538(.data_in(wire_d35_37),.data_out(wire_d35_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363539(.data_in(wire_d35_38),.data_out(wire_d35_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363540(.data_in(wire_d35_39),.data_out(wire_d35_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363541(.data_in(wire_d35_40),.data_out(wire_d35_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363542(.data_in(wire_d35_41),.data_out(wire_d35_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363543(.data_in(wire_d35_42),.data_out(wire_d35_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363544(.data_in(wire_d35_43),.data_out(wire_d35_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363545(.data_in(wire_d35_44),.data_out(wire_d35_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363546(.data_in(wire_d35_45),.data_out(wire_d35_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363547(.data_in(wire_d35_46),.data_out(wire_d35_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363548(.data_in(wire_d35_47),.data_out(wire_d35_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363549(.data_in(wire_d35_48),.data_out(wire_d35_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363550(.data_in(wire_d35_49),.data_out(wire_d35_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363551(.data_in(wire_d35_50),.data_out(wire_d35_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363552(.data_in(wire_d35_51),.data_out(wire_d35_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363553(.data_in(wire_d35_52),.data_out(wire_d35_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363554(.data_in(wire_d35_53),.data_out(wire_d35_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363555(.data_in(wire_d35_54),.data_out(wire_d35_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363556(.data_in(wire_d35_55),.data_out(wire_d35_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363557(.data_in(wire_d35_56),.data_out(wire_d35_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363558(.data_in(wire_d35_57),.data_out(wire_d35_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363559(.data_in(wire_d35_58),.data_out(wire_d35_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363560(.data_in(wire_d35_59),.data_out(wire_d35_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363561(.data_in(wire_d35_60),.data_out(wire_d35_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance363562(.data_in(wire_d35_61),.data_out(wire_d35_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363563(.data_in(wire_d35_62),.data_out(wire_d35_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363564(.data_in(wire_d35_63),.data_out(wire_d35_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363565(.data_in(wire_d35_64),.data_out(wire_d35_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance363566(.data_in(wire_d35_65),.data_out(wire_d35_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363567(.data_in(wire_d35_66),.data_out(wire_d35_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance363568(.data_in(wire_d35_67),.data_out(wire_d35_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance363569(.data_in(wire_d35_68),.data_out(d_out35),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance37360(.data_in(d_in36),.data_out(wire_d36_0),.clk(clk),.rst(rst));            //channel 37
	encoder #(.WIDTH(WIDTH)) encoder_instance37361(.data_in(wire_d36_0),.data_out(wire_d36_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance37362(.data_in(wire_d36_1),.data_out(wire_d36_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance37363(.data_in(wire_d36_2),.data_out(wire_d36_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance37364(.data_in(wire_d36_3),.data_out(wire_d36_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance37365(.data_in(wire_d36_4),.data_out(wire_d36_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance37366(.data_in(wire_d36_5),.data_out(wire_d36_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance37367(.data_in(wire_d36_6),.data_out(wire_d36_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance37368(.data_in(wire_d36_7),.data_out(wire_d36_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance37369(.data_in(wire_d36_8),.data_out(wire_d36_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373610(.data_in(wire_d36_9),.data_out(wire_d36_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373611(.data_in(wire_d36_10),.data_out(wire_d36_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373612(.data_in(wire_d36_11),.data_out(wire_d36_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373613(.data_in(wire_d36_12),.data_out(wire_d36_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373614(.data_in(wire_d36_13),.data_out(wire_d36_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373615(.data_in(wire_d36_14),.data_out(wire_d36_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373616(.data_in(wire_d36_15),.data_out(wire_d36_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373617(.data_in(wire_d36_16),.data_out(wire_d36_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373618(.data_in(wire_d36_17),.data_out(wire_d36_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373619(.data_in(wire_d36_18),.data_out(wire_d36_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373620(.data_in(wire_d36_19),.data_out(wire_d36_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373621(.data_in(wire_d36_20),.data_out(wire_d36_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373622(.data_in(wire_d36_21),.data_out(wire_d36_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373623(.data_in(wire_d36_22),.data_out(wire_d36_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373624(.data_in(wire_d36_23),.data_out(wire_d36_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373625(.data_in(wire_d36_24),.data_out(wire_d36_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373626(.data_in(wire_d36_25),.data_out(wire_d36_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373627(.data_in(wire_d36_26),.data_out(wire_d36_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373628(.data_in(wire_d36_27),.data_out(wire_d36_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373629(.data_in(wire_d36_28),.data_out(wire_d36_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373630(.data_in(wire_d36_29),.data_out(wire_d36_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373631(.data_in(wire_d36_30),.data_out(wire_d36_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373632(.data_in(wire_d36_31),.data_out(wire_d36_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373633(.data_in(wire_d36_32),.data_out(wire_d36_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373634(.data_in(wire_d36_33),.data_out(wire_d36_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373635(.data_in(wire_d36_34),.data_out(wire_d36_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373636(.data_in(wire_d36_35),.data_out(wire_d36_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373637(.data_in(wire_d36_36),.data_out(wire_d36_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373638(.data_in(wire_d36_37),.data_out(wire_d36_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373639(.data_in(wire_d36_38),.data_out(wire_d36_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373640(.data_in(wire_d36_39),.data_out(wire_d36_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373641(.data_in(wire_d36_40),.data_out(wire_d36_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373642(.data_in(wire_d36_41),.data_out(wire_d36_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373643(.data_in(wire_d36_42),.data_out(wire_d36_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373644(.data_in(wire_d36_43),.data_out(wire_d36_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373645(.data_in(wire_d36_44),.data_out(wire_d36_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373646(.data_in(wire_d36_45),.data_out(wire_d36_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373647(.data_in(wire_d36_46),.data_out(wire_d36_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373648(.data_in(wire_d36_47),.data_out(wire_d36_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373649(.data_in(wire_d36_48),.data_out(wire_d36_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373650(.data_in(wire_d36_49),.data_out(wire_d36_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373651(.data_in(wire_d36_50),.data_out(wire_d36_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373652(.data_in(wire_d36_51),.data_out(wire_d36_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373653(.data_in(wire_d36_52),.data_out(wire_d36_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373654(.data_in(wire_d36_53),.data_out(wire_d36_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373655(.data_in(wire_d36_54),.data_out(wire_d36_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373656(.data_in(wire_d36_55),.data_out(wire_d36_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373657(.data_in(wire_d36_56),.data_out(wire_d36_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance373658(.data_in(wire_d36_57),.data_out(wire_d36_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373659(.data_in(wire_d36_58),.data_out(wire_d36_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373660(.data_in(wire_d36_59),.data_out(wire_d36_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373661(.data_in(wire_d36_60),.data_out(wire_d36_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373662(.data_in(wire_d36_61),.data_out(wire_d36_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373663(.data_in(wire_d36_62),.data_out(wire_d36_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373664(.data_in(wire_d36_63),.data_out(wire_d36_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance373665(.data_in(wire_d36_64),.data_out(wire_d36_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373666(.data_in(wire_d36_65),.data_out(wire_d36_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373667(.data_in(wire_d36_66),.data_out(wire_d36_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance373668(.data_in(wire_d36_67),.data_out(wire_d36_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance373669(.data_in(wire_d36_68),.data_out(d_out36),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance38370(.data_in(d_in37),.data_out(wire_d37_0),.clk(clk),.rst(rst));            //channel 38
	encoder #(.WIDTH(WIDTH)) encoder_instance38371(.data_in(wire_d37_0),.data_out(wire_d37_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance38372(.data_in(wire_d37_1),.data_out(wire_d37_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance38373(.data_in(wire_d37_2),.data_out(wire_d37_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance38374(.data_in(wire_d37_3),.data_out(wire_d37_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance38375(.data_in(wire_d37_4),.data_out(wire_d37_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance38376(.data_in(wire_d37_5),.data_out(wire_d37_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance38377(.data_in(wire_d37_6),.data_out(wire_d37_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance38378(.data_in(wire_d37_7),.data_out(wire_d37_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance38379(.data_in(wire_d37_8),.data_out(wire_d37_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383710(.data_in(wire_d37_9),.data_out(wire_d37_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383711(.data_in(wire_d37_10),.data_out(wire_d37_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383712(.data_in(wire_d37_11),.data_out(wire_d37_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383713(.data_in(wire_d37_12),.data_out(wire_d37_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383714(.data_in(wire_d37_13),.data_out(wire_d37_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383715(.data_in(wire_d37_14),.data_out(wire_d37_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383716(.data_in(wire_d37_15),.data_out(wire_d37_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383717(.data_in(wire_d37_16),.data_out(wire_d37_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383718(.data_in(wire_d37_17),.data_out(wire_d37_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383719(.data_in(wire_d37_18),.data_out(wire_d37_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383720(.data_in(wire_d37_19),.data_out(wire_d37_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383721(.data_in(wire_d37_20),.data_out(wire_d37_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383722(.data_in(wire_d37_21),.data_out(wire_d37_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383723(.data_in(wire_d37_22),.data_out(wire_d37_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383724(.data_in(wire_d37_23),.data_out(wire_d37_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383725(.data_in(wire_d37_24),.data_out(wire_d37_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383726(.data_in(wire_d37_25),.data_out(wire_d37_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383727(.data_in(wire_d37_26),.data_out(wire_d37_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383728(.data_in(wire_d37_27),.data_out(wire_d37_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383729(.data_in(wire_d37_28),.data_out(wire_d37_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383730(.data_in(wire_d37_29),.data_out(wire_d37_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383731(.data_in(wire_d37_30),.data_out(wire_d37_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383732(.data_in(wire_d37_31),.data_out(wire_d37_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383733(.data_in(wire_d37_32),.data_out(wire_d37_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383734(.data_in(wire_d37_33),.data_out(wire_d37_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383735(.data_in(wire_d37_34),.data_out(wire_d37_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383736(.data_in(wire_d37_35),.data_out(wire_d37_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383737(.data_in(wire_d37_36),.data_out(wire_d37_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383738(.data_in(wire_d37_37),.data_out(wire_d37_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383739(.data_in(wire_d37_38),.data_out(wire_d37_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383740(.data_in(wire_d37_39),.data_out(wire_d37_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383741(.data_in(wire_d37_40),.data_out(wire_d37_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383742(.data_in(wire_d37_41),.data_out(wire_d37_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383743(.data_in(wire_d37_42),.data_out(wire_d37_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383744(.data_in(wire_d37_43),.data_out(wire_d37_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383745(.data_in(wire_d37_44),.data_out(wire_d37_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383746(.data_in(wire_d37_45),.data_out(wire_d37_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383747(.data_in(wire_d37_46),.data_out(wire_d37_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383748(.data_in(wire_d37_47),.data_out(wire_d37_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383749(.data_in(wire_d37_48),.data_out(wire_d37_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383750(.data_in(wire_d37_49),.data_out(wire_d37_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383751(.data_in(wire_d37_50),.data_out(wire_d37_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383752(.data_in(wire_d37_51),.data_out(wire_d37_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383753(.data_in(wire_d37_52),.data_out(wire_d37_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383754(.data_in(wire_d37_53),.data_out(wire_d37_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383755(.data_in(wire_d37_54),.data_out(wire_d37_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383756(.data_in(wire_d37_55),.data_out(wire_d37_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383757(.data_in(wire_d37_56),.data_out(wire_d37_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383758(.data_in(wire_d37_57),.data_out(wire_d37_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383759(.data_in(wire_d37_58),.data_out(wire_d37_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383760(.data_in(wire_d37_59),.data_out(wire_d37_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance383761(.data_in(wire_d37_60),.data_out(wire_d37_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383762(.data_in(wire_d37_61),.data_out(wire_d37_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383763(.data_in(wire_d37_62),.data_out(wire_d37_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance383764(.data_in(wire_d37_63),.data_out(wire_d37_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383765(.data_in(wire_d37_64),.data_out(wire_d37_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383766(.data_in(wire_d37_65),.data_out(wire_d37_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383767(.data_in(wire_d37_66),.data_out(wire_d37_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance383768(.data_in(wire_d37_67),.data_out(wire_d37_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance383769(.data_in(wire_d37_68),.data_out(d_out37),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance39380(.data_in(d_in38),.data_out(wire_d38_0),.clk(clk),.rst(rst));            //channel 39
	invertion #(.WIDTH(WIDTH)) invertion_instance39381(.data_in(wire_d38_0),.data_out(wire_d38_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance39382(.data_in(wire_d38_1),.data_out(wire_d38_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance39383(.data_in(wire_d38_2),.data_out(wire_d38_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance39384(.data_in(wire_d38_3),.data_out(wire_d38_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance39385(.data_in(wire_d38_4),.data_out(wire_d38_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance39386(.data_in(wire_d38_5),.data_out(wire_d38_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance39387(.data_in(wire_d38_6),.data_out(wire_d38_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance39388(.data_in(wire_d38_7),.data_out(wire_d38_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance39389(.data_in(wire_d38_8),.data_out(wire_d38_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393810(.data_in(wire_d38_9),.data_out(wire_d38_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393811(.data_in(wire_d38_10),.data_out(wire_d38_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393812(.data_in(wire_d38_11),.data_out(wire_d38_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393813(.data_in(wire_d38_12),.data_out(wire_d38_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393814(.data_in(wire_d38_13),.data_out(wire_d38_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393815(.data_in(wire_d38_14),.data_out(wire_d38_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393816(.data_in(wire_d38_15),.data_out(wire_d38_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393817(.data_in(wire_d38_16),.data_out(wire_d38_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393818(.data_in(wire_d38_17),.data_out(wire_d38_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393819(.data_in(wire_d38_18),.data_out(wire_d38_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393820(.data_in(wire_d38_19),.data_out(wire_d38_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393821(.data_in(wire_d38_20),.data_out(wire_d38_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393822(.data_in(wire_d38_21),.data_out(wire_d38_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393823(.data_in(wire_d38_22),.data_out(wire_d38_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393824(.data_in(wire_d38_23),.data_out(wire_d38_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393825(.data_in(wire_d38_24),.data_out(wire_d38_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393826(.data_in(wire_d38_25),.data_out(wire_d38_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393827(.data_in(wire_d38_26),.data_out(wire_d38_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393828(.data_in(wire_d38_27),.data_out(wire_d38_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393829(.data_in(wire_d38_28),.data_out(wire_d38_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393830(.data_in(wire_d38_29),.data_out(wire_d38_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393831(.data_in(wire_d38_30),.data_out(wire_d38_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393832(.data_in(wire_d38_31),.data_out(wire_d38_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393833(.data_in(wire_d38_32),.data_out(wire_d38_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393834(.data_in(wire_d38_33),.data_out(wire_d38_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393835(.data_in(wire_d38_34),.data_out(wire_d38_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393836(.data_in(wire_d38_35),.data_out(wire_d38_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393837(.data_in(wire_d38_36),.data_out(wire_d38_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393838(.data_in(wire_d38_37),.data_out(wire_d38_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393839(.data_in(wire_d38_38),.data_out(wire_d38_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393840(.data_in(wire_d38_39),.data_out(wire_d38_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393841(.data_in(wire_d38_40),.data_out(wire_d38_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393842(.data_in(wire_d38_41),.data_out(wire_d38_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393843(.data_in(wire_d38_42),.data_out(wire_d38_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393844(.data_in(wire_d38_43),.data_out(wire_d38_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393845(.data_in(wire_d38_44),.data_out(wire_d38_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393846(.data_in(wire_d38_45),.data_out(wire_d38_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393847(.data_in(wire_d38_46),.data_out(wire_d38_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393848(.data_in(wire_d38_47),.data_out(wire_d38_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393849(.data_in(wire_d38_48),.data_out(wire_d38_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393850(.data_in(wire_d38_49),.data_out(wire_d38_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393851(.data_in(wire_d38_50),.data_out(wire_d38_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393852(.data_in(wire_d38_51),.data_out(wire_d38_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393853(.data_in(wire_d38_52),.data_out(wire_d38_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393854(.data_in(wire_d38_53),.data_out(wire_d38_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393855(.data_in(wire_d38_54),.data_out(wire_d38_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance393856(.data_in(wire_d38_55),.data_out(wire_d38_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393857(.data_in(wire_d38_56),.data_out(wire_d38_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393858(.data_in(wire_d38_57),.data_out(wire_d38_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393859(.data_in(wire_d38_58),.data_out(wire_d38_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393860(.data_in(wire_d38_59),.data_out(wire_d38_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393861(.data_in(wire_d38_60),.data_out(wire_d38_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393862(.data_in(wire_d38_61),.data_out(wire_d38_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance393863(.data_in(wire_d38_62),.data_out(wire_d38_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393864(.data_in(wire_d38_63),.data_out(wire_d38_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393865(.data_in(wire_d38_64),.data_out(wire_d38_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393866(.data_in(wire_d38_65),.data_out(wire_d38_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393867(.data_in(wire_d38_66),.data_out(wire_d38_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance393868(.data_in(wire_d38_67),.data_out(wire_d38_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance393869(.data_in(wire_d38_68),.data_out(d_out38),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance40390(.data_in(d_in39),.data_out(wire_d39_0),.clk(clk),.rst(rst));            //channel 40
	encoder #(.WIDTH(WIDTH)) encoder_instance40391(.data_in(wire_d39_0),.data_out(wire_d39_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance40392(.data_in(wire_d39_1),.data_out(wire_d39_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance40393(.data_in(wire_d39_2),.data_out(wire_d39_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance40394(.data_in(wire_d39_3),.data_out(wire_d39_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance40395(.data_in(wire_d39_4),.data_out(wire_d39_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance40396(.data_in(wire_d39_5),.data_out(wire_d39_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance40397(.data_in(wire_d39_6),.data_out(wire_d39_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance40398(.data_in(wire_d39_7),.data_out(wire_d39_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance40399(.data_in(wire_d39_8),.data_out(wire_d39_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403910(.data_in(wire_d39_9),.data_out(wire_d39_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403911(.data_in(wire_d39_10),.data_out(wire_d39_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403912(.data_in(wire_d39_11),.data_out(wire_d39_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403913(.data_in(wire_d39_12),.data_out(wire_d39_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403914(.data_in(wire_d39_13),.data_out(wire_d39_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403915(.data_in(wire_d39_14),.data_out(wire_d39_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403916(.data_in(wire_d39_15),.data_out(wire_d39_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403917(.data_in(wire_d39_16),.data_out(wire_d39_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403918(.data_in(wire_d39_17),.data_out(wire_d39_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403919(.data_in(wire_d39_18),.data_out(wire_d39_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403920(.data_in(wire_d39_19),.data_out(wire_d39_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403921(.data_in(wire_d39_20),.data_out(wire_d39_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403922(.data_in(wire_d39_21),.data_out(wire_d39_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403923(.data_in(wire_d39_22),.data_out(wire_d39_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403924(.data_in(wire_d39_23),.data_out(wire_d39_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403925(.data_in(wire_d39_24),.data_out(wire_d39_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403926(.data_in(wire_d39_25),.data_out(wire_d39_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403927(.data_in(wire_d39_26),.data_out(wire_d39_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403928(.data_in(wire_d39_27),.data_out(wire_d39_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403929(.data_in(wire_d39_28),.data_out(wire_d39_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403930(.data_in(wire_d39_29),.data_out(wire_d39_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403931(.data_in(wire_d39_30),.data_out(wire_d39_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403932(.data_in(wire_d39_31),.data_out(wire_d39_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403933(.data_in(wire_d39_32),.data_out(wire_d39_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403934(.data_in(wire_d39_33),.data_out(wire_d39_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403935(.data_in(wire_d39_34),.data_out(wire_d39_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403936(.data_in(wire_d39_35),.data_out(wire_d39_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403937(.data_in(wire_d39_36),.data_out(wire_d39_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403938(.data_in(wire_d39_37),.data_out(wire_d39_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403939(.data_in(wire_d39_38),.data_out(wire_d39_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403940(.data_in(wire_d39_39),.data_out(wire_d39_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403941(.data_in(wire_d39_40),.data_out(wire_d39_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403942(.data_in(wire_d39_41),.data_out(wire_d39_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403943(.data_in(wire_d39_42),.data_out(wire_d39_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403944(.data_in(wire_d39_43),.data_out(wire_d39_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403945(.data_in(wire_d39_44),.data_out(wire_d39_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403946(.data_in(wire_d39_45),.data_out(wire_d39_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403947(.data_in(wire_d39_46),.data_out(wire_d39_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403948(.data_in(wire_d39_47),.data_out(wire_d39_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403949(.data_in(wire_d39_48),.data_out(wire_d39_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403950(.data_in(wire_d39_49),.data_out(wire_d39_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403951(.data_in(wire_d39_50),.data_out(wire_d39_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403952(.data_in(wire_d39_51),.data_out(wire_d39_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403953(.data_in(wire_d39_52),.data_out(wire_d39_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403954(.data_in(wire_d39_53),.data_out(wire_d39_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403955(.data_in(wire_d39_54),.data_out(wire_d39_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403956(.data_in(wire_d39_55),.data_out(wire_d39_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403957(.data_in(wire_d39_56),.data_out(wire_d39_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403958(.data_in(wire_d39_57),.data_out(wire_d39_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403959(.data_in(wire_d39_58),.data_out(wire_d39_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403960(.data_in(wire_d39_59),.data_out(wire_d39_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403961(.data_in(wire_d39_60),.data_out(wire_d39_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403962(.data_in(wire_d39_61),.data_out(wire_d39_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance403963(.data_in(wire_d39_62),.data_out(wire_d39_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance403964(.data_in(wire_d39_63),.data_out(wire_d39_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403965(.data_in(wire_d39_64),.data_out(wire_d39_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403966(.data_in(wire_d39_65),.data_out(wire_d39_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403967(.data_in(wire_d39_66),.data_out(wire_d39_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance403968(.data_in(wire_d39_67),.data_out(wire_d39_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance403969(.data_in(wire_d39_68),.data_out(d_out39),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance41400(.data_in(d_in40),.data_out(wire_d40_0),.clk(clk),.rst(rst));            //channel 41
	invertion #(.WIDTH(WIDTH)) invertion_instance41401(.data_in(wire_d40_0),.data_out(wire_d40_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance41402(.data_in(wire_d40_1),.data_out(wire_d40_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance41403(.data_in(wire_d40_2),.data_out(wire_d40_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance41404(.data_in(wire_d40_3),.data_out(wire_d40_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance41405(.data_in(wire_d40_4),.data_out(wire_d40_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance41406(.data_in(wire_d40_5),.data_out(wire_d40_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance41407(.data_in(wire_d40_6),.data_out(wire_d40_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance41408(.data_in(wire_d40_7),.data_out(wire_d40_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance41409(.data_in(wire_d40_8),.data_out(wire_d40_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414010(.data_in(wire_d40_9),.data_out(wire_d40_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414011(.data_in(wire_d40_10),.data_out(wire_d40_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414012(.data_in(wire_d40_11),.data_out(wire_d40_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414013(.data_in(wire_d40_12),.data_out(wire_d40_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414014(.data_in(wire_d40_13),.data_out(wire_d40_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414015(.data_in(wire_d40_14),.data_out(wire_d40_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414016(.data_in(wire_d40_15),.data_out(wire_d40_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414017(.data_in(wire_d40_16),.data_out(wire_d40_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414018(.data_in(wire_d40_17),.data_out(wire_d40_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414019(.data_in(wire_d40_18),.data_out(wire_d40_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414020(.data_in(wire_d40_19),.data_out(wire_d40_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414021(.data_in(wire_d40_20),.data_out(wire_d40_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414022(.data_in(wire_d40_21),.data_out(wire_d40_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414023(.data_in(wire_d40_22),.data_out(wire_d40_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414024(.data_in(wire_d40_23),.data_out(wire_d40_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414025(.data_in(wire_d40_24),.data_out(wire_d40_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414026(.data_in(wire_d40_25),.data_out(wire_d40_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414027(.data_in(wire_d40_26),.data_out(wire_d40_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414028(.data_in(wire_d40_27),.data_out(wire_d40_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414029(.data_in(wire_d40_28),.data_out(wire_d40_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414030(.data_in(wire_d40_29),.data_out(wire_d40_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414031(.data_in(wire_d40_30),.data_out(wire_d40_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414032(.data_in(wire_d40_31),.data_out(wire_d40_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414033(.data_in(wire_d40_32),.data_out(wire_d40_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414034(.data_in(wire_d40_33),.data_out(wire_d40_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414035(.data_in(wire_d40_34),.data_out(wire_d40_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414036(.data_in(wire_d40_35),.data_out(wire_d40_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414037(.data_in(wire_d40_36),.data_out(wire_d40_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414038(.data_in(wire_d40_37),.data_out(wire_d40_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414039(.data_in(wire_d40_38),.data_out(wire_d40_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414040(.data_in(wire_d40_39),.data_out(wire_d40_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414041(.data_in(wire_d40_40),.data_out(wire_d40_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414042(.data_in(wire_d40_41),.data_out(wire_d40_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414043(.data_in(wire_d40_42),.data_out(wire_d40_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414044(.data_in(wire_d40_43),.data_out(wire_d40_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414045(.data_in(wire_d40_44),.data_out(wire_d40_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414046(.data_in(wire_d40_45),.data_out(wire_d40_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414047(.data_in(wire_d40_46),.data_out(wire_d40_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414048(.data_in(wire_d40_47),.data_out(wire_d40_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414049(.data_in(wire_d40_48),.data_out(wire_d40_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414050(.data_in(wire_d40_49),.data_out(wire_d40_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414051(.data_in(wire_d40_50),.data_out(wire_d40_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414052(.data_in(wire_d40_51),.data_out(wire_d40_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414053(.data_in(wire_d40_52),.data_out(wire_d40_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414054(.data_in(wire_d40_53),.data_out(wire_d40_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414055(.data_in(wire_d40_54),.data_out(wire_d40_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414056(.data_in(wire_d40_55),.data_out(wire_d40_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414057(.data_in(wire_d40_56),.data_out(wire_d40_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414058(.data_in(wire_d40_57),.data_out(wire_d40_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414059(.data_in(wire_d40_58),.data_out(wire_d40_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414060(.data_in(wire_d40_59),.data_out(wire_d40_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414061(.data_in(wire_d40_60),.data_out(wire_d40_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414062(.data_in(wire_d40_61),.data_out(wire_d40_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance414063(.data_in(wire_d40_62),.data_out(wire_d40_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414064(.data_in(wire_d40_63),.data_out(wire_d40_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance414065(.data_in(wire_d40_64),.data_out(wire_d40_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414066(.data_in(wire_d40_65),.data_out(wire_d40_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414067(.data_in(wire_d40_66),.data_out(wire_d40_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance414068(.data_in(wire_d40_67),.data_out(wire_d40_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance414069(.data_in(wire_d40_68),.data_out(d_out40),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance42410(.data_in(d_in41),.data_out(wire_d41_0),.clk(clk),.rst(rst));            //channel 42
	invertion #(.WIDTH(WIDTH)) invertion_instance42411(.data_in(wire_d41_0),.data_out(wire_d41_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance42412(.data_in(wire_d41_1),.data_out(wire_d41_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance42413(.data_in(wire_d41_2),.data_out(wire_d41_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance42414(.data_in(wire_d41_3),.data_out(wire_d41_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance42415(.data_in(wire_d41_4),.data_out(wire_d41_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance42416(.data_in(wire_d41_5),.data_out(wire_d41_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance42417(.data_in(wire_d41_6),.data_out(wire_d41_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance42418(.data_in(wire_d41_7),.data_out(wire_d41_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance42419(.data_in(wire_d41_8),.data_out(wire_d41_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424110(.data_in(wire_d41_9),.data_out(wire_d41_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424111(.data_in(wire_d41_10),.data_out(wire_d41_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424112(.data_in(wire_d41_11),.data_out(wire_d41_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424113(.data_in(wire_d41_12),.data_out(wire_d41_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424114(.data_in(wire_d41_13),.data_out(wire_d41_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424115(.data_in(wire_d41_14),.data_out(wire_d41_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424116(.data_in(wire_d41_15),.data_out(wire_d41_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424117(.data_in(wire_d41_16),.data_out(wire_d41_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424118(.data_in(wire_d41_17),.data_out(wire_d41_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424119(.data_in(wire_d41_18),.data_out(wire_d41_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424120(.data_in(wire_d41_19),.data_out(wire_d41_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424121(.data_in(wire_d41_20),.data_out(wire_d41_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424122(.data_in(wire_d41_21),.data_out(wire_d41_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424123(.data_in(wire_d41_22),.data_out(wire_d41_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424124(.data_in(wire_d41_23),.data_out(wire_d41_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424125(.data_in(wire_d41_24),.data_out(wire_d41_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424126(.data_in(wire_d41_25),.data_out(wire_d41_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424127(.data_in(wire_d41_26),.data_out(wire_d41_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424128(.data_in(wire_d41_27),.data_out(wire_d41_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424129(.data_in(wire_d41_28),.data_out(wire_d41_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424130(.data_in(wire_d41_29),.data_out(wire_d41_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424131(.data_in(wire_d41_30),.data_out(wire_d41_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424132(.data_in(wire_d41_31),.data_out(wire_d41_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424133(.data_in(wire_d41_32),.data_out(wire_d41_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424134(.data_in(wire_d41_33),.data_out(wire_d41_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424135(.data_in(wire_d41_34),.data_out(wire_d41_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424136(.data_in(wire_d41_35),.data_out(wire_d41_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424137(.data_in(wire_d41_36),.data_out(wire_d41_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424138(.data_in(wire_d41_37),.data_out(wire_d41_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424139(.data_in(wire_d41_38),.data_out(wire_d41_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424140(.data_in(wire_d41_39),.data_out(wire_d41_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424141(.data_in(wire_d41_40),.data_out(wire_d41_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424142(.data_in(wire_d41_41),.data_out(wire_d41_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424143(.data_in(wire_d41_42),.data_out(wire_d41_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424144(.data_in(wire_d41_43),.data_out(wire_d41_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424145(.data_in(wire_d41_44),.data_out(wire_d41_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424146(.data_in(wire_d41_45),.data_out(wire_d41_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424147(.data_in(wire_d41_46),.data_out(wire_d41_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424148(.data_in(wire_d41_47),.data_out(wire_d41_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424149(.data_in(wire_d41_48),.data_out(wire_d41_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424150(.data_in(wire_d41_49),.data_out(wire_d41_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424151(.data_in(wire_d41_50),.data_out(wire_d41_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424152(.data_in(wire_d41_51),.data_out(wire_d41_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424153(.data_in(wire_d41_52),.data_out(wire_d41_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424154(.data_in(wire_d41_53),.data_out(wire_d41_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424155(.data_in(wire_d41_54),.data_out(wire_d41_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance424156(.data_in(wire_d41_55),.data_out(wire_d41_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424157(.data_in(wire_d41_56),.data_out(wire_d41_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424158(.data_in(wire_d41_57),.data_out(wire_d41_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424159(.data_in(wire_d41_58),.data_out(wire_d41_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424160(.data_in(wire_d41_59),.data_out(wire_d41_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424161(.data_in(wire_d41_60),.data_out(wire_d41_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424162(.data_in(wire_d41_61),.data_out(wire_d41_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424163(.data_in(wire_d41_62),.data_out(wire_d41_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance424164(.data_in(wire_d41_63),.data_out(wire_d41_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424165(.data_in(wire_d41_64),.data_out(wire_d41_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424166(.data_in(wire_d41_65),.data_out(wire_d41_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424167(.data_in(wire_d41_66),.data_out(wire_d41_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance424168(.data_in(wire_d41_67),.data_out(wire_d41_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance424169(.data_in(wire_d41_68),.data_out(d_out41),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance43420(.data_in(d_in42),.data_out(wire_d42_0),.clk(clk),.rst(rst));            //channel 43
	invertion #(.WIDTH(WIDTH)) invertion_instance43421(.data_in(wire_d42_0),.data_out(wire_d42_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance43422(.data_in(wire_d42_1),.data_out(wire_d42_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance43423(.data_in(wire_d42_2),.data_out(wire_d42_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance43424(.data_in(wire_d42_3),.data_out(wire_d42_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance43425(.data_in(wire_d42_4),.data_out(wire_d42_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance43426(.data_in(wire_d42_5),.data_out(wire_d42_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance43427(.data_in(wire_d42_6),.data_out(wire_d42_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance43428(.data_in(wire_d42_7),.data_out(wire_d42_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43429(.data_in(wire_d42_8),.data_out(wire_d42_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434210(.data_in(wire_d42_9),.data_out(wire_d42_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434211(.data_in(wire_d42_10),.data_out(wire_d42_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434212(.data_in(wire_d42_11),.data_out(wire_d42_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434213(.data_in(wire_d42_12),.data_out(wire_d42_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434214(.data_in(wire_d42_13),.data_out(wire_d42_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434215(.data_in(wire_d42_14),.data_out(wire_d42_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434216(.data_in(wire_d42_15),.data_out(wire_d42_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434217(.data_in(wire_d42_16),.data_out(wire_d42_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434218(.data_in(wire_d42_17),.data_out(wire_d42_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434219(.data_in(wire_d42_18),.data_out(wire_d42_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434220(.data_in(wire_d42_19),.data_out(wire_d42_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434221(.data_in(wire_d42_20),.data_out(wire_d42_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434222(.data_in(wire_d42_21),.data_out(wire_d42_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434223(.data_in(wire_d42_22),.data_out(wire_d42_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434224(.data_in(wire_d42_23),.data_out(wire_d42_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434225(.data_in(wire_d42_24),.data_out(wire_d42_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434226(.data_in(wire_d42_25),.data_out(wire_d42_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434227(.data_in(wire_d42_26),.data_out(wire_d42_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434228(.data_in(wire_d42_27),.data_out(wire_d42_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434229(.data_in(wire_d42_28),.data_out(wire_d42_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434230(.data_in(wire_d42_29),.data_out(wire_d42_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434231(.data_in(wire_d42_30),.data_out(wire_d42_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434232(.data_in(wire_d42_31),.data_out(wire_d42_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434233(.data_in(wire_d42_32),.data_out(wire_d42_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434234(.data_in(wire_d42_33),.data_out(wire_d42_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434235(.data_in(wire_d42_34),.data_out(wire_d42_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434236(.data_in(wire_d42_35),.data_out(wire_d42_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434237(.data_in(wire_d42_36),.data_out(wire_d42_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434238(.data_in(wire_d42_37),.data_out(wire_d42_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434239(.data_in(wire_d42_38),.data_out(wire_d42_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434240(.data_in(wire_d42_39),.data_out(wire_d42_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434241(.data_in(wire_d42_40),.data_out(wire_d42_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434242(.data_in(wire_d42_41),.data_out(wire_d42_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434243(.data_in(wire_d42_42),.data_out(wire_d42_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434244(.data_in(wire_d42_43),.data_out(wire_d42_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434245(.data_in(wire_d42_44),.data_out(wire_d42_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434246(.data_in(wire_d42_45),.data_out(wire_d42_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434247(.data_in(wire_d42_46),.data_out(wire_d42_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434248(.data_in(wire_d42_47),.data_out(wire_d42_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434249(.data_in(wire_d42_48),.data_out(wire_d42_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434250(.data_in(wire_d42_49),.data_out(wire_d42_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434251(.data_in(wire_d42_50),.data_out(wire_d42_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434252(.data_in(wire_d42_51),.data_out(wire_d42_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434253(.data_in(wire_d42_52),.data_out(wire_d42_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434254(.data_in(wire_d42_53),.data_out(wire_d42_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434255(.data_in(wire_d42_54),.data_out(wire_d42_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434256(.data_in(wire_d42_55),.data_out(wire_d42_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434257(.data_in(wire_d42_56),.data_out(wire_d42_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434258(.data_in(wire_d42_57),.data_out(wire_d42_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434259(.data_in(wire_d42_58),.data_out(wire_d42_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434260(.data_in(wire_d42_59),.data_out(wire_d42_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434261(.data_in(wire_d42_60),.data_out(wire_d42_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434262(.data_in(wire_d42_61),.data_out(wire_d42_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434263(.data_in(wire_d42_62),.data_out(wire_d42_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434264(.data_in(wire_d42_63),.data_out(wire_d42_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434265(.data_in(wire_d42_64),.data_out(wire_d42_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance434266(.data_in(wire_d42_65),.data_out(wire_d42_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434267(.data_in(wire_d42_66),.data_out(wire_d42_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance434268(.data_in(wire_d42_67),.data_out(wire_d42_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434269(.data_in(wire_d42_68),.data_out(d_out42),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance44430(.data_in(d_in43),.data_out(wire_d43_0),.clk(clk),.rst(rst));            //channel 44
	encoder #(.WIDTH(WIDTH)) encoder_instance44431(.data_in(wire_d43_0),.data_out(wire_d43_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance44432(.data_in(wire_d43_1),.data_out(wire_d43_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance44433(.data_in(wire_d43_2),.data_out(wire_d43_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance44434(.data_in(wire_d43_3),.data_out(wire_d43_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance44435(.data_in(wire_d43_4),.data_out(wire_d43_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance44436(.data_in(wire_d43_5),.data_out(wire_d43_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance44437(.data_in(wire_d43_6),.data_out(wire_d43_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance44438(.data_in(wire_d43_7),.data_out(wire_d43_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance44439(.data_in(wire_d43_8),.data_out(wire_d43_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444310(.data_in(wire_d43_9),.data_out(wire_d43_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444311(.data_in(wire_d43_10),.data_out(wire_d43_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444312(.data_in(wire_d43_11),.data_out(wire_d43_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444313(.data_in(wire_d43_12),.data_out(wire_d43_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444314(.data_in(wire_d43_13),.data_out(wire_d43_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444315(.data_in(wire_d43_14),.data_out(wire_d43_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444316(.data_in(wire_d43_15),.data_out(wire_d43_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444317(.data_in(wire_d43_16),.data_out(wire_d43_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444318(.data_in(wire_d43_17),.data_out(wire_d43_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444319(.data_in(wire_d43_18),.data_out(wire_d43_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444320(.data_in(wire_d43_19),.data_out(wire_d43_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444321(.data_in(wire_d43_20),.data_out(wire_d43_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444322(.data_in(wire_d43_21),.data_out(wire_d43_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444323(.data_in(wire_d43_22),.data_out(wire_d43_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444324(.data_in(wire_d43_23),.data_out(wire_d43_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444325(.data_in(wire_d43_24),.data_out(wire_d43_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444326(.data_in(wire_d43_25),.data_out(wire_d43_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444327(.data_in(wire_d43_26),.data_out(wire_d43_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444328(.data_in(wire_d43_27),.data_out(wire_d43_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444329(.data_in(wire_d43_28),.data_out(wire_d43_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444330(.data_in(wire_d43_29),.data_out(wire_d43_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444331(.data_in(wire_d43_30),.data_out(wire_d43_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444332(.data_in(wire_d43_31),.data_out(wire_d43_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444333(.data_in(wire_d43_32),.data_out(wire_d43_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444334(.data_in(wire_d43_33),.data_out(wire_d43_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444335(.data_in(wire_d43_34),.data_out(wire_d43_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444336(.data_in(wire_d43_35),.data_out(wire_d43_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444337(.data_in(wire_d43_36),.data_out(wire_d43_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444338(.data_in(wire_d43_37),.data_out(wire_d43_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444339(.data_in(wire_d43_38),.data_out(wire_d43_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444340(.data_in(wire_d43_39),.data_out(wire_d43_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444341(.data_in(wire_d43_40),.data_out(wire_d43_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444342(.data_in(wire_d43_41),.data_out(wire_d43_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444343(.data_in(wire_d43_42),.data_out(wire_d43_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444344(.data_in(wire_d43_43),.data_out(wire_d43_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444345(.data_in(wire_d43_44),.data_out(wire_d43_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444346(.data_in(wire_d43_45),.data_out(wire_d43_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444347(.data_in(wire_d43_46),.data_out(wire_d43_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444348(.data_in(wire_d43_47),.data_out(wire_d43_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444349(.data_in(wire_d43_48),.data_out(wire_d43_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444350(.data_in(wire_d43_49),.data_out(wire_d43_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444351(.data_in(wire_d43_50),.data_out(wire_d43_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444352(.data_in(wire_d43_51),.data_out(wire_d43_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444353(.data_in(wire_d43_52),.data_out(wire_d43_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance444354(.data_in(wire_d43_53),.data_out(wire_d43_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444355(.data_in(wire_d43_54),.data_out(wire_d43_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444356(.data_in(wire_d43_55),.data_out(wire_d43_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444357(.data_in(wire_d43_56),.data_out(wire_d43_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444358(.data_in(wire_d43_57),.data_out(wire_d43_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444359(.data_in(wire_d43_58),.data_out(wire_d43_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444360(.data_in(wire_d43_59),.data_out(wire_d43_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444361(.data_in(wire_d43_60),.data_out(wire_d43_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444362(.data_in(wire_d43_61),.data_out(wire_d43_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444363(.data_in(wire_d43_62),.data_out(wire_d43_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444364(.data_in(wire_d43_63),.data_out(wire_d43_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444365(.data_in(wire_d43_64),.data_out(wire_d43_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444366(.data_in(wire_d43_65),.data_out(wire_d43_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance444367(.data_in(wire_d43_66),.data_out(wire_d43_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance444368(.data_in(wire_d43_67),.data_out(wire_d43_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance444369(.data_in(wire_d43_68),.data_out(d_out43),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance45440(.data_in(d_in44),.data_out(wire_d44_0),.clk(clk),.rst(rst));            //channel 45
	invertion #(.WIDTH(WIDTH)) invertion_instance45441(.data_in(wire_d44_0),.data_out(wire_d44_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance45442(.data_in(wire_d44_1),.data_out(wire_d44_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance45443(.data_in(wire_d44_2),.data_out(wire_d44_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance45444(.data_in(wire_d44_3),.data_out(wire_d44_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance45445(.data_in(wire_d44_4),.data_out(wire_d44_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance45446(.data_in(wire_d44_5),.data_out(wire_d44_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance45447(.data_in(wire_d44_6),.data_out(wire_d44_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance45448(.data_in(wire_d44_7),.data_out(wire_d44_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance45449(.data_in(wire_d44_8),.data_out(wire_d44_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454410(.data_in(wire_d44_9),.data_out(wire_d44_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454411(.data_in(wire_d44_10),.data_out(wire_d44_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454412(.data_in(wire_d44_11),.data_out(wire_d44_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454413(.data_in(wire_d44_12),.data_out(wire_d44_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454414(.data_in(wire_d44_13),.data_out(wire_d44_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454415(.data_in(wire_d44_14),.data_out(wire_d44_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454416(.data_in(wire_d44_15),.data_out(wire_d44_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454417(.data_in(wire_d44_16),.data_out(wire_d44_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454418(.data_in(wire_d44_17),.data_out(wire_d44_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454419(.data_in(wire_d44_18),.data_out(wire_d44_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454420(.data_in(wire_d44_19),.data_out(wire_d44_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454421(.data_in(wire_d44_20),.data_out(wire_d44_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454422(.data_in(wire_d44_21),.data_out(wire_d44_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454423(.data_in(wire_d44_22),.data_out(wire_d44_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454424(.data_in(wire_d44_23),.data_out(wire_d44_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454425(.data_in(wire_d44_24),.data_out(wire_d44_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454426(.data_in(wire_d44_25),.data_out(wire_d44_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454427(.data_in(wire_d44_26),.data_out(wire_d44_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454428(.data_in(wire_d44_27),.data_out(wire_d44_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454429(.data_in(wire_d44_28),.data_out(wire_d44_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454430(.data_in(wire_d44_29),.data_out(wire_d44_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454431(.data_in(wire_d44_30),.data_out(wire_d44_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454432(.data_in(wire_d44_31),.data_out(wire_d44_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454433(.data_in(wire_d44_32),.data_out(wire_d44_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454434(.data_in(wire_d44_33),.data_out(wire_d44_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454435(.data_in(wire_d44_34),.data_out(wire_d44_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454436(.data_in(wire_d44_35),.data_out(wire_d44_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454437(.data_in(wire_d44_36),.data_out(wire_d44_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454438(.data_in(wire_d44_37),.data_out(wire_d44_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454439(.data_in(wire_d44_38),.data_out(wire_d44_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454440(.data_in(wire_d44_39),.data_out(wire_d44_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454441(.data_in(wire_d44_40),.data_out(wire_d44_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454442(.data_in(wire_d44_41),.data_out(wire_d44_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454443(.data_in(wire_d44_42),.data_out(wire_d44_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454444(.data_in(wire_d44_43),.data_out(wire_d44_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454445(.data_in(wire_d44_44),.data_out(wire_d44_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454446(.data_in(wire_d44_45),.data_out(wire_d44_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454447(.data_in(wire_d44_46),.data_out(wire_d44_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454448(.data_in(wire_d44_47),.data_out(wire_d44_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454449(.data_in(wire_d44_48),.data_out(wire_d44_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454450(.data_in(wire_d44_49),.data_out(wire_d44_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454451(.data_in(wire_d44_50),.data_out(wire_d44_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454452(.data_in(wire_d44_51),.data_out(wire_d44_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454453(.data_in(wire_d44_52),.data_out(wire_d44_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454454(.data_in(wire_d44_53),.data_out(wire_d44_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454455(.data_in(wire_d44_54),.data_out(wire_d44_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454456(.data_in(wire_d44_55),.data_out(wire_d44_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454457(.data_in(wire_d44_56),.data_out(wire_d44_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance454458(.data_in(wire_d44_57),.data_out(wire_d44_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454459(.data_in(wire_d44_58),.data_out(wire_d44_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454460(.data_in(wire_d44_59),.data_out(wire_d44_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454461(.data_in(wire_d44_60),.data_out(wire_d44_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454462(.data_in(wire_d44_61),.data_out(wire_d44_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454463(.data_in(wire_d44_62),.data_out(wire_d44_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance454464(.data_in(wire_d44_63),.data_out(wire_d44_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454465(.data_in(wire_d44_64),.data_out(wire_d44_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454466(.data_in(wire_d44_65),.data_out(wire_d44_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454467(.data_in(wire_d44_66),.data_out(wire_d44_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance454468(.data_in(wire_d44_67),.data_out(wire_d44_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance454469(.data_in(wire_d44_68),.data_out(d_out44),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance46450(.data_in(d_in45),.data_out(wire_d45_0),.clk(clk),.rst(rst));            //channel 46
	encoder #(.WIDTH(WIDTH)) encoder_instance46451(.data_in(wire_d45_0),.data_out(wire_d45_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance46452(.data_in(wire_d45_1),.data_out(wire_d45_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance46453(.data_in(wire_d45_2),.data_out(wire_d45_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance46454(.data_in(wire_d45_3),.data_out(wire_d45_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance46455(.data_in(wire_d45_4),.data_out(wire_d45_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance46456(.data_in(wire_d45_5),.data_out(wire_d45_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance46457(.data_in(wire_d45_6),.data_out(wire_d45_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance46458(.data_in(wire_d45_7),.data_out(wire_d45_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance46459(.data_in(wire_d45_8),.data_out(wire_d45_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464510(.data_in(wire_d45_9),.data_out(wire_d45_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464511(.data_in(wire_d45_10),.data_out(wire_d45_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464512(.data_in(wire_d45_11),.data_out(wire_d45_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464513(.data_in(wire_d45_12),.data_out(wire_d45_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464514(.data_in(wire_d45_13),.data_out(wire_d45_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464515(.data_in(wire_d45_14),.data_out(wire_d45_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464516(.data_in(wire_d45_15),.data_out(wire_d45_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464517(.data_in(wire_d45_16),.data_out(wire_d45_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464518(.data_in(wire_d45_17),.data_out(wire_d45_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464519(.data_in(wire_d45_18),.data_out(wire_d45_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464520(.data_in(wire_d45_19),.data_out(wire_d45_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464521(.data_in(wire_d45_20),.data_out(wire_d45_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464522(.data_in(wire_d45_21),.data_out(wire_d45_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464523(.data_in(wire_d45_22),.data_out(wire_d45_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464524(.data_in(wire_d45_23),.data_out(wire_d45_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464525(.data_in(wire_d45_24),.data_out(wire_d45_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464526(.data_in(wire_d45_25),.data_out(wire_d45_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464527(.data_in(wire_d45_26),.data_out(wire_d45_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464528(.data_in(wire_d45_27),.data_out(wire_d45_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464529(.data_in(wire_d45_28),.data_out(wire_d45_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464530(.data_in(wire_d45_29),.data_out(wire_d45_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464531(.data_in(wire_d45_30),.data_out(wire_d45_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464532(.data_in(wire_d45_31),.data_out(wire_d45_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464533(.data_in(wire_d45_32),.data_out(wire_d45_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464534(.data_in(wire_d45_33),.data_out(wire_d45_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464535(.data_in(wire_d45_34),.data_out(wire_d45_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464536(.data_in(wire_d45_35),.data_out(wire_d45_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464537(.data_in(wire_d45_36),.data_out(wire_d45_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464538(.data_in(wire_d45_37),.data_out(wire_d45_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464539(.data_in(wire_d45_38),.data_out(wire_d45_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464540(.data_in(wire_d45_39),.data_out(wire_d45_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464541(.data_in(wire_d45_40),.data_out(wire_d45_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464542(.data_in(wire_d45_41),.data_out(wire_d45_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464543(.data_in(wire_d45_42),.data_out(wire_d45_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464544(.data_in(wire_d45_43),.data_out(wire_d45_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464545(.data_in(wire_d45_44),.data_out(wire_d45_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464546(.data_in(wire_d45_45),.data_out(wire_d45_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464547(.data_in(wire_d45_46),.data_out(wire_d45_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464548(.data_in(wire_d45_47),.data_out(wire_d45_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464549(.data_in(wire_d45_48),.data_out(wire_d45_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464550(.data_in(wire_d45_49),.data_out(wire_d45_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464551(.data_in(wire_d45_50),.data_out(wire_d45_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464552(.data_in(wire_d45_51),.data_out(wire_d45_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464553(.data_in(wire_d45_52),.data_out(wire_d45_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464554(.data_in(wire_d45_53),.data_out(wire_d45_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464555(.data_in(wire_d45_54),.data_out(wire_d45_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464556(.data_in(wire_d45_55),.data_out(wire_d45_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464557(.data_in(wire_d45_56),.data_out(wire_d45_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464558(.data_in(wire_d45_57),.data_out(wire_d45_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464559(.data_in(wire_d45_58),.data_out(wire_d45_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464560(.data_in(wire_d45_59),.data_out(wire_d45_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464561(.data_in(wire_d45_60),.data_out(wire_d45_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance464562(.data_in(wire_d45_61),.data_out(wire_d45_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464563(.data_in(wire_d45_62),.data_out(wire_d45_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464564(.data_in(wire_d45_63),.data_out(wire_d45_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance464565(.data_in(wire_d45_64),.data_out(wire_d45_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464566(.data_in(wire_d45_65),.data_out(wire_d45_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464567(.data_in(wire_d45_66),.data_out(wire_d45_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance464568(.data_in(wire_d45_67),.data_out(wire_d45_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance464569(.data_in(wire_d45_68),.data_out(d_out45),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance47460(.data_in(d_in46),.data_out(wire_d46_0),.clk(clk),.rst(rst));            //channel 47
	encoder #(.WIDTH(WIDTH)) encoder_instance47461(.data_in(wire_d46_0),.data_out(wire_d46_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance47462(.data_in(wire_d46_1),.data_out(wire_d46_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance47463(.data_in(wire_d46_2),.data_out(wire_d46_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance47464(.data_in(wire_d46_3),.data_out(wire_d46_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance47465(.data_in(wire_d46_4),.data_out(wire_d46_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance47466(.data_in(wire_d46_5),.data_out(wire_d46_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance47467(.data_in(wire_d46_6),.data_out(wire_d46_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance47468(.data_in(wire_d46_7),.data_out(wire_d46_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance47469(.data_in(wire_d46_8),.data_out(wire_d46_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474610(.data_in(wire_d46_9),.data_out(wire_d46_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474611(.data_in(wire_d46_10),.data_out(wire_d46_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474612(.data_in(wire_d46_11),.data_out(wire_d46_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474613(.data_in(wire_d46_12),.data_out(wire_d46_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474614(.data_in(wire_d46_13),.data_out(wire_d46_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474615(.data_in(wire_d46_14),.data_out(wire_d46_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474616(.data_in(wire_d46_15),.data_out(wire_d46_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474617(.data_in(wire_d46_16),.data_out(wire_d46_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474618(.data_in(wire_d46_17),.data_out(wire_d46_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474619(.data_in(wire_d46_18),.data_out(wire_d46_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474620(.data_in(wire_d46_19),.data_out(wire_d46_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474621(.data_in(wire_d46_20),.data_out(wire_d46_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474622(.data_in(wire_d46_21),.data_out(wire_d46_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474623(.data_in(wire_d46_22),.data_out(wire_d46_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474624(.data_in(wire_d46_23),.data_out(wire_d46_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474625(.data_in(wire_d46_24),.data_out(wire_d46_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474626(.data_in(wire_d46_25),.data_out(wire_d46_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474627(.data_in(wire_d46_26),.data_out(wire_d46_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474628(.data_in(wire_d46_27),.data_out(wire_d46_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474629(.data_in(wire_d46_28),.data_out(wire_d46_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474630(.data_in(wire_d46_29),.data_out(wire_d46_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474631(.data_in(wire_d46_30),.data_out(wire_d46_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474632(.data_in(wire_d46_31),.data_out(wire_d46_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474633(.data_in(wire_d46_32),.data_out(wire_d46_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474634(.data_in(wire_d46_33),.data_out(wire_d46_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474635(.data_in(wire_d46_34),.data_out(wire_d46_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474636(.data_in(wire_d46_35),.data_out(wire_d46_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474637(.data_in(wire_d46_36),.data_out(wire_d46_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474638(.data_in(wire_d46_37),.data_out(wire_d46_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474639(.data_in(wire_d46_38),.data_out(wire_d46_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474640(.data_in(wire_d46_39),.data_out(wire_d46_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474641(.data_in(wire_d46_40),.data_out(wire_d46_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474642(.data_in(wire_d46_41),.data_out(wire_d46_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474643(.data_in(wire_d46_42),.data_out(wire_d46_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474644(.data_in(wire_d46_43),.data_out(wire_d46_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474645(.data_in(wire_d46_44),.data_out(wire_d46_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474646(.data_in(wire_d46_45),.data_out(wire_d46_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474647(.data_in(wire_d46_46),.data_out(wire_d46_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474648(.data_in(wire_d46_47),.data_out(wire_d46_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474649(.data_in(wire_d46_48),.data_out(wire_d46_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474650(.data_in(wire_d46_49),.data_out(wire_d46_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474651(.data_in(wire_d46_50),.data_out(wire_d46_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474652(.data_in(wire_d46_51),.data_out(wire_d46_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474653(.data_in(wire_d46_52),.data_out(wire_d46_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474654(.data_in(wire_d46_53),.data_out(wire_d46_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474655(.data_in(wire_d46_54),.data_out(wire_d46_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474656(.data_in(wire_d46_55),.data_out(wire_d46_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474657(.data_in(wire_d46_56),.data_out(wire_d46_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474658(.data_in(wire_d46_57),.data_out(wire_d46_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474659(.data_in(wire_d46_58),.data_out(wire_d46_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474660(.data_in(wire_d46_59),.data_out(wire_d46_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474661(.data_in(wire_d46_60),.data_out(wire_d46_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474662(.data_in(wire_d46_61),.data_out(wire_d46_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance474663(.data_in(wire_d46_62),.data_out(wire_d46_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474664(.data_in(wire_d46_63),.data_out(wire_d46_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance474665(.data_in(wire_d46_64),.data_out(wire_d46_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474666(.data_in(wire_d46_65),.data_out(wire_d46_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474667(.data_in(wire_d46_66),.data_out(wire_d46_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance474668(.data_in(wire_d46_67),.data_out(wire_d46_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance474669(.data_in(wire_d46_68),.data_out(d_out46),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance48470(.data_in(d_in47),.data_out(wire_d47_0),.clk(clk),.rst(rst));            //channel 48
	register #(.WIDTH(WIDTH)) register_instance48471(.data_in(wire_d47_0),.data_out(wire_d47_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance48472(.data_in(wire_d47_1),.data_out(wire_d47_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance48473(.data_in(wire_d47_2),.data_out(wire_d47_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance48474(.data_in(wire_d47_3),.data_out(wire_d47_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance48475(.data_in(wire_d47_4),.data_out(wire_d47_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance48476(.data_in(wire_d47_5),.data_out(wire_d47_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance48477(.data_in(wire_d47_6),.data_out(wire_d47_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance48478(.data_in(wire_d47_7),.data_out(wire_d47_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance48479(.data_in(wire_d47_8),.data_out(wire_d47_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484710(.data_in(wire_d47_9),.data_out(wire_d47_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484711(.data_in(wire_d47_10),.data_out(wire_d47_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484712(.data_in(wire_d47_11),.data_out(wire_d47_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484713(.data_in(wire_d47_12),.data_out(wire_d47_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484714(.data_in(wire_d47_13),.data_out(wire_d47_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484715(.data_in(wire_d47_14),.data_out(wire_d47_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484716(.data_in(wire_d47_15),.data_out(wire_d47_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484717(.data_in(wire_d47_16),.data_out(wire_d47_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484718(.data_in(wire_d47_17),.data_out(wire_d47_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484719(.data_in(wire_d47_18),.data_out(wire_d47_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484720(.data_in(wire_d47_19),.data_out(wire_d47_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484721(.data_in(wire_d47_20),.data_out(wire_d47_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484722(.data_in(wire_d47_21),.data_out(wire_d47_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484723(.data_in(wire_d47_22),.data_out(wire_d47_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484724(.data_in(wire_d47_23),.data_out(wire_d47_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484725(.data_in(wire_d47_24),.data_out(wire_d47_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484726(.data_in(wire_d47_25),.data_out(wire_d47_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484727(.data_in(wire_d47_26),.data_out(wire_d47_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484728(.data_in(wire_d47_27),.data_out(wire_d47_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484729(.data_in(wire_d47_28),.data_out(wire_d47_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484730(.data_in(wire_d47_29),.data_out(wire_d47_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484731(.data_in(wire_d47_30),.data_out(wire_d47_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484732(.data_in(wire_d47_31),.data_out(wire_d47_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484733(.data_in(wire_d47_32),.data_out(wire_d47_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484734(.data_in(wire_d47_33),.data_out(wire_d47_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484735(.data_in(wire_d47_34),.data_out(wire_d47_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484736(.data_in(wire_d47_35),.data_out(wire_d47_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484737(.data_in(wire_d47_36),.data_out(wire_d47_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484738(.data_in(wire_d47_37),.data_out(wire_d47_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484739(.data_in(wire_d47_38),.data_out(wire_d47_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484740(.data_in(wire_d47_39),.data_out(wire_d47_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484741(.data_in(wire_d47_40),.data_out(wire_d47_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484742(.data_in(wire_d47_41),.data_out(wire_d47_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484743(.data_in(wire_d47_42),.data_out(wire_d47_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484744(.data_in(wire_d47_43),.data_out(wire_d47_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484745(.data_in(wire_d47_44),.data_out(wire_d47_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484746(.data_in(wire_d47_45),.data_out(wire_d47_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484747(.data_in(wire_d47_46),.data_out(wire_d47_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484748(.data_in(wire_d47_47),.data_out(wire_d47_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484749(.data_in(wire_d47_48),.data_out(wire_d47_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484750(.data_in(wire_d47_49),.data_out(wire_d47_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484751(.data_in(wire_d47_50),.data_out(wire_d47_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484752(.data_in(wire_d47_51),.data_out(wire_d47_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484753(.data_in(wire_d47_52),.data_out(wire_d47_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484754(.data_in(wire_d47_53),.data_out(wire_d47_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484755(.data_in(wire_d47_54),.data_out(wire_d47_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484756(.data_in(wire_d47_55),.data_out(wire_d47_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484757(.data_in(wire_d47_56),.data_out(wire_d47_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484758(.data_in(wire_d47_57),.data_out(wire_d47_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484759(.data_in(wire_d47_58),.data_out(wire_d47_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484760(.data_in(wire_d47_59),.data_out(wire_d47_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance484761(.data_in(wire_d47_60),.data_out(wire_d47_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484762(.data_in(wire_d47_61),.data_out(wire_d47_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484763(.data_in(wire_d47_62),.data_out(wire_d47_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484764(.data_in(wire_d47_63),.data_out(wire_d47_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484765(.data_in(wire_d47_64),.data_out(wire_d47_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484766(.data_in(wire_d47_65),.data_out(wire_d47_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance484767(.data_in(wire_d47_66),.data_out(wire_d47_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance484768(.data_in(wire_d47_67),.data_out(wire_d47_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance484769(.data_in(wire_d47_68),.data_out(d_out47),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance49480(.data_in(d_in48),.data_out(wire_d48_0),.clk(clk),.rst(rst));            //channel 49
	large_mux #(.WIDTH(WIDTH)) large_mux_instance49481(.data_in(wire_d48_0),.data_out(wire_d48_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance49482(.data_in(wire_d48_1),.data_out(wire_d48_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance49483(.data_in(wire_d48_2),.data_out(wire_d48_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance49484(.data_in(wire_d48_3),.data_out(wire_d48_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance49485(.data_in(wire_d48_4),.data_out(wire_d48_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance49486(.data_in(wire_d48_5),.data_out(wire_d48_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance49487(.data_in(wire_d48_6),.data_out(wire_d48_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance49488(.data_in(wire_d48_7),.data_out(wire_d48_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance49489(.data_in(wire_d48_8),.data_out(wire_d48_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494810(.data_in(wire_d48_9),.data_out(wire_d48_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494811(.data_in(wire_d48_10),.data_out(wire_d48_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494812(.data_in(wire_d48_11),.data_out(wire_d48_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494813(.data_in(wire_d48_12),.data_out(wire_d48_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494814(.data_in(wire_d48_13),.data_out(wire_d48_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494815(.data_in(wire_d48_14),.data_out(wire_d48_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494816(.data_in(wire_d48_15),.data_out(wire_d48_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494817(.data_in(wire_d48_16),.data_out(wire_d48_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494818(.data_in(wire_d48_17),.data_out(wire_d48_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494819(.data_in(wire_d48_18),.data_out(wire_d48_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494820(.data_in(wire_d48_19),.data_out(wire_d48_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494821(.data_in(wire_d48_20),.data_out(wire_d48_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494822(.data_in(wire_d48_21),.data_out(wire_d48_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494823(.data_in(wire_d48_22),.data_out(wire_d48_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494824(.data_in(wire_d48_23),.data_out(wire_d48_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494825(.data_in(wire_d48_24),.data_out(wire_d48_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494826(.data_in(wire_d48_25),.data_out(wire_d48_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494827(.data_in(wire_d48_26),.data_out(wire_d48_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494828(.data_in(wire_d48_27),.data_out(wire_d48_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494829(.data_in(wire_d48_28),.data_out(wire_d48_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494830(.data_in(wire_d48_29),.data_out(wire_d48_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494831(.data_in(wire_d48_30),.data_out(wire_d48_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494832(.data_in(wire_d48_31),.data_out(wire_d48_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494833(.data_in(wire_d48_32),.data_out(wire_d48_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494834(.data_in(wire_d48_33),.data_out(wire_d48_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494835(.data_in(wire_d48_34),.data_out(wire_d48_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494836(.data_in(wire_d48_35),.data_out(wire_d48_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494837(.data_in(wire_d48_36),.data_out(wire_d48_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494838(.data_in(wire_d48_37),.data_out(wire_d48_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494839(.data_in(wire_d48_38),.data_out(wire_d48_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494840(.data_in(wire_d48_39),.data_out(wire_d48_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494841(.data_in(wire_d48_40),.data_out(wire_d48_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494842(.data_in(wire_d48_41),.data_out(wire_d48_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494843(.data_in(wire_d48_42),.data_out(wire_d48_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494844(.data_in(wire_d48_43),.data_out(wire_d48_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494845(.data_in(wire_d48_44),.data_out(wire_d48_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494846(.data_in(wire_d48_45),.data_out(wire_d48_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494847(.data_in(wire_d48_46),.data_out(wire_d48_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494848(.data_in(wire_d48_47),.data_out(wire_d48_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494849(.data_in(wire_d48_48),.data_out(wire_d48_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494850(.data_in(wire_d48_49),.data_out(wire_d48_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494851(.data_in(wire_d48_50),.data_out(wire_d48_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494852(.data_in(wire_d48_51),.data_out(wire_d48_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494853(.data_in(wire_d48_52),.data_out(wire_d48_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494854(.data_in(wire_d48_53),.data_out(wire_d48_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494855(.data_in(wire_d48_54),.data_out(wire_d48_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494856(.data_in(wire_d48_55),.data_out(wire_d48_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494857(.data_in(wire_d48_56),.data_out(wire_d48_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494858(.data_in(wire_d48_57),.data_out(wire_d48_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494859(.data_in(wire_d48_58),.data_out(wire_d48_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494860(.data_in(wire_d48_59),.data_out(wire_d48_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494861(.data_in(wire_d48_60),.data_out(wire_d48_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494862(.data_in(wire_d48_61),.data_out(wire_d48_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance494863(.data_in(wire_d48_62),.data_out(wire_d48_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494864(.data_in(wire_d48_63),.data_out(wire_d48_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance494865(.data_in(wire_d48_64),.data_out(wire_d48_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494866(.data_in(wire_d48_65),.data_out(wire_d48_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494867(.data_in(wire_d48_66),.data_out(wire_d48_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance494868(.data_in(wire_d48_67),.data_out(wire_d48_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance494869(.data_in(wire_d48_68),.data_out(d_out48),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance50490(.data_in(d_in49),.data_out(wire_d49_0),.clk(clk),.rst(rst));            //channel 50
	invertion #(.WIDTH(WIDTH)) invertion_instance50491(.data_in(wire_d49_0),.data_out(wire_d49_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance50492(.data_in(wire_d49_1),.data_out(wire_d49_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance50493(.data_in(wire_d49_2),.data_out(wire_d49_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance50494(.data_in(wire_d49_3),.data_out(wire_d49_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance50495(.data_in(wire_d49_4),.data_out(wire_d49_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance50496(.data_in(wire_d49_5),.data_out(wire_d49_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance50497(.data_in(wire_d49_6),.data_out(wire_d49_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance50498(.data_in(wire_d49_7),.data_out(wire_d49_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance50499(.data_in(wire_d49_8),.data_out(wire_d49_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504910(.data_in(wire_d49_9),.data_out(wire_d49_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504911(.data_in(wire_d49_10),.data_out(wire_d49_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504912(.data_in(wire_d49_11),.data_out(wire_d49_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504913(.data_in(wire_d49_12),.data_out(wire_d49_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504914(.data_in(wire_d49_13),.data_out(wire_d49_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504915(.data_in(wire_d49_14),.data_out(wire_d49_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504916(.data_in(wire_d49_15),.data_out(wire_d49_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504917(.data_in(wire_d49_16),.data_out(wire_d49_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504918(.data_in(wire_d49_17),.data_out(wire_d49_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504919(.data_in(wire_d49_18),.data_out(wire_d49_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504920(.data_in(wire_d49_19),.data_out(wire_d49_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504921(.data_in(wire_d49_20),.data_out(wire_d49_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504922(.data_in(wire_d49_21),.data_out(wire_d49_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504923(.data_in(wire_d49_22),.data_out(wire_d49_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504924(.data_in(wire_d49_23),.data_out(wire_d49_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504925(.data_in(wire_d49_24),.data_out(wire_d49_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504926(.data_in(wire_d49_25),.data_out(wire_d49_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504927(.data_in(wire_d49_26),.data_out(wire_d49_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504928(.data_in(wire_d49_27),.data_out(wire_d49_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504929(.data_in(wire_d49_28),.data_out(wire_d49_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504930(.data_in(wire_d49_29),.data_out(wire_d49_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504931(.data_in(wire_d49_30),.data_out(wire_d49_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504932(.data_in(wire_d49_31),.data_out(wire_d49_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504933(.data_in(wire_d49_32),.data_out(wire_d49_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504934(.data_in(wire_d49_33),.data_out(wire_d49_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504935(.data_in(wire_d49_34),.data_out(wire_d49_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504936(.data_in(wire_d49_35),.data_out(wire_d49_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504937(.data_in(wire_d49_36),.data_out(wire_d49_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504938(.data_in(wire_d49_37),.data_out(wire_d49_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504939(.data_in(wire_d49_38),.data_out(wire_d49_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504940(.data_in(wire_d49_39),.data_out(wire_d49_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504941(.data_in(wire_d49_40),.data_out(wire_d49_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504942(.data_in(wire_d49_41),.data_out(wire_d49_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504943(.data_in(wire_d49_42),.data_out(wire_d49_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504944(.data_in(wire_d49_43),.data_out(wire_d49_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504945(.data_in(wire_d49_44),.data_out(wire_d49_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504946(.data_in(wire_d49_45),.data_out(wire_d49_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504947(.data_in(wire_d49_46),.data_out(wire_d49_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504948(.data_in(wire_d49_47),.data_out(wire_d49_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504949(.data_in(wire_d49_48),.data_out(wire_d49_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504950(.data_in(wire_d49_49),.data_out(wire_d49_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504951(.data_in(wire_d49_50),.data_out(wire_d49_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504952(.data_in(wire_d49_51),.data_out(wire_d49_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504953(.data_in(wire_d49_52),.data_out(wire_d49_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504954(.data_in(wire_d49_53),.data_out(wire_d49_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504955(.data_in(wire_d49_54),.data_out(wire_d49_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504956(.data_in(wire_d49_55),.data_out(wire_d49_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504957(.data_in(wire_d49_56),.data_out(wire_d49_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504958(.data_in(wire_d49_57),.data_out(wire_d49_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504959(.data_in(wire_d49_58),.data_out(wire_d49_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504960(.data_in(wire_d49_59),.data_out(wire_d49_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504961(.data_in(wire_d49_60),.data_out(wire_d49_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504962(.data_in(wire_d49_61),.data_out(wire_d49_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance504963(.data_in(wire_d49_62),.data_out(wire_d49_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504964(.data_in(wire_d49_63),.data_out(wire_d49_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504965(.data_in(wire_d49_64),.data_out(wire_d49_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance504966(.data_in(wire_d49_65),.data_out(wire_d49_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance504967(.data_in(wire_d49_66),.data_out(wire_d49_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504968(.data_in(wire_d49_67),.data_out(wire_d49_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance504969(.data_in(wire_d49_68),.data_out(d_out49),.clk(clk),.rst(rst));


endmodule