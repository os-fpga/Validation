// `include "encoder.v"
// `include "invertion.v"
// `include "large_adder.v"
// `include "large_mux.v"
// `include "memory_cntrl.v"
// `include "register.v"
// `include "full_adder.v"
// `include "d_latch.v"
// `include "shift_reg.v"
// `include "mod_n_counter.v"
// `include "decoder.v"
// `include "parity_generator.v"

module design210_100_120_top #(parameter WIDTH=32,CHANNEL=100) (clk, rst, in, out);

	localparam OUT_BUS=CHANNEL*WIDTH;
	input clk,rst;
	input [WIDTH-1:0] in;
	output [WIDTH-1:0] out;

	reg [WIDTH-1:0] d_in0;
	reg [WIDTH-1:0] d_in1;
	reg [WIDTH-1:0] d_in2;
	reg [WIDTH-1:0] d_in3;
	reg [WIDTH-1:0] d_in4;
	reg [WIDTH-1:0] d_in5;
	reg [WIDTH-1:0] d_in6;
	reg [WIDTH-1:0] d_in7;
	reg [WIDTH-1:0] d_in8;
	reg [WIDTH-1:0] d_in9;
	reg [WIDTH-1:0] d_in10;
	reg [WIDTH-1:0] d_in11;
	reg [WIDTH-1:0] d_in12;
	reg [WIDTH-1:0] d_in13;
	reg [WIDTH-1:0] d_in14;
	reg [WIDTH-1:0] d_in15;
	reg [WIDTH-1:0] d_in16;
	reg [WIDTH-1:0] d_in17;
	reg [WIDTH-1:0] d_in18;
	reg [WIDTH-1:0] d_in19;
	reg [WIDTH-1:0] d_in20;
	reg [WIDTH-1:0] d_in21;
	reg [WIDTH-1:0] d_in22;
	reg [WIDTH-1:0] d_in23;
	reg [WIDTH-1:0] d_in24;
	reg [WIDTH-1:0] d_in25;
	reg [WIDTH-1:0] d_in26;
	reg [WIDTH-1:0] d_in27;
	reg [WIDTH-1:0] d_in28;
	reg [WIDTH-1:0] d_in29;
	reg [WIDTH-1:0] d_in30;
	reg [WIDTH-1:0] d_in31;
	reg [WIDTH-1:0] d_in32;
	reg [WIDTH-1:0] d_in33;
	reg [WIDTH-1:0] d_in34;
	reg [WIDTH-1:0] d_in35;
	reg [WIDTH-1:0] d_in36;
	reg [WIDTH-1:0] d_in37;
	reg [WIDTH-1:0] d_in38;
	reg [WIDTH-1:0] d_in39;
	reg [WIDTH-1:0] d_in40;
	reg [WIDTH-1:0] d_in41;
	reg [WIDTH-1:0] d_in42;
	reg [WIDTH-1:0] d_in43;
	reg [WIDTH-1:0] d_in44;
	reg [WIDTH-1:0] d_in45;
	reg [WIDTH-1:0] d_in46;
	reg [WIDTH-1:0] d_in47;
	reg [WIDTH-1:0] d_in48;
	reg [WIDTH-1:0] d_in49;
	reg [WIDTH-1:0] d_in50;
	reg [WIDTH-1:0] d_in51;
	reg [WIDTH-1:0] d_in52;
	reg [WIDTH-1:0] d_in53;
	reg [WIDTH-1:0] d_in54;
	reg [WIDTH-1:0] d_in55;
	reg [WIDTH-1:0] d_in56;
	reg [WIDTH-1:0] d_in57;
	reg [WIDTH-1:0] d_in58;
	reg [WIDTH-1:0] d_in59;
	reg [WIDTH-1:0] d_in60;
	reg [WIDTH-1:0] d_in61;
	reg [WIDTH-1:0] d_in62;
	reg [WIDTH-1:0] d_in63;
	reg [WIDTH-1:0] d_in64;
	reg [WIDTH-1:0] d_in65;
	reg [WIDTH-1:0] d_in66;
	reg [WIDTH-1:0] d_in67;
	reg [WIDTH-1:0] d_in68;
	reg [WIDTH-1:0] d_in69;
	reg [WIDTH-1:0] d_in70;
	reg [WIDTH-1:0] d_in71;
	reg [WIDTH-1:0] d_in72;
	reg [WIDTH-1:0] d_in73;
	reg [WIDTH-1:0] d_in74;
	reg [WIDTH-1:0] d_in75;
	reg [WIDTH-1:0] d_in76;
	reg [WIDTH-1:0] d_in77;
	reg [WIDTH-1:0] d_in78;
	reg [WIDTH-1:0] d_in79;
	reg [WIDTH-1:0] d_in80;
	reg [WIDTH-1:0] d_in81;
	reg [WIDTH-1:0] d_in82;
	reg [WIDTH-1:0] d_in83;
	reg [WIDTH-1:0] d_in84;
	reg [WIDTH-1:0] d_in85;
	reg [WIDTH-1:0] d_in86;
	reg [WIDTH-1:0] d_in87;
	reg [WIDTH-1:0] d_in88;
	reg [WIDTH-1:0] d_in89;
	reg [WIDTH-1:0] d_in90;
	reg [WIDTH-1:0] d_in91;
	reg [WIDTH-1:0] d_in92;
	reg [WIDTH-1:0] d_in93;
	reg [WIDTH-1:0] d_in94;
	reg [WIDTH-1:0] d_in95;
	reg [WIDTH-1:0] d_in96;
	reg [WIDTH-1:0] d_in97;
	reg [WIDTH-1:0] d_in98;
	reg [WIDTH-1:0] d_in99;
	wire [WIDTH-1:0] d_out0;
	wire [WIDTH-1:0] d_out1;
	wire [WIDTH-1:0] d_out2;
	wire [WIDTH-1:0] d_out3;
	wire [WIDTH-1:0] d_out4;
	wire [WIDTH-1:0] d_out5;
	wire [WIDTH-1:0] d_out6;
	wire [WIDTH-1:0] d_out7;
	wire [WIDTH-1:0] d_out8;
	wire [WIDTH-1:0] d_out9;
	wire [WIDTH-1:0] d_out10;
	wire [WIDTH-1:0] d_out11;
	wire [WIDTH-1:0] d_out12;
	wire [WIDTH-1:0] d_out13;
	wire [WIDTH-1:0] d_out14;
	wire [WIDTH-1:0] d_out15;
	wire [WIDTH-1:0] d_out16;
	wire [WIDTH-1:0] d_out17;
	wire [WIDTH-1:0] d_out18;
	wire [WIDTH-1:0] d_out19;
	wire [WIDTH-1:0] d_out20;
	wire [WIDTH-1:0] d_out21;
	wire [WIDTH-1:0] d_out22;
	wire [WIDTH-1:0] d_out23;
	wire [WIDTH-1:0] d_out24;
	wire [WIDTH-1:0] d_out25;
	wire [WIDTH-1:0] d_out26;
	wire [WIDTH-1:0] d_out27;
	wire [WIDTH-1:0] d_out28;
	wire [WIDTH-1:0] d_out29;
	wire [WIDTH-1:0] d_out30;
	wire [WIDTH-1:0] d_out31;
	wire [WIDTH-1:0] d_out32;
	wire [WIDTH-1:0] d_out33;
	wire [WIDTH-1:0] d_out34;
	wire [WIDTH-1:0] d_out35;
	wire [WIDTH-1:0] d_out36;
	wire [WIDTH-1:0] d_out37;
	wire [WIDTH-1:0] d_out38;
	wire [WIDTH-1:0] d_out39;
	wire [WIDTH-1:0] d_out40;
	wire [WIDTH-1:0] d_out41;
	wire [WIDTH-1:0] d_out42;
	wire [WIDTH-1:0] d_out43;
	wire [WIDTH-1:0] d_out44;
	wire [WIDTH-1:0] d_out45;
	wire [WIDTH-1:0] d_out46;
	wire [WIDTH-1:0] d_out47;
	wire [WIDTH-1:0] d_out48;
	wire [WIDTH-1:0] d_out49;
	wire [WIDTH-1:0] d_out50;
	wire [WIDTH-1:0] d_out51;
	wire [WIDTH-1:0] d_out52;
	wire [WIDTH-1:0] d_out53;
	wire [WIDTH-1:0] d_out54;
	wire [WIDTH-1:0] d_out55;
	wire [WIDTH-1:0] d_out56;
	wire [WIDTH-1:0] d_out57;
	wire [WIDTH-1:0] d_out58;
	wire [WIDTH-1:0] d_out59;
	wire [WIDTH-1:0] d_out60;
	wire [WIDTH-1:0] d_out61;
	wire [WIDTH-1:0] d_out62;
	wire [WIDTH-1:0] d_out63;
	wire [WIDTH-1:0] d_out64;
	wire [WIDTH-1:0] d_out65;
	wire [WIDTH-1:0] d_out66;
	wire [WIDTH-1:0] d_out67;
	wire [WIDTH-1:0] d_out68;
	wire [WIDTH-1:0] d_out69;
	wire [WIDTH-1:0] d_out70;
	wire [WIDTH-1:0] d_out71;
	wire [WIDTH-1:0] d_out72;
	wire [WIDTH-1:0] d_out73;
	wire [WIDTH-1:0] d_out74;
	wire [WIDTH-1:0] d_out75;
	wire [WIDTH-1:0] d_out76;
	wire [WIDTH-1:0] d_out77;
	wire [WIDTH-1:0] d_out78;
	wire [WIDTH-1:0] d_out79;
	wire [WIDTH-1:0] d_out80;
	wire [WIDTH-1:0] d_out81;
	wire [WIDTH-1:0] d_out82;
	wire [WIDTH-1:0] d_out83;
	wire [WIDTH-1:0] d_out84;
	wire [WIDTH-1:0] d_out85;
	wire [WIDTH-1:0] d_out86;
	wire [WIDTH-1:0] d_out87;
	wire [WIDTH-1:0] d_out88;
	wire [WIDTH-1:0] d_out89;
	wire [WIDTH-1:0] d_out90;
	wire [WIDTH-1:0] d_out91;
	wire [WIDTH-1:0] d_out92;
	wire [WIDTH-1:0] d_out93;
	wire [WIDTH-1:0] d_out94;
	wire [WIDTH-1:0] d_out95;
	wire [WIDTH-1:0] d_out96;
	wire [WIDTH-1:0] d_out97;
	wire [WIDTH-1:0] d_out98;
	wire [WIDTH-1:0] d_out99;

	reg [OUT_BUS-1:0] tmp;

	always @ (posedge clk or posedge rst) begin
		if (rst)
			tmp <= 0;
		else
			tmp <= {tmp[OUT_BUS-(WIDTH-1):0],in};
	end

	always @ (posedge clk) begin
		d_in0 <= tmp[WIDTH-1:0];
		d_in1 <= tmp[(WIDTH*2)-1:WIDTH*1];
		d_in2 <= tmp[(WIDTH*3)-1:WIDTH*2];
		d_in3 <= tmp[(WIDTH*4)-1:WIDTH*3];
		d_in4 <= tmp[(WIDTH*5)-1:WIDTH*4];
		d_in5 <= tmp[(WIDTH*6)-1:WIDTH*5];
		d_in6 <= tmp[(WIDTH*7)-1:WIDTH*6];
		d_in7 <= tmp[(WIDTH*8)-1:WIDTH*7];
		d_in8 <= tmp[(WIDTH*9)-1:WIDTH*8];
		d_in9 <= tmp[(WIDTH*10)-1:WIDTH*9];
		d_in10 <= tmp[(WIDTH*11)-1:WIDTH*10];
		d_in11 <= tmp[(WIDTH*12)-1:WIDTH*11];
		d_in12 <= tmp[(WIDTH*13)-1:WIDTH*12];
		d_in13 <= tmp[(WIDTH*14)-1:WIDTH*13];
		d_in14 <= tmp[(WIDTH*15)-1:WIDTH*14];
		d_in15 <= tmp[(WIDTH*16)-1:WIDTH*15];
		d_in16 <= tmp[(WIDTH*17)-1:WIDTH*16];
		d_in17 <= tmp[(WIDTH*18)-1:WIDTH*17];
		d_in18 <= tmp[(WIDTH*19)-1:WIDTH*18];
		d_in19 <= tmp[(WIDTH*20)-1:WIDTH*19];
		d_in20 <= tmp[(WIDTH*21)-1:WIDTH*20];
		d_in21 <= tmp[(WIDTH*22)-1:WIDTH*21];
		d_in22 <= tmp[(WIDTH*23)-1:WIDTH*22];
		d_in23 <= tmp[(WIDTH*24)-1:WIDTH*23];
		d_in24 <= tmp[(WIDTH*25)-1:WIDTH*24];
		d_in25 <= tmp[(WIDTH*26)-1:WIDTH*25];
		d_in26 <= tmp[(WIDTH*27)-1:WIDTH*26];
		d_in27 <= tmp[(WIDTH*28)-1:WIDTH*27];
		d_in28 <= tmp[(WIDTH*29)-1:WIDTH*28];
		d_in29 <= tmp[(WIDTH*30)-1:WIDTH*29];
		d_in30 <= tmp[(WIDTH*31)-1:WIDTH*30];
		d_in31 <= tmp[(WIDTH*32)-1:WIDTH*31];
		d_in32 <= tmp[(WIDTH*33)-1:WIDTH*32];
		d_in33 <= tmp[(WIDTH*34)-1:WIDTH*33];
		d_in34 <= tmp[(WIDTH*35)-1:WIDTH*34];
		d_in35 <= tmp[(WIDTH*36)-1:WIDTH*35];
		d_in36 <= tmp[(WIDTH*37)-1:WIDTH*36];
		d_in37 <= tmp[(WIDTH*38)-1:WIDTH*37];
		d_in38 <= tmp[(WIDTH*39)-1:WIDTH*38];
		d_in39 <= tmp[(WIDTH*40)-1:WIDTH*39];
		d_in40 <= tmp[(WIDTH*41)-1:WIDTH*40];
		d_in41 <= tmp[(WIDTH*42)-1:WIDTH*41];
		d_in42 <= tmp[(WIDTH*43)-1:WIDTH*42];
		d_in43 <= tmp[(WIDTH*44)-1:WIDTH*43];
		d_in44 <= tmp[(WIDTH*45)-1:WIDTH*44];
		d_in45 <= tmp[(WIDTH*46)-1:WIDTH*45];
		d_in46 <= tmp[(WIDTH*47)-1:WIDTH*46];
		d_in47 <= tmp[(WIDTH*48)-1:WIDTH*47];
		d_in48 <= tmp[(WIDTH*49)-1:WIDTH*48];
		d_in49 <= tmp[(WIDTH*50)-1:WIDTH*49];
		d_in50 <= tmp[(WIDTH*51)-1:WIDTH*50];
		d_in51 <= tmp[(WIDTH*52)-1:WIDTH*51];
		d_in52 <= tmp[(WIDTH*53)-1:WIDTH*52];
		d_in53 <= tmp[(WIDTH*54)-1:WIDTH*53];
		d_in54 <= tmp[(WIDTH*55)-1:WIDTH*54];
		d_in55 <= tmp[(WIDTH*56)-1:WIDTH*55];
		d_in56 <= tmp[(WIDTH*57)-1:WIDTH*56];
		d_in57 <= tmp[(WIDTH*58)-1:WIDTH*57];
		d_in58 <= tmp[(WIDTH*59)-1:WIDTH*58];
		d_in59 <= tmp[(WIDTH*60)-1:WIDTH*59];
		d_in60 <= tmp[(WIDTH*61)-1:WIDTH*60];
		d_in61 <= tmp[(WIDTH*62)-1:WIDTH*61];
		d_in62 <= tmp[(WIDTH*63)-1:WIDTH*62];
		d_in63 <= tmp[(WIDTH*64)-1:WIDTH*63];
		d_in64 <= tmp[(WIDTH*65)-1:WIDTH*64];
		d_in65 <= tmp[(WIDTH*66)-1:WIDTH*65];
		d_in66 <= tmp[(WIDTH*67)-1:WIDTH*66];
		d_in67 <= tmp[(WIDTH*68)-1:WIDTH*67];
		d_in68 <= tmp[(WIDTH*69)-1:WIDTH*68];
		d_in69 <= tmp[(WIDTH*70)-1:WIDTH*69];
		d_in70 <= tmp[(WIDTH*71)-1:WIDTH*70];
		d_in71 <= tmp[(WIDTH*72)-1:WIDTH*71];
		d_in72 <= tmp[(WIDTH*73)-1:WIDTH*72];
		d_in73 <= tmp[(WIDTH*74)-1:WIDTH*73];
		d_in74 <= tmp[(WIDTH*75)-1:WIDTH*74];
		d_in75 <= tmp[(WIDTH*76)-1:WIDTH*75];
		d_in76 <= tmp[(WIDTH*77)-1:WIDTH*76];
		d_in77 <= tmp[(WIDTH*78)-1:WIDTH*77];
		d_in78 <= tmp[(WIDTH*79)-1:WIDTH*78];
		d_in79 <= tmp[(WIDTH*80)-1:WIDTH*79];
		d_in80 <= tmp[(WIDTH*81)-1:WIDTH*80];
		d_in81 <= tmp[(WIDTH*82)-1:WIDTH*81];
		d_in82 <= tmp[(WIDTH*83)-1:WIDTH*82];
		d_in83 <= tmp[(WIDTH*84)-1:WIDTH*83];
		d_in84 <= tmp[(WIDTH*85)-1:WIDTH*84];
		d_in85 <= tmp[(WIDTH*86)-1:WIDTH*85];
		d_in86 <= tmp[(WIDTH*87)-1:WIDTH*86];
		d_in87 <= tmp[(WIDTH*88)-1:WIDTH*87];
		d_in88 <= tmp[(WIDTH*89)-1:WIDTH*88];
		d_in89 <= tmp[(WIDTH*90)-1:WIDTH*89];
		d_in90 <= tmp[(WIDTH*91)-1:WIDTH*90];
		d_in91 <= tmp[(WIDTH*92)-1:WIDTH*91];
		d_in92 <= tmp[(WIDTH*93)-1:WIDTH*92];
		d_in93 <= tmp[(WIDTH*94)-1:WIDTH*93];
		d_in94 <= tmp[(WIDTH*95)-1:WIDTH*94];
		d_in95 <= tmp[(WIDTH*96)-1:WIDTH*95];
		d_in96 <= tmp[(WIDTH*97)-1:WIDTH*96];
		d_in97 <= tmp[(WIDTH*98)-1:WIDTH*97];
		d_in98 <= tmp[(WIDTH*99)-1:WIDTH*98];
		d_in99 <= tmp[(WIDTH*100)-1:WIDTH*99];
	end

	design210_100_120 #(.WIDTH(WIDTH)) design210_100_120_inst(.d_in0(d_in0),.d_in1(d_in1),.d_in2(d_in2),.d_in3(d_in3),.d_in4(d_in4),.d_in5(d_in5),.d_in6(d_in6),.d_in7(d_in7),.d_in8(d_in8),.d_in9(d_in9),.d_in10(d_in10),.d_in11(d_in11),.d_in12(d_in12),.d_in13(d_in13),.d_in14(d_in14),.d_in15(d_in15),.d_in16(d_in16),.d_in17(d_in17),.d_in18(d_in18),.d_in19(d_in19),.d_in20(d_in20),.d_in21(d_in21),.d_in22(d_in22),.d_in23(d_in23),.d_in24(d_in24),.d_in25(d_in25),.d_in26(d_in26),.d_in27(d_in27),.d_in28(d_in28),.d_in29(d_in29),.d_in30(d_in30),.d_in31(d_in31),.d_in32(d_in32),.d_in33(d_in33),.d_in34(d_in34),.d_in35(d_in35),.d_in36(d_in36),.d_in37(d_in37),.d_in38(d_in38),.d_in39(d_in39),.d_in40(d_in40),.d_in41(d_in41),.d_in42(d_in42),.d_in43(d_in43),.d_in44(d_in44),.d_in45(d_in45),.d_in46(d_in46),.d_in47(d_in47),.d_in48(d_in48),.d_in49(d_in49),.d_in50(d_in50),.d_in51(d_in51),.d_in52(d_in52),.d_in53(d_in53),.d_in54(d_in54),.d_in55(d_in55),.d_in56(d_in56),.d_in57(d_in57),.d_in58(d_in58),.d_in59(d_in59),.d_in60(d_in60),.d_in61(d_in61),.d_in62(d_in62),.d_in63(d_in63),.d_in64(d_in64),.d_in65(d_in65),.d_in66(d_in66),.d_in67(d_in67),.d_in68(d_in68),.d_in69(d_in69),.d_in70(d_in70),.d_in71(d_in71),.d_in72(d_in72),.d_in73(d_in73),.d_in74(d_in74),.d_in75(d_in75),.d_in76(d_in76),.d_in77(d_in77),.d_in78(d_in78),.d_in79(d_in79),.d_in80(d_in80),.d_in81(d_in81),.d_in82(d_in82),.d_in83(d_in83),.d_in84(d_in84),.d_in85(d_in85),.d_in86(d_in86),.d_in87(d_in87),.d_in88(d_in88),.d_in89(d_in89),.d_in90(d_in90),.d_in91(d_in91),.d_in92(d_in92),.d_in93(d_in93),.d_in94(d_in94),.d_in95(d_in95),.d_in96(d_in96),.d_in97(d_in97),.d_in98(d_in98),.d_in99(d_in99),.d_out0(d_out0),.d_out1(d_out1),.d_out2(d_out2),.d_out3(d_out3),.d_out4(d_out4),.d_out5(d_out5),.d_out6(d_out6),.d_out7(d_out7),.d_out8(d_out8),.d_out9(d_out9),.d_out10(d_out10),.d_out11(d_out11),.d_out12(d_out12),.d_out13(d_out13),.d_out14(d_out14),.d_out15(d_out15),.d_out16(d_out16),.d_out17(d_out17),.d_out18(d_out18),.d_out19(d_out19),.d_out20(d_out20),.d_out21(d_out21),.d_out22(d_out22),.d_out23(d_out23),.d_out24(d_out24),.d_out25(d_out25),.d_out26(d_out26),.d_out27(d_out27),.d_out28(d_out28),.d_out29(d_out29),.d_out30(d_out30),.d_out31(d_out31),.d_out32(d_out32),.d_out33(d_out33),.d_out34(d_out34),.d_out35(d_out35),.d_out36(d_out36),.d_out37(d_out37),.d_out38(d_out38),.d_out39(d_out39),.d_out40(d_out40),.d_out41(d_out41),.d_out42(d_out42),.d_out43(d_out43),.d_out44(d_out44),.d_out45(d_out45),.d_out46(d_out46),.d_out47(d_out47),.d_out48(d_out48),.d_out49(d_out49),.d_out50(d_out50),.d_out51(d_out51),.d_out52(d_out52),.d_out53(d_out53),.d_out54(d_out54),.d_out55(d_out55),.d_out56(d_out56),.d_out57(d_out57),.d_out58(d_out58),.d_out59(d_out59),.d_out60(d_out60),.d_out61(d_out61),.d_out62(d_out62),.d_out63(d_out63),.d_out64(d_out64),.d_out65(d_out65),.d_out66(d_out66),.d_out67(d_out67),.d_out68(d_out68),.d_out69(d_out69),.d_out70(d_out70),.d_out71(d_out71),.d_out72(d_out72),.d_out73(d_out73),.d_out74(d_out74),.d_out75(d_out75),.d_out76(d_out76),.d_out77(d_out77),.d_out78(d_out78),.d_out79(d_out79),.d_out80(d_out80),.d_out81(d_out81),.d_out82(d_out82),.d_out83(d_out83),.d_out84(d_out84),.d_out85(d_out85),.d_out86(d_out86),.d_out87(d_out87),.d_out88(d_out88),.d_out89(d_out89),.d_out90(d_out90),.d_out91(d_out91),.d_out92(d_out92),.d_out93(d_out93),.d_out94(d_out94),.d_out95(d_out95),.d_out96(d_out96),.d_out97(d_out97),.d_out98(d_out98),.d_out99(d_out99),.clk(clk),.rst(rst));

	assign out = d_out0^d_out1^d_out2^d_out3^d_out4^d_out5^d_out6^d_out7^d_out8^d_out9^d_out10^d_out11^d_out12^d_out13^d_out14^d_out15^d_out16^d_out17^d_out18^d_out19^d_out20^d_out21^d_out22^d_out23^d_out24^d_out25^d_out26^d_out27^d_out28^d_out29^d_out30^d_out31^d_out32^d_out33^d_out34^d_out35^d_out36^d_out37^d_out38^d_out39^d_out40^d_out41^d_out42^d_out43^d_out44^d_out45^d_out46^d_out47^d_out48^d_out49^d_out50^d_out51^d_out52^d_out53^d_out54^d_out55^d_out56^d_out57^d_out58^d_out59^d_out60^d_out61^d_out62^d_out63^d_out64^d_out65^d_out66^d_out67^d_out68^d_out69^d_out70^d_out71^d_out72^d_out73^d_out74^d_out75^d_out76^d_out77^d_out78^d_out79^d_out80^d_out81^d_out82^d_out83^d_out84^d_out85^d_out86^d_out87^d_out88^d_out89^d_out90^d_out91^d_out92^d_out93^d_out94^d_out95^d_out96^d_out97^d_out98^d_out99;

endmodule

module design210_100_120 #(parameter WIDTH=32) (d_in0, d_in1, d_in2, d_in3, d_in4, d_in5, d_in6, d_in7, d_in8, d_in9, d_in10, d_in11, d_in12, d_in13, d_in14, d_in15, d_in16, d_in17, d_in18, d_in19, d_in20, d_in21, d_in22, d_in23, d_in24, d_in25, d_in26, d_in27, d_in28, d_in29, d_in30, d_in31, d_in32, d_in33, d_in34, d_in35, d_in36, d_in37, d_in38, d_in39, d_in40, d_in41, d_in42, d_in43, d_in44, d_in45, d_in46, d_in47, d_in48, d_in49, d_in50, d_in51, d_in52, d_in53, d_in54, d_in55, d_in56, d_in57, d_in58, d_in59, d_in60, d_in61, d_in62, d_in63, d_in64, d_in65, d_in66, d_in67, d_in68, d_in69, d_in70, d_in71, d_in72, d_in73, d_in74, d_in75, d_in76, d_in77, d_in78, d_in79, d_in80, d_in81, d_in82, d_in83, d_in84, d_in85, d_in86, d_in87, d_in88, d_in89, d_in90, d_in91, d_in92, d_in93, d_in94, d_in95, d_in96, d_in97, d_in98, d_in99, d_out0, d_out1, d_out2, d_out3, d_out4, d_out5, d_out6, d_out7, d_out8, d_out9, d_out10, d_out11, d_out12, d_out13, d_out14, d_out15, d_out16, d_out17, d_out18, d_out19, d_out20, d_out21, d_out22, d_out23, d_out24, d_out25, d_out26, d_out27, d_out28, d_out29, d_out30, d_out31, d_out32, d_out33, d_out34, d_out35, d_out36, d_out37, d_out38, d_out39, d_out40, d_out41, d_out42, d_out43, d_out44, d_out45, d_out46, d_out47, d_out48, d_out49, d_out50, d_out51, d_out52, d_out53, d_out54, d_out55, d_out56, d_out57, d_out58, d_out59, d_out60, d_out61, d_out62, d_out63, d_out64, d_out65, d_out66, d_out67, d_out68, d_out69, d_out70, d_out71, d_out72, d_out73, d_out74, d_out75, d_out76, d_out77, d_out78, d_out79, d_out80, d_out81, d_out82, d_out83, d_out84, d_out85, d_out86, d_out87, d_out88, d_out89, d_out90, d_out91, d_out92, d_out93, d_out94, d_out95, d_out96, d_out97, d_out98, d_out99, clk, rst);
	input clk;
	input rst;
	input [WIDTH-1:0] d_in0; 
	input [WIDTH-1:0] d_in1; 
	input [WIDTH-1:0] d_in2; 
	input [WIDTH-1:0] d_in3; 
	input [WIDTH-1:0] d_in4; 
	input [WIDTH-1:0] d_in5; 
	input [WIDTH-1:0] d_in6; 
	input [WIDTH-1:0] d_in7; 
	input [WIDTH-1:0] d_in8; 
	input [WIDTH-1:0] d_in9; 
	input [WIDTH-1:0] d_in10; 
	input [WIDTH-1:0] d_in11; 
	input [WIDTH-1:0] d_in12; 
	input [WIDTH-1:0] d_in13; 
	input [WIDTH-1:0] d_in14; 
	input [WIDTH-1:0] d_in15; 
	input [WIDTH-1:0] d_in16; 
	input [WIDTH-1:0] d_in17; 
	input [WIDTH-1:0] d_in18; 
	input [WIDTH-1:0] d_in19; 
	input [WIDTH-1:0] d_in20; 
	input [WIDTH-1:0] d_in21; 
	input [WIDTH-1:0] d_in22; 
	input [WIDTH-1:0] d_in23; 
	input [WIDTH-1:0] d_in24; 
	input [WIDTH-1:0] d_in25; 
	input [WIDTH-1:0] d_in26; 
	input [WIDTH-1:0] d_in27; 
	input [WIDTH-1:0] d_in28; 
	input [WIDTH-1:0] d_in29; 
	input [WIDTH-1:0] d_in30; 
	input [WIDTH-1:0] d_in31; 
	input [WIDTH-1:0] d_in32; 
	input [WIDTH-1:0] d_in33; 
	input [WIDTH-1:0] d_in34; 
	input [WIDTH-1:0] d_in35; 
	input [WIDTH-1:0] d_in36; 
	input [WIDTH-1:0] d_in37; 
	input [WIDTH-1:0] d_in38; 
	input [WIDTH-1:0] d_in39; 
	input [WIDTH-1:0] d_in40; 
	input [WIDTH-1:0] d_in41; 
	input [WIDTH-1:0] d_in42; 
	input [WIDTH-1:0] d_in43; 
	input [WIDTH-1:0] d_in44; 
	input [WIDTH-1:0] d_in45; 
	input [WIDTH-1:0] d_in46; 
	input [WIDTH-1:0] d_in47; 
	input [WIDTH-1:0] d_in48; 
	input [WIDTH-1:0] d_in49; 
	input [WIDTH-1:0] d_in50; 
	input [WIDTH-1:0] d_in51; 
	input [WIDTH-1:0] d_in52; 
	input [WIDTH-1:0] d_in53; 
	input [WIDTH-1:0] d_in54; 
	input [WIDTH-1:0] d_in55; 
	input [WIDTH-1:0] d_in56; 
	input [WIDTH-1:0] d_in57; 
	input [WIDTH-1:0] d_in58; 
	input [WIDTH-1:0] d_in59; 
	input [WIDTH-1:0] d_in60; 
	input [WIDTH-1:0] d_in61; 
	input [WIDTH-1:0] d_in62; 
	input [WIDTH-1:0] d_in63; 
	input [WIDTH-1:0] d_in64; 
	input [WIDTH-1:0] d_in65; 
	input [WIDTH-1:0] d_in66; 
	input [WIDTH-1:0] d_in67; 
	input [WIDTH-1:0] d_in68; 
	input [WIDTH-1:0] d_in69; 
	input [WIDTH-1:0] d_in70; 
	input [WIDTH-1:0] d_in71; 
	input [WIDTH-1:0] d_in72; 
	input [WIDTH-1:0] d_in73; 
	input [WIDTH-1:0] d_in74; 
	input [WIDTH-1:0] d_in75; 
	input [WIDTH-1:0] d_in76; 
	input [WIDTH-1:0] d_in77; 
	input [WIDTH-1:0] d_in78; 
	input [WIDTH-1:0] d_in79; 
	input [WIDTH-1:0] d_in80; 
	input [WIDTH-1:0] d_in81; 
	input [WIDTH-1:0] d_in82; 
	input [WIDTH-1:0] d_in83; 
	input [WIDTH-1:0] d_in84; 
	input [WIDTH-1:0] d_in85; 
	input [WIDTH-1:0] d_in86; 
	input [WIDTH-1:0] d_in87; 
	input [WIDTH-1:0] d_in88; 
	input [WIDTH-1:0] d_in89; 
	input [WIDTH-1:0] d_in90; 
	input [WIDTH-1:0] d_in91; 
	input [WIDTH-1:0] d_in92; 
	input [WIDTH-1:0] d_in93; 
	input [WIDTH-1:0] d_in94; 
	input [WIDTH-1:0] d_in95; 
	input [WIDTH-1:0] d_in96; 
	input [WIDTH-1:0] d_in97; 
	input [WIDTH-1:0] d_in98; 
	input [WIDTH-1:0] d_in99; 
	output [WIDTH-1:0] d_out0; 
	output [WIDTH-1:0] d_out1; 
	output [WIDTH-1:0] d_out2; 
	output [WIDTH-1:0] d_out3; 
	output [WIDTH-1:0] d_out4; 
	output [WIDTH-1:0] d_out5; 
	output [WIDTH-1:0] d_out6; 
	output [WIDTH-1:0] d_out7; 
	output [WIDTH-1:0] d_out8; 
	output [WIDTH-1:0] d_out9; 
	output [WIDTH-1:0] d_out10; 
	output [WIDTH-1:0] d_out11; 
	output [WIDTH-1:0] d_out12; 
	output [WIDTH-1:0] d_out13; 
	output [WIDTH-1:0] d_out14; 
	output [WIDTH-1:0] d_out15; 
	output [WIDTH-1:0] d_out16; 
	output [WIDTH-1:0] d_out17; 
	output [WIDTH-1:0] d_out18; 
	output [WIDTH-1:0] d_out19; 
	output [WIDTH-1:0] d_out20; 
	output [WIDTH-1:0] d_out21; 
	output [WIDTH-1:0] d_out22; 
	output [WIDTH-1:0] d_out23; 
	output [WIDTH-1:0] d_out24; 
	output [WIDTH-1:0] d_out25; 
	output [WIDTH-1:0] d_out26; 
	output [WIDTH-1:0] d_out27; 
	output [WIDTH-1:0] d_out28; 
	output [WIDTH-1:0] d_out29; 
	output [WIDTH-1:0] d_out30; 
	output [WIDTH-1:0] d_out31; 
	output [WIDTH-1:0] d_out32; 
	output [WIDTH-1:0] d_out33; 
	output [WIDTH-1:0] d_out34; 
	output [WIDTH-1:0] d_out35; 
	output [WIDTH-1:0] d_out36; 
	output [WIDTH-1:0] d_out37; 
	output [WIDTH-1:0] d_out38; 
	output [WIDTH-1:0] d_out39; 
	output [WIDTH-1:0] d_out40; 
	output [WIDTH-1:0] d_out41; 
	output [WIDTH-1:0] d_out42; 
	output [WIDTH-1:0] d_out43; 
	output [WIDTH-1:0] d_out44; 
	output [WIDTH-1:0] d_out45; 
	output [WIDTH-1:0] d_out46; 
	output [WIDTH-1:0] d_out47; 
	output [WIDTH-1:0] d_out48; 
	output [WIDTH-1:0] d_out49; 
	output [WIDTH-1:0] d_out50; 
	output [WIDTH-1:0] d_out51; 
	output [WIDTH-1:0] d_out52; 
	output [WIDTH-1:0] d_out53; 
	output [WIDTH-1:0] d_out54; 
	output [WIDTH-1:0] d_out55; 
	output [WIDTH-1:0] d_out56; 
	output [WIDTH-1:0] d_out57; 
	output [WIDTH-1:0] d_out58; 
	output [WIDTH-1:0] d_out59; 
	output [WIDTH-1:0] d_out60; 
	output [WIDTH-1:0] d_out61; 
	output [WIDTH-1:0] d_out62; 
	output [WIDTH-1:0] d_out63; 
	output [WIDTH-1:0] d_out64; 
	output [WIDTH-1:0] d_out65; 
	output [WIDTH-1:0] d_out66; 
	output [WIDTH-1:0] d_out67; 
	output [WIDTH-1:0] d_out68; 
	output [WIDTH-1:0] d_out69; 
	output [WIDTH-1:0] d_out70; 
	output [WIDTH-1:0] d_out71; 
	output [WIDTH-1:0] d_out72; 
	output [WIDTH-1:0] d_out73; 
	output [WIDTH-1:0] d_out74; 
	output [WIDTH-1:0] d_out75; 
	output [WIDTH-1:0] d_out76; 
	output [WIDTH-1:0] d_out77; 
	output [WIDTH-1:0] d_out78; 
	output [WIDTH-1:0] d_out79; 
	output [WIDTH-1:0] d_out80; 
	output [WIDTH-1:0] d_out81; 
	output [WIDTH-1:0] d_out82; 
	output [WIDTH-1:0] d_out83; 
	output [WIDTH-1:0] d_out84; 
	output [WIDTH-1:0] d_out85; 
	output [WIDTH-1:0] d_out86; 
	output [WIDTH-1:0] d_out87; 
	output [WIDTH-1:0] d_out88; 
	output [WIDTH-1:0] d_out89; 
	output [WIDTH-1:0] d_out90; 
	output [WIDTH-1:0] d_out91; 
	output [WIDTH-1:0] d_out92; 
	output [WIDTH-1:0] d_out93; 
	output [WIDTH-1:0] d_out94; 
	output [WIDTH-1:0] d_out95; 
	output [WIDTH-1:0] d_out96; 
	output [WIDTH-1:0] d_out97; 
	output [WIDTH-1:0] d_out98; 
	output [WIDTH-1:0] d_out99; 

	wire [WIDTH-1:0] wire_d0_0;
	wire [WIDTH-1:0] wire_d0_1;
	wire [WIDTH-1:0] wire_d0_2;
	wire [WIDTH-1:0] wire_d0_3;
	wire [WIDTH-1:0] wire_d0_4;
	wire [WIDTH-1:0] wire_d0_5;
	wire [WIDTH-1:0] wire_d0_6;
	wire [WIDTH-1:0] wire_d0_7;
	wire [WIDTH-1:0] wire_d0_8;
	wire [WIDTH-1:0] wire_d0_9;
	wire [WIDTH-1:0] wire_d0_10;
	wire [WIDTH-1:0] wire_d0_11;
	wire [WIDTH-1:0] wire_d0_12;
	wire [WIDTH-1:0] wire_d0_13;
	wire [WIDTH-1:0] wire_d0_14;
	wire [WIDTH-1:0] wire_d0_15;
	wire [WIDTH-1:0] wire_d0_16;
	wire [WIDTH-1:0] wire_d0_17;
	wire [WIDTH-1:0] wire_d0_18;
	wire [WIDTH-1:0] wire_d0_19;
	wire [WIDTH-1:0] wire_d0_20;
	wire [WIDTH-1:0] wire_d0_21;
	wire [WIDTH-1:0] wire_d0_22;
	wire [WIDTH-1:0] wire_d0_23;
	wire [WIDTH-1:0] wire_d0_24;
	wire [WIDTH-1:0] wire_d0_25;
	wire [WIDTH-1:0] wire_d0_26;
	wire [WIDTH-1:0] wire_d0_27;
	wire [WIDTH-1:0] wire_d0_28;
	wire [WIDTH-1:0] wire_d0_29;
	wire [WIDTH-1:0] wire_d0_30;
	wire [WIDTH-1:0] wire_d0_31;
	wire [WIDTH-1:0] wire_d0_32;
	wire [WIDTH-1:0] wire_d0_33;
	wire [WIDTH-1:0] wire_d0_34;
	wire [WIDTH-1:0] wire_d0_35;
	wire [WIDTH-1:0] wire_d0_36;
	wire [WIDTH-1:0] wire_d0_37;
	wire [WIDTH-1:0] wire_d0_38;
	wire [WIDTH-1:0] wire_d0_39;
	wire [WIDTH-1:0] wire_d0_40;
	wire [WIDTH-1:0] wire_d0_41;
	wire [WIDTH-1:0] wire_d0_42;
	wire [WIDTH-1:0] wire_d0_43;
	wire [WIDTH-1:0] wire_d0_44;
	wire [WIDTH-1:0] wire_d0_45;
	wire [WIDTH-1:0] wire_d0_46;
	wire [WIDTH-1:0] wire_d0_47;
	wire [WIDTH-1:0] wire_d0_48;
	wire [WIDTH-1:0] wire_d0_49;
	wire [WIDTH-1:0] wire_d0_50;
	wire [WIDTH-1:0] wire_d0_51;
	wire [WIDTH-1:0] wire_d0_52;
	wire [WIDTH-1:0] wire_d0_53;
	wire [WIDTH-1:0] wire_d0_54;
	wire [WIDTH-1:0] wire_d0_55;
	wire [WIDTH-1:0] wire_d0_56;
	wire [WIDTH-1:0] wire_d0_57;
	wire [WIDTH-1:0] wire_d0_58;
	wire [WIDTH-1:0] wire_d0_59;
	wire [WIDTH-1:0] wire_d0_60;
	wire [WIDTH-1:0] wire_d0_61;
	wire [WIDTH-1:0] wire_d0_62;
	wire [WIDTH-1:0] wire_d0_63;
	wire [WIDTH-1:0] wire_d0_64;
	wire [WIDTH-1:0] wire_d0_65;
	wire [WIDTH-1:0] wire_d0_66;
	wire [WIDTH-1:0] wire_d0_67;
	wire [WIDTH-1:0] wire_d0_68;
	wire [WIDTH-1:0] wire_d0_69;
	wire [WIDTH-1:0] wire_d0_70;
	wire [WIDTH-1:0] wire_d0_71;
	wire [WIDTH-1:0] wire_d0_72;
	wire [WIDTH-1:0] wire_d0_73;
	wire [WIDTH-1:0] wire_d0_74;
	wire [WIDTH-1:0] wire_d0_75;
	wire [WIDTH-1:0] wire_d0_76;
	wire [WIDTH-1:0] wire_d0_77;
	wire [WIDTH-1:0] wire_d0_78;
	wire [WIDTH-1:0] wire_d0_79;
	wire [WIDTH-1:0] wire_d0_80;
	wire [WIDTH-1:0] wire_d0_81;
	wire [WIDTH-1:0] wire_d0_82;
	wire [WIDTH-1:0] wire_d0_83;
	wire [WIDTH-1:0] wire_d0_84;
	wire [WIDTH-1:0] wire_d0_85;
	wire [WIDTH-1:0] wire_d0_86;
	wire [WIDTH-1:0] wire_d0_87;
	wire [WIDTH-1:0] wire_d0_88;
	wire [WIDTH-1:0] wire_d0_89;
	wire [WIDTH-1:0] wire_d0_90;
	wire [WIDTH-1:0] wire_d0_91;
	wire [WIDTH-1:0] wire_d0_92;
	wire [WIDTH-1:0] wire_d0_93;
	wire [WIDTH-1:0] wire_d0_94;
	wire [WIDTH-1:0] wire_d0_95;
	wire [WIDTH-1:0] wire_d0_96;
	wire [WIDTH-1:0] wire_d0_97;
	wire [WIDTH-1:0] wire_d0_98;
	wire [WIDTH-1:0] wire_d0_99;
	wire [WIDTH-1:0] wire_d0_100;
	wire [WIDTH-1:0] wire_d0_101;
	wire [WIDTH-1:0] wire_d0_102;
	wire [WIDTH-1:0] wire_d0_103;
	wire [WIDTH-1:0] wire_d0_104;
	wire [WIDTH-1:0] wire_d0_105;
	wire [WIDTH-1:0] wire_d0_106;
	wire [WIDTH-1:0] wire_d0_107;
	wire [WIDTH-1:0] wire_d0_108;
	wire [WIDTH-1:0] wire_d0_109;
	wire [WIDTH-1:0] wire_d0_110;
	wire [WIDTH-1:0] wire_d0_111;
	wire [WIDTH-1:0] wire_d0_112;
	wire [WIDTH-1:0] wire_d0_113;
	wire [WIDTH-1:0] wire_d0_114;
	wire [WIDTH-1:0] wire_d0_115;
	wire [WIDTH-1:0] wire_d0_116;
	wire [WIDTH-1:0] wire_d0_117;
	wire [WIDTH-1:0] wire_d0_118;
	wire [WIDTH-1:0] wire_d1_0;
	wire [WIDTH-1:0] wire_d1_1;
	wire [WIDTH-1:0] wire_d1_2;
	wire [WIDTH-1:0] wire_d1_3;
	wire [WIDTH-1:0] wire_d1_4;
	wire [WIDTH-1:0] wire_d1_5;
	wire [WIDTH-1:0] wire_d1_6;
	wire [WIDTH-1:0] wire_d1_7;
	wire [WIDTH-1:0] wire_d1_8;
	wire [WIDTH-1:0] wire_d1_9;
	wire [WIDTH-1:0] wire_d1_10;
	wire [WIDTH-1:0] wire_d1_11;
	wire [WIDTH-1:0] wire_d1_12;
	wire [WIDTH-1:0] wire_d1_13;
	wire [WIDTH-1:0] wire_d1_14;
	wire [WIDTH-1:0] wire_d1_15;
	wire [WIDTH-1:0] wire_d1_16;
	wire [WIDTH-1:0] wire_d1_17;
	wire [WIDTH-1:0] wire_d1_18;
	wire [WIDTH-1:0] wire_d1_19;
	wire [WIDTH-1:0] wire_d1_20;
	wire [WIDTH-1:0] wire_d1_21;
	wire [WIDTH-1:0] wire_d1_22;
	wire [WIDTH-1:0] wire_d1_23;
	wire [WIDTH-1:0] wire_d1_24;
	wire [WIDTH-1:0] wire_d1_25;
	wire [WIDTH-1:0] wire_d1_26;
	wire [WIDTH-1:0] wire_d1_27;
	wire [WIDTH-1:0] wire_d1_28;
	wire [WIDTH-1:0] wire_d1_29;
	wire [WIDTH-1:0] wire_d1_30;
	wire [WIDTH-1:0] wire_d1_31;
	wire [WIDTH-1:0] wire_d1_32;
	wire [WIDTH-1:0] wire_d1_33;
	wire [WIDTH-1:0] wire_d1_34;
	wire [WIDTH-1:0] wire_d1_35;
	wire [WIDTH-1:0] wire_d1_36;
	wire [WIDTH-1:0] wire_d1_37;
	wire [WIDTH-1:0] wire_d1_38;
	wire [WIDTH-1:0] wire_d1_39;
	wire [WIDTH-1:0] wire_d1_40;
	wire [WIDTH-1:0] wire_d1_41;
	wire [WIDTH-1:0] wire_d1_42;
	wire [WIDTH-1:0] wire_d1_43;
	wire [WIDTH-1:0] wire_d1_44;
	wire [WIDTH-1:0] wire_d1_45;
	wire [WIDTH-1:0] wire_d1_46;
	wire [WIDTH-1:0] wire_d1_47;
	wire [WIDTH-1:0] wire_d1_48;
	wire [WIDTH-1:0] wire_d1_49;
	wire [WIDTH-1:0] wire_d1_50;
	wire [WIDTH-1:0] wire_d1_51;
	wire [WIDTH-1:0] wire_d1_52;
	wire [WIDTH-1:0] wire_d1_53;
	wire [WIDTH-1:0] wire_d1_54;
	wire [WIDTH-1:0] wire_d1_55;
	wire [WIDTH-1:0] wire_d1_56;
	wire [WIDTH-1:0] wire_d1_57;
	wire [WIDTH-1:0] wire_d1_58;
	wire [WIDTH-1:0] wire_d1_59;
	wire [WIDTH-1:0] wire_d1_60;
	wire [WIDTH-1:0] wire_d1_61;
	wire [WIDTH-1:0] wire_d1_62;
	wire [WIDTH-1:0] wire_d1_63;
	wire [WIDTH-1:0] wire_d1_64;
	wire [WIDTH-1:0] wire_d1_65;
	wire [WIDTH-1:0] wire_d1_66;
	wire [WIDTH-1:0] wire_d1_67;
	wire [WIDTH-1:0] wire_d1_68;
	wire [WIDTH-1:0] wire_d1_69;
	wire [WIDTH-1:0] wire_d1_70;
	wire [WIDTH-1:0] wire_d1_71;
	wire [WIDTH-1:0] wire_d1_72;
	wire [WIDTH-1:0] wire_d1_73;
	wire [WIDTH-1:0] wire_d1_74;
	wire [WIDTH-1:0] wire_d1_75;
	wire [WIDTH-1:0] wire_d1_76;
	wire [WIDTH-1:0] wire_d1_77;
	wire [WIDTH-1:0] wire_d1_78;
	wire [WIDTH-1:0] wire_d1_79;
	wire [WIDTH-1:0] wire_d1_80;
	wire [WIDTH-1:0] wire_d1_81;
	wire [WIDTH-1:0] wire_d1_82;
	wire [WIDTH-1:0] wire_d1_83;
	wire [WIDTH-1:0] wire_d1_84;
	wire [WIDTH-1:0] wire_d1_85;
	wire [WIDTH-1:0] wire_d1_86;
	wire [WIDTH-1:0] wire_d1_87;
	wire [WIDTH-1:0] wire_d1_88;
	wire [WIDTH-1:0] wire_d1_89;
	wire [WIDTH-1:0] wire_d1_90;
	wire [WIDTH-1:0] wire_d1_91;
	wire [WIDTH-1:0] wire_d1_92;
	wire [WIDTH-1:0] wire_d1_93;
	wire [WIDTH-1:0] wire_d1_94;
	wire [WIDTH-1:0] wire_d1_95;
	wire [WIDTH-1:0] wire_d1_96;
	wire [WIDTH-1:0] wire_d1_97;
	wire [WIDTH-1:0] wire_d1_98;
	wire [WIDTH-1:0] wire_d1_99;
	wire [WIDTH-1:0] wire_d1_100;
	wire [WIDTH-1:0] wire_d1_101;
	wire [WIDTH-1:0] wire_d1_102;
	wire [WIDTH-1:0] wire_d1_103;
	wire [WIDTH-1:0] wire_d1_104;
	wire [WIDTH-1:0] wire_d1_105;
	wire [WIDTH-1:0] wire_d1_106;
	wire [WIDTH-1:0] wire_d1_107;
	wire [WIDTH-1:0] wire_d1_108;
	wire [WIDTH-1:0] wire_d1_109;
	wire [WIDTH-1:0] wire_d1_110;
	wire [WIDTH-1:0] wire_d1_111;
	wire [WIDTH-1:0] wire_d1_112;
	wire [WIDTH-1:0] wire_d1_113;
	wire [WIDTH-1:0] wire_d1_114;
	wire [WIDTH-1:0] wire_d1_115;
	wire [WIDTH-1:0] wire_d1_116;
	wire [WIDTH-1:0] wire_d1_117;
	wire [WIDTH-1:0] wire_d1_118;
	wire [WIDTH-1:0] wire_d2_0;
	wire [WIDTH-1:0] wire_d2_1;
	wire [WIDTH-1:0] wire_d2_2;
	wire [WIDTH-1:0] wire_d2_3;
	wire [WIDTH-1:0] wire_d2_4;
	wire [WIDTH-1:0] wire_d2_5;
	wire [WIDTH-1:0] wire_d2_6;
	wire [WIDTH-1:0] wire_d2_7;
	wire [WIDTH-1:0] wire_d2_8;
	wire [WIDTH-1:0] wire_d2_9;
	wire [WIDTH-1:0] wire_d2_10;
	wire [WIDTH-1:0] wire_d2_11;
	wire [WIDTH-1:0] wire_d2_12;
	wire [WIDTH-1:0] wire_d2_13;
	wire [WIDTH-1:0] wire_d2_14;
	wire [WIDTH-1:0] wire_d2_15;
	wire [WIDTH-1:0] wire_d2_16;
	wire [WIDTH-1:0] wire_d2_17;
	wire [WIDTH-1:0] wire_d2_18;
	wire [WIDTH-1:0] wire_d2_19;
	wire [WIDTH-1:0] wire_d2_20;
	wire [WIDTH-1:0] wire_d2_21;
	wire [WIDTH-1:0] wire_d2_22;
	wire [WIDTH-1:0] wire_d2_23;
	wire [WIDTH-1:0] wire_d2_24;
	wire [WIDTH-1:0] wire_d2_25;
	wire [WIDTH-1:0] wire_d2_26;
	wire [WIDTH-1:0] wire_d2_27;
	wire [WIDTH-1:0] wire_d2_28;
	wire [WIDTH-1:0] wire_d2_29;
	wire [WIDTH-1:0] wire_d2_30;
	wire [WIDTH-1:0] wire_d2_31;
	wire [WIDTH-1:0] wire_d2_32;
	wire [WIDTH-1:0] wire_d2_33;
	wire [WIDTH-1:0] wire_d2_34;
	wire [WIDTH-1:0] wire_d2_35;
	wire [WIDTH-1:0] wire_d2_36;
	wire [WIDTH-1:0] wire_d2_37;
	wire [WIDTH-1:0] wire_d2_38;
	wire [WIDTH-1:0] wire_d2_39;
	wire [WIDTH-1:0] wire_d2_40;
	wire [WIDTH-1:0] wire_d2_41;
	wire [WIDTH-1:0] wire_d2_42;
	wire [WIDTH-1:0] wire_d2_43;
	wire [WIDTH-1:0] wire_d2_44;
	wire [WIDTH-1:0] wire_d2_45;
	wire [WIDTH-1:0] wire_d2_46;
	wire [WIDTH-1:0] wire_d2_47;
	wire [WIDTH-1:0] wire_d2_48;
	wire [WIDTH-1:0] wire_d2_49;
	wire [WIDTH-1:0] wire_d2_50;
	wire [WIDTH-1:0] wire_d2_51;
	wire [WIDTH-1:0] wire_d2_52;
	wire [WIDTH-1:0] wire_d2_53;
	wire [WIDTH-1:0] wire_d2_54;
	wire [WIDTH-1:0] wire_d2_55;
	wire [WIDTH-1:0] wire_d2_56;
	wire [WIDTH-1:0] wire_d2_57;
	wire [WIDTH-1:0] wire_d2_58;
	wire [WIDTH-1:0] wire_d2_59;
	wire [WIDTH-1:0] wire_d2_60;
	wire [WIDTH-1:0] wire_d2_61;
	wire [WIDTH-1:0] wire_d2_62;
	wire [WIDTH-1:0] wire_d2_63;
	wire [WIDTH-1:0] wire_d2_64;
	wire [WIDTH-1:0] wire_d2_65;
	wire [WIDTH-1:0] wire_d2_66;
	wire [WIDTH-1:0] wire_d2_67;
	wire [WIDTH-1:0] wire_d2_68;
	wire [WIDTH-1:0] wire_d2_69;
	wire [WIDTH-1:0] wire_d2_70;
	wire [WIDTH-1:0] wire_d2_71;
	wire [WIDTH-1:0] wire_d2_72;
	wire [WIDTH-1:0] wire_d2_73;
	wire [WIDTH-1:0] wire_d2_74;
	wire [WIDTH-1:0] wire_d2_75;
	wire [WIDTH-1:0] wire_d2_76;
	wire [WIDTH-1:0] wire_d2_77;
	wire [WIDTH-1:0] wire_d2_78;
	wire [WIDTH-1:0] wire_d2_79;
	wire [WIDTH-1:0] wire_d2_80;
	wire [WIDTH-1:0] wire_d2_81;
	wire [WIDTH-1:0] wire_d2_82;
	wire [WIDTH-1:0] wire_d2_83;
	wire [WIDTH-1:0] wire_d2_84;
	wire [WIDTH-1:0] wire_d2_85;
	wire [WIDTH-1:0] wire_d2_86;
	wire [WIDTH-1:0] wire_d2_87;
	wire [WIDTH-1:0] wire_d2_88;
	wire [WIDTH-1:0] wire_d2_89;
	wire [WIDTH-1:0] wire_d2_90;
	wire [WIDTH-1:0] wire_d2_91;
	wire [WIDTH-1:0] wire_d2_92;
	wire [WIDTH-1:0] wire_d2_93;
	wire [WIDTH-1:0] wire_d2_94;
	wire [WIDTH-1:0] wire_d2_95;
	wire [WIDTH-1:0] wire_d2_96;
	wire [WIDTH-1:0] wire_d2_97;
	wire [WIDTH-1:0] wire_d2_98;
	wire [WIDTH-1:0] wire_d2_99;
	wire [WIDTH-1:0] wire_d2_100;
	wire [WIDTH-1:0] wire_d2_101;
	wire [WIDTH-1:0] wire_d2_102;
	wire [WIDTH-1:0] wire_d2_103;
	wire [WIDTH-1:0] wire_d2_104;
	wire [WIDTH-1:0] wire_d2_105;
	wire [WIDTH-1:0] wire_d2_106;
	wire [WIDTH-1:0] wire_d2_107;
	wire [WIDTH-1:0] wire_d2_108;
	wire [WIDTH-1:0] wire_d2_109;
	wire [WIDTH-1:0] wire_d2_110;
	wire [WIDTH-1:0] wire_d2_111;
	wire [WIDTH-1:0] wire_d2_112;
	wire [WIDTH-1:0] wire_d2_113;
	wire [WIDTH-1:0] wire_d2_114;
	wire [WIDTH-1:0] wire_d2_115;
	wire [WIDTH-1:0] wire_d2_116;
	wire [WIDTH-1:0] wire_d2_117;
	wire [WIDTH-1:0] wire_d2_118;
	wire [WIDTH-1:0] wire_d3_0;
	wire [WIDTH-1:0] wire_d3_1;
	wire [WIDTH-1:0] wire_d3_2;
	wire [WIDTH-1:0] wire_d3_3;
	wire [WIDTH-1:0] wire_d3_4;
	wire [WIDTH-1:0] wire_d3_5;
	wire [WIDTH-1:0] wire_d3_6;
	wire [WIDTH-1:0] wire_d3_7;
	wire [WIDTH-1:0] wire_d3_8;
	wire [WIDTH-1:0] wire_d3_9;
	wire [WIDTH-1:0] wire_d3_10;
	wire [WIDTH-1:0] wire_d3_11;
	wire [WIDTH-1:0] wire_d3_12;
	wire [WIDTH-1:0] wire_d3_13;
	wire [WIDTH-1:0] wire_d3_14;
	wire [WIDTH-1:0] wire_d3_15;
	wire [WIDTH-1:0] wire_d3_16;
	wire [WIDTH-1:0] wire_d3_17;
	wire [WIDTH-1:0] wire_d3_18;
	wire [WIDTH-1:0] wire_d3_19;
	wire [WIDTH-1:0] wire_d3_20;
	wire [WIDTH-1:0] wire_d3_21;
	wire [WIDTH-1:0] wire_d3_22;
	wire [WIDTH-1:0] wire_d3_23;
	wire [WIDTH-1:0] wire_d3_24;
	wire [WIDTH-1:0] wire_d3_25;
	wire [WIDTH-1:0] wire_d3_26;
	wire [WIDTH-1:0] wire_d3_27;
	wire [WIDTH-1:0] wire_d3_28;
	wire [WIDTH-1:0] wire_d3_29;
	wire [WIDTH-1:0] wire_d3_30;
	wire [WIDTH-1:0] wire_d3_31;
	wire [WIDTH-1:0] wire_d3_32;
	wire [WIDTH-1:0] wire_d3_33;
	wire [WIDTH-1:0] wire_d3_34;
	wire [WIDTH-1:0] wire_d3_35;
	wire [WIDTH-1:0] wire_d3_36;
	wire [WIDTH-1:0] wire_d3_37;
	wire [WIDTH-1:0] wire_d3_38;
	wire [WIDTH-1:0] wire_d3_39;
	wire [WIDTH-1:0] wire_d3_40;
	wire [WIDTH-1:0] wire_d3_41;
	wire [WIDTH-1:0] wire_d3_42;
	wire [WIDTH-1:0] wire_d3_43;
	wire [WIDTH-1:0] wire_d3_44;
	wire [WIDTH-1:0] wire_d3_45;
	wire [WIDTH-1:0] wire_d3_46;
	wire [WIDTH-1:0] wire_d3_47;
	wire [WIDTH-1:0] wire_d3_48;
	wire [WIDTH-1:0] wire_d3_49;
	wire [WIDTH-1:0] wire_d3_50;
	wire [WIDTH-1:0] wire_d3_51;
	wire [WIDTH-1:0] wire_d3_52;
	wire [WIDTH-1:0] wire_d3_53;
	wire [WIDTH-1:0] wire_d3_54;
	wire [WIDTH-1:0] wire_d3_55;
	wire [WIDTH-1:0] wire_d3_56;
	wire [WIDTH-1:0] wire_d3_57;
	wire [WIDTH-1:0] wire_d3_58;
	wire [WIDTH-1:0] wire_d3_59;
	wire [WIDTH-1:0] wire_d3_60;
	wire [WIDTH-1:0] wire_d3_61;
	wire [WIDTH-1:0] wire_d3_62;
	wire [WIDTH-1:0] wire_d3_63;
	wire [WIDTH-1:0] wire_d3_64;
	wire [WIDTH-1:0] wire_d3_65;
	wire [WIDTH-1:0] wire_d3_66;
	wire [WIDTH-1:0] wire_d3_67;
	wire [WIDTH-1:0] wire_d3_68;
	wire [WIDTH-1:0] wire_d3_69;
	wire [WIDTH-1:0] wire_d3_70;
	wire [WIDTH-1:0] wire_d3_71;
	wire [WIDTH-1:0] wire_d3_72;
	wire [WIDTH-1:0] wire_d3_73;
	wire [WIDTH-1:0] wire_d3_74;
	wire [WIDTH-1:0] wire_d3_75;
	wire [WIDTH-1:0] wire_d3_76;
	wire [WIDTH-1:0] wire_d3_77;
	wire [WIDTH-1:0] wire_d3_78;
	wire [WIDTH-1:0] wire_d3_79;
	wire [WIDTH-1:0] wire_d3_80;
	wire [WIDTH-1:0] wire_d3_81;
	wire [WIDTH-1:0] wire_d3_82;
	wire [WIDTH-1:0] wire_d3_83;
	wire [WIDTH-1:0] wire_d3_84;
	wire [WIDTH-1:0] wire_d3_85;
	wire [WIDTH-1:0] wire_d3_86;
	wire [WIDTH-1:0] wire_d3_87;
	wire [WIDTH-1:0] wire_d3_88;
	wire [WIDTH-1:0] wire_d3_89;
	wire [WIDTH-1:0] wire_d3_90;
	wire [WIDTH-1:0] wire_d3_91;
	wire [WIDTH-1:0] wire_d3_92;
	wire [WIDTH-1:0] wire_d3_93;
	wire [WIDTH-1:0] wire_d3_94;
	wire [WIDTH-1:0] wire_d3_95;
	wire [WIDTH-1:0] wire_d3_96;
	wire [WIDTH-1:0] wire_d3_97;
	wire [WIDTH-1:0] wire_d3_98;
	wire [WIDTH-1:0] wire_d3_99;
	wire [WIDTH-1:0] wire_d3_100;
	wire [WIDTH-1:0] wire_d3_101;
	wire [WIDTH-1:0] wire_d3_102;
	wire [WIDTH-1:0] wire_d3_103;
	wire [WIDTH-1:0] wire_d3_104;
	wire [WIDTH-1:0] wire_d3_105;
	wire [WIDTH-1:0] wire_d3_106;
	wire [WIDTH-1:0] wire_d3_107;
	wire [WIDTH-1:0] wire_d3_108;
	wire [WIDTH-1:0] wire_d3_109;
	wire [WIDTH-1:0] wire_d3_110;
	wire [WIDTH-1:0] wire_d3_111;
	wire [WIDTH-1:0] wire_d3_112;
	wire [WIDTH-1:0] wire_d3_113;
	wire [WIDTH-1:0] wire_d3_114;
	wire [WIDTH-1:0] wire_d3_115;
	wire [WIDTH-1:0] wire_d3_116;
	wire [WIDTH-1:0] wire_d3_117;
	wire [WIDTH-1:0] wire_d3_118;
	wire [WIDTH-1:0] wire_d4_0;
	wire [WIDTH-1:0] wire_d4_1;
	wire [WIDTH-1:0] wire_d4_2;
	wire [WIDTH-1:0] wire_d4_3;
	wire [WIDTH-1:0] wire_d4_4;
	wire [WIDTH-1:0] wire_d4_5;
	wire [WIDTH-1:0] wire_d4_6;
	wire [WIDTH-1:0] wire_d4_7;
	wire [WIDTH-1:0] wire_d4_8;
	wire [WIDTH-1:0] wire_d4_9;
	wire [WIDTH-1:0] wire_d4_10;
	wire [WIDTH-1:0] wire_d4_11;
	wire [WIDTH-1:0] wire_d4_12;
	wire [WIDTH-1:0] wire_d4_13;
	wire [WIDTH-1:0] wire_d4_14;
	wire [WIDTH-1:0] wire_d4_15;
	wire [WIDTH-1:0] wire_d4_16;
	wire [WIDTH-1:0] wire_d4_17;
	wire [WIDTH-1:0] wire_d4_18;
	wire [WIDTH-1:0] wire_d4_19;
	wire [WIDTH-1:0] wire_d4_20;
	wire [WIDTH-1:0] wire_d4_21;
	wire [WIDTH-1:0] wire_d4_22;
	wire [WIDTH-1:0] wire_d4_23;
	wire [WIDTH-1:0] wire_d4_24;
	wire [WIDTH-1:0] wire_d4_25;
	wire [WIDTH-1:0] wire_d4_26;
	wire [WIDTH-1:0] wire_d4_27;
	wire [WIDTH-1:0] wire_d4_28;
	wire [WIDTH-1:0] wire_d4_29;
	wire [WIDTH-1:0] wire_d4_30;
	wire [WIDTH-1:0] wire_d4_31;
	wire [WIDTH-1:0] wire_d4_32;
	wire [WIDTH-1:0] wire_d4_33;
	wire [WIDTH-1:0] wire_d4_34;
	wire [WIDTH-1:0] wire_d4_35;
	wire [WIDTH-1:0] wire_d4_36;
	wire [WIDTH-1:0] wire_d4_37;
	wire [WIDTH-1:0] wire_d4_38;
	wire [WIDTH-1:0] wire_d4_39;
	wire [WIDTH-1:0] wire_d4_40;
	wire [WIDTH-1:0] wire_d4_41;
	wire [WIDTH-1:0] wire_d4_42;
	wire [WIDTH-1:0] wire_d4_43;
	wire [WIDTH-1:0] wire_d4_44;
	wire [WIDTH-1:0] wire_d4_45;
	wire [WIDTH-1:0] wire_d4_46;
	wire [WIDTH-1:0] wire_d4_47;
	wire [WIDTH-1:0] wire_d4_48;
	wire [WIDTH-1:0] wire_d4_49;
	wire [WIDTH-1:0] wire_d4_50;
	wire [WIDTH-1:0] wire_d4_51;
	wire [WIDTH-1:0] wire_d4_52;
	wire [WIDTH-1:0] wire_d4_53;
	wire [WIDTH-1:0] wire_d4_54;
	wire [WIDTH-1:0] wire_d4_55;
	wire [WIDTH-1:0] wire_d4_56;
	wire [WIDTH-1:0] wire_d4_57;
	wire [WIDTH-1:0] wire_d4_58;
	wire [WIDTH-1:0] wire_d4_59;
	wire [WIDTH-1:0] wire_d4_60;
	wire [WIDTH-1:0] wire_d4_61;
	wire [WIDTH-1:0] wire_d4_62;
	wire [WIDTH-1:0] wire_d4_63;
	wire [WIDTH-1:0] wire_d4_64;
	wire [WIDTH-1:0] wire_d4_65;
	wire [WIDTH-1:0] wire_d4_66;
	wire [WIDTH-1:0] wire_d4_67;
	wire [WIDTH-1:0] wire_d4_68;
	wire [WIDTH-1:0] wire_d4_69;
	wire [WIDTH-1:0] wire_d4_70;
	wire [WIDTH-1:0] wire_d4_71;
	wire [WIDTH-1:0] wire_d4_72;
	wire [WIDTH-1:0] wire_d4_73;
	wire [WIDTH-1:0] wire_d4_74;
	wire [WIDTH-1:0] wire_d4_75;
	wire [WIDTH-1:0] wire_d4_76;
	wire [WIDTH-1:0] wire_d4_77;
	wire [WIDTH-1:0] wire_d4_78;
	wire [WIDTH-1:0] wire_d4_79;
	wire [WIDTH-1:0] wire_d4_80;
	wire [WIDTH-1:0] wire_d4_81;
	wire [WIDTH-1:0] wire_d4_82;
	wire [WIDTH-1:0] wire_d4_83;
	wire [WIDTH-1:0] wire_d4_84;
	wire [WIDTH-1:0] wire_d4_85;
	wire [WIDTH-1:0] wire_d4_86;
	wire [WIDTH-1:0] wire_d4_87;
	wire [WIDTH-1:0] wire_d4_88;
	wire [WIDTH-1:0] wire_d4_89;
	wire [WIDTH-1:0] wire_d4_90;
	wire [WIDTH-1:0] wire_d4_91;
	wire [WIDTH-1:0] wire_d4_92;
	wire [WIDTH-1:0] wire_d4_93;
	wire [WIDTH-1:0] wire_d4_94;
	wire [WIDTH-1:0] wire_d4_95;
	wire [WIDTH-1:0] wire_d4_96;
	wire [WIDTH-1:0] wire_d4_97;
	wire [WIDTH-1:0] wire_d4_98;
	wire [WIDTH-1:0] wire_d4_99;
	wire [WIDTH-1:0] wire_d4_100;
	wire [WIDTH-1:0] wire_d4_101;
	wire [WIDTH-1:0] wire_d4_102;
	wire [WIDTH-1:0] wire_d4_103;
	wire [WIDTH-1:0] wire_d4_104;
	wire [WIDTH-1:0] wire_d4_105;
	wire [WIDTH-1:0] wire_d4_106;
	wire [WIDTH-1:0] wire_d4_107;
	wire [WIDTH-1:0] wire_d4_108;
	wire [WIDTH-1:0] wire_d4_109;
	wire [WIDTH-1:0] wire_d4_110;
	wire [WIDTH-1:0] wire_d4_111;
	wire [WIDTH-1:0] wire_d4_112;
	wire [WIDTH-1:0] wire_d4_113;
	wire [WIDTH-1:0] wire_d4_114;
	wire [WIDTH-1:0] wire_d4_115;
	wire [WIDTH-1:0] wire_d4_116;
	wire [WIDTH-1:0] wire_d4_117;
	wire [WIDTH-1:0] wire_d4_118;
	wire [WIDTH-1:0] wire_d5_0;
	wire [WIDTH-1:0] wire_d5_1;
	wire [WIDTH-1:0] wire_d5_2;
	wire [WIDTH-1:0] wire_d5_3;
	wire [WIDTH-1:0] wire_d5_4;
	wire [WIDTH-1:0] wire_d5_5;
	wire [WIDTH-1:0] wire_d5_6;
	wire [WIDTH-1:0] wire_d5_7;
	wire [WIDTH-1:0] wire_d5_8;
	wire [WIDTH-1:0] wire_d5_9;
	wire [WIDTH-1:0] wire_d5_10;
	wire [WIDTH-1:0] wire_d5_11;
	wire [WIDTH-1:0] wire_d5_12;
	wire [WIDTH-1:0] wire_d5_13;
	wire [WIDTH-1:0] wire_d5_14;
	wire [WIDTH-1:0] wire_d5_15;
	wire [WIDTH-1:0] wire_d5_16;
	wire [WIDTH-1:0] wire_d5_17;
	wire [WIDTH-1:0] wire_d5_18;
	wire [WIDTH-1:0] wire_d5_19;
	wire [WIDTH-1:0] wire_d5_20;
	wire [WIDTH-1:0] wire_d5_21;
	wire [WIDTH-1:0] wire_d5_22;
	wire [WIDTH-1:0] wire_d5_23;
	wire [WIDTH-1:0] wire_d5_24;
	wire [WIDTH-1:0] wire_d5_25;
	wire [WIDTH-1:0] wire_d5_26;
	wire [WIDTH-1:0] wire_d5_27;
	wire [WIDTH-1:0] wire_d5_28;
	wire [WIDTH-1:0] wire_d5_29;
	wire [WIDTH-1:0] wire_d5_30;
	wire [WIDTH-1:0] wire_d5_31;
	wire [WIDTH-1:0] wire_d5_32;
	wire [WIDTH-1:0] wire_d5_33;
	wire [WIDTH-1:0] wire_d5_34;
	wire [WIDTH-1:0] wire_d5_35;
	wire [WIDTH-1:0] wire_d5_36;
	wire [WIDTH-1:0] wire_d5_37;
	wire [WIDTH-1:0] wire_d5_38;
	wire [WIDTH-1:0] wire_d5_39;
	wire [WIDTH-1:0] wire_d5_40;
	wire [WIDTH-1:0] wire_d5_41;
	wire [WIDTH-1:0] wire_d5_42;
	wire [WIDTH-1:0] wire_d5_43;
	wire [WIDTH-1:0] wire_d5_44;
	wire [WIDTH-1:0] wire_d5_45;
	wire [WIDTH-1:0] wire_d5_46;
	wire [WIDTH-1:0] wire_d5_47;
	wire [WIDTH-1:0] wire_d5_48;
	wire [WIDTH-1:0] wire_d5_49;
	wire [WIDTH-1:0] wire_d5_50;
	wire [WIDTH-1:0] wire_d5_51;
	wire [WIDTH-1:0] wire_d5_52;
	wire [WIDTH-1:0] wire_d5_53;
	wire [WIDTH-1:0] wire_d5_54;
	wire [WIDTH-1:0] wire_d5_55;
	wire [WIDTH-1:0] wire_d5_56;
	wire [WIDTH-1:0] wire_d5_57;
	wire [WIDTH-1:0] wire_d5_58;
	wire [WIDTH-1:0] wire_d5_59;
	wire [WIDTH-1:0] wire_d5_60;
	wire [WIDTH-1:0] wire_d5_61;
	wire [WIDTH-1:0] wire_d5_62;
	wire [WIDTH-1:0] wire_d5_63;
	wire [WIDTH-1:0] wire_d5_64;
	wire [WIDTH-1:0] wire_d5_65;
	wire [WIDTH-1:0] wire_d5_66;
	wire [WIDTH-1:0] wire_d5_67;
	wire [WIDTH-1:0] wire_d5_68;
	wire [WIDTH-1:0] wire_d5_69;
	wire [WIDTH-1:0] wire_d5_70;
	wire [WIDTH-1:0] wire_d5_71;
	wire [WIDTH-1:0] wire_d5_72;
	wire [WIDTH-1:0] wire_d5_73;
	wire [WIDTH-1:0] wire_d5_74;
	wire [WIDTH-1:0] wire_d5_75;
	wire [WIDTH-1:0] wire_d5_76;
	wire [WIDTH-1:0] wire_d5_77;
	wire [WIDTH-1:0] wire_d5_78;
	wire [WIDTH-1:0] wire_d5_79;
	wire [WIDTH-1:0] wire_d5_80;
	wire [WIDTH-1:0] wire_d5_81;
	wire [WIDTH-1:0] wire_d5_82;
	wire [WIDTH-1:0] wire_d5_83;
	wire [WIDTH-1:0] wire_d5_84;
	wire [WIDTH-1:0] wire_d5_85;
	wire [WIDTH-1:0] wire_d5_86;
	wire [WIDTH-1:0] wire_d5_87;
	wire [WIDTH-1:0] wire_d5_88;
	wire [WIDTH-1:0] wire_d5_89;
	wire [WIDTH-1:0] wire_d5_90;
	wire [WIDTH-1:0] wire_d5_91;
	wire [WIDTH-1:0] wire_d5_92;
	wire [WIDTH-1:0] wire_d5_93;
	wire [WIDTH-1:0] wire_d5_94;
	wire [WIDTH-1:0] wire_d5_95;
	wire [WIDTH-1:0] wire_d5_96;
	wire [WIDTH-1:0] wire_d5_97;
	wire [WIDTH-1:0] wire_d5_98;
	wire [WIDTH-1:0] wire_d5_99;
	wire [WIDTH-1:0] wire_d5_100;
	wire [WIDTH-1:0] wire_d5_101;
	wire [WIDTH-1:0] wire_d5_102;
	wire [WIDTH-1:0] wire_d5_103;
	wire [WIDTH-1:0] wire_d5_104;
	wire [WIDTH-1:0] wire_d5_105;
	wire [WIDTH-1:0] wire_d5_106;
	wire [WIDTH-1:0] wire_d5_107;
	wire [WIDTH-1:0] wire_d5_108;
	wire [WIDTH-1:0] wire_d5_109;
	wire [WIDTH-1:0] wire_d5_110;
	wire [WIDTH-1:0] wire_d5_111;
	wire [WIDTH-1:0] wire_d5_112;
	wire [WIDTH-1:0] wire_d5_113;
	wire [WIDTH-1:0] wire_d5_114;
	wire [WIDTH-1:0] wire_d5_115;
	wire [WIDTH-1:0] wire_d5_116;
	wire [WIDTH-1:0] wire_d5_117;
	wire [WIDTH-1:0] wire_d5_118;
	wire [WIDTH-1:0] wire_d6_0;
	wire [WIDTH-1:0] wire_d6_1;
	wire [WIDTH-1:0] wire_d6_2;
	wire [WIDTH-1:0] wire_d6_3;
	wire [WIDTH-1:0] wire_d6_4;
	wire [WIDTH-1:0] wire_d6_5;
	wire [WIDTH-1:0] wire_d6_6;
	wire [WIDTH-1:0] wire_d6_7;
	wire [WIDTH-1:0] wire_d6_8;
	wire [WIDTH-1:0] wire_d6_9;
	wire [WIDTH-1:0] wire_d6_10;
	wire [WIDTH-1:0] wire_d6_11;
	wire [WIDTH-1:0] wire_d6_12;
	wire [WIDTH-1:0] wire_d6_13;
	wire [WIDTH-1:0] wire_d6_14;
	wire [WIDTH-1:0] wire_d6_15;
	wire [WIDTH-1:0] wire_d6_16;
	wire [WIDTH-1:0] wire_d6_17;
	wire [WIDTH-1:0] wire_d6_18;
	wire [WIDTH-1:0] wire_d6_19;
	wire [WIDTH-1:0] wire_d6_20;
	wire [WIDTH-1:0] wire_d6_21;
	wire [WIDTH-1:0] wire_d6_22;
	wire [WIDTH-1:0] wire_d6_23;
	wire [WIDTH-1:0] wire_d6_24;
	wire [WIDTH-1:0] wire_d6_25;
	wire [WIDTH-1:0] wire_d6_26;
	wire [WIDTH-1:0] wire_d6_27;
	wire [WIDTH-1:0] wire_d6_28;
	wire [WIDTH-1:0] wire_d6_29;
	wire [WIDTH-1:0] wire_d6_30;
	wire [WIDTH-1:0] wire_d6_31;
	wire [WIDTH-1:0] wire_d6_32;
	wire [WIDTH-1:0] wire_d6_33;
	wire [WIDTH-1:0] wire_d6_34;
	wire [WIDTH-1:0] wire_d6_35;
	wire [WIDTH-1:0] wire_d6_36;
	wire [WIDTH-1:0] wire_d6_37;
	wire [WIDTH-1:0] wire_d6_38;
	wire [WIDTH-1:0] wire_d6_39;
	wire [WIDTH-1:0] wire_d6_40;
	wire [WIDTH-1:0] wire_d6_41;
	wire [WIDTH-1:0] wire_d6_42;
	wire [WIDTH-1:0] wire_d6_43;
	wire [WIDTH-1:0] wire_d6_44;
	wire [WIDTH-1:0] wire_d6_45;
	wire [WIDTH-1:0] wire_d6_46;
	wire [WIDTH-1:0] wire_d6_47;
	wire [WIDTH-1:0] wire_d6_48;
	wire [WIDTH-1:0] wire_d6_49;
	wire [WIDTH-1:0] wire_d6_50;
	wire [WIDTH-1:0] wire_d6_51;
	wire [WIDTH-1:0] wire_d6_52;
	wire [WIDTH-1:0] wire_d6_53;
	wire [WIDTH-1:0] wire_d6_54;
	wire [WIDTH-1:0] wire_d6_55;
	wire [WIDTH-1:0] wire_d6_56;
	wire [WIDTH-1:0] wire_d6_57;
	wire [WIDTH-1:0] wire_d6_58;
	wire [WIDTH-1:0] wire_d6_59;
	wire [WIDTH-1:0] wire_d6_60;
	wire [WIDTH-1:0] wire_d6_61;
	wire [WIDTH-1:0] wire_d6_62;
	wire [WIDTH-1:0] wire_d6_63;
	wire [WIDTH-1:0] wire_d6_64;
	wire [WIDTH-1:0] wire_d6_65;
	wire [WIDTH-1:0] wire_d6_66;
	wire [WIDTH-1:0] wire_d6_67;
	wire [WIDTH-1:0] wire_d6_68;
	wire [WIDTH-1:0] wire_d6_69;
	wire [WIDTH-1:0] wire_d6_70;
	wire [WIDTH-1:0] wire_d6_71;
	wire [WIDTH-1:0] wire_d6_72;
	wire [WIDTH-1:0] wire_d6_73;
	wire [WIDTH-1:0] wire_d6_74;
	wire [WIDTH-1:0] wire_d6_75;
	wire [WIDTH-1:0] wire_d6_76;
	wire [WIDTH-1:0] wire_d6_77;
	wire [WIDTH-1:0] wire_d6_78;
	wire [WIDTH-1:0] wire_d6_79;
	wire [WIDTH-1:0] wire_d6_80;
	wire [WIDTH-1:0] wire_d6_81;
	wire [WIDTH-1:0] wire_d6_82;
	wire [WIDTH-1:0] wire_d6_83;
	wire [WIDTH-1:0] wire_d6_84;
	wire [WIDTH-1:0] wire_d6_85;
	wire [WIDTH-1:0] wire_d6_86;
	wire [WIDTH-1:0] wire_d6_87;
	wire [WIDTH-1:0] wire_d6_88;
	wire [WIDTH-1:0] wire_d6_89;
	wire [WIDTH-1:0] wire_d6_90;
	wire [WIDTH-1:0] wire_d6_91;
	wire [WIDTH-1:0] wire_d6_92;
	wire [WIDTH-1:0] wire_d6_93;
	wire [WIDTH-1:0] wire_d6_94;
	wire [WIDTH-1:0] wire_d6_95;
	wire [WIDTH-1:0] wire_d6_96;
	wire [WIDTH-1:0] wire_d6_97;
	wire [WIDTH-1:0] wire_d6_98;
	wire [WIDTH-1:0] wire_d6_99;
	wire [WIDTH-1:0] wire_d6_100;
	wire [WIDTH-1:0] wire_d6_101;
	wire [WIDTH-1:0] wire_d6_102;
	wire [WIDTH-1:0] wire_d6_103;
	wire [WIDTH-1:0] wire_d6_104;
	wire [WIDTH-1:0] wire_d6_105;
	wire [WIDTH-1:0] wire_d6_106;
	wire [WIDTH-1:0] wire_d6_107;
	wire [WIDTH-1:0] wire_d6_108;
	wire [WIDTH-1:0] wire_d6_109;
	wire [WIDTH-1:0] wire_d6_110;
	wire [WIDTH-1:0] wire_d6_111;
	wire [WIDTH-1:0] wire_d6_112;
	wire [WIDTH-1:0] wire_d6_113;
	wire [WIDTH-1:0] wire_d6_114;
	wire [WIDTH-1:0] wire_d6_115;
	wire [WIDTH-1:0] wire_d6_116;
	wire [WIDTH-1:0] wire_d6_117;
	wire [WIDTH-1:0] wire_d6_118;
	wire [WIDTH-1:0] wire_d7_0;
	wire [WIDTH-1:0] wire_d7_1;
	wire [WIDTH-1:0] wire_d7_2;
	wire [WIDTH-1:0] wire_d7_3;
	wire [WIDTH-1:0] wire_d7_4;
	wire [WIDTH-1:0] wire_d7_5;
	wire [WIDTH-1:0] wire_d7_6;
	wire [WIDTH-1:0] wire_d7_7;
	wire [WIDTH-1:0] wire_d7_8;
	wire [WIDTH-1:0] wire_d7_9;
	wire [WIDTH-1:0] wire_d7_10;
	wire [WIDTH-1:0] wire_d7_11;
	wire [WIDTH-1:0] wire_d7_12;
	wire [WIDTH-1:0] wire_d7_13;
	wire [WIDTH-1:0] wire_d7_14;
	wire [WIDTH-1:0] wire_d7_15;
	wire [WIDTH-1:0] wire_d7_16;
	wire [WIDTH-1:0] wire_d7_17;
	wire [WIDTH-1:0] wire_d7_18;
	wire [WIDTH-1:0] wire_d7_19;
	wire [WIDTH-1:0] wire_d7_20;
	wire [WIDTH-1:0] wire_d7_21;
	wire [WIDTH-1:0] wire_d7_22;
	wire [WIDTH-1:0] wire_d7_23;
	wire [WIDTH-1:0] wire_d7_24;
	wire [WIDTH-1:0] wire_d7_25;
	wire [WIDTH-1:0] wire_d7_26;
	wire [WIDTH-1:0] wire_d7_27;
	wire [WIDTH-1:0] wire_d7_28;
	wire [WIDTH-1:0] wire_d7_29;
	wire [WIDTH-1:0] wire_d7_30;
	wire [WIDTH-1:0] wire_d7_31;
	wire [WIDTH-1:0] wire_d7_32;
	wire [WIDTH-1:0] wire_d7_33;
	wire [WIDTH-1:0] wire_d7_34;
	wire [WIDTH-1:0] wire_d7_35;
	wire [WIDTH-1:0] wire_d7_36;
	wire [WIDTH-1:0] wire_d7_37;
	wire [WIDTH-1:0] wire_d7_38;
	wire [WIDTH-1:0] wire_d7_39;
	wire [WIDTH-1:0] wire_d7_40;
	wire [WIDTH-1:0] wire_d7_41;
	wire [WIDTH-1:0] wire_d7_42;
	wire [WIDTH-1:0] wire_d7_43;
	wire [WIDTH-1:0] wire_d7_44;
	wire [WIDTH-1:0] wire_d7_45;
	wire [WIDTH-1:0] wire_d7_46;
	wire [WIDTH-1:0] wire_d7_47;
	wire [WIDTH-1:0] wire_d7_48;
	wire [WIDTH-1:0] wire_d7_49;
	wire [WIDTH-1:0] wire_d7_50;
	wire [WIDTH-1:0] wire_d7_51;
	wire [WIDTH-1:0] wire_d7_52;
	wire [WIDTH-1:0] wire_d7_53;
	wire [WIDTH-1:0] wire_d7_54;
	wire [WIDTH-1:0] wire_d7_55;
	wire [WIDTH-1:0] wire_d7_56;
	wire [WIDTH-1:0] wire_d7_57;
	wire [WIDTH-1:0] wire_d7_58;
	wire [WIDTH-1:0] wire_d7_59;
	wire [WIDTH-1:0] wire_d7_60;
	wire [WIDTH-1:0] wire_d7_61;
	wire [WIDTH-1:0] wire_d7_62;
	wire [WIDTH-1:0] wire_d7_63;
	wire [WIDTH-1:0] wire_d7_64;
	wire [WIDTH-1:0] wire_d7_65;
	wire [WIDTH-1:0] wire_d7_66;
	wire [WIDTH-1:0] wire_d7_67;
	wire [WIDTH-1:0] wire_d7_68;
	wire [WIDTH-1:0] wire_d7_69;
	wire [WIDTH-1:0] wire_d7_70;
	wire [WIDTH-1:0] wire_d7_71;
	wire [WIDTH-1:0] wire_d7_72;
	wire [WIDTH-1:0] wire_d7_73;
	wire [WIDTH-1:0] wire_d7_74;
	wire [WIDTH-1:0] wire_d7_75;
	wire [WIDTH-1:0] wire_d7_76;
	wire [WIDTH-1:0] wire_d7_77;
	wire [WIDTH-1:0] wire_d7_78;
	wire [WIDTH-1:0] wire_d7_79;
	wire [WIDTH-1:0] wire_d7_80;
	wire [WIDTH-1:0] wire_d7_81;
	wire [WIDTH-1:0] wire_d7_82;
	wire [WIDTH-1:0] wire_d7_83;
	wire [WIDTH-1:0] wire_d7_84;
	wire [WIDTH-1:0] wire_d7_85;
	wire [WIDTH-1:0] wire_d7_86;
	wire [WIDTH-1:0] wire_d7_87;
	wire [WIDTH-1:0] wire_d7_88;
	wire [WIDTH-1:0] wire_d7_89;
	wire [WIDTH-1:0] wire_d7_90;
	wire [WIDTH-1:0] wire_d7_91;
	wire [WIDTH-1:0] wire_d7_92;
	wire [WIDTH-1:0] wire_d7_93;
	wire [WIDTH-1:0] wire_d7_94;
	wire [WIDTH-1:0] wire_d7_95;
	wire [WIDTH-1:0] wire_d7_96;
	wire [WIDTH-1:0] wire_d7_97;
	wire [WIDTH-1:0] wire_d7_98;
	wire [WIDTH-1:0] wire_d7_99;
	wire [WIDTH-1:0] wire_d7_100;
	wire [WIDTH-1:0] wire_d7_101;
	wire [WIDTH-1:0] wire_d7_102;
	wire [WIDTH-1:0] wire_d7_103;
	wire [WIDTH-1:0] wire_d7_104;
	wire [WIDTH-1:0] wire_d7_105;
	wire [WIDTH-1:0] wire_d7_106;
	wire [WIDTH-1:0] wire_d7_107;
	wire [WIDTH-1:0] wire_d7_108;
	wire [WIDTH-1:0] wire_d7_109;
	wire [WIDTH-1:0] wire_d7_110;
	wire [WIDTH-1:0] wire_d7_111;
	wire [WIDTH-1:0] wire_d7_112;
	wire [WIDTH-1:0] wire_d7_113;
	wire [WIDTH-1:0] wire_d7_114;
	wire [WIDTH-1:0] wire_d7_115;
	wire [WIDTH-1:0] wire_d7_116;
	wire [WIDTH-1:0] wire_d7_117;
	wire [WIDTH-1:0] wire_d7_118;
	wire [WIDTH-1:0] wire_d8_0;
	wire [WIDTH-1:0] wire_d8_1;
	wire [WIDTH-1:0] wire_d8_2;
	wire [WIDTH-1:0] wire_d8_3;
	wire [WIDTH-1:0] wire_d8_4;
	wire [WIDTH-1:0] wire_d8_5;
	wire [WIDTH-1:0] wire_d8_6;
	wire [WIDTH-1:0] wire_d8_7;
	wire [WIDTH-1:0] wire_d8_8;
	wire [WIDTH-1:0] wire_d8_9;
	wire [WIDTH-1:0] wire_d8_10;
	wire [WIDTH-1:0] wire_d8_11;
	wire [WIDTH-1:0] wire_d8_12;
	wire [WIDTH-1:0] wire_d8_13;
	wire [WIDTH-1:0] wire_d8_14;
	wire [WIDTH-1:0] wire_d8_15;
	wire [WIDTH-1:0] wire_d8_16;
	wire [WIDTH-1:0] wire_d8_17;
	wire [WIDTH-1:0] wire_d8_18;
	wire [WIDTH-1:0] wire_d8_19;
	wire [WIDTH-1:0] wire_d8_20;
	wire [WIDTH-1:0] wire_d8_21;
	wire [WIDTH-1:0] wire_d8_22;
	wire [WIDTH-1:0] wire_d8_23;
	wire [WIDTH-1:0] wire_d8_24;
	wire [WIDTH-1:0] wire_d8_25;
	wire [WIDTH-1:0] wire_d8_26;
	wire [WIDTH-1:0] wire_d8_27;
	wire [WIDTH-1:0] wire_d8_28;
	wire [WIDTH-1:0] wire_d8_29;
	wire [WIDTH-1:0] wire_d8_30;
	wire [WIDTH-1:0] wire_d8_31;
	wire [WIDTH-1:0] wire_d8_32;
	wire [WIDTH-1:0] wire_d8_33;
	wire [WIDTH-1:0] wire_d8_34;
	wire [WIDTH-1:0] wire_d8_35;
	wire [WIDTH-1:0] wire_d8_36;
	wire [WIDTH-1:0] wire_d8_37;
	wire [WIDTH-1:0] wire_d8_38;
	wire [WIDTH-1:0] wire_d8_39;
	wire [WIDTH-1:0] wire_d8_40;
	wire [WIDTH-1:0] wire_d8_41;
	wire [WIDTH-1:0] wire_d8_42;
	wire [WIDTH-1:0] wire_d8_43;
	wire [WIDTH-1:0] wire_d8_44;
	wire [WIDTH-1:0] wire_d8_45;
	wire [WIDTH-1:0] wire_d8_46;
	wire [WIDTH-1:0] wire_d8_47;
	wire [WIDTH-1:0] wire_d8_48;
	wire [WIDTH-1:0] wire_d8_49;
	wire [WIDTH-1:0] wire_d8_50;
	wire [WIDTH-1:0] wire_d8_51;
	wire [WIDTH-1:0] wire_d8_52;
	wire [WIDTH-1:0] wire_d8_53;
	wire [WIDTH-1:0] wire_d8_54;
	wire [WIDTH-1:0] wire_d8_55;
	wire [WIDTH-1:0] wire_d8_56;
	wire [WIDTH-1:0] wire_d8_57;
	wire [WIDTH-1:0] wire_d8_58;
	wire [WIDTH-1:0] wire_d8_59;
	wire [WIDTH-1:0] wire_d8_60;
	wire [WIDTH-1:0] wire_d8_61;
	wire [WIDTH-1:0] wire_d8_62;
	wire [WIDTH-1:0] wire_d8_63;
	wire [WIDTH-1:0] wire_d8_64;
	wire [WIDTH-1:0] wire_d8_65;
	wire [WIDTH-1:0] wire_d8_66;
	wire [WIDTH-1:0] wire_d8_67;
	wire [WIDTH-1:0] wire_d8_68;
	wire [WIDTH-1:0] wire_d8_69;
	wire [WIDTH-1:0] wire_d8_70;
	wire [WIDTH-1:0] wire_d8_71;
	wire [WIDTH-1:0] wire_d8_72;
	wire [WIDTH-1:0] wire_d8_73;
	wire [WIDTH-1:0] wire_d8_74;
	wire [WIDTH-1:0] wire_d8_75;
	wire [WIDTH-1:0] wire_d8_76;
	wire [WIDTH-1:0] wire_d8_77;
	wire [WIDTH-1:0] wire_d8_78;
	wire [WIDTH-1:0] wire_d8_79;
	wire [WIDTH-1:0] wire_d8_80;
	wire [WIDTH-1:0] wire_d8_81;
	wire [WIDTH-1:0] wire_d8_82;
	wire [WIDTH-1:0] wire_d8_83;
	wire [WIDTH-1:0] wire_d8_84;
	wire [WIDTH-1:0] wire_d8_85;
	wire [WIDTH-1:0] wire_d8_86;
	wire [WIDTH-1:0] wire_d8_87;
	wire [WIDTH-1:0] wire_d8_88;
	wire [WIDTH-1:0] wire_d8_89;
	wire [WIDTH-1:0] wire_d8_90;
	wire [WIDTH-1:0] wire_d8_91;
	wire [WIDTH-1:0] wire_d8_92;
	wire [WIDTH-1:0] wire_d8_93;
	wire [WIDTH-1:0] wire_d8_94;
	wire [WIDTH-1:0] wire_d8_95;
	wire [WIDTH-1:0] wire_d8_96;
	wire [WIDTH-1:0] wire_d8_97;
	wire [WIDTH-1:0] wire_d8_98;
	wire [WIDTH-1:0] wire_d8_99;
	wire [WIDTH-1:0] wire_d8_100;
	wire [WIDTH-1:0] wire_d8_101;
	wire [WIDTH-1:0] wire_d8_102;
	wire [WIDTH-1:0] wire_d8_103;
	wire [WIDTH-1:0] wire_d8_104;
	wire [WIDTH-1:0] wire_d8_105;
	wire [WIDTH-1:0] wire_d8_106;
	wire [WIDTH-1:0] wire_d8_107;
	wire [WIDTH-1:0] wire_d8_108;
	wire [WIDTH-1:0] wire_d8_109;
	wire [WIDTH-1:0] wire_d8_110;
	wire [WIDTH-1:0] wire_d8_111;
	wire [WIDTH-1:0] wire_d8_112;
	wire [WIDTH-1:0] wire_d8_113;
	wire [WIDTH-1:0] wire_d8_114;
	wire [WIDTH-1:0] wire_d8_115;
	wire [WIDTH-1:0] wire_d8_116;
	wire [WIDTH-1:0] wire_d8_117;
	wire [WIDTH-1:0] wire_d8_118;
	wire [WIDTH-1:0] wire_d9_0;
	wire [WIDTH-1:0] wire_d9_1;
	wire [WIDTH-1:0] wire_d9_2;
	wire [WIDTH-1:0] wire_d9_3;
	wire [WIDTH-1:0] wire_d9_4;
	wire [WIDTH-1:0] wire_d9_5;
	wire [WIDTH-1:0] wire_d9_6;
	wire [WIDTH-1:0] wire_d9_7;
	wire [WIDTH-1:0] wire_d9_8;
	wire [WIDTH-1:0] wire_d9_9;
	wire [WIDTH-1:0] wire_d9_10;
	wire [WIDTH-1:0] wire_d9_11;
	wire [WIDTH-1:0] wire_d9_12;
	wire [WIDTH-1:0] wire_d9_13;
	wire [WIDTH-1:0] wire_d9_14;
	wire [WIDTH-1:0] wire_d9_15;
	wire [WIDTH-1:0] wire_d9_16;
	wire [WIDTH-1:0] wire_d9_17;
	wire [WIDTH-1:0] wire_d9_18;
	wire [WIDTH-1:0] wire_d9_19;
	wire [WIDTH-1:0] wire_d9_20;
	wire [WIDTH-1:0] wire_d9_21;
	wire [WIDTH-1:0] wire_d9_22;
	wire [WIDTH-1:0] wire_d9_23;
	wire [WIDTH-1:0] wire_d9_24;
	wire [WIDTH-1:0] wire_d9_25;
	wire [WIDTH-1:0] wire_d9_26;
	wire [WIDTH-1:0] wire_d9_27;
	wire [WIDTH-1:0] wire_d9_28;
	wire [WIDTH-1:0] wire_d9_29;
	wire [WIDTH-1:0] wire_d9_30;
	wire [WIDTH-1:0] wire_d9_31;
	wire [WIDTH-1:0] wire_d9_32;
	wire [WIDTH-1:0] wire_d9_33;
	wire [WIDTH-1:0] wire_d9_34;
	wire [WIDTH-1:0] wire_d9_35;
	wire [WIDTH-1:0] wire_d9_36;
	wire [WIDTH-1:0] wire_d9_37;
	wire [WIDTH-1:0] wire_d9_38;
	wire [WIDTH-1:0] wire_d9_39;
	wire [WIDTH-1:0] wire_d9_40;
	wire [WIDTH-1:0] wire_d9_41;
	wire [WIDTH-1:0] wire_d9_42;
	wire [WIDTH-1:0] wire_d9_43;
	wire [WIDTH-1:0] wire_d9_44;
	wire [WIDTH-1:0] wire_d9_45;
	wire [WIDTH-1:0] wire_d9_46;
	wire [WIDTH-1:0] wire_d9_47;
	wire [WIDTH-1:0] wire_d9_48;
	wire [WIDTH-1:0] wire_d9_49;
	wire [WIDTH-1:0] wire_d9_50;
	wire [WIDTH-1:0] wire_d9_51;
	wire [WIDTH-1:0] wire_d9_52;
	wire [WIDTH-1:0] wire_d9_53;
	wire [WIDTH-1:0] wire_d9_54;
	wire [WIDTH-1:0] wire_d9_55;
	wire [WIDTH-1:0] wire_d9_56;
	wire [WIDTH-1:0] wire_d9_57;
	wire [WIDTH-1:0] wire_d9_58;
	wire [WIDTH-1:0] wire_d9_59;
	wire [WIDTH-1:0] wire_d9_60;
	wire [WIDTH-1:0] wire_d9_61;
	wire [WIDTH-1:0] wire_d9_62;
	wire [WIDTH-1:0] wire_d9_63;
	wire [WIDTH-1:0] wire_d9_64;
	wire [WIDTH-1:0] wire_d9_65;
	wire [WIDTH-1:0] wire_d9_66;
	wire [WIDTH-1:0] wire_d9_67;
	wire [WIDTH-1:0] wire_d9_68;
	wire [WIDTH-1:0] wire_d9_69;
	wire [WIDTH-1:0] wire_d9_70;
	wire [WIDTH-1:0] wire_d9_71;
	wire [WIDTH-1:0] wire_d9_72;
	wire [WIDTH-1:0] wire_d9_73;
	wire [WIDTH-1:0] wire_d9_74;
	wire [WIDTH-1:0] wire_d9_75;
	wire [WIDTH-1:0] wire_d9_76;
	wire [WIDTH-1:0] wire_d9_77;
	wire [WIDTH-1:0] wire_d9_78;
	wire [WIDTH-1:0] wire_d9_79;
	wire [WIDTH-1:0] wire_d9_80;
	wire [WIDTH-1:0] wire_d9_81;
	wire [WIDTH-1:0] wire_d9_82;
	wire [WIDTH-1:0] wire_d9_83;
	wire [WIDTH-1:0] wire_d9_84;
	wire [WIDTH-1:0] wire_d9_85;
	wire [WIDTH-1:0] wire_d9_86;
	wire [WIDTH-1:0] wire_d9_87;
	wire [WIDTH-1:0] wire_d9_88;
	wire [WIDTH-1:0] wire_d9_89;
	wire [WIDTH-1:0] wire_d9_90;
	wire [WIDTH-1:0] wire_d9_91;
	wire [WIDTH-1:0] wire_d9_92;
	wire [WIDTH-1:0] wire_d9_93;
	wire [WIDTH-1:0] wire_d9_94;
	wire [WIDTH-1:0] wire_d9_95;
	wire [WIDTH-1:0] wire_d9_96;
	wire [WIDTH-1:0] wire_d9_97;
	wire [WIDTH-1:0] wire_d9_98;
	wire [WIDTH-1:0] wire_d9_99;
	wire [WIDTH-1:0] wire_d9_100;
	wire [WIDTH-1:0] wire_d9_101;
	wire [WIDTH-1:0] wire_d9_102;
	wire [WIDTH-1:0] wire_d9_103;
	wire [WIDTH-1:0] wire_d9_104;
	wire [WIDTH-1:0] wire_d9_105;
	wire [WIDTH-1:0] wire_d9_106;
	wire [WIDTH-1:0] wire_d9_107;
	wire [WIDTH-1:0] wire_d9_108;
	wire [WIDTH-1:0] wire_d9_109;
	wire [WIDTH-1:0] wire_d9_110;
	wire [WIDTH-1:0] wire_d9_111;
	wire [WIDTH-1:0] wire_d9_112;
	wire [WIDTH-1:0] wire_d9_113;
	wire [WIDTH-1:0] wire_d9_114;
	wire [WIDTH-1:0] wire_d9_115;
	wire [WIDTH-1:0] wire_d9_116;
	wire [WIDTH-1:0] wire_d9_117;
	wire [WIDTH-1:0] wire_d9_118;
	wire [WIDTH-1:0] wire_d10_0;
	wire [WIDTH-1:0] wire_d10_1;
	wire [WIDTH-1:0] wire_d10_2;
	wire [WIDTH-1:0] wire_d10_3;
	wire [WIDTH-1:0] wire_d10_4;
	wire [WIDTH-1:0] wire_d10_5;
	wire [WIDTH-1:0] wire_d10_6;
	wire [WIDTH-1:0] wire_d10_7;
	wire [WIDTH-1:0] wire_d10_8;
	wire [WIDTH-1:0] wire_d10_9;
	wire [WIDTH-1:0] wire_d10_10;
	wire [WIDTH-1:0] wire_d10_11;
	wire [WIDTH-1:0] wire_d10_12;
	wire [WIDTH-1:0] wire_d10_13;
	wire [WIDTH-1:0] wire_d10_14;
	wire [WIDTH-1:0] wire_d10_15;
	wire [WIDTH-1:0] wire_d10_16;
	wire [WIDTH-1:0] wire_d10_17;
	wire [WIDTH-1:0] wire_d10_18;
	wire [WIDTH-1:0] wire_d10_19;
	wire [WIDTH-1:0] wire_d10_20;
	wire [WIDTH-1:0] wire_d10_21;
	wire [WIDTH-1:0] wire_d10_22;
	wire [WIDTH-1:0] wire_d10_23;
	wire [WIDTH-1:0] wire_d10_24;
	wire [WIDTH-1:0] wire_d10_25;
	wire [WIDTH-1:0] wire_d10_26;
	wire [WIDTH-1:0] wire_d10_27;
	wire [WIDTH-1:0] wire_d10_28;
	wire [WIDTH-1:0] wire_d10_29;
	wire [WIDTH-1:0] wire_d10_30;
	wire [WIDTH-1:0] wire_d10_31;
	wire [WIDTH-1:0] wire_d10_32;
	wire [WIDTH-1:0] wire_d10_33;
	wire [WIDTH-1:0] wire_d10_34;
	wire [WIDTH-1:0] wire_d10_35;
	wire [WIDTH-1:0] wire_d10_36;
	wire [WIDTH-1:0] wire_d10_37;
	wire [WIDTH-1:0] wire_d10_38;
	wire [WIDTH-1:0] wire_d10_39;
	wire [WIDTH-1:0] wire_d10_40;
	wire [WIDTH-1:0] wire_d10_41;
	wire [WIDTH-1:0] wire_d10_42;
	wire [WIDTH-1:0] wire_d10_43;
	wire [WIDTH-1:0] wire_d10_44;
	wire [WIDTH-1:0] wire_d10_45;
	wire [WIDTH-1:0] wire_d10_46;
	wire [WIDTH-1:0] wire_d10_47;
	wire [WIDTH-1:0] wire_d10_48;
	wire [WIDTH-1:0] wire_d10_49;
	wire [WIDTH-1:0] wire_d10_50;
	wire [WIDTH-1:0] wire_d10_51;
	wire [WIDTH-1:0] wire_d10_52;
	wire [WIDTH-1:0] wire_d10_53;
	wire [WIDTH-1:0] wire_d10_54;
	wire [WIDTH-1:0] wire_d10_55;
	wire [WIDTH-1:0] wire_d10_56;
	wire [WIDTH-1:0] wire_d10_57;
	wire [WIDTH-1:0] wire_d10_58;
	wire [WIDTH-1:0] wire_d10_59;
	wire [WIDTH-1:0] wire_d10_60;
	wire [WIDTH-1:0] wire_d10_61;
	wire [WIDTH-1:0] wire_d10_62;
	wire [WIDTH-1:0] wire_d10_63;
	wire [WIDTH-1:0] wire_d10_64;
	wire [WIDTH-1:0] wire_d10_65;
	wire [WIDTH-1:0] wire_d10_66;
	wire [WIDTH-1:0] wire_d10_67;
	wire [WIDTH-1:0] wire_d10_68;
	wire [WIDTH-1:0] wire_d10_69;
	wire [WIDTH-1:0] wire_d10_70;
	wire [WIDTH-1:0] wire_d10_71;
	wire [WIDTH-1:0] wire_d10_72;
	wire [WIDTH-1:0] wire_d10_73;
	wire [WIDTH-1:0] wire_d10_74;
	wire [WIDTH-1:0] wire_d10_75;
	wire [WIDTH-1:0] wire_d10_76;
	wire [WIDTH-1:0] wire_d10_77;
	wire [WIDTH-1:0] wire_d10_78;
	wire [WIDTH-1:0] wire_d10_79;
	wire [WIDTH-1:0] wire_d10_80;
	wire [WIDTH-1:0] wire_d10_81;
	wire [WIDTH-1:0] wire_d10_82;
	wire [WIDTH-1:0] wire_d10_83;
	wire [WIDTH-1:0] wire_d10_84;
	wire [WIDTH-1:0] wire_d10_85;
	wire [WIDTH-1:0] wire_d10_86;
	wire [WIDTH-1:0] wire_d10_87;
	wire [WIDTH-1:0] wire_d10_88;
	wire [WIDTH-1:0] wire_d10_89;
	wire [WIDTH-1:0] wire_d10_90;
	wire [WIDTH-1:0] wire_d10_91;
	wire [WIDTH-1:0] wire_d10_92;
	wire [WIDTH-1:0] wire_d10_93;
	wire [WIDTH-1:0] wire_d10_94;
	wire [WIDTH-1:0] wire_d10_95;
	wire [WIDTH-1:0] wire_d10_96;
	wire [WIDTH-1:0] wire_d10_97;
	wire [WIDTH-1:0] wire_d10_98;
	wire [WIDTH-1:0] wire_d10_99;
	wire [WIDTH-1:0] wire_d10_100;
	wire [WIDTH-1:0] wire_d10_101;
	wire [WIDTH-1:0] wire_d10_102;
	wire [WIDTH-1:0] wire_d10_103;
	wire [WIDTH-1:0] wire_d10_104;
	wire [WIDTH-1:0] wire_d10_105;
	wire [WIDTH-1:0] wire_d10_106;
	wire [WIDTH-1:0] wire_d10_107;
	wire [WIDTH-1:0] wire_d10_108;
	wire [WIDTH-1:0] wire_d10_109;
	wire [WIDTH-1:0] wire_d10_110;
	wire [WIDTH-1:0] wire_d10_111;
	wire [WIDTH-1:0] wire_d10_112;
	wire [WIDTH-1:0] wire_d10_113;
	wire [WIDTH-1:0] wire_d10_114;
	wire [WIDTH-1:0] wire_d10_115;
	wire [WIDTH-1:0] wire_d10_116;
	wire [WIDTH-1:0] wire_d10_117;
	wire [WIDTH-1:0] wire_d10_118;
	wire [WIDTH-1:0] wire_d11_0;
	wire [WIDTH-1:0] wire_d11_1;
	wire [WIDTH-1:0] wire_d11_2;
	wire [WIDTH-1:0] wire_d11_3;
	wire [WIDTH-1:0] wire_d11_4;
	wire [WIDTH-1:0] wire_d11_5;
	wire [WIDTH-1:0] wire_d11_6;
	wire [WIDTH-1:0] wire_d11_7;
	wire [WIDTH-1:0] wire_d11_8;
	wire [WIDTH-1:0] wire_d11_9;
	wire [WIDTH-1:0] wire_d11_10;
	wire [WIDTH-1:0] wire_d11_11;
	wire [WIDTH-1:0] wire_d11_12;
	wire [WIDTH-1:0] wire_d11_13;
	wire [WIDTH-1:0] wire_d11_14;
	wire [WIDTH-1:0] wire_d11_15;
	wire [WIDTH-1:0] wire_d11_16;
	wire [WIDTH-1:0] wire_d11_17;
	wire [WIDTH-1:0] wire_d11_18;
	wire [WIDTH-1:0] wire_d11_19;
	wire [WIDTH-1:0] wire_d11_20;
	wire [WIDTH-1:0] wire_d11_21;
	wire [WIDTH-1:0] wire_d11_22;
	wire [WIDTH-1:0] wire_d11_23;
	wire [WIDTH-1:0] wire_d11_24;
	wire [WIDTH-1:0] wire_d11_25;
	wire [WIDTH-1:0] wire_d11_26;
	wire [WIDTH-1:0] wire_d11_27;
	wire [WIDTH-1:0] wire_d11_28;
	wire [WIDTH-1:0] wire_d11_29;
	wire [WIDTH-1:0] wire_d11_30;
	wire [WIDTH-1:0] wire_d11_31;
	wire [WIDTH-1:0] wire_d11_32;
	wire [WIDTH-1:0] wire_d11_33;
	wire [WIDTH-1:0] wire_d11_34;
	wire [WIDTH-1:0] wire_d11_35;
	wire [WIDTH-1:0] wire_d11_36;
	wire [WIDTH-1:0] wire_d11_37;
	wire [WIDTH-1:0] wire_d11_38;
	wire [WIDTH-1:0] wire_d11_39;
	wire [WIDTH-1:0] wire_d11_40;
	wire [WIDTH-1:0] wire_d11_41;
	wire [WIDTH-1:0] wire_d11_42;
	wire [WIDTH-1:0] wire_d11_43;
	wire [WIDTH-1:0] wire_d11_44;
	wire [WIDTH-1:0] wire_d11_45;
	wire [WIDTH-1:0] wire_d11_46;
	wire [WIDTH-1:0] wire_d11_47;
	wire [WIDTH-1:0] wire_d11_48;
	wire [WIDTH-1:0] wire_d11_49;
	wire [WIDTH-1:0] wire_d11_50;
	wire [WIDTH-1:0] wire_d11_51;
	wire [WIDTH-1:0] wire_d11_52;
	wire [WIDTH-1:0] wire_d11_53;
	wire [WIDTH-1:0] wire_d11_54;
	wire [WIDTH-1:0] wire_d11_55;
	wire [WIDTH-1:0] wire_d11_56;
	wire [WIDTH-1:0] wire_d11_57;
	wire [WIDTH-1:0] wire_d11_58;
	wire [WIDTH-1:0] wire_d11_59;
	wire [WIDTH-1:0] wire_d11_60;
	wire [WIDTH-1:0] wire_d11_61;
	wire [WIDTH-1:0] wire_d11_62;
	wire [WIDTH-1:0] wire_d11_63;
	wire [WIDTH-1:0] wire_d11_64;
	wire [WIDTH-1:0] wire_d11_65;
	wire [WIDTH-1:0] wire_d11_66;
	wire [WIDTH-1:0] wire_d11_67;
	wire [WIDTH-1:0] wire_d11_68;
	wire [WIDTH-1:0] wire_d11_69;
	wire [WIDTH-1:0] wire_d11_70;
	wire [WIDTH-1:0] wire_d11_71;
	wire [WIDTH-1:0] wire_d11_72;
	wire [WIDTH-1:0] wire_d11_73;
	wire [WIDTH-1:0] wire_d11_74;
	wire [WIDTH-1:0] wire_d11_75;
	wire [WIDTH-1:0] wire_d11_76;
	wire [WIDTH-1:0] wire_d11_77;
	wire [WIDTH-1:0] wire_d11_78;
	wire [WIDTH-1:0] wire_d11_79;
	wire [WIDTH-1:0] wire_d11_80;
	wire [WIDTH-1:0] wire_d11_81;
	wire [WIDTH-1:0] wire_d11_82;
	wire [WIDTH-1:0] wire_d11_83;
	wire [WIDTH-1:0] wire_d11_84;
	wire [WIDTH-1:0] wire_d11_85;
	wire [WIDTH-1:0] wire_d11_86;
	wire [WIDTH-1:0] wire_d11_87;
	wire [WIDTH-1:0] wire_d11_88;
	wire [WIDTH-1:0] wire_d11_89;
	wire [WIDTH-1:0] wire_d11_90;
	wire [WIDTH-1:0] wire_d11_91;
	wire [WIDTH-1:0] wire_d11_92;
	wire [WIDTH-1:0] wire_d11_93;
	wire [WIDTH-1:0] wire_d11_94;
	wire [WIDTH-1:0] wire_d11_95;
	wire [WIDTH-1:0] wire_d11_96;
	wire [WIDTH-1:0] wire_d11_97;
	wire [WIDTH-1:0] wire_d11_98;
	wire [WIDTH-1:0] wire_d11_99;
	wire [WIDTH-1:0] wire_d11_100;
	wire [WIDTH-1:0] wire_d11_101;
	wire [WIDTH-1:0] wire_d11_102;
	wire [WIDTH-1:0] wire_d11_103;
	wire [WIDTH-1:0] wire_d11_104;
	wire [WIDTH-1:0] wire_d11_105;
	wire [WIDTH-1:0] wire_d11_106;
	wire [WIDTH-1:0] wire_d11_107;
	wire [WIDTH-1:0] wire_d11_108;
	wire [WIDTH-1:0] wire_d11_109;
	wire [WIDTH-1:0] wire_d11_110;
	wire [WIDTH-1:0] wire_d11_111;
	wire [WIDTH-1:0] wire_d11_112;
	wire [WIDTH-1:0] wire_d11_113;
	wire [WIDTH-1:0] wire_d11_114;
	wire [WIDTH-1:0] wire_d11_115;
	wire [WIDTH-1:0] wire_d11_116;
	wire [WIDTH-1:0] wire_d11_117;
	wire [WIDTH-1:0] wire_d11_118;
	wire [WIDTH-1:0] wire_d12_0;
	wire [WIDTH-1:0] wire_d12_1;
	wire [WIDTH-1:0] wire_d12_2;
	wire [WIDTH-1:0] wire_d12_3;
	wire [WIDTH-1:0] wire_d12_4;
	wire [WIDTH-1:0] wire_d12_5;
	wire [WIDTH-1:0] wire_d12_6;
	wire [WIDTH-1:0] wire_d12_7;
	wire [WIDTH-1:0] wire_d12_8;
	wire [WIDTH-1:0] wire_d12_9;
	wire [WIDTH-1:0] wire_d12_10;
	wire [WIDTH-1:0] wire_d12_11;
	wire [WIDTH-1:0] wire_d12_12;
	wire [WIDTH-1:0] wire_d12_13;
	wire [WIDTH-1:0] wire_d12_14;
	wire [WIDTH-1:0] wire_d12_15;
	wire [WIDTH-1:0] wire_d12_16;
	wire [WIDTH-1:0] wire_d12_17;
	wire [WIDTH-1:0] wire_d12_18;
	wire [WIDTH-1:0] wire_d12_19;
	wire [WIDTH-1:0] wire_d12_20;
	wire [WIDTH-1:0] wire_d12_21;
	wire [WIDTH-1:0] wire_d12_22;
	wire [WIDTH-1:0] wire_d12_23;
	wire [WIDTH-1:0] wire_d12_24;
	wire [WIDTH-1:0] wire_d12_25;
	wire [WIDTH-1:0] wire_d12_26;
	wire [WIDTH-1:0] wire_d12_27;
	wire [WIDTH-1:0] wire_d12_28;
	wire [WIDTH-1:0] wire_d12_29;
	wire [WIDTH-1:0] wire_d12_30;
	wire [WIDTH-1:0] wire_d12_31;
	wire [WIDTH-1:0] wire_d12_32;
	wire [WIDTH-1:0] wire_d12_33;
	wire [WIDTH-1:0] wire_d12_34;
	wire [WIDTH-1:0] wire_d12_35;
	wire [WIDTH-1:0] wire_d12_36;
	wire [WIDTH-1:0] wire_d12_37;
	wire [WIDTH-1:0] wire_d12_38;
	wire [WIDTH-1:0] wire_d12_39;
	wire [WIDTH-1:0] wire_d12_40;
	wire [WIDTH-1:0] wire_d12_41;
	wire [WIDTH-1:0] wire_d12_42;
	wire [WIDTH-1:0] wire_d12_43;
	wire [WIDTH-1:0] wire_d12_44;
	wire [WIDTH-1:0] wire_d12_45;
	wire [WIDTH-1:0] wire_d12_46;
	wire [WIDTH-1:0] wire_d12_47;
	wire [WIDTH-1:0] wire_d12_48;
	wire [WIDTH-1:0] wire_d12_49;
	wire [WIDTH-1:0] wire_d12_50;
	wire [WIDTH-1:0] wire_d12_51;
	wire [WIDTH-1:0] wire_d12_52;
	wire [WIDTH-1:0] wire_d12_53;
	wire [WIDTH-1:0] wire_d12_54;
	wire [WIDTH-1:0] wire_d12_55;
	wire [WIDTH-1:0] wire_d12_56;
	wire [WIDTH-1:0] wire_d12_57;
	wire [WIDTH-1:0] wire_d12_58;
	wire [WIDTH-1:0] wire_d12_59;
	wire [WIDTH-1:0] wire_d12_60;
	wire [WIDTH-1:0] wire_d12_61;
	wire [WIDTH-1:0] wire_d12_62;
	wire [WIDTH-1:0] wire_d12_63;
	wire [WIDTH-1:0] wire_d12_64;
	wire [WIDTH-1:0] wire_d12_65;
	wire [WIDTH-1:0] wire_d12_66;
	wire [WIDTH-1:0] wire_d12_67;
	wire [WIDTH-1:0] wire_d12_68;
	wire [WIDTH-1:0] wire_d12_69;
	wire [WIDTH-1:0] wire_d12_70;
	wire [WIDTH-1:0] wire_d12_71;
	wire [WIDTH-1:0] wire_d12_72;
	wire [WIDTH-1:0] wire_d12_73;
	wire [WIDTH-1:0] wire_d12_74;
	wire [WIDTH-1:0] wire_d12_75;
	wire [WIDTH-1:0] wire_d12_76;
	wire [WIDTH-1:0] wire_d12_77;
	wire [WIDTH-1:0] wire_d12_78;
	wire [WIDTH-1:0] wire_d12_79;
	wire [WIDTH-1:0] wire_d12_80;
	wire [WIDTH-1:0] wire_d12_81;
	wire [WIDTH-1:0] wire_d12_82;
	wire [WIDTH-1:0] wire_d12_83;
	wire [WIDTH-1:0] wire_d12_84;
	wire [WIDTH-1:0] wire_d12_85;
	wire [WIDTH-1:0] wire_d12_86;
	wire [WIDTH-1:0] wire_d12_87;
	wire [WIDTH-1:0] wire_d12_88;
	wire [WIDTH-1:0] wire_d12_89;
	wire [WIDTH-1:0] wire_d12_90;
	wire [WIDTH-1:0] wire_d12_91;
	wire [WIDTH-1:0] wire_d12_92;
	wire [WIDTH-1:0] wire_d12_93;
	wire [WIDTH-1:0] wire_d12_94;
	wire [WIDTH-1:0] wire_d12_95;
	wire [WIDTH-1:0] wire_d12_96;
	wire [WIDTH-1:0] wire_d12_97;
	wire [WIDTH-1:0] wire_d12_98;
	wire [WIDTH-1:0] wire_d12_99;
	wire [WIDTH-1:0] wire_d12_100;
	wire [WIDTH-1:0] wire_d12_101;
	wire [WIDTH-1:0] wire_d12_102;
	wire [WIDTH-1:0] wire_d12_103;
	wire [WIDTH-1:0] wire_d12_104;
	wire [WIDTH-1:0] wire_d12_105;
	wire [WIDTH-1:0] wire_d12_106;
	wire [WIDTH-1:0] wire_d12_107;
	wire [WIDTH-1:0] wire_d12_108;
	wire [WIDTH-1:0] wire_d12_109;
	wire [WIDTH-1:0] wire_d12_110;
	wire [WIDTH-1:0] wire_d12_111;
	wire [WIDTH-1:0] wire_d12_112;
	wire [WIDTH-1:0] wire_d12_113;
	wire [WIDTH-1:0] wire_d12_114;
	wire [WIDTH-1:0] wire_d12_115;
	wire [WIDTH-1:0] wire_d12_116;
	wire [WIDTH-1:0] wire_d12_117;
	wire [WIDTH-1:0] wire_d12_118;
	wire [WIDTH-1:0] wire_d13_0;
	wire [WIDTH-1:0] wire_d13_1;
	wire [WIDTH-1:0] wire_d13_2;
	wire [WIDTH-1:0] wire_d13_3;
	wire [WIDTH-1:0] wire_d13_4;
	wire [WIDTH-1:0] wire_d13_5;
	wire [WIDTH-1:0] wire_d13_6;
	wire [WIDTH-1:0] wire_d13_7;
	wire [WIDTH-1:0] wire_d13_8;
	wire [WIDTH-1:0] wire_d13_9;
	wire [WIDTH-1:0] wire_d13_10;
	wire [WIDTH-1:0] wire_d13_11;
	wire [WIDTH-1:0] wire_d13_12;
	wire [WIDTH-1:0] wire_d13_13;
	wire [WIDTH-1:0] wire_d13_14;
	wire [WIDTH-1:0] wire_d13_15;
	wire [WIDTH-1:0] wire_d13_16;
	wire [WIDTH-1:0] wire_d13_17;
	wire [WIDTH-1:0] wire_d13_18;
	wire [WIDTH-1:0] wire_d13_19;
	wire [WIDTH-1:0] wire_d13_20;
	wire [WIDTH-1:0] wire_d13_21;
	wire [WIDTH-1:0] wire_d13_22;
	wire [WIDTH-1:0] wire_d13_23;
	wire [WIDTH-1:0] wire_d13_24;
	wire [WIDTH-1:0] wire_d13_25;
	wire [WIDTH-1:0] wire_d13_26;
	wire [WIDTH-1:0] wire_d13_27;
	wire [WIDTH-1:0] wire_d13_28;
	wire [WIDTH-1:0] wire_d13_29;
	wire [WIDTH-1:0] wire_d13_30;
	wire [WIDTH-1:0] wire_d13_31;
	wire [WIDTH-1:0] wire_d13_32;
	wire [WIDTH-1:0] wire_d13_33;
	wire [WIDTH-1:0] wire_d13_34;
	wire [WIDTH-1:0] wire_d13_35;
	wire [WIDTH-1:0] wire_d13_36;
	wire [WIDTH-1:0] wire_d13_37;
	wire [WIDTH-1:0] wire_d13_38;
	wire [WIDTH-1:0] wire_d13_39;
	wire [WIDTH-1:0] wire_d13_40;
	wire [WIDTH-1:0] wire_d13_41;
	wire [WIDTH-1:0] wire_d13_42;
	wire [WIDTH-1:0] wire_d13_43;
	wire [WIDTH-1:0] wire_d13_44;
	wire [WIDTH-1:0] wire_d13_45;
	wire [WIDTH-1:0] wire_d13_46;
	wire [WIDTH-1:0] wire_d13_47;
	wire [WIDTH-1:0] wire_d13_48;
	wire [WIDTH-1:0] wire_d13_49;
	wire [WIDTH-1:0] wire_d13_50;
	wire [WIDTH-1:0] wire_d13_51;
	wire [WIDTH-1:0] wire_d13_52;
	wire [WIDTH-1:0] wire_d13_53;
	wire [WIDTH-1:0] wire_d13_54;
	wire [WIDTH-1:0] wire_d13_55;
	wire [WIDTH-1:0] wire_d13_56;
	wire [WIDTH-1:0] wire_d13_57;
	wire [WIDTH-1:0] wire_d13_58;
	wire [WIDTH-1:0] wire_d13_59;
	wire [WIDTH-1:0] wire_d13_60;
	wire [WIDTH-1:0] wire_d13_61;
	wire [WIDTH-1:0] wire_d13_62;
	wire [WIDTH-1:0] wire_d13_63;
	wire [WIDTH-1:0] wire_d13_64;
	wire [WIDTH-1:0] wire_d13_65;
	wire [WIDTH-1:0] wire_d13_66;
	wire [WIDTH-1:0] wire_d13_67;
	wire [WIDTH-1:0] wire_d13_68;
	wire [WIDTH-1:0] wire_d13_69;
	wire [WIDTH-1:0] wire_d13_70;
	wire [WIDTH-1:0] wire_d13_71;
	wire [WIDTH-1:0] wire_d13_72;
	wire [WIDTH-1:0] wire_d13_73;
	wire [WIDTH-1:0] wire_d13_74;
	wire [WIDTH-1:0] wire_d13_75;
	wire [WIDTH-1:0] wire_d13_76;
	wire [WIDTH-1:0] wire_d13_77;
	wire [WIDTH-1:0] wire_d13_78;
	wire [WIDTH-1:0] wire_d13_79;
	wire [WIDTH-1:0] wire_d13_80;
	wire [WIDTH-1:0] wire_d13_81;
	wire [WIDTH-1:0] wire_d13_82;
	wire [WIDTH-1:0] wire_d13_83;
	wire [WIDTH-1:0] wire_d13_84;
	wire [WIDTH-1:0] wire_d13_85;
	wire [WIDTH-1:0] wire_d13_86;
	wire [WIDTH-1:0] wire_d13_87;
	wire [WIDTH-1:0] wire_d13_88;
	wire [WIDTH-1:0] wire_d13_89;
	wire [WIDTH-1:0] wire_d13_90;
	wire [WIDTH-1:0] wire_d13_91;
	wire [WIDTH-1:0] wire_d13_92;
	wire [WIDTH-1:0] wire_d13_93;
	wire [WIDTH-1:0] wire_d13_94;
	wire [WIDTH-1:0] wire_d13_95;
	wire [WIDTH-1:0] wire_d13_96;
	wire [WIDTH-1:0] wire_d13_97;
	wire [WIDTH-1:0] wire_d13_98;
	wire [WIDTH-1:0] wire_d13_99;
	wire [WIDTH-1:0] wire_d13_100;
	wire [WIDTH-1:0] wire_d13_101;
	wire [WIDTH-1:0] wire_d13_102;
	wire [WIDTH-1:0] wire_d13_103;
	wire [WIDTH-1:0] wire_d13_104;
	wire [WIDTH-1:0] wire_d13_105;
	wire [WIDTH-1:0] wire_d13_106;
	wire [WIDTH-1:0] wire_d13_107;
	wire [WIDTH-1:0] wire_d13_108;
	wire [WIDTH-1:0] wire_d13_109;
	wire [WIDTH-1:0] wire_d13_110;
	wire [WIDTH-1:0] wire_d13_111;
	wire [WIDTH-1:0] wire_d13_112;
	wire [WIDTH-1:0] wire_d13_113;
	wire [WIDTH-1:0] wire_d13_114;
	wire [WIDTH-1:0] wire_d13_115;
	wire [WIDTH-1:0] wire_d13_116;
	wire [WIDTH-1:0] wire_d13_117;
	wire [WIDTH-1:0] wire_d13_118;
	wire [WIDTH-1:0] wire_d14_0;
	wire [WIDTH-1:0] wire_d14_1;
	wire [WIDTH-1:0] wire_d14_2;
	wire [WIDTH-1:0] wire_d14_3;
	wire [WIDTH-1:0] wire_d14_4;
	wire [WIDTH-1:0] wire_d14_5;
	wire [WIDTH-1:0] wire_d14_6;
	wire [WIDTH-1:0] wire_d14_7;
	wire [WIDTH-1:0] wire_d14_8;
	wire [WIDTH-1:0] wire_d14_9;
	wire [WIDTH-1:0] wire_d14_10;
	wire [WIDTH-1:0] wire_d14_11;
	wire [WIDTH-1:0] wire_d14_12;
	wire [WIDTH-1:0] wire_d14_13;
	wire [WIDTH-1:0] wire_d14_14;
	wire [WIDTH-1:0] wire_d14_15;
	wire [WIDTH-1:0] wire_d14_16;
	wire [WIDTH-1:0] wire_d14_17;
	wire [WIDTH-1:0] wire_d14_18;
	wire [WIDTH-1:0] wire_d14_19;
	wire [WIDTH-1:0] wire_d14_20;
	wire [WIDTH-1:0] wire_d14_21;
	wire [WIDTH-1:0] wire_d14_22;
	wire [WIDTH-1:0] wire_d14_23;
	wire [WIDTH-1:0] wire_d14_24;
	wire [WIDTH-1:0] wire_d14_25;
	wire [WIDTH-1:0] wire_d14_26;
	wire [WIDTH-1:0] wire_d14_27;
	wire [WIDTH-1:0] wire_d14_28;
	wire [WIDTH-1:0] wire_d14_29;
	wire [WIDTH-1:0] wire_d14_30;
	wire [WIDTH-1:0] wire_d14_31;
	wire [WIDTH-1:0] wire_d14_32;
	wire [WIDTH-1:0] wire_d14_33;
	wire [WIDTH-1:0] wire_d14_34;
	wire [WIDTH-1:0] wire_d14_35;
	wire [WIDTH-1:0] wire_d14_36;
	wire [WIDTH-1:0] wire_d14_37;
	wire [WIDTH-1:0] wire_d14_38;
	wire [WIDTH-1:0] wire_d14_39;
	wire [WIDTH-1:0] wire_d14_40;
	wire [WIDTH-1:0] wire_d14_41;
	wire [WIDTH-1:0] wire_d14_42;
	wire [WIDTH-1:0] wire_d14_43;
	wire [WIDTH-1:0] wire_d14_44;
	wire [WIDTH-1:0] wire_d14_45;
	wire [WIDTH-1:0] wire_d14_46;
	wire [WIDTH-1:0] wire_d14_47;
	wire [WIDTH-1:0] wire_d14_48;
	wire [WIDTH-1:0] wire_d14_49;
	wire [WIDTH-1:0] wire_d14_50;
	wire [WIDTH-1:0] wire_d14_51;
	wire [WIDTH-1:0] wire_d14_52;
	wire [WIDTH-1:0] wire_d14_53;
	wire [WIDTH-1:0] wire_d14_54;
	wire [WIDTH-1:0] wire_d14_55;
	wire [WIDTH-1:0] wire_d14_56;
	wire [WIDTH-1:0] wire_d14_57;
	wire [WIDTH-1:0] wire_d14_58;
	wire [WIDTH-1:0] wire_d14_59;
	wire [WIDTH-1:0] wire_d14_60;
	wire [WIDTH-1:0] wire_d14_61;
	wire [WIDTH-1:0] wire_d14_62;
	wire [WIDTH-1:0] wire_d14_63;
	wire [WIDTH-1:0] wire_d14_64;
	wire [WIDTH-1:0] wire_d14_65;
	wire [WIDTH-1:0] wire_d14_66;
	wire [WIDTH-1:0] wire_d14_67;
	wire [WIDTH-1:0] wire_d14_68;
	wire [WIDTH-1:0] wire_d14_69;
	wire [WIDTH-1:0] wire_d14_70;
	wire [WIDTH-1:0] wire_d14_71;
	wire [WIDTH-1:0] wire_d14_72;
	wire [WIDTH-1:0] wire_d14_73;
	wire [WIDTH-1:0] wire_d14_74;
	wire [WIDTH-1:0] wire_d14_75;
	wire [WIDTH-1:0] wire_d14_76;
	wire [WIDTH-1:0] wire_d14_77;
	wire [WIDTH-1:0] wire_d14_78;
	wire [WIDTH-1:0] wire_d14_79;
	wire [WIDTH-1:0] wire_d14_80;
	wire [WIDTH-1:0] wire_d14_81;
	wire [WIDTH-1:0] wire_d14_82;
	wire [WIDTH-1:0] wire_d14_83;
	wire [WIDTH-1:0] wire_d14_84;
	wire [WIDTH-1:0] wire_d14_85;
	wire [WIDTH-1:0] wire_d14_86;
	wire [WIDTH-1:0] wire_d14_87;
	wire [WIDTH-1:0] wire_d14_88;
	wire [WIDTH-1:0] wire_d14_89;
	wire [WIDTH-1:0] wire_d14_90;
	wire [WIDTH-1:0] wire_d14_91;
	wire [WIDTH-1:0] wire_d14_92;
	wire [WIDTH-1:0] wire_d14_93;
	wire [WIDTH-1:0] wire_d14_94;
	wire [WIDTH-1:0] wire_d14_95;
	wire [WIDTH-1:0] wire_d14_96;
	wire [WIDTH-1:0] wire_d14_97;
	wire [WIDTH-1:0] wire_d14_98;
	wire [WIDTH-1:0] wire_d14_99;
	wire [WIDTH-1:0] wire_d14_100;
	wire [WIDTH-1:0] wire_d14_101;
	wire [WIDTH-1:0] wire_d14_102;
	wire [WIDTH-1:0] wire_d14_103;
	wire [WIDTH-1:0] wire_d14_104;
	wire [WIDTH-1:0] wire_d14_105;
	wire [WIDTH-1:0] wire_d14_106;
	wire [WIDTH-1:0] wire_d14_107;
	wire [WIDTH-1:0] wire_d14_108;
	wire [WIDTH-1:0] wire_d14_109;
	wire [WIDTH-1:0] wire_d14_110;
	wire [WIDTH-1:0] wire_d14_111;
	wire [WIDTH-1:0] wire_d14_112;
	wire [WIDTH-1:0] wire_d14_113;
	wire [WIDTH-1:0] wire_d14_114;
	wire [WIDTH-1:0] wire_d14_115;
	wire [WIDTH-1:0] wire_d14_116;
	wire [WIDTH-1:0] wire_d14_117;
	wire [WIDTH-1:0] wire_d14_118;
	wire [WIDTH-1:0] wire_d15_0;
	wire [WIDTH-1:0] wire_d15_1;
	wire [WIDTH-1:0] wire_d15_2;
	wire [WIDTH-1:0] wire_d15_3;
	wire [WIDTH-1:0] wire_d15_4;
	wire [WIDTH-1:0] wire_d15_5;
	wire [WIDTH-1:0] wire_d15_6;
	wire [WIDTH-1:0] wire_d15_7;
	wire [WIDTH-1:0] wire_d15_8;
	wire [WIDTH-1:0] wire_d15_9;
	wire [WIDTH-1:0] wire_d15_10;
	wire [WIDTH-1:0] wire_d15_11;
	wire [WIDTH-1:0] wire_d15_12;
	wire [WIDTH-1:0] wire_d15_13;
	wire [WIDTH-1:0] wire_d15_14;
	wire [WIDTH-1:0] wire_d15_15;
	wire [WIDTH-1:0] wire_d15_16;
	wire [WIDTH-1:0] wire_d15_17;
	wire [WIDTH-1:0] wire_d15_18;
	wire [WIDTH-1:0] wire_d15_19;
	wire [WIDTH-1:0] wire_d15_20;
	wire [WIDTH-1:0] wire_d15_21;
	wire [WIDTH-1:0] wire_d15_22;
	wire [WIDTH-1:0] wire_d15_23;
	wire [WIDTH-1:0] wire_d15_24;
	wire [WIDTH-1:0] wire_d15_25;
	wire [WIDTH-1:0] wire_d15_26;
	wire [WIDTH-1:0] wire_d15_27;
	wire [WIDTH-1:0] wire_d15_28;
	wire [WIDTH-1:0] wire_d15_29;
	wire [WIDTH-1:0] wire_d15_30;
	wire [WIDTH-1:0] wire_d15_31;
	wire [WIDTH-1:0] wire_d15_32;
	wire [WIDTH-1:0] wire_d15_33;
	wire [WIDTH-1:0] wire_d15_34;
	wire [WIDTH-1:0] wire_d15_35;
	wire [WIDTH-1:0] wire_d15_36;
	wire [WIDTH-1:0] wire_d15_37;
	wire [WIDTH-1:0] wire_d15_38;
	wire [WIDTH-1:0] wire_d15_39;
	wire [WIDTH-1:0] wire_d15_40;
	wire [WIDTH-1:0] wire_d15_41;
	wire [WIDTH-1:0] wire_d15_42;
	wire [WIDTH-1:0] wire_d15_43;
	wire [WIDTH-1:0] wire_d15_44;
	wire [WIDTH-1:0] wire_d15_45;
	wire [WIDTH-1:0] wire_d15_46;
	wire [WIDTH-1:0] wire_d15_47;
	wire [WIDTH-1:0] wire_d15_48;
	wire [WIDTH-1:0] wire_d15_49;
	wire [WIDTH-1:0] wire_d15_50;
	wire [WIDTH-1:0] wire_d15_51;
	wire [WIDTH-1:0] wire_d15_52;
	wire [WIDTH-1:0] wire_d15_53;
	wire [WIDTH-1:0] wire_d15_54;
	wire [WIDTH-1:0] wire_d15_55;
	wire [WIDTH-1:0] wire_d15_56;
	wire [WIDTH-1:0] wire_d15_57;
	wire [WIDTH-1:0] wire_d15_58;
	wire [WIDTH-1:0] wire_d15_59;
	wire [WIDTH-1:0] wire_d15_60;
	wire [WIDTH-1:0] wire_d15_61;
	wire [WIDTH-1:0] wire_d15_62;
	wire [WIDTH-1:0] wire_d15_63;
	wire [WIDTH-1:0] wire_d15_64;
	wire [WIDTH-1:0] wire_d15_65;
	wire [WIDTH-1:0] wire_d15_66;
	wire [WIDTH-1:0] wire_d15_67;
	wire [WIDTH-1:0] wire_d15_68;
	wire [WIDTH-1:0] wire_d15_69;
	wire [WIDTH-1:0] wire_d15_70;
	wire [WIDTH-1:0] wire_d15_71;
	wire [WIDTH-1:0] wire_d15_72;
	wire [WIDTH-1:0] wire_d15_73;
	wire [WIDTH-1:0] wire_d15_74;
	wire [WIDTH-1:0] wire_d15_75;
	wire [WIDTH-1:0] wire_d15_76;
	wire [WIDTH-1:0] wire_d15_77;
	wire [WIDTH-1:0] wire_d15_78;
	wire [WIDTH-1:0] wire_d15_79;
	wire [WIDTH-1:0] wire_d15_80;
	wire [WIDTH-1:0] wire_d15_81;
	wire [WIDTH-1:0] wire_d15_82;
	wire [WIDTH-1:0] wire_d15_83;
	wire [WIDTH-1:0] wire_d15_84;
	wire [WIDTH-1:0] wire_d15_85;
	wire [WIDTH-1:0] wire_d15_86;
	wire [WIDTH-1:0] wire_d15_87;
	wire [WIDTH-1:0] wire_d15_88;
	wire [WIDTH-1:0] wire_d15_89;
	wire [WIDTH-1:0] wire_d15_90;
	wire [WIDTH-1:0] wire_d15_91;
	wire [WIDTH-1:0] wire_d15_92;
	wire [WIDTH-1:0] wire_d15_93;
	wire [WIDTH-1:0] wire_d15_94;
	wire [WIDTH-1:0] wire_d15_95;
	wire [WIDTH-1:0] wire_d15_96;
	wire [WIDTH-1:0] wire_d15_97;
	wire [WIDTH-1:0] wire_d15_98;
	wire [WIDTH-1:0] wire_d15_99;
	wire [WIDTH-1:0] wire_d15_100;
	wire [WIDTH-1:0] wire_d15_101;
	wire [WIDTH-1:0] wire_d15_102;
	wire [WIDTH-1:0] wire_d15_103;
	wire [WIDTH-1:0] wire_d15_104;
	wire [WIDTH-1:0] wire_d15_105;
	wire [WIDTH-1:0] wire_d15_106;
	wire [WIDTH-1:0] wire_d15_107;
	wire [WIDTH-1:0] wire_d15_108;
	wire [WIDTH-1:0] wire_d15_109;
	wire [WIDTH-1:0] wire_d15_110;
	wire [WIDTH-1:0] wire_d15_111;
	wire [WIDTH-1:0] wire_d15_112;
	wire [WIDTH-1:0] wire_d15_113;
	wire [WIDTH-1:0] wire_d15_114;
	wire [WIDTH-1:0] wire_d15_115;
	wire [WIDTH-1:0] wire_d15_116;
	wire [WIDTH-1:0] wire_d15_117;
	wire [WIDTH-1:0] wire_d15_118;
	wire [WIDTH-1:0] wire_d16_0;
	wire [WIDTH-1:0] wire_d16_1;
	wire [WIDTH-1:0] wire_d16_2;
	wire [WIDTH-1:0] wire_d16_3;
	wire [WIDTH-1:0] wire_d16_4;
	wire [WIDTH-1:0] wire_d16_5;
	wire [WIDTH-1:0] wire_d16_6;
	wire [WIDTH-1:0] wire_d16_7;
	wire [WIDTH-1:0] wire_d16_8;
	wire [WIDTH-1:0] wire_d16_9;
	wire [WIDTH-1:0] wire_d16_10;
	wire [WIDTH-1:0] wire_d16_11;
	wire [WIDTH-1:0] wire_d16_12;
	wire [WIDTH-1:0] wire_d16_13;
	wire [WIDTH-1:0] wire_d16_14;
	wire [WIDTH-1:0] wire_d16_15;
	wire [WIDTH-1:0] wire_d16_16;
	wire [WIDTH-1:0] wire_d16_17;
	wire [WIDTH-1:0] wire_d16_18;
	wire [WIDTH-1:0] wire_d16_19;
	wire [WIDTH-1:0] wire_d16_20;
	wire [WIDTH-1:0] wire_d16_21;
	wire [WIDTH-1:0] wire_d16_22;
	wire [WIDTH-1:0] wire_d16_23;
	wire [WIDTH-1:0] wire_d16_24;
	wire [WIDTH-1:0] wire_d16_25;
	wire [WIDTH-1:0] wire_d16_26;
	wire [WIDTH-1:0] wire_d16_27;
	wire [WIDTH-1:0] wire_d16_28;
	wire [WIDTH-1:0] wire_d16_29;
	wire [WIDTH-1:0] wire_d16_30;
	wire [WIDTH-1:0] wire_d16_31;
	wire [WIDTH-1:0] wire_d16_32;
	wire [WIDTH-1:0] wire_d16_33;
	wire [WIDTH-1:0] wire_d16_34;
	wire [WIDTH-1:0] wire_d16_35;
	wire [WIDTH-1:0] wire_d16_36;
	wire [WIDTH-1:0] wire_d16_37;
	wire [WIDTH-1:0] wire_d16_38;
	wire [WIDTH-1:0] wire_d16_39;
	wire [WIDTH-1:0] wire_d16_40;
	wire [WIDTH-1:0] wire_d16_41;
	wire [WIDTH-1:0] wire_d16_42;
	wire [WIDTH-1:0] wire_d16_43;
	wire [WIDTH-1:0] wire_d16_44;
	wire [WIDTH-1:0] wire_d16_45;
	wire [WIDTH-1:0] wire_d16_46;
	wire [WIDTH-1:0] wire_d16_47;
	wire [WIDTH-1:0] wire_d16_48;
	wire [WIDTH-1:0] wire_d16_49;
	wire [WIDTH-1:0] wire_d16_50;
	wire [WIDTH-1:0] wire_d16_51;
	wire [WIDTH-1:0] wire_d16_52;
	wire [WIDTH-1:0] wire_d16_53;
	wire [WIDTH-1:0] wire_d16_54;
	wire [WIDTH-1:0] wire_d16_55;
	wire [WIDTH-1:0] wire_d16_56;
	wire [WIDTH-1:0] wire_d16_57;
	wire [WIDTH-1:0] wire_d16_58;
	wire [WIDTH-1:0] wire_d16_59;
	wire [WIDTH-1:0] wire_d16_60;
	wire [WIDTH-1:0] wire_d16_61;
	wire [WIDTH-1:0] wire_d16_62;
	wire [WIDTH-1:0] wire_d16_63;
	wire [WIDTH-1:0] wire_d16_64;
	wire [WIDTH-1:0] wire_d16_65;
	wire [WIDTH-1:0] wire_d16_66;
	wire [WIDTH-1:0] wire_d16_67;
	wire [WIDTH-1:0] wire_d16_68;
	wire [WIDTH-1:0] wire_d16_69;
	wire [WIDTH-1:0] wire_d16_70;
	wire [WIDTH-1:0] wire_d16_71;
	wire [WIDTH-1:0] wire_d16_72;
	wire [WIDTH-1:0] wire_d16_73;
	wire [WIDTH-1:0] wire_d16_74;
	wire [WIDTH-1:0] wire_d16_75;
	wire [WIDTH-1:0] wire_d16_76;
	wire [WIDTH-1:0] wire_d16_77;
	wire [WIDTH-1:0] wire_d16_78;
	wire [WIDTH-1:0] wire_d16_79;
	wire [WIDTH-1:0] wire_d16_80;
	wire [WIDTH-1:0] wire_d16_81;
	wire [WIDTH-1:0] wire_d16_82;
	wire [WIDTH-1:0] wire_d16_83;
	wire [WIDTH-1:0] wire_d16_84;
	wire [WIDTH-1:0] wire_d16_85;
	wire [WIDTH-1:0] wire_d16_86;
	wire [WIDTH-1:0] wire_d16_87;
	wire [WIDTH-1:0] wire_d16_88;
	wire [WIDTH-1:0] wire_d16_89;
	wire [WIDTH-1:0] wire_d16_90;
	wire [WIDTH-1:0] wire_d16_91;
	wire [WIDTH-1:0] wire_d16_92;
	wire [WIDTH-1:0] wire_d16_93;
	wire [WIDTH-1:0] wire_d16_94;
	wire [WIDTH-1:0] wire_d16_95;
	wire [WIDTH-1:0] wire_d16_96;
	wire [WIDTH-1:0] wire_d16_97;
	wire [WIDTH-1:0] wire_d16_98;
	wire [WIDTH-1:0] wire_d16_99;
	wire [WIDTH-1:0] wire_d16_100;
	wire [WIDTH-1:0] wire_d16_101;
	wire [WIDTH-1:0] wire_d16_102;
	wire [WIDTH-1:0] wire_d16_103;
	wire [WIDTH-1:0] wire_d16_104;
	wire [WIDTH-1:0] wire_d16_105;
	wire [WIDTH-1:0] wire_d16_106;
	wire [WIDTH-1:0] wire_d16_107;
	wire [WIDTH-1:0] wire_d16_108;
	wire [WIDTH-1:0] wire_d16_109;
	wire [WIDTH-1:0] wire_d16_110;
	wire [WIDTH-1:0] wire_d16_111;
	wire [WIDTH-1:0] wire_d16_112;
	wire [WIDTH-1:0] wire_d16_113;
	wire [WIDTH-1:0] wire_d16_114;
	wire [WIDTH-1:0] wire_d16_115;
	wire [WIDTH-1:0] wire_d16_116;
	wire [WIDTH-1:0] wire_d16_117;
	wire [WIDTH-1:0] wire_d16_118;
	wire [WIDTH-1:0] wire_d17_0;
	wire [WIDTH-1:0] wire_d17_1;
	wire [WIDTH-1:0] wire_d17_2;
	wire [WIDTH-1:0] wire_d17_3;
	wire [WIDTH-1:0] wire_d17_4;
	wire [WIDTH-1:0] wire_d17_5;
	wire [WIDTH-1:0] wire_d17_6;
	wire [WIDTH-1:0] wire_d17_7;
	wire [WIDTH-1:0] wire_d17_8;
	wire [WIDTH-1:0] wire_d17_9;
	wire [WIDTH-1:0] wire_d17_10;
	wire [WIDTH-1:0] wire_d17_11;
	wire [WIDTH-1:0] wire_d17_12;
	wire [WIDTH-1:0] wire_d17_13;
	wire [WIDTH-1:0] wire_d17_14;
	wire [WIDTH-1:0] wire_d17_15;
	wire [WIDTH-1:0] wire_d17_16;
	wire [WIDTH-1:0] wire_d17_17;
	wire [WIDTH-1:0] wire_d17_18;
	wire [WIDTH-1:0] wire_d17_19;
	wire [WIDTH-1:0] wire_d17_20;
	wire [WIDTH-1:0] wire_d17_21;
	wire [WIDTH-1:0] wire_d17_22;
	wire [WIDTH-1:0] wire_d17_23;
	wire [WIDTH-1:0] wire_d17_24;
	wire [WIDTH-1:0] wire_d17_25;
	wire [WIDTH-1:0] wire_d17_26;
	wire [WIDTH-1:0] wire_d17_27;
	wire [WIDTH-1:0] wire_d17_28;
	wire [WIDTH-1:0] wire_d17_29;
	wire [WIDTH-1:0] wire_d17_30;
	wire [WIDTH-1:0] wire_d17_31;
	wire [WIDTH-1:0] wire_d17_32;
	wire [WIDTH-1:0] wire_d17_33;
	wire [WIDTH-1:0] wire_d17_34;
	wire [WIDTH-1:0] wire_d17_35;
	wire [WIDTH-1:0] wire_d17_36;
	wire [WIDTH-1:0] wire_d17_37;
	wire [WIDTH-1:0] wire_d17_38;
	wire [WIDTH-1:0] wire_d17_39;
	wire [WIDTH-1:0] wire_d17_40;
	wire [WIDTH-1:0] wire_d17_41;
	wire [WIDTH-1:0] wire_d17_42;
	wire [WIDTH-1:0] wire_d17_43;
	wire [WIDTH-1:0] wire_d17_44;
	wire [WIDTH-1:0] wire_d17_45;
	wire [WIDTH-1:0] wire_d17_46;
	wire [WIDTH-1:0] wire_d17_47;
	wire [WIDTH-1:0] wire_d17_48;
	wire [WIDTH-1:0] wire_d17_49;
	wire [WIDTH-1:0] wire_d17_50;
	wire [WIDTH-1:0] wire_d17_51;
	wire [WIDTH-1:0] wire_d17_52;
	wire [WIDTH-1:0] wire_d17_53;
	wire [WIDTH-1:0] wire_d17_54;
	wire [WIDTH-1:0] wire_d17_55;
	wire [WIDTH-1:0] wire_d17_56;
	wire [WIDTH-1:0] wire_d17_57;
	wire [WIDTH-1:0] wire_d17_58;
	wire [WIDTH-1:0] wire_d17_59;
	wire [WIDTH-1:0] wire_d17_60;
	wire [WIDTH-1:0] wire_d17_61;
	wire [WIDTH-1:0] wire_d17_62;
	wire [WIDTH-1:0] wire_d17_63;
	wire [WIDTH-1:0] wire_d17_64;
	wire [WIDTH-1:0] wire_d17_65;
	wire [WIDTH-1:0] wire_d17_66;
	wire [WIDTH-1:0] wire_d17_67;
	wire [WIDTH-1:0] wire_d17_68;
	wire [WIDTH-1:0] wire_d17_69;
	wire [WIDTH-1:0] wire_d17_70;
	wire [WIDTH-1:0] wire_d17_71;
	wire [WIDTH-1:0] wire_d17_72;
	wire [WIDTH-1:0] wire_d17_73;
	wire [WIDTH-1:0] wire_d17_74;
	wire [WIDTH-1:0] wire_d17_75;
	wire [WIDTH-1:0] wire_d17_76;
	wire [WIDTH-1:0] wire_d17_77;
	wire [WIDTH-1:0] wire_d17_78;
	wire [WIDTH-1:0] wire_d17_79;
	wire [WIDTH-1:0] wire_d17_80;
	wire [WIDTH-1:0] wire_d17_81;
	wire [WIDTH-1:0] wire_d17_82;
	wire [WIDTH-1:0] wire_d17_83;
	wire [WIDTH-1:0] wire_d17_84;
	wire [WIDTH-1:0] wire_d17_85;
	wire [WIDTH-1:0] wire_d17_86;
	wire [WIDTH-1:0] wire_d17_87;
	wire [WIDTH-1:0] wire_d17_88;
	wire [WIDTH-1:0] wire_d17_89;
	wire [WIDTH-1:0] wire_d17_90;
	wire [WIDTH-1:0] wire_d17_91;
	wire [WIDTH-1:0] wire_d17_92;
	wire [WIDTH-1:0] wire_d17_93;
	wire [WIDTH-1:0] wire_d17_94;
	wire [WIDTH-1:0] wire_d17_95;
	wire [WIDTH-1:0] wire_d17_96;
	wire [WIDTH-1:0] wire_d17_97;
	wire [WIDTH-1:0] wire_d17_98;
	wire [WIDTH-1:0] wire_d17_99;
	wire [WIDTH-1:0] wire_d17_100;
	wire [WIDTH-1:0] wire_d17_101;
	wire [WIDTH-1:0] wire_d17_102;
	wire [WIDTH-1:0] wire_d17_103;
	wire [WIDTH-1:0] wire_d17_104;
	wire [WIDTH-1:0] wire_d17_105;
	wire [WIDTH-1:0] wire_d17_106;
	wire [WIDTH-1:0] wire_d17_107;
	wire [WIDTH-1:0] wire_d17_108;
	wire [WIDTH-1:0] wire_d17_109;
	wire [WIDTH-1:0] wire_d17_110;
	wire [WIDTH-1:0] wire_d17_111;
	wire [WIDTH-1:0] wire_d17_112;
	wire [WIDTH-1:0] wire_d17_113;
	wire [WIDTH-1:0] wire_d17_114;
	wire [WIDTH-1:0] wire_d17_115;
	wire [WIDTH-1:0] wire_d17_116;
	wire [WIDTH-1:0] wire_d17_117;
	wire [WIDTH-1:0] wire_d17_118;
	wire [WIDTH-1:0] wire_d18_0;
	wire [WIDTH-1:0] wire_d18_1;
	wire [WIDTH-1:0] wire_d18_2;
	wire [WIDTH-1:0] wire_d18_3;
	wire [WIDTH-1:0] wire_d18_4;
	wire [WIDTH-1:0] wire_d18_5;
	wire [WIDTH-1:0] wire_d18_6;
	wire [WIDTH-1:0] wire_d18_7;
	wire [WIDTH-1:0] wire_d18_8;
	wire [WIDTH-1:0] wire_d18_9;
	wire [WIDTH-1:0] wire_d18_10;
	wire [WIDTH-1:0] wire_d18_11;
	wire [WIDTH-1:0] wire_d18_12;
	wire [WIDTH-1:0] wire_d18_13;
	wire [WIDTH-1:0] wire_d18_14;
	wire [WIDTH-1:0] wire_d18_15;
	wire [WIDTH-1:0] wire_d18_16;
	wire [WIDTH-1:0] wire_d18_17;
	wire [WIDTH-1:0] wire_d18_18;
	wire [WIDTH-1:0] wire_d18_19;
	wire [WIDTH-1:0] wire_d18_20;
	wire [WIDTH-1:0] wire_d18_21;
	wire [WIDTH-1:0] wire_d18_22;
	wire [WIDTH-1:0] wire_d18_23;
	wire [WIDTH-1:0] wire_d18_24;
	wire [WIDTH-1:0] wire_d18_25;
	wire [WIDTH-1:0] wire_d18_26;
	wire [WIDTH-1:0] wire_d18_27;
	wire [WIDTH-1:0] wire_d18_28;
	wire [WIDTH-1:0] wire_d18_29;
	wire [WIDTH-1:0] wire_d18_30;
	wire [WIDTH-1:0] wire_d18_31;
	wire [WIDTH-1:0] wire_d18_32;
	wire [WIDTH-1:0] wire_d18_33;
	wire [WIDTH-1:0] wire_d18_34;
	wire [WIDTH-1:0] wire_d18_35;
	wire [WIDTH-1:0] wire_d18_36;
	wire [WIDTH-1:0] wire_d18_37;
	wire [WIDTH-1:0] wire_d18_38;
	wire [WIDTH-1:0] wire_d18_39;
	wire [WIDTH-1:0] wire_d18_40;
	wire [WIDTH-1:0] wire_d18_41;
	wire [WIDTH-1:0] wire_d18_42;
	wire [WIDTH-1:0] wire_d18_43;
	wire [WIDTH-1:0] wire_d18_44;
	wire [WIDTH-1:0] wire_d18_45;
	wire [WIDTH-1:0] wire_d18_46;
	wire [WIDTH-1:0] wire_d18_47;
	wire [WIDTH-1:0] wire_d18_48;
	wire [WIDTH-1:0] wire_d18_49;
	wire [WIDTH-1:0] wire_d18_50;
	wire [WIDTH-1:0] wire_d18_51;
	wire [WIDTH-1:0] wire_d18_52;
	wire [WIDTH-1:0] wire_d18_53;
	wire [WIDTH-1:0] wire_d18_54;
	wire [WIDTH-1:0] wire_d18_55;
	wire [WIDTH-1:0] wire_d18_56;
	wire [WIDTH-1:0] wire_d18_57;
	wire [WIDTH-1:0] wire_d18_58;
	wire [WIDTH-1:0] wire_d18_59;
	wire [WIDTH-1:0] wire_d18_60;
	wire [WIDTH-1:0] wire_d18_61;
	wire [WIDTH-1:0] wire_d18_62;
	wire [WIDTH-1:0] wire_d18_63;
	wire [WIDTH-1:0] wire_d18_64;
	wire [WIDTH-1:0] wire_d18_65;
	wire [WIDTH-1:0] wire_d18_66;
	wire [WIDTH-1:0] wire_d18_67;
	wire [WIDTH-1:0] wire_d18_68;
	wire [WIDTH-1:0] wire_d18_69;
	wire [WIDTH-1:0] wire_d18_70;
	wire [WIDTH-1:0] wire_d18_71;
	wire [WIDTH-1:0] wire_d18_72;
	wire [WIDTH-1:0] wire_d18_73;
	wire [WIDTH-1:0] wire_d18_74;
	wire [WIDTH-1:0] wire_d18_75;
	wire [WIDTH-1:0] wire_d18_76;
	wire [WIDTH-1:0] wire_d18_77;
	wire [WIDTH-1:0] wire_d18_78;
	wire [WIDTH-1:0] wire_d18_79;
	wire [WIDTH-1:0] wire_d18_80;
	wire [WIDTH-1:0] wire_d18_81;
	wire [WIDTH-1:0] wire_d18_82;
	wire [WIDTH-1:0] wire_d18_83;
	wire [WIDTH-1:0] wire_d18_84;
	wire [WIDTH-1:0] wire_d18_85;
	wire [WIDTH-1:0] wire_d18_86;
	wire [WIDTH-1:0] wire_d18_87;
	wire [WIDTH-1:0] wire_d18_88;
	wire [WIDTH-1:0] wire_d18_89;
	wire [WIDTH-1:0] wire_d18_90;
	wire [WIDTH-1:0] wire_d18_91;
	wire [WIDTH-1:0] wire_d18_92;
	wire [WIDTH-1:0] wire_d18_93;
	wire [WIDTH-1:0] wire_d18_94;
	wire [WIDTH-1:0] wire_d18_95;
	wire [WIDTH-1:0] wire_d18_96;
	wire [WIDTH-1:0] wire_d18_97;
	wire [WIDTH-1:0] wire_d18_98;
	wire [WIDTH-1:0] wire_d18_99;
	wire [WIDTH-1:0] wire_d18_100;
	wire [WIDTH-1:0] wire_d18_101;
	wire [WIDTH-1:0] wire_d18_102;
	wire [WIDTH-1:0] wire_d18_103;
	wire [WIDTH-1:0] wire_d18_104;
	wire [WIDTH-1:0] wire_d18_105;
	wire [WIDTH-1:0] wire_d18_106;
	wire [WIDTH-1:0] wire_d18_107;
	wire [WIDTH-1:0] wire_d18_108;
	wire [WIDTH-1:0] wire_d18_109;
	wire [WIDTH-1:0] wire_d18_110;
	wire [WIDTH-1:0] wire_d18_111;
	wire [WIDTH-1:0] wire_d18_112;
	wire [WIDTH-1:0] wire_d18_113;
	wire [WIDTH-1:0] wire_d18_114;
	wire [WIDTH-1:0] wire_d18_115;
	wire [WIDTH-1:0] wire_d18_116;
	wire [WIDTH-1:0] wire_d18_117;
	wire [WIDTH-1:0] wire_d18_118;
	wire [WIDTH-1:0] wire_d19_0;
	wire [WIDTH-1:0] wire_d19_1;
	wire [WIDTH-1:0] wire_d19_2;
	wire [WIDTH-1:0] wire_d19_3;
	wire [WIDTH-1:0] wire_d19_4;
	wire [WIDTH-1:0] wire_d19_5;
	wire [WIDTH-1:0] wire_d19_6;
	wire [WIDTH-1:0] wire_d19_7;
	wire [WIDTH-1:0] wire_d19_8;
	wire [WIDTH-1:0] wire_d19_9;
	wire [WIDTH-1:0] wire_d19_10;
	wire [WIDTH-1:0] wire_d19_11;
	wire [WIDTH-1:0] wire_d19_12;
	wire [WIDTH-1:0] wire_d19_13;
	wire [WIDTH-1:0] wire_d19_14;
	wire [WIDTH-1:0] wire_d19_15;
	wire [WIDTH-1:0] wire_d19_16;
	wire [WIDTH-1:0] wire_d19_17;
	wire [WIDTH-1:0] wire_d19_18;
	wire [WIDTH-1:0] wire_d19_19;
	wire [WIDTH-1:0] wire_d19_20;
	wire [WIDTH-1:0] wire_d19_21;
	wire [WIDTH-1:0] wire_d19_22;
	wire [WIDTH-1:0] wire_d19_23;
	wire [WIDTH-1:0] wire_d19_24;
	wire [WIDTH-1:0] wire_d19_25;
	wire [WIDTH-1:0] wire_d19_26;
	wire [WIDTH-1:0] wire_d19_27;
	wire [WIDTH-1:0] wire_d19_28;
	wire [WIDTH-1:0] wire_d19_29;
	wire [WIDTH-1:0] wire_d19_30;
	wire [WIDTH-1:0] wire_d19_31;
	wire [WIDTH-1:0] wire_d19_32;
	wire [WIDTH-1:0] wire_d19_33;
	wire [WIDTH-1:0] wire_d19_34;
	wire [WIDTH-1:0] wire_d19_35;
	wire [WIDTH-1:0] wire_d19_36;
	wire [WIDTH-1:0] wire_d19_37;
	wire [WIDTH-1:0] wire_d19_38;
	wire [WIDTH-1:0] wire_d19_39;
	wire [WIDTH-1:0] wire_d19_40;
	wire [WIDTH-1:0] wire_d19_41;
	wire [WIDTH-1:0] wire_d19_42;
	wire [WIDTH-1:0] wire_d19_43;
	wire [WIDTH-1:0] wire_d19_44;
	wire [WIDTH-1:0] wire_d19_45;
	wire [WIDTH-1:0] wire_d19_46;
	wire [WIDTH-1:0] wire_d19_47;
	wire [WIDTH-1:0] wire_d19_48;
	wire [WIDTH-1:0] wire_d19_49;
	wire [WIDTH-1:0] wire_d19_50;
	wire [WIDTH-1:0] wire_d19_51;
	wire [WIDTH-1:0] wire_d19_52;
	wire [WIDTH-1:0] wire_d19_53;
	wire [WIDTH-1:0] wire_d19_54;
	wire [WIDTH-1:0] wire_d19_55;
	wire [WIDTH-1:0] wire_d19_56;
	wire [WIDTH-1:0] wire_d19_57;
	wire [WIDTH-1:0] wire_d19_58;
	wire [WIDTH-1:0] wire_d19_59;
	wire [WIDTH-1:0] wire_d19_60;
	wire [WIDTH-1:0] wire_d19_61;
	wire [WIDTH-1:0] wire_d19_62;
	wire [WIDTH-1:0] wire_d19_63;
	wire [WIDTH-1:0] wire_d19_64;
	wire [WIDTH-1:0] wire_d19_65;
	wire [WIDTH-1:0] wire_d19_66;
	wire [WIDTH-1:0] wire_d19_67;
	wire [WIDTH-1:0] wire_d19_68;
	wire [WIDTH-1:0] wire_d19_69;
	wire [WIDTH-1:0] wire_d19_70;
	wire [WIDTH-1:0] wire_d19_71;
	wire [WIDTH-1:0] wire_d19_72;
	wire [WIDTH-1:0] wire_d19_73;
	wire [WIDTH-1:0] wire_d19_74;
	wire [WIDTH-1:0] wire_d19_75;
	wire [WIDTH-1:0] wire_d19_76;
	wire [WIDTH-1:0] wire_d19_77;
	wire [WIDTH-1:0] wire_d19_78;
	wire [WIDTH-1:0] wire_d19_79;
	wire [WIDTH-1:0] wire_d19_80;
	wire [WIDTH-1:0] wire_d19_81;
	wire [WIDTH-1:0] wire_d19_82;
	wire [WIDTH-1:0] wire_d19_83;
	wire [WIDTH-1:0] wire_d19_84;
	wire [WIDTH-1:0] wire_d19_85;
	wire [WIDTH-1:0] wire_d19_86;
	wire [WIDTH-1:0] wire_d19_87;
	wire [WIDTH-1:0] wire_d19_88;
	wire [WIDTH-1:0] wire_d19_89;
	wire [WIDTH-1:0] wire_d19_90;
	wire [WIDTH-1:0] wire_d19_91;
	wire [WIDTH-1:0] wire_d19_92;
	wire [WIDTH-1:0] wire_d19_93;
	wire [WIDTH-1:0] wire_d19_94;
	wire [WIDTH-1:0] wire_d19_95;
	wire [WIDTH-1:0] wire_d19_96;
	wire [WIDTH-1:0] wire_d19_97;
	wire [WIDTH-1:0] wire_d19_98;
	wire [WIDTH-1:0] wire_d19_99;
	wire [WIDTH-1:0] wire_d19_100;
	wire [WIDTH-1:0] wire_d19_101;
	wire [WIDTH-1:0] wire_d19_102;
	wire [WIDTH-1:0] wire_d19_103;
	wire [WIDTH-1:0] wire_d19_104;
	wire [WIDTH-1:0] wire_d19_105;
	wire [WIDTH-1:0] wire_d19_106;
	wire [WIDTH-1:0] wire_d19_107;
	wire [WIDTH-1:0] wire_d19_108;
	wire [WIDTH-1:0] wire_d19_109;
	wire [WIDTH-1:0] wire_d19_110;
	wire [WIDTH-1:0] wire_d19_111;
	wire [WIDTH-1:0] wire_d19_112;
	wire [WIDTH-1:0] wire_d19_113;
	wire [WIDTH-1:0] wire_d19_114;
	wire [WIDTH-1:0] wire_d19_115;
	wire [WIDTH-1:0] wire_d19_116;
	wire [WIDTH-1:0] wire_d19_117;
	wire [WIDTH-1:0] wire_d19_118;
	wire [WIDTH-1:0] wire_d20_0;
	wire [WIDTH-1:0] wire_d20_1;
	wire [WIDTH-1:0] wire_d20_2;
	wire [WIDTH-1:0] wire_d20_3;
	wire [WIDTH-1:0] wire_d20_4;
	wire [WIDTH-1:0] wire_d20_5;
	wire [WIDTH-1:0] wire_d20_6;
	wire [WIDTH-1:0] wire_d20_7;
	wire [WIDTH-1:0] wire_d20_8;
	wire [WIDTH-1:0] wire_d20_9;
	wire [WIDTH-1:0] wire_d20_10;
	wire [WIDTH-1:0] wire_d20_11;
	wire [WIDTH-1:0] wire_d20_12;
	wire [WIDTH-1:0] wire_d20_13;
	wire [WIDTH-1:0] wire_d20_14;
	wire [WIDTH-1:0] wire_d20_15;
	wire [WIDTH-1:0] wire_d20_16;
	wire [WIDTH-1:0] wire_d20_17;
	wire [WIDTH-1:0] wire_d20_18;
	wire [WIDTH-1:0] wire_d20_19;
	wire [WIDTH-1:0] wire_d20_20;
	wire [WIDTH-1:0] wire_d20_21;
	wire [WIDTH-1:0] wire_d20_22;
	wire [WIDTH-1:0] wire_d20_23;
	wire [WIDTH-1:0] wire_d20_24;
	wire [WIDTH-1:0] wire_d20_25;
	wire [WIDTH-1:0] wire_d20_26;
	wire [WIDTH-1:0] wire_d20_27;
	wire [WIDTH-1:0] wire_d20_28;
	wire [WIDTH-1:0] wire_d20_29;
	wire [WIDTH-1:0] wire_d20_30;
	wire [WIDTH-1:0] wire_d20_31;
	wire [WIDTH-1:0] wire_d20_32;
	wire [WIDTH-1:0] wire_d20_33;
	wire [WIDTH-1:0] wire_d20_34;
	wire [WIDTH-1:0] wire_d20_35;
	wire [WIDTH-1:0] wire_d20_36;
	wire [WIDTH-1:0] wire_d20_37;
	wire [WIDTH-1:0] wire_d20_38;
	wire [WIDTH-1:0] wire_d20_39;
	wire [WIDTH-1:0] wire_d20_40;
	wire [WIDTH-1:0] wire_d20_41;
	wire [WIDTH-1:0] wire_d20_42;
	wire [WIDTH-1:0] wire_d20_43;
	wire [WIDTH-1:0] wire_d20_44;
	wire [WIDTH-1:0] wire_d20_45;
	wire [WIDTH-1:0] wire_d20_46;
	wire [WIDTH-1:0] wire_d20_47;
	wire [WIDTH-1:0] wire_d20_48;
	wire [WIDTH-1:0] wire_d20_49;
	wire [WIDTH-1:0] wire_d20_50;
	wire [WIDTH-1:0] wire_d20_51;
	wire [WIDTH-1:0] wire_d20_52;
	wire [WIDTH-1:0] wire_d20_53;
	wire [WIDTH-1:0] wire_d20_54;
	wire [WIDTH-1:0] wire_d20_55;
	wire [WIDTH-1:0] wire_d20_56;
	wire [WIDTH-1:0] wire_d20_57;
	wire [WIDTH-1:0] wire_d20_58;
	wire [WIDTH-1:0] wire_d20_59;
	wire [WIDTH-1:0] wire_d20_60;
	wire [WIDTH-1:0] wire_d20_61;
	wire [WIDTH-1:0] wire_d20_62;
	wire [WIDTH-1:0] wire_d20_63;
	wire [WIDTH-1:0] wire_d20_64;
	wire [WIDTH-1:0] wire_d20_65;
	wire [WIDTH-1:0] wire_d20_66;
	wire [WIDTH-1:0] wire_d20_67;
	wire [WIDTH-1:0] wire_d20_68;
	wire [WIDTH-1:0] wire_d20_69;
	wire [WIDTH-1:0] wire_d20_70;
	wire [WIDTH-1:0] wire_d20_71;
	wire [WIDTH-1:0] wire_d20_72;
	wire [WIDTH-1:0] wire_d20_73;
	wire [WIDTH-1:0] wire_d20_74;
	wire [WIDTH-1:0] wire_d20_75;
	wire [WIDTH-1:0] wire_d20_76;
	wire [WIDTH-1:0] wire_d20_77;
	wire [WIDTH-1:0] wire_d20_78;
	wire [WIDTH-1:0] wire_d20_79;
	wire [WIDTH-1:0] wire_d20_80;
	wire [WIDTH-1:0] wire_d20_81;
	wire [WIDTH-1:0] wire_d20_82;
	wire [WIDTH-1:0] wire_d20_83;
	wire [WIDTH-1:0] wire_d20_84;
	wire [WIDTH-1:0] wire_d20_85;
	wire [WIDTH-1:0] wire_d20_86;
	wire [WIDTH-1:0] wire_d20_87;
	wire [WIDTH-1:0] wire_d20_88;
	wire [WIDTH-1:0] wire_d20_89;
	wire [WIDTH-1:0] wire_d20_90;
	wire [WIDTH-1:0] wire_d20_91;
	wire [WIDTH-1:0] wire_d20_92;
	wire [WIDTH-1:0] wire_d20_93;
	wire [WIDTH-1:0] wire_d20_94;
	wire [WIDTH-1:0] wire_d20_95;
	wire [WIDTH-1:0] wire_d20_96;
	wire [WIDTH-1:0] wire_d20_97;
	wire [WIDTH-1:0] wire_d20_98;
	wire [WIDTH-1:0] wire_d20_99;
	wire [WIDTH-1:0] wire_d20_100;
	wire [WIDTH-1:0] wire_d20_101;
	wire [WIDTH-1:0] wire_d20_102;
	wire [WIDTH-1:0] wire_d20_103;
	wire [WIDTH-1:0] wire_d20_104;
	wire [WIDTH-1:0] wire_d20_105;
	wire [WIDTH-1:0] wire_d20_106;
	wire [WIDTH-1:0] wire_d20_107;
	wire [WIDTH-1:0] wire_d20_108;
	wire [WIDTH-1:0] wire_d20_109;
	wire [WIDTH-1:0] wire_d20_110;
	wire [WIDTH-1:0] wire_d20_111;
	wire [WIDTH-1:0] wire_d20_112;
	wire [WIDTH-1:0] wire_d20_113;
	wire [WIDTH-1:0] wire_d20_114;
	wire [WIDTH-1:0] wire_d20_115;
	wire [WIDTH-1:0] wire_d20_116;
	wire [WIDTH-1:0] wire_d20_117;
	wire [WIDTH-1:0] wire_d20_118;
	wire [WIDTH-1:0] wire_d21_0;
	wire [WIDTH-1:0] wire_d21_1;
	wire [WIDTH-1:0] wire_d21_2;
	wire [WIDTH-1:0] wire_d21_3;
	wire [WIDTH-1:0] wire_d21_4;
	wire [WIDTH-1:0] wire_d21_5;
	wire [WIDTH-1:0] wire_d21_6;
	wire [WIDTH-1:0] wire_d21_7;
	wire [WIDTH-1:0] wire_d21_8;
	wire [WIDTH-1:0] wire_d21_9;
	wire [WIDTH-1:0] wire_d21_10;
	wire [WIDTH-1:0] wire_d21_11;
	wire [WIDTH-1:0] wire_d21_12;
	wire [WIDTH-1:0] wire_d21_13;
	wire [WIDTH-1:0] wire_d21_14;
	wire [WIDTH-1:0] wire_d21_15;
	wire [WIDTH-1:0] wire_d21_16;
	wire [WIDTH-1:0] wire_d21_17;
	wire [WIDTH-1:0] wire_d21_18;
	wire [WIDTH-1:0] wire_d21_19;
	wire [WIDTH-1:0] wire_d21_20;
	wire [WIDTH-1:0] wire_d21_21;
	wire [WIDTH-1:0] wire_d21_22;
	wire [WIDTH-1:0] wire_d21_23;
	wire [WIDTH-1:0] wire_d21_24;
	wire [WIDTH-1:0] wire_d21_25;
	wire [WIDTH-1:0] wire_d21_26;
	wire [WIDTH-1:0] wire_d21_27;
	wire [WIDTH-1:0] wire_d21_28;
	wire [WIDTH-1:0] wire_d21_29;
	wire [WIDTH-1:0] wire_d21_30;
	wire [WIDTH-1:0] wire_d21_31;
	wire [WIDTH-1:0] wire_d21_32;
	wire [WIDTH-1:0] wire_d21_33;
	wire [WIDTH-1:0] wire_d21_34;
	wire [WIDTH-1:0] wire_d21_35;
	wire [WIDTH-1:0] wire_d21_36;
	wire [WIDTH-1:0] wire_d21_37;
	wire [WIDTH-1:0] wire_d21_38;
	wire [WIDTH-1:0] wire_d21_39;
	wire [WIDTH-1:0] wire_d21_40;
	wire [WIDTH-1:0] wire_d21_41;
	wire [WIDTH-1:0] wire_d21_42;
	wire [WIDTH-1:0] wire_d21_43;
	wire [WIDTH-1:0] wire_d21_44;
	wire [WIDTH-1:0] wire_d21_45;
	wire [WIDTH-1:0] wire_d21_46;
	wire [WIDTH-1:0] wire_d21_47;
	wire [WIDTH-1:0] wire_d21_48;
	wire [WIDTH-1:0] wire_d21_49;
	wire [WIDTH-1:0] wire_d21_50;
	wire [WIDTH-1:0] wire_d21_51;
	wire [WIDTH-1:0] wire_d21_52;
	wire [WIDTH-1:0] wire_d21_53;
	wire [WIDTH-1:0] wire_d21_54;
	wire [WIDTH-1:0] wire_d21_55;
	wire [WIDTH-1:0] wire_d21_56;
	wire [WIDTH-1:0] wire_d21_57;
	wire [WIDTH-1:0] wire_d21_58;
	wire [WIDTH-1:0] wire_d21_59;
	wire [WIDTH-1:0] wire_d21_60;
	wire [WIDTH-1:0] wire_d21_61;
	wire [WIDTH-1:0] wire_d21_62;
	wire [WIDTH-1:0] wire_d21_63;
	wire [WIDTH-1:0] wire_d21_64;
	wire [WIDTH-1:0] wire_d21_65;
	wire [WIDTH-1:0] wire_d21_66;
	wire [WIDTH-1:0] wire_d21_67;
	wire [WIDTH-1:0] wire_d21_68;
	wire [WIDTH-1:0] wire_d21_69;
	wire [WIDTH-1:0] wire_d21_70;
	wire [WIDTH-1:0] wire_d21_71;
	wire [WIDTH-1:0] wire_d21_72;
	wire [WIDTH-1:0] wire_d21_73;
	wire [WIDTH-1:0] wire_d21_74;
	wire [WIDTH-1:0] wire_d21_75;
	wire [WIDTH-1:0] wire_d21_76;
	wire [WIDTH-1:0] wire_d21_77;
	wire [WIDTH-1:0] wire_d21_78;
	wire [WIDTH-1:0] wire_d21_79;
	wire [WIDTH-1:0] wire_d21_80;
	wire [WIDTH-1:0] wire_d21_81;
	wire [WIDTH-1:0] wire_d21_82;
	wire [WIDTH-1:0] wire_d21_83;
	wire [WIDTH-1:0] wire_d21_84;
	wire [WIDTH-1:0] wire_d21_85;
	wire [WIDTH-1:0] wire_d21_86;
	wire [WIDTH-1:0] wire_d21_87;
	wire [WIDTH-1:0] wire_d21_88;
	wire [WIDTH-1:0] wire_d21_89;
	wire [WIDTH-1:0] wire_d21_90;
	wire [WIDTH-1:0] wire_d21_91;
	wire [WIDTH-1:0] wire_d21_92;
	wire [WIDTH-1:0] wire_d21_93;
	wire [WIDTH-1:0] wire_d21_94;
	wire [WIDTH-1:0] wire_d21_95;
	wire [WIDTH-1:0] wire_d21_96;
	wire [WIDTH-1:0] wire_d21_97;
	wire [WIDTH-1:0] wire_d21_98;
	wire [WIDTH-1:0] wire_d21_99;
	wire [WIDTH-1:0] wire_d21_100;
	wire [WIDTH-1:0] wire_d21_101;
	wire [WIDTH-1:0] wire_d21_102;
	wire [WIDTH-1:0] wire_d21_103;
	wire [WIDTH-1:0] wire_d21_104;
	wire [WIDTH-1:0] wire_d21_105;
	wire [WIDTH-1:0] wire_d21_106;
	wire [WIDTH-1:0] wire_d21_107;
	wire [WIDTH-1:0] wire_d21_108;
	wire [WIDTH-1:0] wire_d21_109;
	wire [WIDTH-1:0] wire_d21_110;
	wire [WIDTH-1:0] wire_d21_111;
	wire [WIDTH-1:0] wire_d21_112;
	wire [WIDTH-1:0] wire_d21_113;
	wire [WIDTH-1:0] wire_d21_114;
	wire [WIDTH-1:0] wire_d21_115;
	wire [WIDTH-1:0] wire_d21_116;
	wire [WIDTH-1:0] wire_d21_117;
	wire [WIDTH-1:0] wire_d21_118;
	wire [WIDTH-1:0] wire_d22_0;
	wire [WIDTH-1:0] wire_d22_1;
	wire [WIDTH-1:0] wire_d22_2;
	wire [WIDTH-1:0] wire_d22_3;
	wire [WIDTH-1:0] wire_d22_4;
	wire [WIDTH-1:0] wire_d22_5;
	wire [WIDTH-1:0] wire_d22_6;
	wire [WIDTH-1:0] wire_d22_7;
	wire [WIDTH-1:0] wire_d22_8;
	wire [WIDTH-1:0] wire_d22_9;
	wire [WIDTH-1:0] wire_d22_10;
	wire [WIDTH-1:0] wire_d22_11;
	wire [WIDTH-1:0] wire_d22_12;
	wire [WIDTH-1:0] wire_d22_13;
	wire [WIDTH-1:0] wire_d22_14;
	wire [WIDTH-1:0] wire_d22_15;
	wire [WIDTH-1:0] wire_d22_16;
	wire [WIDTH-1:0] wire_d22_17;
	wire [WIDTH-1:0] wire_d22_18;
	wire [WIDTH-1:0] wire_d22_19;
	wire [WIDTH-1:0] wire_d22_20;
	wire [WIDTH-1:0] wire_d22_21;
	wire [WIDTH-1:0] wire_d22_22;
	wire [WIDTH-1:0] wire_d22_23;
	wire [WIDTH-1:0] wire_d22_24;
	wire [WIDTH-1:0] wire_d22_25;
	wire [WIDTH-1:0] wire_d22_26;
	wire [WIDTH-1:0] wire_d22_27;
	wire [WIDTH-1:0] wire_d22_28;
	wire [WIDTH-1:0] wire_d22_29;
	wire [WIDTH-1:0] wire_d22_30;
	wire [WIDTH-1:0] wire_d22_31;
	wire [WIDTH-1:0] wire_d22_32;
	wire [WIDTH-1:0] wire_d22_33;
	wire [WIDTH-1:0] wire_d22_34;
	wire [WIDTH-1:0] wire_d22_35;
	wire [WIDTH-1:0] wire_d22_36;
	wire [WIDTH-1:0] wire_d22_37;
	wire [WIDTH-1:0] wire_d22_38;
	wire [WIDTH-1:0] wire_d22_39;
	wire [WIDTH-1:0] wire_d22_40;
	wire [WIDTH-1:0] wire_d22_41;
	wire [WIDTH-1:0] wire_d22_42;
	wire [WIDTH-1:0] wire_d22_43;
	wire [WIDTH-1:0] wire_d22_44;
	wire [WIDTH-1:0] wire_d22_45;
	wire [WIDTH-1:0] wire_d22_46;
	wire [WIDTH-1:0] wire_d22_47;
	wire [WIDTH-1:0] wire_d22_48;
	wire [WIDTH-1:0] wire_d22_49;
	wire [WIDTH-1:0] wire_d22_50;
	wire [WIDTH-1:0] wire_d22_51;
	wire [WIDTH-1:0] wire_d22_52;
	wire [WIDTH-1:0] wire_d22_53;
	wire [WIDTH-1:0] wire_d22_54;
	wire [WIDTH-1:0] wire_d22_55;
	wire [WIDTH-1:0] wire_d22_56;
	wire [WIDTH-1:0] wire_d22_57;
	wire [WIDTH-1:0] wire_d22_58;
	wire [WIDTH-1:0] wire_d22_59;
	wire [WIDTH-1:0] wire_d22_60;
	wire [WIDTH-1:0] wire_d22_61;
	wire [WIDTH-1:0] wire_d22_62;
	wire [WIDTH-1:0] wire_d22_63;
	wire [WIDTH-1:0] wire_d22_64;
	wire [WIDTH-1:0] wire_d22_65;
	wire [WIDTH-1:0] wire_d22_66;
	wire [WIDTH-1:0] wire_d22_67;
	wire [WIDTH-1:0] wire_d22_68;
	wire [WIDTH-1:0] wire_d22_69;
	wire [WIDTH-1:0] wire_d22_70;
	wire [WIDTH-1:0] wire_d22_71;
	wire [WIDTH-1:0] wire_d22_72;
	wire [WIDTH-1:0] wire_d22_73;
	wire [WIDTH-1:0] wire_d22_74;
	wire [WIDTH-1:0] wire_d22_75;
	wire [WIDTH-1:0] wire_d22_76;
	wire [WIDTH-1:0] wire_d22_77;
	wire [WIDTH-1:0] wire_d22_78;
	wire [WIDTH-1:0] wire_d22_79;
	wire [WIDTH-1:0] wire_d22_80;
	wire [WIDTH-1:0] wire_d22_81;
	wire [WIDTH-1:0] wire_d22_82;
	wire [WIDTH-1:0] wire_d22_83;
	wire [WIDTH-1:0] wire_d22_84;
	wire [WIDTH-1:0] wire_d22_85;
	wire [WIDTH-1:0] wire_d22_86;
	wire [WIDTH-1:0] wire_d22_87;
	wire [WIDTH-1:0] wire_d22_88;
	wire [WIDTH-1:0] wire_d22_89;
	wire [WIDTH-1:0] wire_d22_90;
	wire [WIDTH-1:0] wire_d22_91;
	wire [WIDTH-1:0] wire_d22_92;
	wire [WIDTH-1:0] wire_d22_93;
	wire [WIDTH-1:0] wire_d22_94;
	wire [WIDTH-1:0] wire_d22_95;
	wire [WIDTH-1:0] wire_d22_96;
	wire [WIDTH-1:0] wire_d22_97;
	wire [WIDTH-1:0] wire_d22_98;
	wire [WIDTH-1:0] wire_d22_99;
	wire [WIDTH-1:0] wire_d22_100;
	wire [WIDTH-1:0] wire_d22_101;
	wire [WIDTH-1:0] wire_d22_102;
	wire [WIDTH-1:0] wire_d22_103;
	wire [WIDTH-1:0] wire_d22_104;
	wire [WIDTH-1:0] wire_d22_105;
	wire [WIDTH-1:0] wire_d22_106;
	wire [WIDTH-1:0] wire_d22_107;
	wire [WIDTH-1:0] wire_d22_108;
	wire [WIDTH-1:0] wire_d22_109;
	wire [WIDTH-1:0] wire_d22_110;
	wire [WIDTH-1:0] wire_d22_111;
	wire [WIDTH-1:0] wire_d22_112;
	wire [WIDTH-1:0] wire_d22_113;
	wire [WIDTH-1:0] wire_d22_114;
	wire [WIDTH-1:0] wire_d22_115;
	wire [WIDTH-1:0] wire_d22_116;
	wire [WIDTH-1:0] wire_d22_117;
	wire [WIDTH-1:0] wire_d22_118;
	wire [WIDTH-1:0] wire_d23_0;
	wire [WIDTH-1:0] wire_d23_1;
	wire [WIDTH-1:0] wire_d23_2;
	wire [WIDTH-1:0] wire_d23_3;
	wire [WIDTH-1:0] wire_d23_4;
	wire [WIDTH-1:0] wire_d23_5;
	wire [WIDTH-1:0] wire_d23_6;
	wire [WIDTH-1:0] wire_d23_7;
	wire [WIDTH-1:0] wire_d23_8;
	wire [WIDTH-1:0] wire_d23_9;
	wire [WIDTH-1:0] wire_d23_10;
	wire [WIDTH-1:0] wire_d23_11;
	wire [WIDTH-1:0] wire_d23_12;
	wire [WIDTH-1:0] wire_d23_13;
	wire [WIDTH-1:0] wire_d23_14;
	wire [WIDTH-1:0] wire_d23_15;
	wire [WIDTH-1:0] wire_d23_16;
	wire [WIDTH-1:0] wire_d23_17;
	wire [WIDTH-1:0] wire_d23_18;
	wire [WIDTH-1:0] wire_d23_19;
	wire [WIDTH-1:0] wire_d23_20;
	wire [WIDTH-1:0] wire_d23_21;
	wire [WIDTH-1:0] wire_d23_22;
	wire [WIDTH-1:0] wire_d23_23;
	wire [WIDTH-1:0] wire_d23_24;
	wire [WIDTH-1:0] wire_d23_25;
	wire [WIDTH-1:0] wire_d23_26;
	wire [WIDTH-1:0] wire_d23_27;
	wire [WIDTH-1:0] wire_d23_28;
	wire [WIDTH-1:0] wire_d23_29;
	wire [WIDTH-1:0] wire_d23_30;
	wire [WIDTH-1:0] wire_d23_31;
	wire [WIDTH-1:0] wire_d23_32;
	wire [WIDTH-1:0] wire_d23_33;
	wire [WIDTH-1:0] wire_d23_34;
	wire [WIDTH-1:0] wire_d23_35;
	wire [WIDTH-1:0] wire_d23_36;
	wire [WIDTH-1:0] wire_d23_37;
	wire [WIDTH-1:0] wire_d23_38;
	wire [WIDTH-1:0] wire_d23_39;
	wire [WIDTH-1:0] wire_d23_40;
	wire [WIDTH-1:0] wire_d23_41;
	wire [WIDTH-1:0] wire_d23_42;
	wire [WIDTH-1:0] wire_d23_43;
	wire [WIDTH-1:0] wire_d23_44;
	wire [WIDTH-1:0] wire_d23_45;
	wire [WIDTH-1:0] wire_d23_46;
	wire [WIDTH-1:0] wire_d23_47;
	wire [WIDTH-1:0] wire_d23_48;
	wire [WIDTH-1:0] wire_d23_49;
	wire [WIDTH-1:0] wire_d23_50;
	wire [WIDTH-1:0] wire_d23_51;
	wire [WIDTH-1:0] wire_d23_52;
	wire [WIDTH-1:0] wire_d23_53;
	wire [WIDTH-1:0] wire_d23_54;
	wire [WIDTH-1:0] wire_d23_55;
	wire [WIDTH-1:0] wire_d23_56;
	wire [WIDTH-1:0] wire_d23_57;
	wire [WIDTH-1:0] wire_d23_58;
	wire [WIDTH-1:0] wire_d23_59;
	wire [WIDTH-1:0] wire_d23_60;
	wire [WIDTH-1:0] wire_d23_61;
	wire [WIDTH-1:0] wire_d23_62;
	wire [WIDTH-1:0] wire_d23_63;
	wire [WIDTH-1:0] wire_d23_64;
	wire [WIDTH-1:0] wire_d23_65;
	wire [WIDTH-1:0] wire_d23_66;
	wire [WIDTH-1:0] wire_d23_67;
	wire [WIDTH-1:0] wire_d23_68;
	wire [WIDTH-1:0] wire_d23_69;
	wire [WIDTH-1:0] wire_d23_70;
	wire [WIDTH-1:0] wire_d23_71;
	wire [WIDTH-1:0] wire_d23_72;
	wire [WIDTH-1:0] wire_d23_73;
	wire [WIDTH-1:0] wire_d23_74;
	wire [WIDTH-1:0] wire_d23_75;
	wire [WIDTH-1:0] wire_d23_76;
	wire [WIDTH-1:0] wire_d23_77;
	wire [WIDTH-1:0] wire_d23_78;
	wire [WIDTH-1:0] wire_d23_79;
	wire [WIDTH-1:0] wire_d23_80;
	wire [WIDTH-1:0] wire_d23_81;
	wire [WIDTH-1:0] wire_d23_82;
	wire [WIDTH-1:0] wire_d23_83;
	wire [WIDTH-1:0] wire_d23_84;
	wire [WIDTH-1:0] wire_d23_85;
	wire [WIDTH-1:0] wire_d23_86;
	wire [WIDTH-1:0] wire_d23_87;
	wire [WIDTH-1:0] wire_d23_88;
	wire [WIDTH-1:0] wire_d23_89;
	wire [WIDTH-1:0] wire_d23_90;
	wire [WIDTH-1:0] wire_d23_91;
	wire [WIDTH-1:0] wire_d23_92;
	wire [WIDTH-1:0] wire_d23_93;
	wire [WIDTH-1:0] wire_d23_94;
	wire [WIDTH-1:0] wire_d23_95;
	wire [WIDTH-1:0] wire_d23_96;
	wire [WIDTH-1:0] wire_d23_97;
	wire [WIDTH-1:0] wire_d23_98;
	wire [WIDTH-1:0] wire_d23_99;
	wire [WIDTH-1:0] wire_d23_100;
	wire [WIDTH-1:0] wire_d23_101;
	wire [WIDTH-1:0] wire_d23_102;
	wire [WIDTH-1:0] wire_d23_103;
	wire [WIDTH-1:0] wire_d23_104;
	wire [WIDTH-1:0] wire_d23_105;
	wire [WIDTH-1:0] wire_d23_106;
	wire [WIDTH-1:0] wire_d23_107;
	wire [WIDTH-1:0] wire_d23_108;
	wire [WIDTH-1:0] wire_d23_109;
	wire [WIDTH-1:0] wire_d23_110;
	wire [WIDTH-1:0] wire_d23_111;
	wire [WIDTH-1:0] wire_d23_112;
	wire [WIDTH-1:0] wire_d23_113;
	wire [WIDTH-1:0] wire_d23_114;
	wire [WIDTH-1:0] wire_d23_115;
	wire [WIDTH-1:0] wire_d23_116;
	wire [WIDTH-1:0] wire_d23_117;
	wire [WIDTH-1:0] wire_d23_118;
	wire [WIDTH-1:0] wire_d24_0;
	wire [WIDTH-1:0] wire_d24_1;
	wire [WIDTH-1:0] wire_d24_2;
	wire [WIDTH-1:0] wire_d24_3;
	wire [WIDTH-1:0] wire_d24_4;
	wire [WIDTH-1:0] wire_d24_5;
	wire [WIDTH-1:0] wire_d24_6;
	wire [WIDTH-1:0] wire_d24_7;
	wire [WIDTH-1:0] wire_d24_8;
	wire [WIDTH-1:0] wire_d24_9;
	wire [WIDTH-1:0] wire_d24_10;
	wire [WIDTH-1:0] wire_d24_11;
	wire [WIDTH-1:0] wire_d24_12;
	wire [WIDTH-1:0] wire_d24_13;
	wire [WIDTH-1:0] wire_d24_14;
	wire [WIDTH-1:0] wire_d24_15;
	wire [WIDTH-1:0] wire_d24_16;
	wire [WIDTH-1:0] wire_d24_17;
	wire [WIDTH-1:0] wire_d24_18;
	wire [WIDTH-1:0] wire_d24_19;
	wire [WIDTH-1:0] wire_d24_20;
	wire [WIDTH-1:0] wire_d24_21;
	wire [WIDTH-1:0] wire_d24_22;
	wire [WIDTH-1:0] wire_d24_23;
	wire [WIDTH-1:0] wire_d24_24;
	wire [WIDTH-1:0] wire_d24_25;
	wire [WIDTH-1:0] wire_d24_26;
	wire [WIDTH-1:0] wire_d24_27;
	wire [WIDTH-1:0] wire_d24_28;
	wire [WIDTH-1:0] wire_d24_29;
	wire [WIDTH-1:0] wire_d24_30;
	wire [WIDTH-1:0] wire_d24_31;
	wire [WIDTH-1:0] wire_d24_32;
	wire [WIDTH-1:0] wire_d24_33;
	wire [WIDTH-1:0] wire_d24_34;
	wire [WIDTH-1:0] wire_d24_35;
	wire [WIDTH-1:0] wire_d24_36;
	wire [WIDTH-1:0] wire_d24_37;
	wire [WIDTH-1:0] wire_d24_38;
	wire [WIDTH-1:0] wire_d24_39;
	wire [WIDTH-1:0] wire_d24_40;
	wire [WIDTH-1:0] wire_d24_41;
	wire [WIDTH-1:0] wire_d24_42;
	wire [WIDTH-1:0] wire_d24_43;
	wire [WIDTH-1:0] wire_d24_44;
	wire [WIDTH-1:0] wire_d24_45;
	wire [WIDTH-1:0] wire_d24_46;
	wire [WIDTH-1:0] wire_d24_47;
	wire [WIDTH-1:0] wire_d24_48;
	wire [WIDTH-1:0] wire_d24_49;
	wire [WIDTH-1:0] wire_d24_50;
	wire [WIDTH-1:0] wire_d24_51;
	wire [WIDTH-1:0] wire_d24_52;
	wire [WIDTH-1:0] wire_d24_53;
	wire [WIDTH-1:0] wire_d24_54;
	wire [WIDTH-1:0] wire_d24_55;
	wire [WIDTH-1:0] wire_d24_56;
	wire [WIDTH-1:0] wire_d24_57;
	wire [WIDTH-1:0] wire_d24_58;
	wire [WIDTH-1:0] wire_d24_59;
	wire [WIDTH-1:0] wire_d24_60;
	wire [WIDTH-1:0] wire_d24_61;
	wire [WIDTH-1:0] wire_d24_62;
	wire [WIDTH-1:0] wire_d24_63;
	wire [WIDTH-1:0] wire_d24_64;
	wire [WIDTH-1:0] wire_d24_65;
	wire [WIDTH-1:0] wire_d24_66;
	wire [WIDTH-1:0] wire_d24_67;
	wire [WIDTH-1:0] wire_d24_68;
	wire [WIDTH-1:0] wire_d24_69;
	wire [WIDTH-1:0] wire_d24_70;
	wire [WIDTH-1:0] wire_d24_71;
	wire [WIDTH-1:0] wire_d24_72;
	wire [WIDTH-1:0] wire_d24_73;
	wire [WIDTH-1:0] wire_d24_74;
	wire [WIDTH-1:0] wire_d24_75;
	wire [WIDTH-1:0] wire_d24_76;
	wire [WIDTH-1:0] wire_d24_77;
	wire [WIDTH-1:0] wire_d24_78;
	wire [WIDTH-1:0] wire_d24_79;
	wire [WIDTH-1:0] wire_d24_80;
	wire [WIDTH-1:0] wire_d24_81;
	wire [WIDTH-1:0] wire_d24_82;
	wire [WIDTH-1:0] wire_d24_83;
	wire [WIDTH-1:0] wire_d24_84;
	wire [WIDTH-1:0] wire_d24_85;
	wire [WIDTH-1:0] wire_d24_86;
	wire [WIDTH-1:0] wire_d24_87;
	wire [WIDTH-1:0] wire_d24_88;
	wire [WIDTH-1:0] wire_d24_89;
	wire [WIDTH-1:0] wire_d24_90;
	wire [WIDTH-1:0] wire_d24_91;
	wire [WIDTH-1:0] wire_d24_92;
	wire [WIDTH-1:0] wire_d24_93;
	wire [WIDTH-1:0] wire_d24_94;
	wire [WIDTH-1:0] wire_d24_95;
	wire [WIDTH-1:0] wire_d24_96;
	wire [WIDTH-1:0] wire_d24_97;
	wire [WIDTH-1:0] wire_d24_98;
	wire [WIDTH-1:0] wire_d24_99;
	wire [WIDTH-1:0] wire_d24_100;
	wire [WIDTH-1:0] wire_d24_101;
	wire [WIDTH-1:0] wire_d24_102;
	wire [WIDTH-1:0] wire_d24_103;
	wire [WIDTH-1:0] wire_d24_104;
	wire [WIDTH-1:0] wire_d24_105;
	wire [WIDTH-1:0] wire_d24_106;
	wire [WIDTH-1:0] wire_d24_107;
	wire [WIDTH-1:0] wire_d24_108;
	wire [WIDTH-1:0] wire_d24_109;
	wire [WIDTH-1:0] wire_d24_110;
	wire [WIDTH-1:0] wire_d24_111;
	wire [WIDTH-1:0] wire_d24_112;
	wire [WIDTH-1:0] wire_d24_113;
	wire [WIDTH-1:0] wire_d24_114;
	wire [WIDTH-1:0] wire_d24_115;
	wire [WIDTH-1:0] wire_d24_116;
	wire [WIDTH-1:0] wire_d24_117;
	wire [WIDTH-1:0] wire_d24_118;
	wire [WIDTH-1:0] wire_d25_0;
	wire [WIDTH-1:0] wire_d25_1;
	wire [WIDTH-1:0] wire_d25_2;
	wire [WIDTH-1:0] wire_d25_3;
	wire [WIDTH-1:0] wire_d25_4;
	wire [WIDTH-1:0] wire_d25_5;
	wire [WIDTH-1:0] wire_d25_6;
	wire [WIDTH-1:0] wire_d25_7;
	wire [WIDTH-1:0] wire_d25_8;
	wire [WIDTH-1:0] wire_d25_9;
	wire [WIDTH-1:0] wire_d25_10;
	wire [WIDTH-1:0] wire_d25_11;
	wire [WIDTH-1:0] wire_d25_12;
	wire [WIDTH-1:0] wire_d25_13;
	wire [WIDTH-1:0] wire_d25_14;
	wire [WIDTH-1:0] wire_d25_15;
	wire [WIDTH-1:0] wire_d25_16;
	wire [WIDTH-1:0] wire_d25_17;
	wire [WIDTH-1:0] wire_d25_18;
	wire [WIDTH-1:0] wire_d25_19;
	wire [WIDTH-1:0] wire_d25_20;
	wire [WIDTH-1:0] wire_d25_21;
	wire [WIDTH-1:0] wire_d25_22;
	wire [WIDTH-1:0] wire_d25_23;
	wire [WIDTH-1:0] wire_d25_24;
	wire [WIDTH-1:0] wire_d25_25;
	wire [WIDTH-1:0] wire_d25_26;
	wire [WIDTH-1:0] wire_d25_27;
	wire [WIDTH-1:0] wire_d25_28;
	wire [WIDTH-1:0] wire_d25_29;
	wire [WIDTH-1:0] wire_d25_30;
	wire [WIDTH-1:0] wire_d25_31;
	wire [WIDTH-1:0] wire_d25_32;
	wire [WIDTH-1:0] wire_d25_33;
	wire [WIDTH-1:0] wire_d25_34;
	wire [WIDTH-1:0] wire_d25_35;
	wire [WIDTH-1:0] wire_d25_36;
	wire [WIDTH-1:0] wire_d25_37;
	wire [WIDTH-1:0] wire_d25_38;
	wire [WIDTH-1:0] wire_d25_39;
	wire [WIDTH-1:0] wire_d25_40;
	wire [WIDTH-1:0] wire_d25_41;
	wire [WIDTH-1:0] wire_d25_42;
	wire [WIDTH-1:0] wire_d25_43;
	wire [WIDTH-1:0] wire_d25_44;
	wire [WIDTH-1:0] wire_d25_45;
	wire [WIDTH-1:0] wire_d25_46;
	wire [WIDTH-1:0] wire_d25_47;
	wire [WIDTH-1:0] wire_d25_48;
	wire [WIDTH-1:0] wire_d25_49;
	wire [WIDTH-1:0] wire_d25_50;
	wire [WIDTH-1:0] wire_d25_51;
	wire [WIDTH-1:0] wire_d25_52;
	wire [WIDTH-1:0] wire_d25_53;
	wire [WIDTH-1:0] wire_d25_54;
	wire [WIDTH-1:0] wire_d25_55;
	wire [WIDTH-1:0] wire_d25_56;
	wire [WIDTH-1:0] wire_d25_57;
	wire [WIDTH-1:0] wire_d25_58;
	wire [WIDTH-1:0] wire_d25_59;
	wire [WIDTH-1:0] wire_d25_60;
	wire [WIDTH-1:0] wire_d25_61;
	wire [WIDTH-1:0] wire_d25_62;
	wire [WIDTH-1:0] wire_d25_63;
	wire [WIDTH-1:0] wire_d25_64;
	wire [WIDTH-1:0] wire_d25_65;
	wire [WIDTH-1:0] wire_d25_66;
	wire [WIDTH-1:0] wire_d25_67;
	wire [WIDTH-1:0] wire_d25_68;
	wire [WIDTH-1:0] wire_d25_69;
	wire [WIDTH-1:0] wire_d25_70;
	wire [WIDTH-1:0] wire_d25_71;
	wire [WIDTH-1:0] wire_d25_72;
	wire [WIDTH-1:0] wire_d25_73;
	wire [WIDTH-1:0] wire_d25_74;
	wire [WIDTH-1:0] wire_d25_75;
	wire [WIDTH-1:0] wire_d25_76;
	wire [WIDTH-1:0] wire_d25_77;
	wire [WIDTH-1:0] wire_d25_78;
	wire [WIDTH-1:0] wire_d25_79;
	wire [WIDTH-1:0] wire_d25_80;
	wire [WIDTH-1:0] wire_d25_81;
	wire [WIDTH-1:0] wire_d25_82;
	wire [WIDTH-1:0] wire_d25_83;
	wire [WIDTH-1:0] wire_d25_84;
	wire [WIDTH-1:0] wire_d25_85;
	wire [WIDTH-1:0] wire_d25_86;
	wire [WIDTH-1:0] wire_d25_87;
	wire [WIDTH-1:0] wire_d25_88;
	wire [WIDTH-1:0] wire_d25_89;
	wire [WIDTH-1:0] wire_d25_90;
	wire [WIDTH-1:0] wire_d25_91;
	wire [WIDTH-1:0] wire_d25_92;
	wire [WIDTH-1:0] wire_d25_93;
	wire [WIDTH-1:0] wire_d25_94;
	wire [WIDTH-1:0] wire_d25_95;
	wire [WIDTH-1:0] wire_d25_96;
	wire [WIDTH-1:0] wire_d25_97;
	wire [WIDTH-1:0] wire_d25_98;
	wire [WIDTH-1:0] wire_d25_99;
	wire [WIDTH-1:0] wire_d25_100;
	wire [WIDTH-1:0] wire_d25_101;
	wire [WIDTH-1:0] wire_d25_102;
	wire [WIDTH-1:0] wire_d25_103;
	wire [WIDTH-1:0] wire_d25_104;
	wire [WIDTH-1:0] wire_d25_105;
	wire [WIDTH-1:0] wire_d25_106;
	wire [WIDTH-1:0] wire_d25_107;
	wire [WIDTH-1:0] wire_d25_108;
	wire [WIDTH-1:0] wire_d25_109;
	wire [WIDTH-1:0] wire_d25_110;
	wire [WIDTH-1:0] wire_d25_111;
	wire [WIDTH-1:0] wire_d25_112;
	wire [WIDTH-1:0] wire_d25_113;
	wire [WIDTH-1:0] wire_d25_114;
	wire [WIDTH-1:0] wire_d25_115;
	wire [WIDTH-1:0] wire_d25_116;
	wire [WIDTH-1:0] wire_d25_117;
	wire [WIDTH-1:0] wire_d25_118;
	wire [WIDTH-1:0] wire_d26_0;
	wire [WIDTH-1:0] wire_d26_1;
	wire [WIDTH-1:0] wire_d26_2;
	wire [WIDTH-1:0] wire_d26_3;
	wire [WIDTH-1:0] wire_d26_4;
	wire [WIDTH-1:0] wire_d26_5;
	wire [WIDTH-1:0] wire_d26_6;
	wire [WIDTH-1:0] wire_d26_7;
	wire [WIDTH-1:0] wire_d26_8;
	wire [WIDTH-1:0] wire_d26_9;
	wire [WIDTH-1:0] wire_d26_10;
	wire [WIDTH-1:0] wire_d26_11;
	wire [WIDTH-1:0] wire_d26_12;
	wire [WIDTH-1:0] wire_d26_13;
	wire [WIDTH-1:0] wire_d26_14;
	wire [WIDTH-1:0] wire_d26_15;
	wire [WIDTH-1:0] wire_d26_16;
	wire [WIDTH-1:0] wire_d26_17;
	wire [WIDTH-1:0] wire_d26_18;
	wire [WIDTH-1:0] wire_d26_19;
	wire [WIDTH-1:0] wire_d26_20;
	wire [WIDTH-1:0] wire_d26_21;
	wire [WIDTH-1:0] wire_d26_22;
	wire [WIDTH-1:0] wire_d26_23;
	wire [WIDTH-1:0] wire_d26_24;
	wire [WIDTH-1:0] wire_d26_25;
	wire [WIDTH-1:0] wire_d26_26;
	wire [WIDTH-1:0] wire_d26_27;
	wire [WIDTH-1:0] wire_d26_28;
	wire [WIDTH-1:0] wire_d26_29;
	wire [WIDTH-1:0] wire_d26_30;
	wire [WIDTH-1:0] wire_d26_31;
	wire [WIDTH-1:0] wire_d26_32;
	wire [WIDTH-1:0] wire_d26_33;
	wire [WIDTH-1:0] wire_d26_34;
	wire [WIDTH-1:0] wire_d26_35;
	wire [WIDTH-1:0] wire_d26_36;
	wire [WIDTH-1:0] wire_d26_37;
	wire [WIDTH-1:0] wire_d26_38;
	wire [WIDTH-1:0] wire_d26_39;
	wire [WIDTH-1:0] wire_d26_40;
	wire [WIDTH-1:0] wire_d26_41;
	wire [WIDTH-1:0] wire_d26_42;
	wire [WIDTH-1:0] wire_d26_43;
	wire [WIDTH-1:0] wire_d26_44;
	wire [WIDTH-1:0] wire_d26_45;
	wire [WIDTH-1:0] wire_d26_46;
	wire [WIDTH-1:0] wire_d26_47;
	wire [WIDTH-1:0] wire_d26_48;
	wire [WIDTH-1:0] wire_d26_49;
	wire [WIDTH-1:0] wire_d26_50;
	wire [WIDTH-1:0] wire_d26_51;
	wire [WIDTH-1:0] wire_d26_52;
	wire [WIDTH-1:0] wire_d26_53;
	wire [WIDTH-1:0] wire_d26_54;
	wire [WIDTH-1:0] wire_d26_55;
	wire [WIDTH-1:0] wire_d26_56;
	wire [WIDTH-1:0] wire_d26_57;
	wire [WIDTH-1:0] wire_d26_58;
	wire [WIDTH-1:0] wire_d26_59;
	wire [WIDTH-1:0] wire_d26_60;
	wire [WIDTH-1:0] wire_d26_61;
	wire [WIDTH-1:0] wire_d26_62;
	wire [WIDTH-1:0] wire_d26_63;
	wire [WIDTH-1:0] wire_d26_64;
	wire [WIDTH-1:0] wire_d26_65;
	wire [WIDTH-1:0] wire_d26_66;
	wire [WIDTH-1:0] wire_d26_67;
	wire [WIDTH-1:0] wire_d26_68;
	wire [WIDTH-1:0] wire_d26_69;
	wire [WIDTH-1:0] wire_d26_70;
	wire [WIDTH-1:0] wire_d26_71;
	wire [WIDTH-1:0] wire_d26_72;
	wire [WIDTH-1:0] wire_d26_73;
	wire [WIDTH-1:0] wire_d26_74;
	wire [WIDTH-1:0] wire_d26_75;
	wire [WIDTH-1:0] wire_d26_76;
	wire [WIDTH-1:0] wire_d26_77;
	wire [WIDTH-1:0] wire_d26_78;
	wire [WIDTH-1:0] wire_d26_79;
	wire [WIDTH-1:0] wire_d26_80;
	wire [WIDTH-1:0] wire_d26_81;
	wire [WIDTH-1:0] wire_d26_82;
	wire [WIDTH-1:0] wire_d26_83;
	wire [WIDTH-1:0] wire_d26_84;
	wire [WIDTH-1:0] wire_d26_85;
	wire [WIDTH-1:0] wire_d26_86;
	wire [WIDTH-1:0] wire_d26_87;
	wire [WIDTH-1:0] wire_d26_88;
	wire [WIDTH-1:0] wire_d26_89;
	wire [WIDTH-1:0] wire_d26_90;
	wire [WIDTH-1:0] wire_d26_91;
	wire [WIDTH-1:0] wire_d26_92;
	wire [WIDTH-1:0] wire_d26_93;
	wire [WIDTH-1:0] wire_d26_94;
	wire [WIDTH-1:0] wire_d26_95;
	wire [WIDTH-1:0] wire_d26_96;
	wire [WIDTH-1:0] wire_d26_97;
	wire [WIDTH-1:0] wire_d26_98;
	wire [WIDTH-1:0] wire_d26_99;
	wire [WIDTH-1:0] wire_d26_100;
	wire [WIDTH-1:0] wire_d26_101;
	wire [WIDTH-1:0] wire_d26_102;
	wire [WIDTH-1:0] wire_d26_103;
	wire [WIDTH-1:0] wire_d26_104;
	wire [WIDTH-1:0] wire_d26_105;
	wire [WIDTH-1:0] wire_d26_106;
	wire [WIDTH-1:0] wire_d26_107;
	wire [WIDTH-1:0] wire_d26_108;
	wire [WIDTH-1:0] wire_d26_109;
	wire [WIDTH-1:0] wire_d26_110;
	wire [WIDTH-1:0] wire_d26_111;
	wire [WIDTH-1:0] wire_d26_112;
	wire [WIDTH-1:0] wire_d26_113;
	wire [WIDTH-1:0] wire_d26_114;
	wire [WIDTH-1:0] wire_d26_115;
	wire [WIDTH-1:0] wire_d26_116;
	wire [WIDTH-1:0] wire_d26_117;
	wire [WIDTH-1:0] wire_d26_118;
	wire [WIDTH-1:0] wire_d27_0;
	wire [WIDTH-1:0] wire_d27_1;
	wire [WIDTH-1:0] wire_d27_2;
	wire [WIDTH-1:0] wire_d27_3;
	wire [WIDTH-1:0] wire_d27_4;
	wire [WIDTH-1:0] wire_d27_5;
	wire [WIDTH-1:0] wire_d27_6;
	wire [WIDTH-1:0] wire_d27_7;
	wire [WIDTH-1:0] wire_d27_8;
	wire [WIDTH-1:0] wire_d27_9;
	wire [WIDTH-1:0] wire_d27_10;
	wire [WIDTH-1:0] wire_d27_11;
	wire [WIDTH-1:0] wire_d27_12;
	wire [WIDTH-1:0] wire_d27_13;
	wire [WIDTH-1:0] wire_d27_14;
	wire [WIDTH-1:0] wire_d27_15;
	wire [WIDTH-1:0] wire_d27_16;
	wire [WIDTH-1:0] wire_d27_17;
	wire [WIDTH-1:0] wire_d27_18;
	wire [WIDTH-1:0] wire_d27_19;
	wire [WIDTH-1:0] wire_d27_20;
	wire [WIDTH-1:0] wire_d27_21;
	wire [WIDTH-1:0] wire_d27_22;
	wire [WIDTH-1:0] wire_d27_23;
	wire [WIDTH-1:0] wire_d27_24;
	wire [WIDTH-1:0] wire_d27_25;
	wire [WIDTH-1:0] wire_d27_26;
	wire [WIDTH-1:0] wire_d27_27;
	wire [WIDTH-1:0] wire_d27_28;
	wire [WIDTH-1:0] wire_d27_29;
	wire [WIDTH-1:0] wire_d27_30;
	wire [WIDTH-1:0] wire_d27_31;
	wire [WIDTH-1:0] wire_d27_32;
	wire [WIDTH-1:0] wire_d27_33;
	wire [WIDTH-1:0] wire_d27_34;
	wire [WIDTH-1:0] wire_d27_35;
	wire [WIDTH-1:0] wire_d27_36;
	wire [WIDTH-1:0] wire_d27_37;
	wire [WIDTH-1:0] wire_d27_38;
	wire [WIDTH-1:0] wire_d27_39;
	wire [WIDTH-1:0] wire_d27_40;
	wire [WIDTH-1:0] wire_d27_41;
	wire [WIDTH-1:0] wire_d27_42;
	wire [WIDTH-1:0] wire_d27_43;
	wire [WIDTH-1:0] wire_d27_44;
	wire [WIDTH-1:0] wire_d27_45;
	wire [WIDTH-1:0] wire_d27_46;
	wire [WIDTH-1:0] wire_d27_47;
	wire [WIDTH-1:0] wire_d27_48;
	wire [WIDTH-1:0] wire_d27_49;
	wire [WIDTH-1:0] wire_d27_50;
	wire [WIDTH-1:0] wire_d27_51;
	wire [WIDTH-1:0] wire_d27_52;
	wire [WIDTH-1:0] wire_d27_53;
	wire [WIDTH-1:0] wire_d27_54;
	wire [WIDTH-1:0] wire_d27_55;
	wire [WIDTH-1:0] wire_d27_56;
	wire [WIDTH-1:0] wire_d27_57;
	wire [WIDTH-1:0] wire_d27_58;
	wire [WIDTH-1:0] wire_d27_59;
	wire [WIDTH-1:0] wire_d27_60;
	wire [WIDTH-1:0] wire_d27_61;
	wire [WIDTH-1:0] wire_d27_62;
	wire [WIDTH-1:0] wire_d27_63;
	wire [WIDTH-1:0] wire_d27_64;
	wire [WIDTH-1:0] wire_d27_65;
	wire [WIDTH-1:0] wire_d27_66;
	wire [WIDTH-1:0] wire_d27_67;
	wire [WIDTH-1:0] wire_d27_68;
	wire [WIDTH-1:0] wire_d27_69;
	wire [WIDTH-1:0] wire_d27_70;
	wire [WIDTH-1:0] wire_d27_71;
	wire [WIDTH-1:0] wire_d27_72;
	wire [WIDTH-1:0] wire_d27_73;
	wire [WIDTH-1:0] wire_d27_74;
	wire [WIDTH-1:0] wire_d27_75;
	wire [WIDTH-1:0] wire_d27_76;
	wire [WIDTH-1:0] wire_d27_77;
	wire [WIDTH-1:0] wire_d27_78;
	wire [WIDTH-1:0] wire_d27_79;
	wire [WIDTH-1:0] wire_d27_80;
	wire [WIDTH-1:0] wire_d27_81;
	wire [WIDTH-1:0] wire_d27_82;
	wire [WIDTH-1:0] wire_d27_83;
	wire [WIDTH-1:0] wire_d27_84;
	wire [WIDTH-1:0] wire_d27_85;
	wire [WIDTH-1:0] wire_d27_86;
	wire [WIDTH-1:0] wire_d27_87;
	wire [WIDTH-1:0] wire_d27_88;
	wire [WIDTH-1:0] wire_d27_89;
	wire [WIDTH-1:0] wire_d27_90;
	wire [WIDTH-1:0] wire_d27_91;
	wire [WIDTH-1:0] wire_d27_92;
	wire [WIDTH-1:0] wire_d27_93;
	wire [WIDTH-1:0] wire_d27_94;
	wire [WIDTH-1:0] wire_d27_95;
	wire [WIDTH-1:0] wire_d27_96;
	wire [WIDTH-1:0] wire_d27_97;
	wire [WIDTH-1:0] wire_d27_98;
	wire [WIDTH-1:0] wire_d27_99;
	wire [WIDTH-1:0] wire_d27_100;
	wire [WIDTH-1:0] wire_d27_101;
	wire [WIDTH-1:0] wire_d27_102;
	wire [WIDTH-1:0] wire_d27_103;
	wire [WIDTH-1:0] wire_d27_104;
	wire [WIDTH-1:0] wire_d27_105;
	wire [WIDTH-1:0] wire_d27_106;
	wire [WIDTH-1:0] wire_d27_107;
	wire [WIDTH-1:0] wire_d27_108;
	wire [WIDTH-1:0] wire_d27_109;
	wire [WIDTH-1:0] wire_d27_110;
	wire [WIDTH-1:0] wire_d27_111;
	wire [WIDTH-1:0] wire_d27_112;
	wire [WIDTH-1:0] wire_d27_113;
	wire [WIDTH-1:0] wire_d27_114;
	wire [WIDTH-1:0] wire_d27_115;
	wire [WIDTH-1:0] wire_d27_116;
	wire [WIDTH-1:0] wire_d27_117;
	wire [WIDTH-1:0] wire_d27_118;
	wire [WIDTH-1:0] wire_d28_0;
	wire [WIDTH-1:0] wire_d28_1;
	wire [WIDTH-1:0] wire_d28_2;
	wire [WIDTH-1:0] wire_d28_3;
	wire [WIDTH-1:0] wire_d28_4;
	wire [WIDTH-1:0] wire_d28_5;
	wire [WIDTH-1:0] wire_d28_6;
	wire [WIDTH-1:0] wire_d28_7;
	wire [WIDTH-1:0] wire_d28_8;
	wire [WIDTH-1:0] wire_d28_9;
	wire [WIDTH-1:0] wire_d28_10;
	wire [WIDTH-1:0] wire_d28_11;
	wire [WIDTH-1:0] wire_d28_12;
	wire [WIDTH-1:0] wire_d28_13;
	wire [WIDTH-1:0] wire_d28_14;
	wire [WIDTH-1:0] wire_d28_15;
	wire [WIDTH-1:0] wire_d28_16;
	wire [WIDTH-1:0] wire_d28_17;
	wire [WIDTH-1:0] wire_d28_18;
	wire [WIDTH-1:0] wire_d28_19;
	wire [WIDTH-1:0] wire_d28_20;
	wire [WIDTH-1:0] wire_d28_21;
	wire [WIDTH-1:0] wire_d28_22;
	wire [WIDTH-1:0] wire_d28_23;
	wire [WIDTH-1:0] wire_d28_24;
	wire [WIDTH-1:0] wire_d28_25;
	wire [WIDTH-1:0] wire_d28_26;
	wire [WIDTH-1:0] wire_d28_27;
	wire [WIDTH-1:0] wire_d28_28;
	wire [WIDTH-1:0] wire_d28_29;
	wire [WIDTH-1:0] wire_d28_30;
	wire [WIDTH-1:0] wire_d28_31;
	wire [WIDTH-1:0] wire_d28_32;
	wire [WIDTH-1:0] wire_d28_33;
	wire [WIDTH-1:0] wire_d28_34;
	wire [WIDTH-1:0] wire_d28_35;
	wire [WIDTH-1:0] wire_d28_36;
	wire [WIDTH-1:0] wire_d28_37;
	wire [WIDTH-1:0] wire_d28_38;
	wire [WIDTH-1:0] wire_d28_39;
	wire [WIDTH-1:0] wire_d28_40;
	wire [WIDTH-1:0] wire_d28_41;
	wire [WIDTH-1:0] wire_d28_42;
	wire [WIDTH-1:0] wire_d28_43;
	wire [WIDTH-1:0] wire_d28_44;
	wire [WIDTH-1:0] wire_d28_45;
	wire [WIDTH-1:0] wire_d28_46;
	wire [WIDTH-1:0] wire_d28_47;
	wire [WIDTH-1:0] wire_d28_48;
	wire [WIDTH-1:0] wire_d28_49;
	wire [WIDTH-1:0] wire_d28_50;
	wire [WIDTH-1:0] wire_d28_51;
	wire [WIDTH-1:0] wire_d28_52;
	wire [WIDTH-1:0] wire_d28_53;
	wire [WIDTH-1:0] wire_d28_54;
	wire [WIDTH-1:0] wire_d28_55;
	wire [WIDTH-1:0] wire_d28_56;
	wire [WIDTH-1:0] wire_d28_57;
	wire [WIDTH-1:0] wire_d28_58;
	wire [WIDTH-1:0] wire_d28_59;
	wire [WIDTH-1:0] wire_d28_60;
	wire [WIDTH-1:0] wire_d28_61;
	wire [WIDTH-1:0] wire_d28_62;
	wire [WIDTH-1:0] wire_d28_63;
	wire [WIDTH-1:0] wire_d28_64;
	wire [WIDTH-1:0] wire_d28_65;
	wire [WIDTH-1:0] wire_d28_66;
	wire [WIDTH-1:0] wire_d28_67;
	wire [WIDTH-1:0] wire_d28_68;
	wire [WIDTH-1:0] wire_d28_69;
	wire [WIDTH-1:0] wire_d28_70;
	wire [WIDTH-1:0] wire_d28_71;
	wire [WIDTH-1:0] wire_d28_72;
	wire [WIDTH-1:0] wire_d28_73;
	wire [WIDTH-1:0] wire_d28_74;
	wire [WIDTH-1:0] wire_d28_75;
	wire [WIDTH-1:0] wire_d28_76;
	wire [WIDTH-1:0] wire_d28_77;
	wire [WIDTH-1:0] wire_d28_78;
	wire [WIDTH-1:0] wire_d28_79;
	wire [WIDTH-1:0] wire_d28_80;
	wire [WIDTH-1:0] wire_d28_81;
	wire [WIDTH-1:0] wire_d28_82;
	wire [WIDTH-1:0] wire_d28_83;
	wire [WIDTH-1:0] wire_d28_84;
	wire [WIDTH-1:0] wire_d28_85;
	wire [WIDTH-1:0] wire_d28_86;
	wire [WIDTH-1:0] wire_d28_87;
	wire [WIDTH-1:0] wire_d28_88;
	wire [WIDTH-1:0] wire_d28_89;
	wire [WIDTH-1:0] wire_d28_90;
	wire [WIDTH-1:0] wire_d28_91;
	wire [WIDTH-1:0] wire_d28_92;
	wire [WIDTH-1:0] wire_d28_93;
	wire [WIDTH-1:0] wire_d28_94;
	wire [WIDTH-1:0] wire_d28_95;
	wire [WIDTH-1:0] wire_d28_96;
	wire [WIDTH-1:0] wire_d28_97;
	wire [WIDTH-1:0] wire_d28_98;
	wire [WIDTH-1:0] wire_d28_99;
	wire [WIDTH-1:0] wire_d28_100;
	wire [WIDTH-1:0] wire_d28_101;
	wire [WIDTH-1:0] wire_d28_102;
	wire [WIDTH-1:0] wire_d28_103;
	wire [WIDTH-1:0] wire_d28_104;
	wire [WIDTH-1:0] wire_d28_105;
	wire [WIDTH-1:0] wire_d28_106;
	wire [WIDTH-1:0] wire_d28_107;
	wire [WIDTH-1:0] wire_d28_108;
	wire [WIDTH-1:0] wire_d28_109;
	wire [WIDTH-1:0] wire_d28_110;
	wire [WIDTH-1:0] wire_d28_111;
	wire [WIDTH-1:0] wire_d28_112;
	wire [WIDTH-1:0] wire_d28_113;
	wire [WIDTH-1:0] wire_d28_114;
	wire [WIDTH-1:0] wire_d28_115;
	wire [WIDTH-1:0] wire_d28_116;
	wire [WIDTH-1:0] wire_d28_117;
	wire [WIDTH-1:0] wire_d28_118;
	wire [WIDTH-1:0] wire_d29_0;
	wire [WIDTH-1:0] wire_d29_1;
	wire [WIDTH-1:0] wire_d29_2;
	wire [WIDTH-1:0] wire_d29_3;
	wire [WIDTH-1:0] wire_d29_4;
	wire [WIDTH-1:0] wire_d29_5;
	wire [WIDTH-1:0] wire_d29_6;
	wire [WIDTH-1:0] wire_d29_7;
	wire [WIDTH-1:0] wire_d29_8;
	wire [WIDTH-1:0] wire_d29_9;
	wire [WIDTH-1:0] wire_d29_10;
	wire [WIDTH-1:0] wire_d29_11;
	wire [WIDTH-1:0] wire_d29_12;
	wire [WIDTH-1:0] wire_d29_13;
	wire [WIDTH-1:0] wire_d29_14;
	wire [WIDTH-1:0] wire_d29_15;
	wire [WIDTH-1:0] wire_d29_16;
	wire [WIDTH-1:0] wire_d29_17;
	wire [WIDTH-1:0] wire_d29_18;
	wire [WIDTH-1:0] wire_d29_19;
	wire [WIDTH-1:0] wire_d29_20;
	wire [WIDTH-1:0] wire_d29_21;
	wire [WIDTH-1:0] wire_d29_22;
	wire [WIDTH-1:0] wire_d29_23;
	wire [WIDTH-1:0] wire_d29_24;
	wire [WIDTH-1:0] wire_d29_25;
	wire [WIDTH-1:0] wire_d29_26;
	wire [WIDTH-1:0] wire_d29_27;
	wire [WIDTH-1:0] wire_d29_28;
	wire [WIDTH-1:0] wire_d29_29;
	wire [WIDTH-1:0] wire_d29_30;
	wire [WIDTH-1:0] wire_d29_31;
	wire [WIDTH-1:0] wire_d29_32;
	wire [WIDTH-1:0] wire_d29_33;
	wire [WIDTH-1:0] wire_d29_34;
	wire [WIDTH-1:0] wire_d29_35;
	wire [WIDTH-1:0] wire_d29_36;
	wire [WIDTH-1:0] wire_d29_37;
	wire [WIDTH-1:0] wire_d29_38;
	wire [WIDTH-1:0] wire_d29_39;
	wire [WIDTH-1:0] wire_d29_40;
	wire [WIDTH-1:0] wire_d29_41;
	wire [WIDTH-1:0] wire_d29_42;
	wire [WIDTH-1:0] wire_d29_43;
	wire [WIDTH-1:0] wire_d29_44;
	wire [WIDTH-1:0] wire_d29_45;
	wire [WIDTH-1:0] wire_d29_46;
	wire [WIDTH-1:0] wire_d29_47;
	wire [WIDTH-1:0] wire_d29_48;
	wire [WIDTH-1:0] wire_d29_49;
	wire [WIDTH-1:0] wire_d29_50;
	wire [WIDTH-1:0] wire_d29_51;
	wire [WIDTH-1:0] wire_d29_52;
	wire [WIDTH-1:0] wire_d29_53;
	wire [WIDTH-1:0] wire_d29_54;
	wire [WIDTH-1:0] wire_d29_55;
	wire [WIDTH-1:0] wire_d29_56;
	wire [WIDTH-1:0] wire_d29_57;
	wire [WIDTH-1:0] wire_d29_58;
	wire [WIDTH-1:0] wire_d29_59;
	wire [WIDTH-1:0] wire_d29_60;
	wire [WIDTH-1:0] wire_d29_61;
	wire [WIDTH-1:0] wire_d29_62;
	wire [WIDTH-1:0] wire_d29_63;
	wire [WIDTH-1:0] wire_d29_64;
	wire [WIDTH-1:0] wire_d29_65;
	wire [WIDTH-1:0] wire_d29_66;
	wire [WIDTH-1:0] wire_d29_67;
	wire [WIDTH-1:0] wire_d29_68;
	wire [WIDTH-1:0] wire_d29_69;
	wire [WIDTH-1:0] wire_d29_70;
	wire [WIDTH-1:0] wire_d29_71;
	wire [WIDTH-1:0] wire_d29_72;
	wire [WIDTH-1:0] wire_d29_73;
	wire [WIDTH-1:0] wire_d29_74;
	wire [WIDTH-1:0] wire_d29_75;
	wire [WIDTH-1:0] wire_d29_76;
	wire [WIDTH-1:0] wire_d29_77;
	wire [WIDTH-1:0] wire_d29_78;
	wire [WIDTH-1:0] wire_d29_79;
	wire [WIDTH-1:0] wire_d29_80;
	wire [WIDTH-1:0] wire_d29_81;
	wire [WIDTH-1:0] wire_d29_82;
	wire [WIDTH-1:0] wire_d29_83;
	wire [WIDTH-1:0] wire_d29_84;
	wire [WIDTH-1:0] wire_d29_85;
	wire [WIDTH-1:0] wire_d29_86;
	wire [WIDTH-1:0] wire_d29_87;
	wire [WIDTH-1:0] wire_d29_88;
	wire [WIDTH-1:0] wire_d29_89;
	wire [WIDTH-1:0] wire_d29_90;
	wire [WIDTH-1:0] wire_d29_91;
	wire [WIDTH-1:0] wire_d29_92;
	wire [WIDTH-1:0] wire_d29_93;
	wire [WIDTH-1:0] wire_d29_94;
	wire [WIDTH-1:0] wire_d29_95;
	wire [WIDTH-1:0] wire_d29_96;
	wire [WIDTH-1:0] wire_d29_97;
	wire [WIDTH-1:0] wire_d29_98;
	wire [WIDTH-1:0] wire_d29_99;
	wire [WIDTH-1:0] wire_d29_100;
	wire [WIDTH-1:0] wire_d29_101;
	wire [WIDTH-1:0] wire_d29_102;
	wire [WIDTH-1:0] wire_d29_103;
	wire [WIDTH-1:0] wire_d29_104;
	wire [WIDTH-1:0] wire_d29_105;
	wire [WIDTH-1:0] wire_d29_106;
	wire [WIDTH-1:0] wire_d29_107;
	wire [WIDTH-1:0] wire_d29_108;
	wire [WIDTH-1:0] wire_d29_109;
	wire [WIDTH-1:0] wire_d29_110;
	wire [WIDTH-1:0] wire_d29_111;
	wire [WIDTH-1:0] wire_d29_112;
	wire [WIDTH-1:0] wire_d29_113;
	wire [WIDTH-1:0] wire_d29_114;
	wire [WIDTH-1:0] wire_d29_115;
	wire [WIDTH-1:0] wire_d29_116;
	wire [WIDTH-1:0] wire_d29_117;
	wire [WIDTH-1:0] wire_d29_118;
	wire [WIDTH-1:0] wire_d30_0;
	wire [WIDTH-1:0] wire_d30_1;
	wire [WIDTH-1:0] wire_d30_2;
	wire [WIDTH-1:0] wire_d30_3;
	wire [WIDTH-1:0] wire_d30_4;
	wire [WIDTH-1:0] wire_d30_5;
	wire [WIDTH-1:0] wire_d30_6;
	wire [WIDTH-1:0] wire_d30_7;
	wire [WIDTH-1:0] wire_d30_8;
	wire [WIDTH-1:0] wire_d30_9;
	wire [WIDTH-1:0] wire_d30_10;
	wire [WIDTH-1:0] wire_d30_11;
	wire [WIDTH-1:0] wire_d30_12;
	wire [WIDTH-1:0] wire_d30_13;
	wire [WIDTH-1:0] wire_d30_14;
	wire [WIDTH-1:0] wire_d30_15;
	wire [WIDTH-1:0] wire_d30_16;
	wire [WIDTH-1:0] wire_d30_17;
	wire [WIDTH-1:0] wire_d30_18;
	wire [WIDTH-1:0] wire_d30_19;
	wire [WIDTH-1:0] wire_d30_20;
	wire [WIDTH-1:0] wire_d30_21;
	wire [WIDTH-1:0] wire_d30_22;
	wire [WIDTH-1:0] wire_d30_23;
	wire [WIDTH-1:0] wire_d30_24;
	wire [WIDTH-1:0] wire_d30_25;
	wire [WIDTH-1:0] wire_d30_26;
	wire [WIDTH-1:0] wire_d30_27;
	wire [WIDTH-1:0] wire_d30_28;
	wire [WIDTH-1:0] wire_d30_29;
	wire [WIDTH-1:0] wire_d30_30;
	wire [WIDTH-1:0] wire_d30_31;
	wire [WIDTH-1:0] wire_d30_32;
	wire [WIDTH-1:0] wire_d30_33;
	wire [WIDTH-1:0] wire_d30_34;
	wire [WIDTH-1:0] wire_d30_35;
	wire [WIDTH-1:0] wire_d30_36;
	wire [WIDTH-1:0] wire_d30_37;
	wire [WIDTH-1:0] wire_d30_38;
	wire [WIDTH-1:0] wire_d30_39;
	wire [WIDTH-1:0] wire_d30_40;
	wire [WIDTH-1:0] wire_d30_41;
	wire [WIDTH-1:0] wire_d30_42;
	wire [WIDTH-1:0] wire_d30_43;
	wire [WIDTH-1:0] wire_d30_44;
	wire [WIDTH-1:0] wire_d30_45;
	wire [WIDTH-1:0] wire_d30_46;
	wire [WIDTH-1:0] wire_d30_47;
	wire [WIDTH-1:0] wire_d30_48;
	wire [WIDTH-1:0] wire_d30_49;
	wire [WIDTH-1:0] wire_d30_50;
	wire [WIDTH-1:0] wire_d30_51;
	wire [WIDTH-1:0] wire_d30_52;
	wire [WIDTH-1:0] wire_d30_53;
	wire [WIDTH-1:0] wire_d30_54;
	wire [WIDTH-1:0] wire_d30_55;
	wire [WIDTH-1:0] wire_d30_56;
	wire [WIDTH-1:0] wire_d30_57;
	wire [WIDTH-1:0] wire_d30_58;
	wire [WIDTH-1:0] wire_d30_59;
	wire [WIDTH-1:0] wire_d30_60;
	wire [WIDTH-1:0] wire_d30_61;
	wire [WIDTH-1:0] wire_d30_62;
	wire [WIDTH-1:0] wire_d30_63;
	wire [WIDTH-1:0] wire_d30_64;
	wire [WIDTH-1:0] wire_d30_65;
	wire [WIDTH-1:0] wire_d30_66;
	wire [WIDTH-1:0] wire_d30_67;
	wire [WIDTH-1:0] wire_d30_68;
	wire [WIDTH-1:0] wire_d30_69;
	wire [WIDTH-1:0] wire_d30_70;
	wire [WIDTH-1:0] wire_d30_71;
	wire [WIDTH-1:0] wire_d30_72;
	wire [WIDTH-1:0] wire_d30_73;
	wire [WIDTH-1:0] wire_d30_74;
	wire [WIDTH-1:0] wire_d30_75;
	wire [WIDTH-1:0] wire_d30_76;
	wire [WIDTH-1:0] wire_d30_77;
	wire [WIDTH-1:0] wire_d30_78;
	wire [WIDTH-1:0] wire_d30_79;
	wire [WIDTH-1:0] wire_d30_80;
	wire [WIDTH-1:0] wire_d30_81;
	wire [WIDTH-1:0] wire_d30_82;
	wire [WIDTH-1:0] wire_d30_83;
	wire [WIDTH-1:0] wire_d30_84;
	wire [WIDTH-1:0] wire_d30_85;
	wire [WIDTH-1:0] wire_d30_86;
	wire [WIDTH-1:0] wire_d30_87;
	wire [WIDTH-1:0] wire_d30_88;
	wire [WIDTH-1:0] wire_d30_89;
	wire [WIDTH-1:0] wire_d30_90;
	wire [WIDTH-1:0] wire_d30_91;
	wire [WIDTH-1:0] wire_d30_92;
	wire [WIDTH-1:0] wire_d30_93;
	wire [WIDTH-1:0] wire_d30_94;
	wire [WIDTH-1:0] wire_d30_95;
	wire [WIDTH-1:0] wire_d30_96;
	wire [WIDTH-1:0] wire_d30_97;
	wire [WIDTH-1:0] wire_d30_98;
	wire [WIDTH-1:0] wire_d30_99;
	wire [WIDTH-1:0] wire_d30_100;
	wire [WIDTH-1:0] wire_d30_101;
	wire [WIDTH-1:0] wire_d30_102;
	wire [WIDTH-1:0] wire_d30_103;
	wire [WIDTH-1:0] wire_d30_104;
	wire [WIDTH-1:0] wire_d30_105;
	wire [WIDTH-1:0] wire_d30_106;
	wire [WIDTH-1:0] wire_d30_107;
	wire [WIDTH-1:0] wire_d30_108;
	wire [WIDTH-1:0] wire_d30_109;
	wire [WIDTH-1:0] wire_d30_110;
	wire [WIDTH-1:0] wire_d30_111;
	wire [WIDTH-1:0] wire_d30_112;
	wire [WIDTH-1:0] wire_d30_113;
	wire [WIDTH-1:0] wire_d30_114;
	wire [WIDTH-1:0] wire_d30_115;
	wire [WIDTH-1:0] wire_d30_116;
	wire [WIDTH-1:0] wire_d30_117;
	wire [WIDTH-1:0] wire_d30_118;
	wire [WIDTH-1:0] wire_d31_0;
	wire [WIDTH-1:0] wire_d31_1;
	wire [WIDTH-1:0] wire_d31_2;
	wire [WIDTH-1:0] wire_d31_3;
	wire [WIDTH-1:0] wire_d31_4;
	wire [WIDTH-1:0] wire_d31_5;
	wire [WIDTH-1:0] wire_d31_6;
	wire [WIDTH-1:0] wire_d31_7;
	wire [WIDTH-1:0] wire_d31_8;
	wire [WIDTH-1:0] wire_d31_9;
	wire [WIDTH-1:0] wire_d31_10;
	wire [WIDTH-1:0] wire_d31_11;
	wire [WIDTH-1:0] wire_d31_12;
	wire [WIDTH-1:0] wire_d31_13;
	wire [WIDTH-1:0] wire_d31_14;
	wire [WIDTH-1:0] wire_d31_15;
	wire [WIDTH-1:0] wire_d31_16;
	wire [WIDTH-1:0] wire_d31_17;
	wire [WIDTH-1:0] wire_d31_18;
	wire [WIDTH-1:0] wire_d31_19;
	wire [WIDTH-1:0] wire_d31_20;
	wire [WIDTH-1:0] wire_d31_21;
	wire [WIDTH-1:0] wire_d31_22;
	wire [WIDTH-1:0] wire_d31_23;
	wire [WIDTH-1:0] wire_d31_24;
	wire [WIDTH-1:0] wire_d31_25;
	wire [WIDTH-1:0] wire_d31_26;
	wire [WIDTH-1:0] wire_d31_27;
	wire [WIDTH-1:0] wire_d31_28;
	wire [WIDTH-1:0] wire_d31_29;
	wire [WIDTH-1:0] wire_d31_30;
	wire [WIDTH-1:0] wire_d31_31;
	wire [WIDTH-1:0] wire_d31_32;
	wire [WIDTH-1:0] wire_d31_33;
	wire [WIDTH-1:0] wire_d31_34;
	wire [WIDTH-1:0] wire_d31_35;
	wire [WIDTH-1:0] wire_d31_36;
	wire [WIDTH-1:0] wire_d31_37;
	wire [WIDTH-1:0] wire_d31_38;
	wire [WIDTH-1:0] wire_d31_39;
	wire [WIDTH-1:0] wire_d31_40;
	wire [WIDTH-1:0] wire_d31_41;
	wire [WIDTH-1:0] wire_d31_42;
	wire [WIDTH-1:0] wire_d31_43;
	wire [WIDTH-1:0] wire_d31_44;
	wire [WIDTH-1:0] wire_d31_45;
	wire [WIDTH-1:0] wire_d31_46;
	wire [WIDTH-1:0] wire_d31_47;
	wire [WIDTH-1:0] wire_d31_48;
	wire [WIDTH-1:0] wire_d31_49;
	wire [WIDTH-1:0] wire_d31_50;
	wire [WIDTH-1:0] wire_d31_51;
	wire [WIDTH-1:0] wire_d31_52;
	wire [WIDTH-1:0] wire_d31_53;
	wire [WIDTH-1:0] wire_d31_54;
	wire [WIDTH-1:0] wire_d31_55;
	wire [WIDTH-1:0] wire_d31_56;
	wire [WIDTH-1:0] wire_d31_57;
	wire [WIDTH-1:0] wire_d31_58;
	wire [WIDTH-1:0] wire_d31_59;
	wire [WIDTH-1:0] wire_d31_60;
	wire [WIDTH-1:0] wire_d31_61;
	wire [WIDTH-1:0] wire_d31_62;
	wire [WIDTH-1:0] wire_d31_63;
	wire [WIDTH-1:0] wire_d31_64;
	wire [WIDTH-1:0] wire_d31_65;
	wire [WIDTH-1:0] wire_d31_66;
	wire [WIDTH-1:0] wire_d31_67;
	wire [WIDTH-1:0] wire_d31_68;
	wire [WIDTH-1:0] wire_d31_69;
	wire [WIDTH-1:0] wire_d31_70;
	wire [WIDTH-1:0] wire_d31_71;
	wire [WIDTH-1:0] wire_d31_72;
	wire [WIDTH-1:0] wire_d31_73;
	wire [WIDTH-1:0] wire_d31_74;
	wire [WIDTH-1:0] wire_d31_75;
	wire [WIDTH-1:0] wire_d31_76;
	wire [WIDTH-1:0] wire_d31_77;
	wire [WIDTH-1:0] wire_d31_78;
	wire [WIDTH-1:0] wire_d31_79;
	wire [WIDTH-1:0] wire_d31_80;
	wire [WIDTH-1:0] wire_d31_81;
	wire [WIDTH-1:0] wire_d31_82;
	wire [WIDTH-1:0] wire_d31_83;
	wire [WIDTH-1:0] wire_d31_84;
	wire [WIDTH-1:0] wire_d31_85;
	wire [WIDTH-1:0] wire_d31_86;
	wire [WIDTH-1:0] wire_d31_87;
	wire [WIDTH-1:0] wire_d31_88;
	wire [WIDTH-1:0] wire_d31_89;
	wire [WIDTH-1:0] wire_d31_90;
	wire [WIDTH-1:0] wire_d31_91;
	wire [WIDTH-1:0] wire_d31_92;
	wire [WIDTH-1:0] wire_d31_93;
	wire [WIDTH-1:0] wire_d31_94;
	wire [WIDTH-1:0] wire_d31_95;
	wire [WIDTH-1:0] wire_d31_96;
	wire [WIDTH-1:0] wire_d31_97;
	wire [WIDTH-1:0] wire_d31_98;
	wire [WIDTH-1:0] wire_d31_99;
	wire [WIDTH-1:0] wire_d31_100;
	wire [WIDTH-1:0] wire_d31_101;
	wire [WIDTH-1:0] wire_d31_102;
	wire [WIDTH-1:0] wire_d31_103;
	wire [WIDTH-1:0] wire_d31_104;
	wire [WIDTH-1:0] wire_d31_105;
	wire [WIDTH-1:0] wire_d31_106;
	wire [WIDTH-1:0] wire_d31_107;
	wire [WIDTH-1:0] wire_d31_108;
	wire [WIDTH-1:0] wire_d31_109;
	wire [WIDTH-1:0] wire_d31_110;
	wire [WIDTH-1:0] wire_d31_111;
	wire [WIDTH-1:0] wire_d31_112;
	wire [WIDTH-1:0] wire_d31_113;
	wire [WIDTH-1:0] wire_d31_114;
	wire [WIDTH-1:0] wire_d31_115;
	wire [WIDTH-1:0] wire_d31_116;
	wire [WIDTH-1:0] wire_d31_117;
	wire [WIDTH-1:0] wire_d31_118;
	wire [WIDTH-1:0] wire_d32_0;
	wire [WIDTH-1:0] wire_d32_1;
	wire [WIDTH-1:0] wire_d32_2;
	wire [WIDTH-1:0] wire_d32_3;
	wire [WIDTH-1:0] wire_d32_4;
	wire [WIDTH-1:0] wire_d32_5;
	wire [WIDTH-1:0] wire_d32_6;
	wire [WIDTH-1:0] wire_d32_7;
	wire [WIDTH-1:0] wire_d32_8;
	wire [WIDTH-1:0] wire_d32_9;
	wire [WIDTH-1:0] wire_d32_10;
	wire [WIDTH-1:0] wire_d32_11;
	wire [WIDTH-1:0] wire_d32_12;
	wire [WIDTH-1:0] wire_d32_13;
	wire [WIDTH-1:0] wire_d32_14;
	wire [WIDTH-1:0] wire_d32_15;
	wire [WIDTH-1:0] wire_d32_16;
	wire [WIDTH-1:0] wire_d32_17;
	wire [WIDTH-1:0] wire_d32_18;
	wire [WIDTH-1:0] wire_d32_19;
	wire [WIDTH-1:0] wire_d32_20;
	wire [WIDTH-1:0] wire_d32_21;
	wire [WIDTH-1:0] wire_d32_22;
	wire [WIDTH-1:0] wire_d32_23;
	wire [WIDTH-1:0] wire_d32_24;
	wire [WIDTH-1:0] wire_d32_25;
	wire [WIDTH-1:0] wire_d32_26;
	wire [WIDTH-1:0] wire_d32_27;
	wire [WIDTH-1:0] wire_d32_28;
	wire [WIDTH-1:0] wire_d32_29;
	wire [WIDTH-1:0] wire_d32_30;
	wire [WIDTH-1:0] wire_d32_31;
	wire [WIDTH-1:0] wire_d32_32;
	wire [WIDTH-1:0] wire_d32_33;
	wire [WIDTH-1:0] wire_d32_34;
	wire [WIDTH-1:0] wire_d32_35;
	wire [WIDTH-1:0] wire_d32_36;
	wire [WIDTH-1:0] wire_d32_37;
	wire [WIDTH-1:0] wire_d32_38;
	wire [WIDTH-1:0] wire_d32_39;
	wire [WIDTH-1:0] wire_d32_40;
	wire [WIDTH-1:0] wire_d32_41;
	wire [WIDTH-1:0] wire_d32_42;
	wire [WIDTH-1:0] wire_d32_43;
	wire [WIDTH-1:0] wire_d32_44;
	wire [WIDTH-1:0] wire_d32_45;
	wire [WIDTH-1:0] wire_d32_46;
	wire [WIDTH-1:0] wire_d32_47;
	wire [WIDTH-1:0] wire_d32_48;
	wire [WIDTH-1:0] wire_d32_49;
	wire [WIDTH-1:0] wire_d32_50;
	wire [WIDTH-1:0] wire_d32_51;
	wire [WIDTH-1:0] wire_d32_52;
	wire [WIDTH-1:0] wire_d32_53;
	wire [WIDTH-1:0] wire_d32_54;
	wire [WIDTH-1:0] wire_d32_55;
	wire [WIDTH-1:0] wire_d32_56;
	wire [WIDTH-1:0] wire_d32_57;
	wire [WIDTH-1:0] wire_d32_58;
	wire [WIDTH-1:0] wire_d32_59;
	wire [WIDTH-1:0] wire_d32_60;
	wire [WIDTH-1:0] wire_d32_61;
	wire [WIDTH-1:0] wire_d32_62;
	wire [WIDTH-1:0] wire_d32_63;
	wire [WIDTH-1:0] wire_d32_64;
	wire [WIDTH-1:0] wire_d32_65;
	wire [WIDTH-1:0] wire_d32_66;
	wire [WIDTH-1:0] wire_d32_67;
	wire [WIDTH-1:0] wire_d32_68;
	wire [WIDTH-1:0] wire_d32_69;
	wire [WIDTH-1:0] wire_d32_70;
	wire [WIDTH-1:0] wire_d32_71;
	wire [WIDTH-1:0] wire_d32_72;
	wire [WIDTH-1:0] wire_d32_73;
	wire [WIDTH-1:0] wire_d32_74;
	wire [WIDTH-1:0] wire_d32_75;
	wire [WIDTH-1:0] wire_d32_76;
	wire [WIDTH-1:0] wire_d32_77;
	wire [WIDTH-1:0] wire_d32_78;
	wire [WIDTH-1:0] wire_d32_79;
	wire [WIDTH-1:0] wire_d32_80;
	wire [WIDTH-1:0] wire_d32_81;
	wire [WIDTH-1:0] wire_d32_82;
	wire [WIDTH-1:0] wire_d32_83;
	wire [WIDTH-1:0] wire_d32_84;
	wire [WIDTH-1:0] wire_d32_85;
	wire [WIDTH-1:0] wire_d32_86;
	wire [WIDTH-1:0] wire_d32_87;
	wire [WIDTH-1:0] wire_d32_88;
	wire [WIDTH-1:0] wire_d32_89;
	wire [WIDTH-1:0] wire_d32_90;
	wire [WIDTH-1:0] wire_d32_91;
	wire [WIDTH-1:0] wire_d32_92;
	wire [WIDTH-1:0] wire_d32_93;
	wire [WIDTH-1:0] wire_d32_94;
	wire [WIDTH-1:0] wire_d32_95;
	wire [WIDTH-1:0] wire_d32_96;
	wire [WIDTH-1:0] wire_d32_97;
	wire [WIDTH-1:0] wire_d32_98;
	wire [WIDTH-1:0] wire_d32_99;
	wire [WIDTH-1:0] wire_d32_100;
	wire [WIDTH-1:0] wire_d32_101;
	wire [WIDTH-1:0] wire_d32_102;
	wire [WIDTH-1:0] wire_d32_103;
	wire [WIDTH-1:0] wire_d32_104;
	wire [WIDTH-1:0] wire_d32_105;
	wire [WIDTH-1:0] wire_d32_106;
	wire [WIDTH-1:0] wire_d32_107;
	wire [WIDTH-1:0] wire_d32_108;
	wire [WIDTH-1:0] wire_d32_109;
	wire [WIDTH-1:0] wire_d32_110;
	wire [WIDTH-1:0] wire_d32_111;
	wire [WIDTH-1:0] wire_d32_112;
	wire [WIDTH-1:0] wire_d32_113;
	wire [WIDTH-1:0] wire_d32_114;
	wire [WIDTH-1:0] wire_d32_115;
	wire [WIDTH-1:0] wire_d32_116;
	wire [WIDTH-1:0] wire_d32_117;
	wire [WIDTH-1:0] wire_d32_118;
	wire [WIDTH-1:0] wire_d33_0;
	wire [WIDTH-1:0] wire_d33_1;
	wire [WIDTH-1:0] wire_d33_2;
	wire [WIDTH-1:0] wire_d33_3;
	wire [WIDTH-1:0] wire_d33_4;
	wire [WIDTH-1:0] wire_d33_5;
	wire [WIDTH-1:0] wire_d33_6;
	wire [WIDTH-1:0] wire_d33_7;
	wire [WIDTH-1:0] wire_d33_8;
	wire [WIDTH-1:0] wire_d33_9;
	wire [WIDTH-1:0] wire_d33_10;
	wire [WIDTH-1:0] wire_d33_11;
	wire [WIDTH-1:0] wire_d33_12;
	wire [WIDTH-1:0] wire_d33_13;
	wire [WIDTH-1:0] wire_d33_14;
	wire [WIDTH-1:0] wire_d33_15;
	wire [WIDTH-1:0] wire_d33_16;
	wire [WIDTH-1:0] wire_d33_17;
	wire [WIDTH-1:0] wire_d33_18;
	wire [WIDTH-1:0] wire_d33_19;
	wire [WIDTH-1:0] wire_d33_20;
	wire [WIDTH-1:0] wire_d33_21;
	wire [WIDTH-1:0] wire_d33_22;
	wire [WIDTH-1:0] wire_d33_23;
	wire [WIDTH-1:0] wire_d33_24;
	wire [WIDTH-1:0] wire_d33_25;
	wire [WIDTH-1:0] wire_d33_26;
	wire [WIDTH-1:0] wire_d33_27;
	wire [WIDTH-1:0] wire_d33_28;
	wire [WIDTH-1:0] wire_d33_29;
	wire [WIDTH-1:0] wire_d33_30;
	wire [WIDTH-1:0] wire_d33_31;
	wire [WIDTH-1:0] wire_d33_32;
	wire [WIDTH-1:0] wire_d33_33;
	wire [WIDTH-1:0] wire_d33_34;
	wire [WIDTH-1:0] wire_d33_35;
	wire [WIDTH-1:0] wire_d33_36;
	wire [WIDTH-1:0] wire_d33_37;
	wire [WIDTH-1:0] wire_d33_38;
	wire [WIDTH-1:0] wire_d33_39;
	wire [WIDTH-1:0] wire_d33_40;
	wire [WIDTH-1:0] wire_d33_41;
	wire [WIDTH-1:0] wire_d33_42;
	wire [WIDTH-1:0] wire_d33_43;
	wire [WIDTH-1:0] wire_d33_44;
	wire [WIDTH-1:0] wire_d33_45;
	wire [WIDTH-1:0] wire_d33_46;
	wire [WIDTH-1:0] wire_d33_47;
	wire [WIDTH-1:0] wire_d33_48;
	wire [WIDTH-1:0] wire_d33_49;
	wire [WIDTH-1:0] wire_d33_50;
	wire [WIDTH-1:0] wire_d33_51;
	wire [WIDTH-1:0] wire_d33_52;
	wire [WIDTH-1:0] wire_d33_53;
	wire [WIDTH-1:0] wire_d33_54;
	wire [WIDTH-1:0] wire_d33_55;
	wire [WIDTH-1:0] wire_d33_56;
	wire [WIDTH-1:0] wire_d33_57;
	wire [WIDTH-1:0] wire_d33_58;
	wire [WIDTH-1:0] wire_d33_59;
	wire [WIDTH-1:0] wire_d33_60;
	wire [WIDTH-1:0] wire_d33_61;
	wire [WIDTH-1:0] wire_d33_62;
	wire [WIDTH-1:0] wire_d33_63;
	wire [WIDTH-1:0] wire_d33_64;
	wire [WIDTH-1:0] wire_d33_65;
	wire [WIDTH-1:0] wire_d33_66;
	wire [WIDTH-1:0] wire_d33_67;
	wire [WIDTH-1:0] wire_d33_68;
	wire [WIDTH-1:0] wire_d33_69;
	wire [WIDTH-1:0] wire_d33_70;
	wire [WIDTH-1:0] wire_d33_71;
	wire [WIDTH-1:0] wire_d33_72;
	wire [WIDTH-1:0] wire_d33_73;
	wire [WIDTH-1:0] wire_d33_74;
	wire [WIDTH-1:0] wire_d33_75;
	wire [WIDTH-1:0] wire_d33_76;
	wire [WIDTH-1:0] wire_d33_77;
	wire [WIDTH-1:0] wire_d33_78;
	wire [WIDTH-1:0] wire_d33_79;
	wire [WIDTH-1:0] wire_d33_80;
	wire [WIDTH-1:0] wire_d33_81;
	wire [WIDTH-1:0] wire_d33_82;
	wire [WIDTH-1:0] wire_d33_83;
	wire [WIDTH-1:0] wire_d33_84;
	wire [WIDTH-1:0] wire_d33_85;
	wire [WIDTH-1:0] wire_d33_86;
	wire [WIDTH-1:0] wire_d33_87;
	wire [WIDTH-1:0] wire_d33_88;
	wire [WIDTH-1:0] wire_d33_89;
	wire [WIDTH-1:0] wire_d33_90;
	wire [WIDTH-1:0] wire_d33_91;
	wire [WIDTH-1:0] wire_d33_92;
	wire [WIDTH-1:0] wire_d33_93;
	wire [WIDTH-1:0] wire_d33_94;
	wire [WIDTH-1:0] wire_d33_95;
	wire [WIDTH-1:0] wire_d33_96;
	wire [WIDTH-1:0] wire_d33_97;
	wire [WIDTH-1:0] wire_d33_98;
	wire [WIDTH-1:0] wire_d33_99;
	wire [WIDTH-1:0] wire_d33_100;
	wire [WIDTH-1:0] wire_d33_101;
	wire [WIDTH-1:0] wire_d33_102;
	wire [WIDTH-1:0] wire_d33_103;
	wire [WIDTH-1:0] wire_d33_104;
	wire [WIDTH-1:0] wire_d33_105;
	wire [WIDTH-1:0] wire_d33_106;
	wire [WIDTH-1:0] wire_d33_107;
	wire [WIDTH-1:0] wire_d33_108;
	wire [WIDTH-1:0] wire_d33_109;
	wire [WIDTH-1:0] wire_d33_110;
	wire [WIDTH-1:0] wire_d33_111;
	wire [WIDTH-1:0] wire_d33_112;
	wire [WIDTH-1:0] wire_d33_113;
	wire [WIDTH-1:0] wire_d33_114;
	wire [WIDTH-1:0] wire_d33_115;
	wire [WIDTH-1:0] wire_d33_116;
	wire [WIDTH-1:0] wire_d33_117;
	wire [WIDTH-1:0] wire_d33_118;
	wire [WIDTH-1:0] wire_d34_0;
	wire [WIDTH-1:0] wire_d34_1;
	wire [WIDTH-1:0] wire_d34_2;
	wire [WIDTH-1:0] wire_d34_3;
	wire [WIDTH-1:0] wire_d34_4;
	wire [WIDTH-1:0] wire_d34_5;
	wire [WIDTH-1:0] wire_d34_6;
	wire [WIDTH-1:0] wire_d34_7;
	wire [WIDTH-1:0] wire_d34_8;
	wire [WIDTH-1:0] wire_d34_9;
	wire [WIDTH-1:0] wire_d34_10;
	wire [WIDTH-1:0] wire_d34_11;
	wire [WIDTH-1:0] wire_d34_12;
	wire [WIDTH-1:0] wire_d34_13;
	wire [WIDTH-1:0] wire_d34_14;
	wire [WIDTH-1:0] wire_d34_15;
	wire [WIDTH-1:0] wire_d34_16;
	wire [WIDTH-1:0] wire_d34_17;
	wire [WIDTH-1:0] wire_d34_18;
	wire [WIDTH-1:0] wire_d34_19;
	wire [WIDTH-1:0] wire_d34_20;
	wire [WIDTH-1:0] wire_d34_21;
	wire [WIDTH-1:0] wire_d34_22;
	wire [WIDTH-1:0] wire_d34_23;
	wire [WIDTH-1:0] wire_d34_24;
	wire [WIDTH-1:0] wire_d34_25;
	wire [WIDTH-1:0] wire_d34_26;
	wire [WIDTH-1:0] wire_d34_27;
	wire [WIDTH-1:0] wire_d34_28;
	wire [WIDTH-1:0] wire_d34_29;
	wire [WIDTH-1:0] wire_d34_30;
	wire [WIDTH-1:0] wire_d34_31;
	wire [WIDTH-1:0] wire_d34_32;
	wire [WIDTH-1:0] wire_d34_33;
	wire [WIDTH-1:0] wire_d34_34;
	wire [WIDTH-1:0] wire_d34_35;
	wire [WIDTH-1:0] wire_d34_36;
	wire [WIDTH-1:0] wire_d34_37;
	wire [WIDTH-1:0] wire_d34_38;
	wire [WIDTH-1:0] wire_d34_39;
	wire [WIDTH-1:0] wire_d34_40;
	wire [WIDTH-1:0] wire_d34_41;
	wire [WIDTH-1:0] wire_d34_42;
	wire [WIDTH-1:0] wire_d34_43;
	wire [WIDTH-1:0] wire_d34_44;
	wire [WIDTH-1:0] wire_d34_45;
	wire [WIDTH-1:0] wire_d34_46;
	wire [WIDTH-1:0] wire_d34_47;
	wire [WIDTH-1:0] wire_d34_48;
	wire [WIDTH-1:0] wire_d34_49;
	wire [WIDTH-1:0] wire_d34_50;
	wire [WIDTH-1:0] wire_d34_51;
	wire [WIDTH-1:0] wire_d34_52;
	wire [WIDTH-1:0] wire_d34_53;
	wire [WIDTH-1:0] wire_d34_54;
	wire [WIDTH-1:0] wire_d34_55;
	wire [WIDTH-1:0] wire_d34_56;
	wire [WIDTH-1:0] wire_d34_57;
	wire [WIDTH-1:0] wire_d34_58;
	wire [WIDTH-1:0] wire_d34_59;
	wire [WIDTH-1:0] wire_d34_60;
	wire [WIDTH-1:0] wire_d34_61;
	wire [WIDTH-1:0] wire_d34_62;
	wire [WIDTH-1:0] wire_d34_63;
	wire [WIDTH-1:0] wire_d34_64;
	wire [WIDTH-1:0] wire_d34_65;
	wire [WIDTH-1:0] wire_d34_66;
	wire [WIDTH-1:0] wire_d34_67;
	wire [WIDTH-1:0] wire_d34_68;
	wire [WIDTH-1:0] wire_d34_69;
	wire [WIDTH-1:0] wire_d34_70;
	wire [WIDTH-1:0] wire_d34_71;
	wire [WIDTH-1:0] wire_d34_72;
	wire [WIDTH-1:0] wire_d34_73;
	wire [WIDTH-1:0] wire_d34_74;
	wire [WIDTH-1:0] wire_d34_75;
	wire [WIDTH-1:0] wire_d34_76;
	wire [WIDTH-1:0] wire_d34_77;
	wire [WIDTH-1:0] wire_d34_78;
	wire [WIDTH-1:0] wire_d34_79;
	wire [WIDTH-1:0] wire_d34_80;
	wire [WIDTH-1:0] wire_d34_81;
	wire [WIDTH-1:0] wire_d34_82;
	wire [WIDTH-1:0] wire_d34_83;
	wire [WIDTH-1:0] wire_d34_84;
	wire [WIDTH-1:0] wire_d34_85;
	wire [WIDTH-1:0] wire_d34_86;
	wire [WIDTH-1:0] wire_d34_87;
	wire [WIDTH-1:0] wire_d34_88;
	wire [WIDTH-1:0] wire_d34_89;
	wire [WIDTH-1:0] wire_d34_90;
	wire [WIDTH-1:0] wire_d34_91;
	wire [WIDTH-1:0] wire_d34_92;
	wire [WIDTH-1:0] wire_d34_93;
	wire [WIDTH-1:0] wire_d34_94;
	wire [WIDTH-1:0] wire_d34_95;
	wire [WIDTH-1:0] wire_d34_96;
	wire [WIDTH-1:0] wire_d34_97;
	wire [WIDTH-1:0] wire_d34_98;
	wire [WIDTH-1:0] wire_d34_99;
	wire [WIDTH-1:0] wire_d34_100;
	wire [WIDTH-1:0] wire_d34_101;
	wire [WIDTH-1:0] wire_d34_102;
	wire [WIDTH-1:0] wire_d34_103;
	wire [WIDTH-1:0] wire_d34_104;
	wire [WIDTH-1:0] wire_d34_105;
	wire [WIDTH-1:0] wire_d34_106;
	wire [WIDTH-1:0] wire_d34_107;
	wire [WIDTH-1:0] wire_d34_108;
	wire [WIDTH-1:0] wire_d34_109;
	wire [WIDTH-1:0] wire_d34_110;
	wire [WIDTH-1:0] wire_d34_111;
	wire [WIDTH-1:0] wire_d34_112;
	wire [WIDTH-1:0] wire_d34_113;
	wire [WIDTH-1:0] wire_d34_114;
	wire [WIDTH-1:0] wire_d34_115;
	wire [WIDTH-1:0] wire_d34_116;
	wire [WIDTH-1:0] wire_d34_117;
	wire [WIDTH-1:0] wire_d34_118;
	wire [WIDTH-1:0] wire_d35_0;
	wire [WIDTH-1:0] wire_d35_1;
	wire [WIDTH-1:0] wire_d35_2;
	wire [WIDTH-1:0] wire_d35_3;
	wire [WIDTH-1:0] wire_d35_4;
	wire [WIDTH-1:0] wire_d35_5;
	wire [WIDTH-1:0] wire_d35_6;
	wire [WIDTH-1:0] wire_d35_7;
	wire [WIDTH-1:0] wire_d35_8;
	wire [WIDTH-1:0] wire_d35_9;
	wire [WIDTH-1:0] wire_d35_10;
	wire [WIDTH-1:0] wire_d35_11;
	wire [WIDTH-1:0] wire_d35_12;
	wire [WIDTH-1:0] wire_d35_13;
	wire [WIDTH-1:0] wire_d35_14;
	wire [WIDTH-1:0] wire_d35_15;
	wire [WIDTH-1:0] wire_d35_16;
	wire [WIDTH-1:0] wire_d35_17;
	wire [WIDTH-1:0] wire_d35_18;
	wire [WIDTH-1:0] wire_d35_19;
	wire [WIDTH-1:0] wire_d35_20;
	wire [WIDTH-1:0] wire_d35_21;
	wire [WIDTH-1:0] wire_d35_22;
	wire [WIDTH-1:0] wire_d35_23;
	wire [WIDTH-1:0] wire_d35_24;
	wire [WIDTH-1:0] wire_d35_25;
	wire [WIDTH-1:0] wire_d35_26;
	wire [WIDTH-1:0] wire_d35_27;
	wire [WIDTH-1:0] wire_d35_28;
	wire [WIDTH-1:0] wire_d35_29;
	wire [WIDTH-1:0] wire_d35_30;
	wire [WIDTH-1:0] wire_d35_31;
	wire [WIDTH-1:0] wire_d35_32;
	wire [WIDTH-1:0] wire_d35_33;
	wire [WIDTH-1:0] wire_d35_34;
	wire [WIDTH-1:0] wire_d35_35;
	wire [WIDTH-1:0] wire_d35_36;
	wire [WIDTH-1:0] wire_d35_37;
	wire [WIDTH-1:0] wire_d35_38;
	wire [WIDTH-1:0] wire_d35_39;
	wire [WIDTH-1:0] wire_d35_40;
	wire [WIDTH-1:0] wire_d35_41;
	wire [WIDTH-1:0] wire_d35_42;
	wire [WIDTH-1:0] wire_d35_43;
	wire [WIDTH-1:0] wire_d35_44;
	wire [WIDTH-1:0] wire_d35_45;
	wire [WIDTH-1:0] wire_d35_46;
	wire [WIDTH-1:0] wire_d35_47;
	wire [WIDTH-1:0] wire_d35_48;
	wire [WIDTH-1:0] wire_d35_49;
	wire [WIDTH-1:0] wire_d35_50;
	wire [WIDTH-1:0] wire_d35_51;
	wire [WIDTH-1:0] wire_d35_52;
	wire [WIDTH-1:0] wire_d35_53;
	wire [WIDTH-1:0] wire_d35_54;
	wire [WIDTH-1:0] wire_d35_55;
	wire [WIDTH-1:0] wire_d35_56;
	wire [WIDTH-1:0] wire_d35_57;
	wire [WIDTH-1:0] wire_d35_58;
	wire [WIDTH-1:0] wire_d35_59;
	wire [WIDTH-1:0] wire_d35_60;
	wire [WIDTH-1:0] wire_d35_61;
	wire [WIDTH-1:0] wire_d35_62;
	wire [WIDTH-1:0] wire_d35_63;
	wire [WIDTH-1:0] wire_d35_64;
	wire [WIDTH-1:0] wire_d35_65;
	wire [WIDTH-1:0] wire_d35_66;
	wire [WIDTH-1:0] wire_d35_67;
	wire [WIDTH-1:0] wire_d35_68;
	wire [WIDTH-1:0] wire_d35_69;
	wire [WIDTH-1:0] wire_d35_70;
	wire [WIDTH-1:0] wire_d35_71;
	wire [WIDTH-1:0] wire_d35_72;
	wire [WIDTH-1:0] wire_d35_73;
	wire [WIDTH-1:0] wire_d35_74;
	wire [WIDTH-1:0] wire_d35_75;
	wire [WIDTH-1:0] wire_d35_76;
	wire [WIDTH-1:0] wire_d35_77;
	wire [WIDTH-1:0] wire_d35_78;
	wire [WIDTH-1:0] wire_d35_79;
	wire [WIDTH-1:0] wire_d35_80;
	wire [WIDTH-1:0] wire_d35_81;
	wire [WIDTH-1:0] wire_d35_82;
	wire [WIDTH-1:0] wire_d35_83;
	wire [WIDTH-1:0] wire_d35_84;
	wire [WIDTH-1:0] wire_d35_85;
	wire [WIDTH-1:0] wire_d35_86;
	wire [WIDTH-1:0] wire_d35_87;
	wire [WIDTH-1:0] wire_d35_88;
	wire [WIDTH-1:0] wire_d35_89;
	wire [WIDTH-1:0] wire_d35_90;
	wire [WIDTH-1:0] wire_d35_91;
	wire [WIDTH-1:0] wire_d35_92;
	wire [WIDTH-1:0] wire_d35_93;
	wire [WIDTH-1:0] wire_d35_94;
	wire [WIDTH-1:0] wire_d35_95;
	wire [WIDTH-1:0] wire_d35_96;
	wire [WIDTH-1:0] wire_d35_97;
	wire [WIDTH-1:0] wire_d35_98;
	wire [WIDTH-1:0] wire_d35_99;
	wire [WIDTH-1:0] wire_d35_100;
	wire [WIDTH-1:0] wire_d35_101;
	wire [WIDTH-1:0] wire_d35_102;
	wire [WIDTH-1:0] wire_d35_103;
	wire [WIDTH-1:0] wire_d35_104;
	wire [WIDTH-1:0] wire_d35_105;
	wire [WIDTH-1:0] wire_d35_106;
	wire [WIDTH-1:0] wire_d35_107;
	wire [WIDTH-1:0] wire_d35_108;
	wire [WIDTH-1:0] wire_d35_109;
	wire [WIDTH-1:0] wire_d35_110;
	wire [WIDTH-1:0] wire_d35_111;
	wire [WIDTH-1:0] wire_d35_112;
	wire [WIDTH-1:0] wire_d35_113;
	wire [WIDTH-1:0] wire_d35_114;
	wire [WIDTH-1:0] wire_d35_115;
	wire [WIDTH-1:0] wire_d35_116;
	wire [WIDTH-1:0] wire_d35_117;
	wire [WIDTH-1:0] wire_d35_118;
	wire [WIDTH-1:0] wire_d36_0;
	wire [WIDTH-1:0] wire_d36_1;
	wire [WIDTH-1:0] wire_d36_2;
	wire [WIDTH-1:0] wire_d36_3;
	wire [WIDTH-1:0] wire_d36_4;
	wire [WIDTH-1:0] wire_d36_5;
	wire [WIDTH-1:0] wire_d36_6;
	wire [WIDTH-1:0] wire_d36_7;
	wire [WIDTH-1:0] wire_d36_8;
	wire [WIDTH-1:0] wire_d36_9;
	wire [WIDTH-1:0] wire_d36_10;
	wire [WIDTH-1:0] wire_d36_11;
	wire [WIDTH-1:0] wire_d36_12;
	wire [WIDTH-1:0] wire_d36_13;
	wire [WIDTH-1:0] wire_d36_14;
	wire [WIDTH-1:0] wire_d36_15;
	wire [WIDTH-1:0] wire_d36_16;
	wire [WIDTH-1:0] wire_d36_17;
	wire [WIDTH-1:0] wire_d36_18;
	wire [WIDTH-1:0] wire_d36_19;
	wire [WIDTH-1:0] wire_d36_20;
	wire [WIDTH-1:0] wire_d36_21;
	wire [WIDTH-1:0] wire_d36_22;
	wire [WIDTH-1:0] wire_d36_23;
	wire [WIDTH-1:0] wire_d36_24;
	wire [WIDTH-1:0] wire_d36_25;
	wire [WIDTH-1:0] wire_d36_26;
	wire [WIDTH-1:0] wire_d36_27;
	wire [WIDTH-1:0] wire_d36_28;
	wire [WIDTH-1:0] wire_d36_29;
	wire [WIDTH-1:0] wire_d36_30;
	wire [WIDTH-1:0] wire_d36_31;
	wire [WIDTH-1:0] wire_d36_32;
	wire [WIDTH-1:0] wire_d36_33;
	wire [WIDTH-1:0] wire_d36_34;
	wire [WIDTH-1:0] wire_d36_35;
	wire [WIDTH-1:0] wire_d36_36;
	wire [WIDTH-1:0] wire_d36_37;
	wire [WIDTH-1:0] wire_d36_38;
	wire [WIDTH-1:0] wire_d36_39;
	wire [WIDTH-1:0] wire_d36_40;
	wire [WIDTH-1:0] wire_d36_41;
	wire [WIDTH-1:0] wire_d36_42;
	wire [WIDTH-1:0] wire_d36_43;
	wire [WIDTH-1:0] wire_d36_44;
	wire [WIDTH-1:0] wire_d36_45;
	wire [WIDTH-1:0] wire_d36_46;
	wire [WIDTH-1:0] wire_d36_47;
	wire [WIDTH-1:0] wire_d36_48;
	wire [WIDTH-1:0] wire_d36_49;
	wire [WIDTH-1:0] wire_d36_50;
	wire [WIDTH-1:0] wire_d36_51;
	wire [WIDTH-1:0] wire_d36_52;
	wire [WIDTH-1:0] wire_d36_53;
	wire [WIDTH-1:0] wire_d36_54;
	wire [WIDTH-1:0] wire_d36_55;
	wire [WIDTH-1:0] wire_d36_56;
	wire [WIDTH-1:0] wire_d36_57;
	wire [WIDTH-1:0] wire_d36_58;
	wire [WIDTH-1:0] wire_d36_59;
	wire [WIDTH-1:0] wire_d36_60;
	wire [WIDTH-1:0] wire_d36_61;
	wire [WIDTH-1:0] wire_d36_62;
	wire [WIDTH-1:0] wire_d36_63;
	wire [WIDTH-1:0] wire_d36_64;
	wire [WIDTH-1:0] wire_d36_65;
	wire [WIDTH-1:0] wire_d36_66;
	wire [WIDTH-1:0] wire_d36_67;
	wire [WIDTH-1:0] wire_d36_68;
	wire [WIDTH-1:0] wire_d36_69;
	wire [WIDTH-1:0] wire_d36_70;
	wire [WIDTH-1:0] wire_d36_71;
	wire [WIDTH-1:0] wire_d36_72;
	wire [WIDTH-1:0] wire_d36_73;
	wire [WIDTH-1:0] wire_d36_74;
	wire [WIDTH-1:0] wire_d36_75;
	wire [WIDTH-1:0] wire_d36_76;
	wire [WIDTH-1:0] wire_d36_77;
	wire [WIDTH-1:0] wire_d36_78;
	wire [WIDTH-1:0] wire_d36_79;
	wire [WIDTH-1:0] wire_d36_80;
	wire [WIDTH-1:0] wire_d36_81;
	wire [WIDTH-1:0] wire_d36_82;
	wire [WIDTH-1:0] wire_d36_83;
	wire [WIDTH-1:0] wire_d36_84;
	wire [WIDTH-1:0] wire_d36_85;
	wire [WIDTH-1:0] wire_d36_86;
	wire [WIDTH-1:0] wire_d36_87;
	wire [WIDTH-1:0] wire_d36_88;
	wire [WIDTH-1:0] wire_d36_89;
	wire [WIDTH-1:0] wire_d36_90;
	wire [WIDTH-1:0] wire_d36_91;
	wire [WIDTH-1:0] wire_d36_92;
	wire [WIDTH-1:0] wire_d36_93;
	wire [WIDTH-1:0] wire_d36_94;
	wire [WIDTH-1:0] wire_d36_95;
	wire [WIDTH-1:0] wire_d36_96;
	wire [WIDTH-1:0] wire_d36_97;
	wire [WIDTH-1:0] wire_d36_98;
	wire [WIDTH-1:0] wire_d36_99;
	wire [WIDTH-1:0] wire_d36_100;
	wire [WIDTH-1:0] wire_d36_101;
	wire [WIDTH-1:0] wire_d36_102;
	wire [WIDTH-1:0] wire_d36_103;
	wire [WIDTH-1:0] wire_d36_104;
	wire [WIDTH-1:0] wire_d36_105;
	wire [WIDTH-1:0] wire_d36_106;
	wire [WIDTH-1:0] wire_d36_107;
	wire [WIDTH-1:0] wire_d36_108;
	wire [WIDTH-1:0] wire_d36_109;
	wire [WIDTH-1:0] wire_d36_110;
	wire [WIDTH-1:0] wire_d36_111;
	wire [WIDTH-1:0] wire_d36_112;
	wire [WIDTH-1:0] wire_d36_113;
	wire [WIDTH-1:0] wire_d36_114;
	wire [WIDTH-1:0] wire_d36_115;
	wire [WIDTH-1:0] wire_d36_116;
	wire [WIDTH-1:0] wire_d36_117;
	wire [WIDTH-1:0] wire_d36_118;
	wire [WIDTH-1:0] wire_d37_0;
	wire [WIDTH-1:0] wire_d37_1;
	wire [WIDTH-1:0] wire_d37_2;
	wire [WIDTH-1:0] wire_d37_3;
	wire [WIDTH-1:0] wire_d37_4;
	wire [WIDTH-1:0] wire_d37_5;
	wire [WIDTH-1:0] wire_d37_6;
	wire [WIDTH-1:0] wire_d37_7;
	wire [WIDTH-1:0] wire_d37_8;
	wire [WIDTH-1:0] wire_d37_9;
	wire [WIDTH-1:0] wire_d37_10;
	wire [WIDTH-1:0] wire_d37_11;
	wire [WIDTH-1:0] wire_d37_12;
	wire [WIDTH-1:0] wire_d37_13;
	wire [WIDTH-1:0] wire_d37_14;
	wire [WIDTH-1:0] wire_d37_15;
	wire [WIDTH-1:0] wire_d37_16;
	wire [WIDTH-1:0] wire_d37_17;
	wire [WIDTH-1:0] wire_d37_18;
	wire [WIDTH-1:0] wire_d37_19;
	wire [WIDTH-1:0] wire_d37_20;
	wire [WIDTH-1:0] wire_d37_21;
	wire [WIDTH-1:0] wire_d37_22;
	wire [WIDTH-1:0] wire_d37_23;
	wire [WIDTH-1:0] wire_d37_24;
	wire [WIDTH-1:0] wire_d37_25;
	wire [WIDTH-1:0] wire_d37_26;
	wire [WIDTH-1:0] wire_d37_27;
	wire [WIDTH-1:0] wire_d37_28;
	wire [WIDTH-1:0] wire_d37_29;
	wire [WIDTH-1:0] wire_d37_30;
	wire [WIDTH-1:0] wire_d37_31;
	wire [WIDTH-1:0] wire_d37_32;
	wire [WIDTH-1:0] wire_d37_33;
	wire [WIDTH-1:0] wire_d37_34;
	wire [WIDTH-1:0] wire_d37_35;
	wire [WIDTH-1:0] wire_d37_36;
	wire [WIDTH-1:0] wire_d37_37;
	wire [WIDTH-1:0] wire_d37_38;
	wire [WIDTH-1:0] wire_d37_39;
	wire [WIDTH-1:0] wire_d37_40;
	wire [WIDTH-1:0] wire_d37_41;
	wire [WIDTH-1:0] wire_d37_42;
	wire [WIDTH-1:0] wire_d37_43;
	wire [WIDTH-1:0] wire_d37_44;
	wire [WIDTH-1:0] wire_d37_45;
	wire [WIDTH-1:0] wire_d37_46;
	wire [WIDTH-1:0] wire_d37_47;
	wire [WIDTH-1:0] wire_d37_48;
	wire [WIDTH-1:0] wire_d37_49;
	wire [WIDTH-1:0] wire_d37_50;
	wire [WIDTH-1:0] wire_d37_51;
	wire [WIDTH-1:0] wire_d37_52;
	wire [WIDTH-1:0] wire_d37_53;
	wire [WIDTH-1:0] wire_d37_54;
	wire [WIDTH-1:0] wire_d37_55;
	wire [WIDTH-1:0] wire_d37_56;
	wire [WIDTH-1:0] wire_d37_57;
	wire [WIDTH-1:0] wire_d37_58;
	wire [WIDTH-1:0] wire_d37_59;
	wire [WIDTH-1:0] wire_d37_60;
	wire [WIDTH-1:0] wire_d37_61;
	wire [WIDTH-1:0] wire_d37_62;
	wire [WIDTH-1:0] wire_d37_63;
	wire [WIDTH-1:0] wire_d37_64;
	wire [WIDTH-1:0] wire_d37_65;
	wire [WIDTH-1:0] wire_d37_66;
	wire [WIDTH-1:0] wire_d37_67;
	wire [WIDTH-1:0] wire_d37_68;
	wire [WIDTH-1:0] wire_d37_69;
	wire [WIDTH-1:0] wire_d37_70;
	wire [WIDTH-1:0] wire_d37_71;
	wire [WIDTH-1:0] wire_d37_72;
	wire [WIDTH-1:0] wire_d37_73;
	wire [WIDTH-1:0] wire_d37_74;
	wire [WIDTH-1:0] wire_d37_75;
	wire [WIDTH-1:0] wire_d37_76;
	wire [WIDTH-1:0] wire_d37_77;
	wire [WIDTH-1:0] wire_d37_78;
	wire [WIDTH-1:0] wire_d37_79;
	wire [WIDTH-1:0] wire_d37_80;
	wire [WIDTH-1:0] wire_d37_81;
	wire [WIDTH-1:0] wire_d37_82;
	wire [WIDTH-1:0] wire_d37_83;
	wire [WIDTH-1:0] wire_d37_84;
	wire [WIDTH-1:0] wire_d37_85;
	wire [WIDTH-1:0] wire_d37_86;
	wire [WIDTH-1:0] wire_d37_87;
	wire [WIDTH-1:0] wire_d37_88;
	wire [WIDTH-1:0] wire_d37_89;
	wire [WIDTH-1:0] wire_d37_90;
	wire [WIDTH-1:0] wire_d37_91;
	wire [WIDTH-1:0] wire_d37_92;
	wire [WIDTH-1:0] wire_d37_93;
	wire [WIDTH-1:0] wire_d37_94;
	wire [WIDTH-1:0] wire_d37_95;
	wire [WIDTH-1:0] wire_d37_96;
	wire [WIDTH-1:0] wire_d37_97;
	wire [WIDTH-1:0] wire_d37_98;
	wire [WIDTH-1:0] wire_d37_99;
	wire [WIDTH-1:0] wire_d37_100;
	wire [WIDTH-1:0] wire_d37_101;
	wire [WIDTH-1:0] wire_d37_102;
	wire [WIDTH-1:0] wire_d37_103;
	wire [WIDTH-1:0] wire_d37_104;
	wire [WIDTH-1:0] wire_d37_105;
	wire [WIDTH-1:0] wire_d37_106;
	wire [WIDTH-1:0] wire_d37_107;
	wire [WIDTH-1:0] wire_d37_108;
	wire [WIDTH-1:0] wire_d37_109;
	wire [WIDTH-1:0] wire_d37_110;
	wire [WIDTH-1:0] wire_d37_111;
	wire [WIDTH-1:0] wire_d37_112;
	wire [WIDTH-1:0] wire_d37_113;
	wire [WIDTH-1:0] wire_d37_114;
	wire [WIDTH-1:0] wire_d37_115;
	wire [WIDTH-1:0] wire_d37_116;
	wire [WIDTH-1:0] wire_d37_117;
	wire [WIDTH-1:0] wire_d37_118;
	wire [WIDTH-1:0] wire_d38_0;
	wire [WIDTH-1:0] wire_d38_1;
	wire [WIDTH-1:0] wire_d38_2;
	wire [WIDTH-1:0] wire_d38_3;
	wire [WIDTH-1:0] wire_d38_4;
	wire [WIDTH-1:0] wire_d38_5;
	wire [WIDTH-1:0] wire_d38_6;
	wire [WIDTH-1:0] wire_d38_7;
	wire [WIDTH-1:0] wire_d38_8;
	wire [WIDTH-1:0] wire_d38_9;
	wire [WIDTH-1:0] wire_d38_10;
	wire [WIDTH-1:0] wire_d38_11;
	wire [WIDTH-1:0] wire_d38_12;
	wire [WIDTH-1:0] wire_d38_13;
	wire [WIDTH-1:0] wire_d38_14;
	wire [WIDTH-1:0] wire_d38_15;
	wire [WIDTH-1:0] wire_d38_16;
	wire [WIDTH-1:0] wire_d38_17;
	wire [WIDTH-1:0] wire_d38_18;
	wire [WIDTH-1:0] wire_d38_19;
	wire [WIDTH-1:0] wire_d38_20;
	wire [WIDTH-1:0] wire_d38_21;
	wire [WIDTH-1:0] wire_d38_22;
	wire [WIDTH-1:0] wire_d38_23;
	wire [WIDTH-1:0] wire_d38_24;
	wire [WIDTH-1:0] wire_d38_25;
	wire [WIDTH-1:0] wire_d38_26;
	wire [WIDTH-1:0] wire_d38_27;
	wire [WIDTH-1:0] wire_d38_28;
	wire [WIDTH-1:0] wire_d38_29;
	wire [WIDTH-1:0] wire_d38_30;
	wire [WIDTH-1:0] wire_d38_31;
	wire [WIDTH-1:0] wire_d38_32;
	wire [WIDTH-1:0] wire_d38_33;
	wire [WIDTH-1:0] wire_d38_34;
	wire [WIDTH-1:0] wire_d38_35;
	wire [WIDTH-1:0] wire_d38_36;
	wire [WIDTH-1:0] wire_d38_37;
	wire [WIDTH-1:0] wire_d38_38;
	wire [WIDTH-1:0] wire_d38_39;
	wire [WIDTH-1:0] wire_d38_40;
	wire [WIDTH-1:0] wire_d38_41;
	wire [WIDTH-1:0] wire_d38_42;
	wire [WIDTH-1:0] wire_d38_43;
	wire [WIDTH-1:0] wire_d38_44;
	wire [WIDTH-1:0] wire_d38_45;
	wire [WIDTH-1:0] wire_d38_46;
	wire [WIDTH-1:0] wire_d38_47;
	wire [WIDTH-1:0] wire_d38_48;
	wire [WIDTH-1:0] wire_d38_49;
	wire [WIDTH-1:0] wire_d38_50;
	wire [WIDTH-1:0] wire_d38_51;
	wire [WIDTH-1:0] wire_d38_52;
	wire [WIDTH-1:0] wire_d38_53;
	wire [WIDTH-1:0] wire_d38_54;
	wire [WIDTH-1:0] wire_d38_55;
	wire [WIDTH-1:0] wire_d38_56;
	wire [WIDTH-1:0] wire_d38_57;
	wire [WIDTH-1:0] wire_d38_58;
	wire [WIDTH-1:0] wire_d38_59;
	wire [WIDTH-1:0] wire_d38_60;
	wire [WIDTH-1:0] wire_d38_61;
	wire [WIDTH-1:0] wire_d38_62;
	wire [WIDTH-1:0] wire_d38_63;
	wire [WIDTH-1:0] wire_d38_64;
	wire [WIDTH-1:0] wire_d38_65;
	wire [WIDTH-1:0] wire_d38_66;
	wire [WIDTH-1:0] wire_d38_67;
	wire [WIDTH-1:0] wire_d38_68;
	wire [WIDTH-1:0] wire_d38_69;
	wire [WIDTH-1:0] wire_d38_70;
	wire [WIDTH-1:0] wire_d38_71;
	wire [WIDTH-1:0] wire_d38_72;
	wire [WIDTH-1:0] wire_d38_73;
	wire [WIDTH-1:0] wire_d38_74;
	wire [WIDTH-1:0] wire_d38_75;
	wire [WIDTH-1:0] wire_d38_76;
	wire [WIDTH-1:0] wire_d38_77;
	wire [WIDTH-1:0] wire_d38_78;
	wire [WIDTH-1:0] wire_d38_79;
	wire [WIDTH-1:0] wire_d38_80;
	wire [WIDTH-1:0] wire_d38_81;
	wire [WIDTH-1:0] wire_d38_82;
	wire [WIDTH-1:0] wire_d38_83;
	wire [WIDTH-1:0] wire_d38_84;
	wire [WIDTH-1:0] wire_d38_85;
	wire [WIDTH-1:0] wire_d38_86;
	wire [WIDTH-1:0] wire_d38_87;
	wire [WIDTH-1:0] wire_d38_88;
	wire [WIDTH-1:0] wire_d38_89;
	wire [WIDTH-1:0] wire_d38_90;
	wire [WIDTH-1:0] wire_d38_91;
	wire [WIDTH-1:0] wire_d38_92;
	wire [WIDTH-1:0] wire_d38_93;
	wire [WIDTH-1:0] wire_d38_94;
	wire [WIDTH-1:0] wire_d38_95;
	wire [WIDTH-1:0] wire_d38_96;
	wire [WIDTH-1:0] wire_d38_97;
	wire [WIDTH-1:0] wire_d38_98;
	wire [WIDTH-1:0] wire_d38_99;
	wire [WIDTH-1:0] wire_d38_100;
	wire [WIDTH-1:0] wire_d38_101;
	wire [WIDTH-1:0] wire_d38_102;
	wire [WIDTH-1:0] wire_d38_103;
	wire [WIDTH-1:0] wire_d38_104;
	wire [WIDTH-1:0] wire_d38_105;
	wire [WIDTH-1:0] wire_d38_106;
	wire [WIDTH-1:0] wire_d38_107;
	wire [WIDTH-1:0] wire_d38_108;
	wire [WIDTH-1:0] wire_d38_109;
	wire [WIDTH-1:0] wire_d38_110;
	wire [WIDTH-1:0] wire_d38_111;
	wire [WIDTH-1:0] wire_d38_112;
	wire [WIDTH-1:0] wire_d38_113;
	wire [WIDTH-1:0] wire_d38_114;
	wire [WIDTH-1:0] wire_d38_115;
	wire [WIDTH-1:0] wire_d38_116;
	wire [WIDTH-1:0] wire_d38_117;
	wire [WIDTH-1:0] wire_d38_118;
	wire [WIDTH-1:0] wire_d39_0;
	wire [WIDTH-1:0] wire_d39_1;
	wire [WIDTH-1:0] wire_d39_2;
	wire [WIDTH-1:0] wire_d39_3;
	wire [WIDTH-1:0] wire_d39_4;
	wire [WIDTH-1:0] wire_d39_5;
	wire [WIDTH-1:0] wire_d39_6;
	wire [WIDTH-1:0] wire_d39_7;
	wire [WIDTH-1:0] wire_d39_8;
	wire [WIDTH-1:0] wire_d39_9;
	wire [WIDTH-1:0] wire_d39_10;
	wire [WIDTH-1:0] wire_d39_11;
	wire [WIDTH-1:0] wire_d39_12;
	wire [WIDTH-1:0] wire_d39_13;
	wire [WIDTH-1:0] wire_d39_14;
	wire [WIDTH-1:0] wire_d39_15;
	wire [WIDTH-1:0] wire_d39_16;
	wire [WIDTH-1:0] wire_d39_17;
	wire [WIDTH-1:0] wire_d39_18;
	wire [WIDTH-1:0] wire_d39_19;
	wire [WIDTH-1:0] wire_d39_20;
	wire [WIDTH-1:0] wire_d39_21;
	wire [WIDTH-1:0] wire_d39_22;
	wire [WIDTH-1:0] wire_d39_23;
	wire [WIDTH-1:0] wire_d39_24;
	wire [WIDTH-1:0] wire_d39_25;
	wire [WIDTH-1:0] wire_d39_26;
	wire [WIDTH-1:0] wire_d39_27;
	wire [WIDTH-1:0] wire_d39_28;
	wire [WIDTH-1:0] wire_d39_29;
	wire [WIDTH-1:0] wire_d39_30;
	wire [WIDTH-1:0] wire_d39_31;
	wire [WIDTH-1:0] wire_d39_32;
	wire [WIDTH-1:0] wire_d39_33;
	wire [WIDTH-1:0] wire_d39_34;
	wire [WIDTH-1:0] wire_d39_35;
	wire [WIDTH-1:0] wire_d39_36;
	wire [WIDTH-1:0] wire_d39_37;
	wire [WIDTH-1:0] wire_d39_38;
	wire [WIDTH-1:0] wire_d39_39;
	wire [WIDTH-1:0] wire_d39_40;
	wire [WIDTH-1:0] wire_d39_41;
	wire [WIDTH-1:0] wire_d39_42;
	wire [WIDTH-1:0] wire_d39_43;
	wire [WIDTH-1:0] wire_d39_44;
	wire [WIDTH-1:0] wire_d39_45;
	wire [WIDTH-1:0] wire_d39_46;
	wire [WIDTH-1:0] wire_d39_47;
	wire [WIDTH-1:0] wire_d39_48;
	wire [WIDTH-1:0] wire_d39_49;
	wire [WIDTH-1:0] wire_d39_50;
	wire [WIDTH-1:0] wire_d39_51;
	wire [WIDTH-1:0] wire_d39_52;
	wire [WIDTH-1:0] wire_d39_53;
	wire [WIDTH-1:0] wire_d39_54;
	wire [WIDTH-1:0] wire_d39_55;
	wire [WIDTH-1:0] wire_d39_56;
	wire [WIDTH-1:0] wire_d39_57;
	wire [WIDTH-1:0] wire_d39_58;
	wire [WIDTH-1:0] wire_d39_59;
	wire [WIDTH-1:0] wire_d39_60;
	wire [WIDTH-1:0] wire_d39_61;
	wire [WIDTH-1:0] wire_d39_62;
	wire [WIDTH-1:0] wire_d39_63;
	wire [WIDTH-1:0] wire_d39_64;
	wire [WIDTH-1:0] wire_d39_65;
	wire [WIDTH-1:0] wire_d39_66;
	wire [WIDTH-1:0] wire_d39_67;
	wire [WIDTH-1:0] wire_d39_68;
	wire [WIDTH-1:0] wire_d39_69;
	wire [WIDTH-1:0] wire_d39_70;
	wire [WIDTH-1:0] wire_d39_71;
	wire [WIDTH-1:0] wire_d39_72;
	wire [WIDTH-1:0] wire_d39_73;
	wire [WIDTH-1:0] wire_d39_74;
	wire [WIDTH-1:0] wire_d39_75;
	wire [WIDTH-1:0] wire_d39_76;
	wire [WIDTH-1:0] wire_d39_77;
	wire [WIDTH-1:0] wire_d39_78;
	wire [WIDTH-1:0] wire_d39_79;
	wire [WIDTH-1:0] wire_d39_80;
	wire [WIDTH-1:0] wire_d39_81;
	wire [WIDTH-1:0] wire_d39_82;
	wire [WIDTH-1:0] wire_d39_83;
	wire [WIDTH-1:0] wire_d39_84;
	wire [WIDTH-1:0] wire_d39_85;
	wire [WIDTH-1:0] wire_d39_86;
	wire [WIDTH-1:0] wire_d39_87;
	wire [WIDTH-1:0] wire_d39_88;
	wire [WIDTH-1:0] wire_d39_89;
	wire [WIDTH-1:0] wire_d39_90;
	wire [WIDTH-1:0] wire_d39_91;
	wire [WIDTH-1:0] wire_d39_92;
	wire [WIDTH-1:0] wire_d39_93;
	wire [WIDTH-1:0] wire_d39_94;
	wire [WIDTH-1:0] wire_d39_95;
	wire [WIDTH-1:0] wire_d39_96;
	wire [WIDTH-1:0] wire_d39_97;
	wire [WIDTH-1:0] wire_d39_98;
	wire [WIDTH-1:0] wire_d39_99;
	wire [WIDTH-1:0] wire_d39_100;
	wire [WIDTH-1:0] wire_d39_101;
	wire [WIDTH-1:0] wire_d39_102;
	wire [WIDTH-1:0] wire_d39_103;
	wire [WIDTH-1:0] wire_d39_104;
	wire [WIDTH-1:0] wire_d39_105;
	wire [WIDTH-1:0] wire_d39_106;
	wire [WIDTH-1:0] wire_d39_107;
	wire [WIDTH-1:0] wire_d39_108;
	wire [WIDTH-1:0] wire_d39_109;
	wire [WIDTH-1:0] wire_d39_110;
	wire [WIDTH-1:0] wire_d39_111;
	wire [WIDTH-1:0] wire_d39_112;
	wire [WIDTH-1:0] wire_d39_113;
	wire [WIDTH-1:0] wire_d39_114;
	wire [WIDTH-1:0] wire_d39_115;
	wire [WIDTH-1:0] wire_d39_116;
	wire [WIDTH-1:0] wire_d39_117;
	wire [WIDTH-1:0] wire_d39_118;
	wire [WIDTH-1:0] wire_d40_0;
	wire [WIDTH-1:0] wire_d40_1;
	wire [WIDTH-1:0] wire_d40_2;
	wire [WIDTH-1:0] wire_d40_3;
	wire [WIDTH-1:0] wire_d40_4;
	wire [WIDTH-1:0] wire_d40_5;
	wire [WIDTH-1:0] wire_d40_6;
	wire [WIDTH-1:0] wire_d40_7;
	wire [WIDTH-1:0] wire_d40_8;
	wire [WIDTH-1:0] wire_d40_9;
	wire [WIDTH-1:0] wire_d40_10;
	wire [WIDTH-1:0] wire_d40_11;
	wire [WIDTH-1:0] wire_d40_12;
	wire [WIDTH-1:0] wire_d40_13;
	wire [WIDTH-1:0] wire_d40_14;
	wire [WIDTH-1:0] wire_d40_15;
	wire [WIDTH-1:0] wire_d40_16;
	wire [WIDTH-1:0] wire_d40_17;
	wire [WIDTH-1:0] wire_d40_18;
	wire [WIDTH-1:0] wire_d40_19;
	wire [WIDTH-1:0] wire_d40_20;
	wire [WIDTH-1:0] wire_d40_21;
	wire [WIDTH-1:0] wire_d40_22;
	wire [WIDTH-1:0] wire_d40_23;
	wire [WIDTH-1:0] wire_d40_24;
	wire [WIDTH-1:0] wire_d40_25;
	wire [WIDTH-1:0] wire_d40_26;
	wire [WIDTH-1:0] wire_d40_27;
	wire [WIDTH-1:0] wire_d40_28;
	wire [WIDTH-1:0] wire_d40_29;
	wire [WIDTH-1:0] wire_d40_30;
	wire [WIDTH-1:0] wire_d40_31;
	wire [WIDTH-1:0] wire_d40_32;
	wire [WIDTH-1:0] wire_d40_33;
	wire [WIDTH-1:0] wire_d40_34;
	wire [WIDTH-1:0] wire_d40_35;
	wire [WIDTH-1:0] wire_d40_36;
	wire [WIDTH-1:0] wire_d40_37;
	wire [WIDTH-1:0] wire_d40_38;
	wire [WIDTH-1:0] wire_d40_39;
	wire [WIDTH-1:0] wire_d40_40;
	wire [WIDTH-1:0] wire_d40_41;
	wire [WIDTH-1:0] wire_d40_42;
	wire [WIDTH-1:0] wire_d40_43;
	wire [WIDTH-1:0] wire_d40_44;
	wire [WIDTH-1:0] wire_d40_45;
	wire [WIDTH-1:0] wire_d40_46;
	wire [WIDTH-1:0] wire_d40_47;
	wire [WIDTH-1:0] wire_d40_48;
	wire [WIDTH-1:0] wire_d40_49;
	wire [WIDTH-1:0] wire_d40_50;
	wire [WIDTH-1:0] wire_d40_51;
	wire [WIDTH-1:0] wire_d40_52;
	wire [WIDTH-1:0] wire_d40_53;
	wire [WIDTH-1:0] wire_d40_54;
	wire [WIDTH-1:0] wire_d40_55;
	wire [WIDTH-1:0] wire_d40_56;
	wire [WIDTH-1:0] wire_d40_57;
	wire [WIDTH-1:0] wire_d40_58;
	wire [WIDTH-1:0] wire_d40_59;
	wire [WIDTH-1:0] wire_d40_60;
	wire [WIDTH-1:0] wire_d40_61;
	wire [WIDTH-1:0] wire_d40_62;
	wire [WIDTH-1:0] wire_d40_63;
	wire [WIDTH-1:0] wire_d40_64;
	wire [WIDTH-1:0] wire_d40_65;
	wire [WIDTH-1:0] wire_d40_66;
	wire [WIDTH-1:0] wire_d40_67;
	wire [WIDTH-1:0] wire_d40_68;
	wire [WIDTH-1:0] wire_d40_69;
	wire [WIDTH-1:0] wire_d40_70;
	wire [WIDTH-1:0] wire_d40_71;
	wire [WIDTH-1:0] wire_d40_72;
	wire [WIDTH-1:0] wire_d40_73;
	wire [WIDTH-1:0] wire_d40_74;
	wire [WIDTH-1:0] wire_d40_75;
	wire [WIDTH-1:0] wire_d40_76;
	wire [WIDTH-1:0] wire_d40_77;
	wire [WIDTH-1:0] wire_d40_78;
	wire [WIDTH-1:0] wire_d40_79;
	wire [WIDTH-1:0] wire_d40_80;
	wire [WIDTH-1:0] wire_d40_81;
	wire [WIDTH-1:0] wire_d40_82;
	wire [WIDTH-1:0] wire_d40_83;
	wire [WIDTH-1:0] wire_d40_84;
	wire [WIDTH-1:0] wire_d40_85;
	wire [WIDTH-1:0] wire_d40_86;
	wire [WIDTH-1:0] wire_d40_87;
	wire [WIDTH-1:0] wire_d40_88;
	wire [WIDTH-1:0] wire_d40_89;
	wire [WIDTH-1:0] wire_d40_90;
	wire [WIDTH-1:0] wire_d40_91;
	wire [WIDTH-1:0] wire_d40_92;
	wire [WIDTH-1:0] wire_d40_93;
	wire [WIDTH-1:0] wire_d40_94;
	wire [WIDTH-1:0] wire_d40_95;
	wire [WIDTH-1:0] wire_d40_96;
	wire [WIDTH-1:0] wire_d40_97;
	wire [WIDTH-1:0] wire_d40_98;
	wire [WIDTH-1:0] wire_d40_99;
	wire [WIDTH-1:0] wire_d40_100;
	wire [WIDTH-1:0] wire_d40_101;
	wire [WIDTH-1:0] wire_d40_102;
	wire [WIDTH-1:0] wire_d40_103;
	wire [WIDTH-1:0] wire_d40_104;
	wire [WIDTH-1:0] wire_d40_105;
	wire [WIDTH-1:0] wire_d40_106;
	wire [WIDTH-1:0] wire_d40_107;
	wire [WIDTH-1:0] wire_d40_108;
	wire [WIDTH-1:0] wire_d40_109;
	wire [WIDTH-1:0] wire_d40_110;
	wire [WIDTH-1:0] wire_d40_111;
	wire [WIDTH-1:0] wire_d40_112;
	wire [WIDTH-1:0] wire_d40_113;
	wire [WIDTH-1:0] wire_d40_114;
	wire [WIDTH-1:0] wire_d40_115;
	wire [WIDTH-1:0] wire_d40_116;
	wire [WIDTH-1:0] wire_d40_117;
	wire [WIDTH-1:0] wire_d40_118;
	wire [WIDTH-1:0] wire_d41_0;
	wire [WIDTH-1:0] wire_d41_1;
	wire [WIDTH-1:0] wire_d41_2;
	wire [WIDTH-1:0] wire_d41_3;
	wire [WIDTH-1:0] wire_d41_4;
	wire [WIDTH-1:0] wire_d41_5;
	wire [WIDTH-1:0] wire_d41_6;
	wire [WIDTH-1:0] wire_d41_7;
	wire [WIDTH-1:0] wire_d41_8;
	wire [WIDTH-1:0] wire_d41_9;
	wire [WIDTH-1:0] wire_d41_10;
	wire [WIDTH-1:0] wire_d41_11;
	wire [WIDTH-1:0] wire_d41_12;
	wire [WIDTH-1:0] wire_d41_13;
	wire [WIDTH-1:0] wire_d41_14;
	wire [WIDTH-1:0] wire_d41_15;
	wire [WIDTH-1:0] wire_d41_16;
	wire [WIDTH-1:0] wire_d41_17;
	wire [WIDTH-1:0] wire_d41_18;
	wire [WIDTH-1:0] wire_d41_19;
	wire [WIDTH-1:0] wire_d41_20;
	wire [WIDTH-1:0] wire_d41_21;
	wire [WIDTH-1:0] wire_d41_22;
	wire [WIDTH-1:0] wire_d41_23;
	wire [WIDTH-1:0] wire_d41_24;
	wire [WIDTH-1:0] wire_d41_25;
	wire [WIDTH-1:0] wire_d41_26;
	wire [WIDTH-1:0] wire_d41_27;
	wire [WIDTH-1:0] wire_d41_28;
	wire [WIDTH-1:0] wire_d41_29;
	wire [WIDTH-1:0] wire_d41_30;
	wire [WIDTH-1:0] wire_d41_31;
	wire [WIDTH-1:0] wire_d41_32;
	wire [WIDTH-1:0] wire_d41_33;
	wire [WIDTH-1:0] wire_d41_34;
	wire [WIDTH-1:0] wire_d41_35;
	wire [WIDTH-1:0] wire_d41_36;
	wire [WIDTH-1:0] wire_d41_37;
	wire [WIDTH-1:0] wire_d41_38;
	wire [WIDTH-1:0] wire_d41_39;
	wire [WIDTH-1:0] wire_d41_40;
	wire [WIDTH-1:0] wire_d41_41;
	wire [WIDTH-1:0] wire_d41_42;
	wire [WIDTH-1:0] wire_d41_43;
	wire [WIDTH-1:0] wire_d41_44;
	wire [WIDTH-1:0] wire_d41_45;
	wire [WIDTH-1:0] wire_d41_46;
	wire [WIDTH-1:0] wire_d41_47;
	wire [WIDTH-1:0] wire_d41_48;
	wire [WIDTH-1:0] wire_d41_49;
	wire [WIDTH-1:0] wire_d41_50;
	wire [WIDTH-1:0] wire_d41_51;
	wire [WIDTH-1:0] wire_d41_52;
	wire [WIDTH-1:0] wire_d41_53;
	wire [WIDTH-1:0] wire_d41_54;
	wire [WIDTH-1:0] wire_d41_55;
	wire [WIDTH-1:0] wire_d41_56;
	wire [WIDTH-1:0] wire_d41_57;
	wire [WIDTH-1:0] wire_d41_58;
	wire [WIDTH-1:0] wire_d41_59;
	wire [WIDTH-1:0] wire_d41_60;
	wire [WIDTH-1:0] wire_d41_61;
	wire [WIDTH-1:0] wire_d41_62;
	wire [WIDTH-1:0] wire_d41_63;
	wire [WIDTH-1:0] wire_d41_64;
	wire [WIDTH-1:0] wire_d41_65;
	wire [WIDTH-1:0] wire_d41_66;
	wire [WIDTH-1:0] wire_d41_67;
	wire [WIDTH-1:0] wire_d41_68;
	wire [WIDTH-1:0] wire_d41_69;
	wire [WIDTH-1:0] wire_d41_70;
	wire [WIDTH-1:0] wire_d41_71;
	wire [WIDTH-1:0] wire_d41_72;
	wire [WIDTH-1:0] wire_d41_73;
	wire [WIDTH-1:0] wire_d41_74;
	wire [WIDTH-1:0] wire_d41_75;
	wire [WIDTH-1:0] wire_d41_76;
	wire [WIDTH-1:0] wire_d41_77;
	wire [WIDTH-1:0] wire_d41_78;
	wire [WIDTH-1:0] wire_d41_79;
	wire [WIDTH-1:0] wire_d41_80;
	wire [WIDTH-1:0] wire_d41_81;
	wire [WIDTH-1:0] wire_d41_82;
	wire [WIDTH-1:0] wire_d41_83;
	wire [WIDTH-1:0] wire_d41_84;
	wire [WIDTH-1:0] wire_d41_85;
	wire [WIDTH-1:0] wire_d41_86;
	wire [WIDTH-1:0] wire_d41_87;
	wire [WIDTH-1:0] wire_d41_88;
	wire [WIDTH-1:0] wire_d41_89;
	wire [WIDTH-1:0] wire_d41_90;
	wire [WIDTH-1:0] wire_d41_91;
	wire [WIDTH-1:0] wire_d41_92;
	wire [WIDTH-1:0] wire_d41_93;
	wire [WIDTH-1:0] wire_d41_94;
	wire [WIDTH-1:0] wire_d41_95;
	wire [WIDTH-1:0] wire_d41_96;
	wire [WIDTH-1:0] wire_d41_97;
	wire [WIDTH-1:0] wire_d41_98;
	wire [WIDTH-1:0] wire_d41_99;
	wire [WIDTH-1:0] wire_d41_100;
	wire [WIDTH-1:0] wire_d41_101;
	wire [WIDTH-1:0] wire_d41_102;
	wire [WIDTH-1:0] wire_d41_103;
	wire [WIDTH-1:0] wire_d41_104;
	wire [WIDTH-1:0] wire_d41_105;
	wire [WIDTH-1:0] wire_d41_106;
	wire [WIDTH-1:0] wire_d41_107;
	wire [WIDTH-1:0] wire_d41_108;
	wire [WIDTH-1:0] wire_d41_109;
	wire [WIDTH-1:0] wire_d41_110;
	wire [WIDTH-1:0] wire_d41_111;
	wire [WIDTH-1:0] wire_d41_112;
	wire [WIDTH-1:0] wire_d41_113;
	wire [WIDTH-1:0] wire_d41_114;
	wire [WIDTH-1:0] wire_d41_115;
	wire [WIDTH-1:0] wire_d41_116;
	wire [WIDTH-1:0] wire_d41_117;
	wire [WIDTH-1:0] wire_d41_118;
	wire [WIDTH-1:0] wire_d42_0;
	wire [WIDTH-1:0] wire_d42_1;
	wire [WIDTH-1:0] wire_d42_2;
	wire [WIDTH-1:0] wire_d42_3;
	wire [WIDTH-1:0] wire_d42_4;
	wire [WIDTH-1:0] wire_d42_5;
	wire [WIDTH-1:0] wire_d42_6;
	wire [WIDTH-1:0] wire_d42_7;
	wire [WIDTH-1:0] wire_d42_8;
	wire [WIDTH-1:0] wire_d42_9;
	wire [WIDTH-1:0] wire_d42_10;
	wire [WIDTH-1:0] wire_d42_11;
	wire [WIDTH-1:0] wire_d42_12;
	wire [WIDTH-1:0] wire_d42_13;
	wire [WIDTH-1:0] wire_d42_14;
	wire [WIDTH-1:0] wire_d42_15;
	wire [WIDTH-1:0] wire_d42_16;
	wire [WIDTH-1:0] wire_d42_17;
	wire [WIDTH-1:0] wire_d42_18;
	wire [WIDTH-1:0] wire_d42_19;
	wire [WIDTH-1:0] wire_d42_20;
	wire [WIDTH-1:0] wire_d42_21;
	wire [WIDTH-1:0] wire_d42_22;
	wire [WIDTH-1:0] wire_d42_23;
	wire [WIDTH-1:0] wire_d42_24;
	wire [WIDTH-1:0] wire_d42_25;
	wire [WIDTH-1:0] wire_d42_26;
	wire [WIDTH-1:0] wire_d42_27;
	wire [WIDTH-1:0] wire_d42_28;
	wire [WIDTH-1:0] wire_d42_29;
	wire [WIDTH-1:0] wire_d42_30;
	wire [WIDTH-1:0] wire_d42_31;
	wire [WIDTH-1:0] wire_d42_32;
	wire [WIDTH-1:0] wire_d42_33;
	wire [WIDTH-1:0] wire_d42_34;
	wire [WIDTH-1:0] wire_d42_35;
	wire [WIDTH-1:0] wire_d42_36;
	wire [WIDTH-1:0] wire_d42_37;
	wire [WIDTH-1:0] wire_d42_38;
	wire [WIDTH-1:0] wire_d42_39;
	wire [WIDTH-1:0] wire_d42_40;
	wire [WIDTH-1:0] wire_d42_41;
	wire [WIDTH-1:0] wire_d42_42;
	wire [WIDTH-1:0] wire_d42_43;
	wire [WIDTH-1:0] wire_d42_44;
	wire [WIDTH-1:0] wire_d42_45;
	wire [WIDTH-1:0] wire_d42_46;
	wire [WIDTH-1:0] wire_d42_47;
	wire [WIDTH-1:0] wire_d42_48;
	wire [WIDTH-1:0] wire_d42_49;
	wire [WIDTH-1:0] wire_d42_50;
	wire [WIDTH-1:0] wire_d42_51;
	wire [WIDTH-1:0] wire_d42_52;
	wire [WIDTH-1:0] wire_d42_53;
	wire [WIDTH-1:0] wire_d42_54;
	wire [WIDTH-1:0] wire_d42_55;
	wire [WIDTH-1:0] wire_d42_56;
	wire [WIDTH-1:0] wire_d42_57;
	wire [WIDTH-1:0] wire_d42_58;
	wire [WIDTH-1:0] wire_d42_59;
	wire [WIDTH-1:0] wire_d42_60;
	wire [WIDTH-1:0] wire_d42_61;
	wire [WIDTH-1:0] wire_d42_62;
	wire [WIDTH-1:0] wire_d42_63;
	wire [WIDTH-1:0] wire_d42_64;
	wire [WIDTH-1:0] wire_d42_65;
	wire [WIDTH-1:0] wire_d42_66;
	wire [WIDTH-1:0] wire_d42_67;
	wire [WIDTH-1:0] wire_d42_68;
	wire [WIDTH-1:0] wire_d42_69;
	wire [WIDTH-1:0] wire_d42_70;
	wire [WIDTH-1:0] wire_d42_71;
	wire [WIDTH-1:0] wire_d42_72;
	wire [WIDTH-1:0] wire_d42_73;
	wire [WIDTH-1:0] wire_d42_74;
	wire [WIDTH-1:0] wire_d42_75;
	wire [WIDTH-1:0] wire_d42_76;
	wire [WIDTH-1:0] wire_d42_77;
	wire [WIDTH-1:0] wire_d42_78;
	wire [WIDTH-1:0] wire_d42_79;
	wire [WIDTH-1:0] wire_d42_80;
	wire [WIDTH-1:0] wire_d42_81;
	wire [WIDTH-1:0] wire_d42_82;
	wire [WIDTH-1:0] wire_d42_83;
	wire [WIDTH-1:0] wire_d42_84;
	wire [WIDTH-1:0] wire_d42_85;
	wire [WIDTH-1:0] wire_d42_86;
	wire [WIDTH-1:0] wire_d42_87;
	wire [WIDTH-1:0] wire_d42_88;
	wire [WIDTH-1:0] wire_d42_89;
	wire [WIDTH-1:0] wire_d42_90;
	wire [WIDTH-1:0] wire_d42_91;
	wire [WIDTH-1:0] wire_d42_92;
	wire [WIDTH-1:0] wire_d42_93;
	wire [WIDTH-1:0] wire_d42_94;
	wire [WIDTH-1:0] wire_d42_95;
	wire [WIDTH-1:0] wire_d42_96;
	wire [WIDTH-1:0] wire_d42_97;
	wire [WIDTH-1:0] wire_d42_98;
	wire [WIDTH-1:0] wire_d42_99;
	wire [WIDTH-1:0] wire_d42_100;
	wire [WIDTH-1:0] wire_d42_101;
	wire [WIDTH-1:0] wire_d42_102;
	wire [WIDTH-1:0] wire_d42_103;
	wire [WIDTH-1:0] wire_d42_104;
	wire [WIDTH-1:0] wire_d42_105;
	wire [WIDTH-1:0] wire_d42_106;
	wire [WIDTH-1:0] wire_d42_107;
	wire [WIDTH-1:0] wire_d42_108;
	wire [WIDTH-1:0] wire_d42_109;
	wire [WIDTH-1:0] wire_d42_110;
	wire [WIDTH-1:0] wire_d42_111;
	wire [WIDTH-1:0] wire_d42_112;
	wire [WIDTH-1:0] wire_d42_113;
	wire [WIDTH-1:0] wire_d42_114;
	wire [WIDTH-1:0] wire_d42_115;
	wire [WIDTH-1:0] wire_d42_116;
	wire [WIDTH-1:0] wire_d42_117;
	wire [WIDTH-1:0] wire_d42_118;
	wire [WIDTH-1:0] wire_d43_0;
	wire [WIDTH-1:0] wire_d43_1;
	wire [WIDTH-1:0] wire_d43_2;
	wire [WIDTH-1:0] wire_d43_3;
	wire [WIDTH-1:0] wire_d43_4;
	wire [WIDTH-1:0] wire_d43_5;
	wire [WIDTH-1:0] wire_d43_6;
	wire [WIDTH-1:0] wire_d43_7;
	wire [WIDTH-1:0] wire_d43_8;
	wire [WIDTH-1:0] wire_d43_9;
	wire [WIDTH-1:0] wire_d43_10;
	wire [WIDTH-1:0] wire_d43_11;
	wire [WIDTH-1:0] wire_d43_12;
	wire [WIDTH-1:0] wire_d43_13;
	wire [WIDTH-1:0] wire_d43_14;
	wire [WIDTH-1:0] wire_d43_15;
	wire [WIDTH-1:0] wire_d43_16;
	wire [WIDTH-1:0] wire_d43_17;
	wire [WIDTH-1:0] wire_d43_18;
	wire [WIDTH-1:0] wire_d43_19;
	wire [WIDTH-1:0] wire_d43_20;
	wire [WIDTH-1:0] wire_d43_21;
	wire [WIDTH-1:0] wire_d43_22;
	wire [WIDTH-1:0] wire_d43_23;
	wire [WIDTH-1:0] wire_d43_24;
	wire [WIDTH-1:0] wire_d43_25;
	wire [WIDTH-1:0] wire_d43_26;
	wire [WIDTH-1:0] wire_d43_27;
	wire [WIDTH-1:0] wire_d43_28;
	wire [WIDTH-1:0] wire_d43_29;
	wire [WIDTH-1:0] wire_d43_30;
	wire [WIDTH-1:0] wire_d43_31;
	wire [WIDTH-1:0] wire_d43_32;
	wire [WIDTH-1:0] wire_d43_33;
	wire [WIDTH-1:0] wire_d43_34;
	wire [WIDTH-1:0] wire_d43_35;
	wire [WIDTH-1:0] wire_d43_36;
	wire [WIDTH-1:0] wire_d43_37;
	wire [WIDTH-1:0] wire_d43_38;
	wire [WIDTH-1:0] wire_d43_39;
	wire [WIDTH-1:0] wire_d43_40;
	wire [WIDTH-1:0] wire_d43_41;
	wire [WIDTH-1:0] wire_d43_42;
	wire [WIDTH-1:0] wire_d43_43;
	wire [WIDTH-1:0] wire_d43_44;
	wire [WIDTH-1:0] wire_d43_45;
	wire [WIDTH-1:0] wire_d43_46;
	wire [WIDTH-1:0] wire_d43_47;
	wire [WIDTH-1:0] wire_d43_48;
	wire [WIDTH-1:0] wire_d43_49;
	wire [WIDTH-1:0] wire_d43_50;
	wire [WIDTH-1:0] wire_d43_51;
	wire [WIDTH-1:0] wire_d43_52;
	wire [WIDTH-1:0] wire_d43_53;
	wire [WIDTH-1:0] wire_d43_54;
	wire [WIDTH-1:0] wire_d43_55;
	wire [WIDTH-1:0] wire_d43_56;
	wire [WIDTH-1:0] wire_d43_57;
	wire [WIDTH-1:0] wire_d43_58;
	wire [WIDTH-1:0] wire_d43_59;
	wire [WIDTH-1:0] wire_d43_60;
	wire [WIDTH-1:0] wire_d43_61;
	wire [WIDTH-1:0] wire_d43_62;
	wire [WIDTH-1:0] wire_d43_63;
	wire [WIDTH-1:0] wire_d43_64;
	wire [WIDTH-1:0] wire_d43_65;
	wire [WIDTH-1:0] wire_d43_66;
	wire [WIDTH-1:0] wire_d43_67;
	wire [WIDTH-1:0] wire_d43_68;
	wire [WIDTH-1:0] wire_d43_69;
	wire [WIDTH-1:0] wire_d43_70;
	wire [WIDTH-1:0] wire_d43_71;
	wire [WIDTH-1:0] wire_d43_72;
	wire [WIDTH-1:0] wire_d43_73;
	wire [WIDTH-1:0] wire_d43_74;
	wire [WIDTH-1:0] wire_d43_75;
	wire [WIDTH-1:0] wire_d43_76;
	wire [WIDTH-1:0] wire_d43_77;
	wire [WIDTH-1:0] wire_d43_78;
	wire [WIDTH-1:0] wire_d43_79;
	wire [WIDTH-1:0] wire_d43_80;
	wire [WIDTH-1:0] wire_d43_81;
	wire [WIDTH-1:0] wire_d43_82;
	wire [WIDTH-1:0] wire_d43_83;
	wire [WIDTH-1:0] wire_d43_84;
	wire [WIDTH-1:0] wire_d43_85;
	wire [WIDTH-1:0] wire_d43_86;
	wire [WIDTH-1:0] wire_d43_87;
	wire [WIDTH-1:0] wire_d43_88;
	wire [WIDTH-1:0] wire_d43_89;
	wire [WIDTH-1:0] wire_d43_90;
	wire [WIDTH-1:0] wire_d43_91;
	wire [WIDTH-1:0] wire_d43_92;
	wire [WIDTH-1:0] wire_d43_93;
	wire [WIDTH-1:0] wire_d43_94;
	wire [WIDTH-1:0] wire_d43_95;
	wire [WIDTH-1:0] wire_d43_96;
	wire [WIDTH-1:0] wire_d43_97;
	wire [WIDTH-1:0] wire_d43_98;
	wire [WIDTH-1:0] wire_d43_99;
	wire [WIDTH-1:0] wire_d43_100;
	wire [WIDTH-1:0] wire_d43_101;
	wire [WIDTH-1:0] wire_d43_102;
	wire [WIDTH-1:0] wire_d43_103;
	wire [WIDTH-1:0] wire_d43_104;
	wire [WIDTH-1:0] wire_d43_105;
	wire [WIDTH-1:0] wire_d43_106;
	wire [WIDTH-1:0] wire_d43_107;
	wire [WIDTH-1:0] wire_d43_108;
	wire [WIDTH-1:0] wire_d43_109;
	wire [WIDTH-1:0] wire_d43_110;
	wire [WIDTH-1:0] wire_d43_111;
	wire [WIDTH-1:0] wire_d43_112;
	wire [WIDTH-1:0] wire_d43_113;
	wire [WIDTH-1:0] wire_d43_114;
	wire [WIDTH-1:0] wire_d43_115;
	wire [WIDTH-1:0] wire_d43_116;
	wire [WIDTH-1:0] wire_d43_117;
	wire [WIDTH-1:0] wire_d43_118;
	wire [WIDTH-1:0] wire_d44_0;
	wire [WIDTH-1:0] wire_d44_1;
	wire [WIDTH-1:0] wire_d44_2;
	wire [WIDTH-1:0] wire_d44_3;
	wire [WIDTH-1:0] wire_d44_4;
	wire [WIDTH-1:0] wire_d44_5;
	wire [WIDTH-1:0] wire_d44_6;
	wire [WIDTH-1:0] wire_d44_7;
	wire [WIDTH-1:0] wire_d44_8;
	wire [WIDTH-1:0] wire_d44_9;
	wire [WIDTH-1:0] wire_d44_10;
	wire [WIDTH-1:0] wire_d44_11;
	wire [WIDTH-1:0] wire_d44_12;
	wire [WIDTH-1:0] wire_d44_13;
	wire [WIDTH-1:0] wire_d44_14;
	wire [WIDTH-1:0] wire_d44_15;
	wire [WIDTH-1:0] wire_d44_16;
	wire [WIDTH-1:0] wire_d44_17;
	wire [WIDTH-1:0] wire_d44_18;
	wire [WIDTH-1:0] wire_d44_19;
	wire [WIDTH-1:0] wire_d44_20;
	wire [WIDTH-1:0] wire_d44_21;
	wire [WIDTH-1:0] wire_d44_22;
	wire [WIDTH-1:0] wire_d44_23;
	wire [WIDTH-1:0] wire_d44_24;
	wire [WIDTH-1:0] wire_d44_25;
	wire [WIDTH-1:0] wire_d44_26;
	wire [WIDTH-1:0] wire_d44_27;
	wire [WIDTH-1:0] wire_d44_28;
	wire [WIDTH-1:0] wire_d44_29;
	wire [WIDTH-1:0] wire_d44_30;
	wire [WIDTH-1:0] wire_d44_31;
	wire [WIDTH-1:0] wire_d44_32;
	wire [WIDTH-1:0] wire_d44_33;
	wire [WIDTH-1:0] wire_d44_34;
	wire [WIDTH-1:0] wire_d44_35;
	wire [WIDTH-1:0] wire_d44_36;
	wire [WIDTH-1:0] wire_d44_37;
	wire [WIDTH-1:0] wire_d44_38;
	wire [WIDTH-1:0] wire_d44_39;
	wire [WIDTH-1:0] wire_d44_40;
	wire [WIDTH-1:0] wire_d44_41;
	wire [WIDTH-1:0] wire_d44_42;
	wire [WIDTH-1:0] wire_d44_43;
	wire [WIDTH-1:0] wire_d44_44;
	wire [WIDTH-1:0] wire_d44_45;
	wire [WIDTH-1:0] wire_d44_46;
	wire [WIDTH-1:0] wire_d44_47;
	wire [WIDTH-1:0] wire_d44_48;
	wire [WIDTH-1:0] wire_d44_49;
	wire [WIDTH-1:0] wire_d44_50;
	wire [WIDTH-1:0] wire_d44_51;
	wire [WIDTH-1:0] wire_d44_52;
	wire [WIDTH-1:0] wire_d44_53;
	wire [WIDTH-1:0] wire_d44_54;
	wire [WIDTH-1:0] wire_d44_55;
	wire [WIDTH-1:0] wire_d44_56;
	wire [WIDTH-1:0] wire_d44_57;
	wire [WIDTH-1:0] wire_d44_58;
	wire [WIDTH-1:0] wire_d44_59;
	wire [WIDTH-1:0] wire_d44_60;
	wire [WIDTH-1:0] wire_d44_61;
	wire [WIDTH-1:0] wire_d44_62;
	wire [WIDTH-1:0] wire_d44_63;
	wire [WIDTH-1:0] wire_d44_64;
	wire [WIDTH-1:0] wire_d44_65;
	wire [WIDTH-1:0] wire_d44_66;
	wire [WIDTH-1:0] wire_d44_67;
	wire [WIDTH-1:0] wire_d44_68;
	wire [WIDTH-1:0] wire_d44_69;
	wire [WIDTH-1:0] wire_d44_70;
	wire [WIDTH-1:0] wire_d44_71;
	wire [WIDTH-1:0] wire_d44_72;
	wire [WIDTH-1:0] wire_d44_73;
	wire [WIDTH-1:0] wire_d44_74;
	wire [WIDTH-1:0] wire_d44_75;
	wire [WIDTH-1:0] wire_d44_76;
	wire [WIDTH-1:0] wire_d44_77;
	wire [WIDTH-1:0] wire_d44_78;
	wire [WIDTH-1:0] wire_d44_79;
	wire [WIDTH-1:0] wire_d44_80;
	wire [WIDTH-1:0] wire_d44_81;
	wire [WIDTH-1:0] wire_d44_82;
	wire [WIDTH-1:0] wire_d44_83;
	wire [WIDTH-1:0] wire_d44_84;
	wire [WIDTH-1:0] wire_d44_85;
	wire [WIDTH-1:0] wire_d44_86;
	wire [WIDTH-1:0] wire_d44_87;
	wire [WIDTH-1:0] wire_d44_88;
	wire [WIDTH-1:0] wire_d44_89;
	wire [WIDTH-1:0] wire_d44_90;
	wire [WIDTH-1:0] wire_d44_91;
	wire [WIDTH-1:0] wire_d44_92;
	wire [WIDTH-1:0] wire_d44_93;
	wire [WIDTH-1:0] wire_d44_94;
	wire [WIDTH-1:0] wire_d44_95;
	wire [WIDTH-1:0] wire_d44_96;
	wire [WIDTH-1:0] wire_d44_97;
	wire [WIDTH-1:0] wire_d44_98;
	wire [WIDTH-1:0] wire_d44_99;
	wire [WIDTH-1:0] wire_d44_100;
	wire [WIDTH-1:0] wire_d44_101;
	wire [WIDTH-1:0] wire_d44_102;
	wire [WIDTH-1:0] wire_d44_103;
	wire [WIDTH-1:0] wire_d44_104;
	wire [WIDTH-1:0] wire_d44_105;
	wire [WIDTH-1:0] wire_d44_106;
	wire [WIDTH-1:0] wire_d44_107;
	wire [WIDTH-1:0] wire_d44_108;
	wire [WIDTH-1:0] wire_d44_109;
	wire [WIDTH-1:0] wire_d44_110;
	wire [WIDTH-1:0] wire_d44_111;
	wire [WIDTH-1:0] wire_d44_112;
	wire [WIDTH-1:0] wire_d44_113;
	wire [WIDTH-1:0] wire_d44_114;
	wire [WIDTH-1:0] wire_d44_115;
	wire [WIDTH-1:0] wire_d44_116;
	wire [WIDTH-1:0] wire_d44_117;
	wire [WIDTH-1:0] wire_d44_118;
	wire [WIDTH-1:0] wire_d45_0;
	wire [WIDTH-1:0] wire_d45_1;
	wire [WIDTH-1:0] wire_d45_2;
	wire [WIDTH-1:0] wire_d45_3;
	wire [WIDTH-1:0] wire_d45_4;
	wire [WIDTH-1:0] wire_d45_5;
	wire [WIDTH-1:0] wire_d45_6;
	wire [WIDTH-1:0] wire_d45_7;
	wire [WIDTH-1:0] wire_d45_8;
	wire [WIDTH-1:0] wire_d45_9;
	wire [WIDTH-1:0] wire_d45_10;
	wire [WIDTH-1:0] wire_d45_11;
	wire [WIDTH-1:0] wire_d45_12;
	wire [WIDTH-1:0] wire_d45_13;
	wire [WIDTH-1:0] wire_d45_14;
	wire [WIDTH-1:0] wire_d45_15;
	wire [WIDTH-1:0] wire_d45_16;
	wire [WIDTH-1:0] wire_d45_17;
	wire [WIDTH-1:0] wire_d45_18;
	wire [WIDTH-1:0] wire_d45_19;
	wire [WIDTH-1:0] wire_d45_20;
	wire [WIDTH-1:0] wire_d45_21;
	wire [WIDTH-1:0] wire_d45_22;
	wire [WIDTH-1:0] wire_d45_23;
	wire [WIDTH-1:0] wire_d45_24;
	wire [WIDTH-1:0] wire_d45_25;
	wire [WIDTH-1:0] wire_d45_26;
	wire [WIDTH-1:0] wire_d45_27;
	wire [WIDTH-1:0] wire_d45_28;
	wire [WIDTH-1:0] wire_d45_29;
	wire [WIDTH-1:0] wire_d45_30;
	wire [WIDTH-1:0] wire_d45_31;
	wire [WIDTH-1:0] wire_d45_32;
	wire [WIDTH-1:0] wire_d45_33;
	wire [WIDTH-1:0] wire_d45_34;
	wire [WIDTH-1:0] wire_d45_35;
	wire [WIDTH-1:0] wire_d45_36;
	wire [WIDTH-1:0] wire_d45_37;
	wire [WIDTH-1:0] wire_d45_38;
	wire [WIDTH-1:0] wire_d45_39;
	wire [WIDTH-1:0] wire_d45_40;
	wire [WIDTH-1:0] wire_d45_41;
	wire [WIDTH-1:0] wire_d45_42;
	wire [WIDTH-1:0] wire_d45_43;
	wire [WIDTH-1:0] wire_d45_44;
	wire [WIDTH-1:0] wire_d45_45;
	wire [WIDTH-1:0] wire_d45_46;
	wire [WIDTH-1:0] wire_d45_47;
	wire [WIDTH-1:0] wire_d45_48;
	wire [WIDTH-1:0] wire_d45_49;
	wire [WIDTH-1:0] wire_d45_50;
	wire [WIDTH-1:0] wire_d45_51;
	wire [WIDTH-1:0] wire_d45_52;
	wire [WIDTH-1:0] wire_d45_53;
	wire [WIDTH-1:0] wire_d45_54;
	wire [WIDTH-1:0] wire_d45_55;
	wire [WIDTH-1:0] wire_d45_56;
	wire [WIDTH-1:0] wire_d45_57;
	wire [WIDTH-1:0] wire_d45_58;
	wire [WIDTH-1:0] wire_d45_59;
	wire [WIDTH-1:0] wire_d45_60;
	wire [WIDTH-1:0] wire_d45_61;
	wire [WIDTH-1:0] wire_d45_62;
	wire [WIDTH-1:0] wire_d45_63;
	wire [WIDTH-1:0] wire_d45_64;
	wire [WIDTH-1:0] wire_d45_65;
	wire [WIDTH-1:0] wire_d45_66;
	wire [WIDTH-1:0] wire_d45_67;
	wire [WIDTH-1:0] wire_d45_68;
	wire [WIDTH-1:0] wire_d45_69;
	wire [WIDTH-1:0] wire_d45_70;
	wire [WIDTH-1:0] wire_d45_71;
	wire [WIDTH-1:0] wire_d45_72;
	wire [WIDTH-1:0] wire_d45_73;
	wire [WIDTH-1:0] wire_d45_74;
	wire [WIDTH-1:0] wire_d45_75;
	wire [WIDTH-1:0] wire_d45_76;
	wire [WIDTH-1:0] wire_d45_77;
	wire [WIDTH-1:0] wire_d45_78;
	wire [WIDTH-1:0] wire_d45_79;
	wire [WIDTH-1:0] wire_d45_80;
	wire [WIDTH-1:0] wire_d45_81;
	wire [WIDTH-1:0] wire_d45_82;
	wire [WIDTH-1:0] wire_d45_83;
	wire [WIDTH-1:0] wire_d45_84;
	wire [WIDTH-1:0] wire_d45_85;
	wire [WIDTH-1:0] wire_d45_86;
	wire [WIDTH-1:0] wire_d45_87;
	wire [WIDTH-1:0] wire_d45_88;
	wire [WIDTH-1:0] wire_d45_89;
	wire [WIDTH-1:0] wire_d45_90;
	wire [WIDTH-1:0] wire_d45_91;
	wire [WIDTH-1:0] wire_d45_92;
	wire [WIDTH-1:0] wire_d45_93;
	wire [WIDTH-1:0] wire_d45_94;
	wire [WIDTH-1:0] wire_d45_95;
	wire [WIDTH-1:0] wire_d45_96;
	wire [WIDTH-1:0] wire_d45_97;
	wire [WIDTH-1:0] wire_d45_98;
	wire [WIDTH-1:0] wire_d45_99;
	wire [WIDTH-1:0] wire_d45_100;
	wire [WIDTH-1:0] wire_d45_101;
	wire [WIDTH-1:0] wire_d45_102;
	wire [WIDTH-1:0] wire_d45_103;
	wire [WIDTH-1:0] wire_d45_104;
	wire [WIDTH-1:0] wire_d45_105;
	wire [WIDTH-1:0] wire_d45_106;
	wire [WIDTH-1:0] wire_d45_107;
	wire [WIDTH-1:0] wire_d45_108;
	wire [WIDTH-1:0] wire_d45_109;
	wire [WIDTH-1:0] wire_d45_110;
	wire [WIDTH-1:0] wire_d45_111;
	wire [WIDTH-1:0] wire_d45_112;
	wire [WIDTH-1:0] wire_d45_113;
	wire [WIDTH-1:0] wire_d45_114;
	wire [WIDTH-1:0] wire_d45_115;
	wire [WIDTH-1:0] wire_d45_116;
	wire [WIDTH-1:0] wire_d45_117;
	wire [WIDTH-1:0] wire_d45_118;
	wire [WIDTH-1:0] wire_d46_0;
	wire [WIDTH-1:0] wire_d46_1;
	wire [WIDTH-1:0] wire_d46_2;
	wire [WIDTH-1:0] wire_d46_3;
	wire [WIDTH-1:0] wire_d46_4;
	wire [WIDTH-1:0] wire_d46_5;
	wire [WIDTH-1:0] wire_d46_6;
	wire [WIDTH-1:0] wire_d46_7;
	wire [WIDTH-1:0] wire_d46_8;
	wire [WIDTH-1:0] wire_d46_9;
	wire [WIDTH-1:0] wire_d46_10;
	wire [WIDTH-1:0] wire_d46_11;
	wire [WIDTH-1:0] wire_d46_12;
	wire [WIDTH-1:0] wire_d46_13;
	wire [WIDTH-1:0] wire_d46_14;
	wire [WIDTH-1:0] wire_d46_15;
	wire [WIDTH-1:0] wire_d46_16;
	wire [WIDTH-1:0] wire_d46_17;
	wire [WIDTH-1:0] wire_d46_18;
	wire [WIDTH-1:0] wire_d46_19;
	wire [WIDTH-1:0] wire_d46_20;
	wire [WIDTH-1:0] wire_d46_21;
	wire [WIDTH-1:0] wire_d46_22;
	wire [WIDTH-1:0] wire_d46_23;
	wire [WIDTH-1:0] wire_d46_24;
	wire [WIDTH-1:0] wire_d46_25;
	wire [WIDTH-1:0] wire_d46_26;
	wire [WIDTH-1:0] wire_d46_27;
	wire [WIDTH-1:0] wire_d46_28;
	wire [WIDTH-1:0] wire_d46_29;
	wire [WIDTH-1:0] wire_d46_30;
	wire [WIDTH-1:0] wire_d46_31;
	wire [WIDTH-1:0] wire_d46_32;
	wire [WIDTH-1:0] wire_d46_33;
	wire [WIDTH-1:0] wire_d46_34;
	wire [WIDTH-1:0] wire_d46_35;
	wire [WIDTH-1:0] wire_d46_36;
	wire [WIDTH-1:0] wire_d46_37;
	wire [WIDTH-1:0] wire_d46_38;
	wire [WIDTH-1:0] wire_d46_39;
	wire [WIDTH-1:0] wire_d46_40;
	wire [WIDTH-1:0] wire_d46_41;
	wire [WIDTH-1:0] wire_d46_42;
	wire [WIDTH-1:0] wire_d46_43;
	wire [WIDTH-1:0] wire_d46_44;
	wire [WIDTH-1:0] wire_d46_45;
	wire [WIDTH-1:0] wire_d46_46;
	wire [WIDTH-1:0] wire_d46_47;
	wire [WIDTH-1:0] wire_d46_48;
	wire [WIDTH-1:0] wire_d46_49;
	wire [WIDTH-1:0] wire_d46_50;
	wire [WIDTH-1:0] wire_d46_51;
	wire [WIDTH-1:0] wire_d46_52;
	wire [WIDTH-1:0] wire_d46_53;
	wire [WIDTH-1:0] wire_d46_54;
	wire [WIDTH-1:0] wire_d46_55;
	wire [WIDTH-1:0] wire_d46_56;
	wire [WIDTH-1:0] wire_d46_57;
	wire [WIDTH-1:0] wire_d46_58;
	wire [WIDTH-1:0] wire_d46_59;
	wire [WIDTH-1:0] wire_d46_60;
	wire [WIDTH-1:0] wire_d46_61;
	wire [WIDTH-1:0] wire_d46_62;
	wire [WIDTH-1:0] wire_d46_63;
	wire [WIDTH-1:0] wire_d46_64;
	wire [WIDTH-1:0] wire_d46_65;
	wire [WIDTH-1:0] wire_d46_66;
	wire [WIDTH-1:0] wire_d46_67;
	wire [WIDTH-1:0] wire_d46_68;
	wire [WIDTH-1:0] wire_d46_69;
	wire [WIDTH-1:0] wire_d46_70;
	wire [WIDTH-1:0] wire_d46_71;
	wire [WIDTH-1:0] wire_d46_72;
	wire [WIDTH-1:0] wire_d46_73;
	wire [WIDTH-1:0] wire_d46_74;
	wire [WIDTH-1:0] wire_d46_75;
	wire [WIDTH-1:0] wire_d46_76;
	wire [WIDTH-1:0] wire_d46_77;
	wire [WIDTH-1:0] wire_d46_78;
	wire [WIDTH-1:0] wire_d46_79;
	wire [WIDTH-1:0] wire_d46_80;
	wire [WIDTH-1:0] wire_d46_81;
	wire [WIDTH-1:0] wire_d46_82;
	wire [WIDTH-1:0] wire_d46_83;
	wire [WIDTH-1:0] wire_d46_84;
	wire [WIDTH-1:0] wire_d46_85;
	wire [WIDTH-1:0] wire_d46_86;
	wire [WIDTH-1:0] wire_d46_87;
	wire [WIDTH-1:0] wire_d46_88;
	wire [WIDTH-1:0] wire_d46_89;
	wire [WIDTH-1:0] wire_d46_90;
	wire [WIDTH-1:0] wire_d46_91;
	wire [WIDTH-1:0] wire_d46_92;
	wire [WIDTH-1:0] wire_d46_93;
	wire [WIDTH-1:0] wire_d46_94;
	wire [WIDTH-1:0] wire_d46_95;
	wire [WIDTH-1:0] wire_d46_96;
	wire [WIDTH-1:0] wire_d46_97;
	wire [WIDTH-1:0] wire_d46_98;
	wire [WIDTH-1:0] wire_d46_99;
	wire [WIDTH-1:0] wire_d46_100;
	wire [WIDTH-1:0] wire_d46_101;
	wire [WIDTH-1:0] wire_d46_102;
	wire [WIDTH-1:0] wire_d46_103;
	wire [WIDTH-1:0] wire_d46_104;
	wire [WIDTH-1:0] wire_d46_105;
	wire [WIDTH-1:0] wire_d46_106;
	wire [WIDTH-1:0] wire_d46_107;
	wire [WIDTH-1:0] wire_d46_108;
	wire [WIDTH-1:0] wire_d46_109;
	wire [WIDTH-1:0] wire_d46_110;
	wire [WIDTH-1:0] wire_d46_111;
	wire [WIDTH-1:0] wire_d46_112;
	wire [WIDTH-1:0] wire_d46_113;
	wire [WIDTH-1:0] wire_d46_114;
	wire [WIDTH-1:0] wire_d46_115;
	wire [WIDTH-1:0] wire_d46_116;
	wire [WIDTH-1:0] wire_d46_117;
	wire [WIDTH-1:0] wire_d46_118;
	wire [WIDTH-1:0] wire_d47_0;
	wire [WIDTH-1:0] wire_d47_1;
	wire [WIDTH-1:0] wire_d47_2;
	wire [WIDTH-1:0] wire_d47_3;
	wire [WIDTH-1:0] wire_d47_4;
	wire [WIDTH-1:0] wire_d47_5;
	wire [WIDTH-1:0] wire_d47_6;
	wire [WIDTH-1:0] wire_d47_7;
	wire [WIDTH-1:0] wire_d47_8;
	wire [WIDTH-1:0] wire_d47_9;
	wire [WIDTH-1:0] wire_d47_10;
	wire [WIDTH-1:0] wire_d47_11;
	wire [WIDTH-1:0] wire_d47_12;
	wire [WIDTH-1:0] wire_d47_13;
	wire [WIDTH-1:0] wire_d47_14;
	wire [WIDTH-1:0] wire_d47_15;
	wire [WIDTH-1:0] wire_d47_16;
	wire [WIDTH-1:0] wire_d47_17;
	wire [WIDTH-1:0] wire_d47_18;
	wire [WIDTH-1:0] wire_d47_19;
	wire [WIDTH-1:0] wire_d47_20;
	wire [WIDTH-1:0] wire_d47_21;
	wire [WIDTH-1:0] wire_d47_22;
	wire [WIDTH-1:0] wire_d47_23;
	wire [WIDTH-1:0] wire_d47_24;
	wire [WIDTH-1:0] wire_d47_25;
	wire [WIDTH-1:0] wire_d47_26;
	wire [WIDTH-1:0] wire_d47_27;
	wire [WIDTH-1:0] wire_d47_28;
	wire [WIDTH-1:0] wire_d47_29;
	wire [WIDTH-1:0] wire_d47_30;
	wire [WIDTH-1:0] wire_d47_31;
	wire [WIDTH-1:0] wire_d47_32;
	wire [WIDTH-1:0] wire_d47_33;
	wire [WIDTH-1:0] wire_d47_34;
	wire [WIDTH-1:0] wire_d47_35;
	wire [WIDTH-1:0] wire_d47_36;
	wire [WIDTH-1:0] wire_d47_37;
	wire [WIDTH-1:0] wire_d47_38;
	wire [WIDTH-1:0] wire_d47_39;
	wire [WIDTH-1:0] wire_d47_40;
	wire [WIDTH-1:0] wire_d47_41;
	wire [WIDTH-1:0] wire_d47_42;
	wire [WIDTH-1:0] wire_d47_43;
	wire [WIDTH-1:0] wire_d47_44;
	wire [WIDTH-1:0] wire_d47_45;
	wire [WIDTH-1:0] wire_d47_46;
	wire [WIDTH-1:0] wire_d47_47;
	wire [WIDTH-1:0] wire_d47_48;
	wire [WIDTH-1:0] wire_d47_49;
	wire [WIDTH-1:0] wire_d47_50;
	wire [WIDTH-1:0] wire_d47_51;
	wire [WIDTH-1:0] wire_d47_52;
	wire [WIDTH-1:0] wire_d47_53;
	wire [WIDTH-1:0] wire_d47_54;
	wire [WIDTH-1:0] wire_d47_55;
	wire [WIDTH-1:0] wire_d47_56;
	wire [WIDTH-1:0] wire_d47_57;
	wire [WIDTH-1:0] wire_d47_58;
	wire [WIDTH-1:0] wire_d47_59;
	wire [WIDTH-1:0] wire_d47_60;
	wire [WIDTH-1:0] wire_d47_61;
	wire [WIDTH-1:0] wire_d47_62;
	wire [WIDTH-1:0] wire_d47_63;
	wire [WIDTH-1:0] wire_d47_64;
	wire [WIDTH-1:0] wire_d47_65;
	wire [WIDTH-1:0] wire_d47_66;
	wire [WIDTH-1:0] wire_d47_67;
	wire [WIDTH-1:0] wire_d47_68;
	wire [WIDTH-1:0] wire_d47_69;
	wire [WIDTH-1:0] wire_d47_70;
	wire [WIDTH-1:0] wire_d47_71;
	wire [WIDTH-1:0] wire_d47_72;
	wire [WIDTH-1:0] wire_d47_73;
	wire [WIDTH-1:0] wire_d47_74;
	wire [WIDTH-1:0] wire_d47_75;
	wire [WIDTH-1:0] wire_d47_76;
	wire [WIDTH-1:0] wire_d47_77;
	wire [WIDTH-1:0] wire_d47_78;
	wire [WIDTH-1:0] wire_d47_79;
	wire [WIDTH-1:0] wire_d47_80;
	wire [WIDTH-1:0] wire_d47_81;
	wire [WIDTH-1:0] wire_d47_82;
	wire [WIDTH-1:0] wire_d47_83;
	wire [WIDTH-1:0] wire_d47_84;
	wire [WIDTH-1:0] wire_d47_85;
	wire [WIDTH-1:0] wire_d47_86;
	wire [WIDTH-1:0] wire_d47_87;
	wire [WIDTH-1:0] wire_d47_88;
	wire [WIDTH-1:0] wire_d47_89;
	wire [WIDTH-1:0] wire_d47_90;
	wire [WIDTH-1:0] wire_d47_91;
	wire [WIDTH-1:0] wire_d47_92;
	wire [WIDTH-1:0] wire_d47_93;
	wire [WIDTH-1:0] wire_d47_94;
	wire [WIDTH-1:0] wire_d47_95;
	wire [WIDTH-1:0] wire_d47_96;
	wire [WIDTH-1:0] wire_d47_97;
	wire [WIDTH-1:0] wire_d47_98;
	wire [WIDTH-1:0] wire_d47_99;
	wire [WIDTH-1:0] wire_d47_100;
	wire [WIDTH-1:0] wire_d47_101;
	wire [WIDTH-1:0] wire_d47_102;
	wire [WIDTH-1:0] wire_d47_103;
	wire [WIDTH-1:0] wire_d47_104;
	wire [WIDTH-1:0] wire_d47_105;
	wire [WIDTH-1:0] wire_d47_106;
	wire [WIDTH-1:0] wire_d47_107;
	wire [WIDTH-1:0] wire_d47_108;
	wire [WIDTH-1:0] wire_d47_109;
	wire [WIDTH-1:0] wire_d47_110;
	wire [WIDTH-1:0] wire_d47_111;
	wire [WIDTH-1:0] wire_d47_112;
	wire [WIDTH-1:0] wire_d47_113;
	wire [WIDTH-1:0] wire_d47_114;
	wire [WIDTH-1:0] wire_d47_115;
	wire [WIDTH-1:0] wire_d47_116;
	wire [WIDTH-1:0] wire_d47_117;
	wire [WIDTH-1:0] wire_d47_118;
	wire [WIDTH-1:0] wire_d48_0;
	wire [WIDTH-1:0] wire_d48_1;
	wire [WIDTH-1:0] wire_d48_2;
	wire [WIDTH-1:0] wire_d48_3;
	wire [WIDTH-1:0] wire_d48_4;
	wire [WIDTH-1:0] wire_d48_5;
	wire [WIDTH-1:0] wire_d48_6;
	wire [WIDTH-1:0] wire_d48_7;
	wire [WIDTH-1:0] wire_d48_8;
	wire [WIDTH-1:0] wire_d48_9;
	wire [WIDTH-1:0] wire_d48_10;
	wire [WIDTH-1:0] wire_d48_11;
	wire [WIDTH-1:0] wire_d48_12;
	wire [WIDTH-1:0] wire_d48_13;
	wire [WIDTH-1:0] wire_d48_14;
	wire [WIDTH-1:0] wire_d48_15;
	wire [WIDTH-1:0] wire_d48_16;
	wire [WIDTH-1:0] wire_d48_17;
	wire [WIDTH-1:0] wire_d48_18;
	wire [WIDTH-1:0] wire_d48_19;
	wire [WIDTH-1:0] wire_d48_20;
	wire [WIDTH-1:0] wire_d48_21;
	wire [WIDTH-1:0] wire_d48_22;
	wire [WIDTH-1:0] wire_d48_23;
	wire [WIDTH-1:0] wire_d48_24;
	wire [WIDTH-1:0] wire_d48_25;
	wire [WIDTH-1:0] wire_d48_26;
	wire [WIDTH-1:0] wire_d48_27;
	wire [WIDTH-1:0] wire_d48_28;
	wire [WIDTH-1:0] wire_d48_29;
	wire [WIDTH-1:0] wire_d48_30;
	wire [WIDTH-1:0] wire_d48_31;
	wire [WIDTH-1:0] wire_d48_32;
	wire [WIDTH-1:0] wire_d48_33;
	wire [WIDTH-1:0] wire_d48_34;
	wire [WIDTH-1:0] wire_d48_35;
	wire [WIDTH-1:0] wire_d48_36;
	wire [WIDTH-1:0] wire_d48_37;
	wire [WIDTH-1:0] wire_d48_38;
	wire [WIDTH-1:0] wire_d48_39;
	wire [WIDTH-1:0] wire_d48_40;
	wire [WIDTH-1:0] wire_d48_41;
	wire [WIDTH-1:0] wire_d48_42;
	wire [WIDTH-1:0] wire_d48_43;
	wire [WIDTH-1:0] wire_d48_44;
	wire [WIDTH-1:0] wire_d48_45;
	wire [WIDTH-1:0] wire_d48_46;
	wire [WIDTH-1:0] wire_d48_47;
	wire [WIDTH-1:0] wire_d48_48;
	wire [WIDTH-1:0] wire_d48_49;
	wire [WIDTH-1:0] wire_d48_50;
	wire [WIDTH-1:0] wire_d48_51;
	wire [WIDTH-1:0] wire_d48_52;
	wire [WIDTH-1:0] wire_d48_53;
	wire [WIDTH-1:0] wire_d48_54;
	wire [WIDTH-1:0] wire_d48_55;
	wire [WIDTH-1:0] wire_d48_56;
	wire [WIDTH-1:0] wire_d48_57;
	wire [WIDTH-1:0] wire_d48_58;
	wire [WIDTH-1:0] wire_d48_59;
	wire [WIDTH-1:0] wire_d48_60;
	wire [WIDTH-1:0] wire_d48_61;
	wire [WIDTH-1:0] wire_d48_62;
	wire [WIDTH-1:0] wire_d48_63;
	wire [WIDTH-1:0] wire_d48_64;
	wire [WIDTH-1:0] wire_d48_65;
	wire [WIDTH-1:0] wire_d48_66;
	wire [WIDTH-1:0] wire_d48_67;
	wire [WIDTH-1:0] wire_d48_68;
	wire [WIDTH-1:0] wire_d48_69;
	wire [WIDTH-1:0] wire_d48_70;
	wire [WIDTH-1:0] wire_d48_71;
	wire [WIDTH-1:0] wire_d48_72;
	wire [WIDTH-1:0] wire_d48_73;
	wire [WIDTH-1:0] wire_d48_74;
	wire [WIDTH-1:0] wire_d48_75;
	wire [WIDTH-1:0] wire_d48_76;
	wire [WIDTH-1:0] wire_d48_77;
	wire [WIDTH-1:0] wire_d48_78;
	wire [WIDTH-1:0] wire_d48_79;
	wire [WIDTH-1:0] wire_d48_80;
	wire [WIDTH-1:0] wire_d48_81;
	wire [WIDTH-1:0] wire_d48_82;
	wire [WIDTH-1:0] wire_d48_83;
	wire [WIDTH-1:0] wire_d48_84;
	wire [WIDTH-1:0] wire_d48_85;
	wire [WIDTH-1:0] wire_d48_86;
	wire [WIDTH-1:0] wire_d48_87;
	wire [WIDTH-1:0] wire_d48_88;
	wire [WIDTH-1:0] wire_d48_89;
	wire [WIDTH-1:0] wire_d48_90;
	wire [WIDTH-1:0] wire_d48_91;
	wire [WIDTH-1:0] wire_d48_92;
	wire [WIDTH-1:0] wire_d48_93;
	wire [WIDTH-1:0] wire_d48_94;
	wire [WIDTH-1:0] wire_d48_95;
	wire [WIDTH-1:0] wire_d48_96;
	wire [WIDTH-1:0] wire_d48_97;
	wire [WIDTH-1:0] wire_d48_98;
	wire [WIDTH-1:0] wire_d48_99;
	wire [WIDTH-1:0] wire_d48_100;
	wire [WIDTH-1:0] wire_d48_101;
	wire [WIDTH-1:0] wire_d48_102;
	wire [WIDTH-1:0] wire_d48_103;
	wire [WIDTH-1:0] wire_d48_104;
	wire [WIDTH-1:0] wire_d48_105;
	wire [WIDTH-1:0] wire_d48_106;
	wire [WIDTH-1:0] wire_d48_107;
	wire [WIDTH-1:0] wire_d48_108;
	wire [WIDTH-1:0] wire_d48_109;
	wire [WIDTH-1:0] wire_d48_110;
	wire [WIDTH-1:0] wire_d48_111;
	wire [WIDTH-1:0] wire_d48_112;
	wire [WIDTH-1:0] wire_d48_113;
	wire [WIDTH-1:0] wire_d48_114;
	wire [WIDTH-1:0] wire_d48_115;
	wire [WIDTH-1:0] wire_d48_116;
	wire [WIDTH-1:0] wire_d48_117;
	wire [WIDTH-1:0] wire_d48_118;
	wire [WIDTH-1:0] wire_d49_0;
	wire [WIDTH-1:0] wire_d49_1;
	wire [WIDTH-1:0] wire_d49_2;
	wire [WIDTH-1:0] wire_d49_3;
	wire [WIDTH-1:0] wire_d49_4;
	wire [WIDTH-1:0] wire_d49_5;
	wire [WIDTH-1:0] wire_d49_6;
	wire [WIDTH-1:0] wire_d49_7;
	wire [WIDTH-1:0] wire_d49_8;
	wire [WIDTH-1:0] wire_d49_9;
	wire [WIDTH-1:0] wire_d49_10;
	wire [WIDTH-1:0] wire_d49_11;
	wire [WIDTH-1:0] wire_d49_12;
	wire [WIDTH-1:0] wire_d49_13;
	wire [WIDTH-1:0] wire_d49_14;
	wire [WIDTH-1:0] wire_d49_15;
	wire [WIDTH-1:0] wire_d49_16;
	wire [WIDTH-1:0] wire_d49_17;
	wire [WIDTH-1:0] wire_d49_18;
	wire [WIDTH-1:0] wire_d49_19;
	wire [WIDTH-1:0] wire_d49_20;
	wire [WIDTH-1:0] wire_d49_21;
	wire [WIDTH-1:0] wire_d49_22;
	wire [WIDTH-1:0] wire_d49_23;
	wire [WIDTH-1:0] wire_d49_24;
	wire [WIDTH-1:0] wire_d49_25;
	wire [WIDTH-1:0] wire_d49_26;
	wire [WIDTH-1:0] wire_d49_27;
	wire [WIDTH-1:0] wire_d49_28;
	wire [WIDTH-1:0] wire_d49_29;
	wire [WIDTH-1:0] wire_d49_30;
	wire [WIDTH-1:0] wire_d49_31;
	wire [WIDTH-1:0] wire_d49_32;
	wire [WIDTH-1:0] wire_d49_33;
	wire [WIDTH-1:0] wire_d49_34;
	wire [WIDTH-1:0] wire_d49_35;
	wire [WIDTH-1:0] wire_d49_36;
	wire [WIDTH-1:0] wire_d49_37;
	wire [WIDTH-1:0] wire_d49_38;
	wire [WIDTH-1:0] wire_d49_39;
	wire [WIDTH-1:0] wire_d49_40;
	wire [WIDTH-1:0] wire_d49_41;
	wire [WIDTH-1:0] wire_d49_42;
	wire [WIDTH-1:0] wire_d49_43;
	wire [WIDTH-1:0] wire_d49_44;
	wire [WIDTH-1:0] wire_d49_45;
	wire [WIDTH-1:0] wire_d49_46;
	wire [WIDTH-1:0] wire_d49_47;
	wire [WIDTH-1:0] wire_d49_48;
	wire [WIDTH-1:0] wire_d49_49;
	wire [WIDTH-1:0] wire_d49_50;
	wire [WIDTH-1:0] wire_d49_51;
	wire [WIDTH-1:0] wire_d49_52;
	wire [WIDTH-1:0] wire_d49_53;
	wire [WIDTH-1:0] wire_d49_54;
	wire [WIDTH-1:0] wire_d49_55;
	wire [WIDTH-1:0] wire_d49_56;
	wire [WIDTH-1:0] wire_d49_57;
	wire [WIDTH-1:0] wire_d49_58;
	wire [WIDTH-1:0] wire_d49_59;
	wire [WIDTH-1:0] wire_d49_60;
	wire [WIDTH-1:0] wire_d49_61;
	wire [WIDTH-1:0] wire_d49_62;
	wire [WIDTH-1:0] wire_d49_63;
	wire [WIDTH-1:0] wire_d49_64;
	wire [WIDTH-1:0] wire_d49_65;
	wire [WIDTH-1:0] wire_d49_66;
	wire [WIDTH-1:0] wire_d49_67;
	wire [WIDTH-1:0] wire_d49_68;
	wire [WIDTH-1:0] wire_d49_69;
	wire [WIDTH-1:0] wire_d49_70;
	wire [WIDTH-1:0] wire_d49_71;
	wire [WIDTH-1:0] wire_d49_72;
	wire [WIDTH-1:0] wire_d49_73;
	wire [WIDTH-1:0] wire_d49_74;
	wire [WIDTH-1:0] wire_d49_75;
	wire [WIDTH-1:0] wire_d49_76;
	wire [WIDTH-1:0] wire_d49_77;
	wire [WIDTH-1:0] wire_d49_78;
	wire [WIDTH-1:0] wire_d49_79;
	wire [WIDTH-1:0] wire_d49_80;
	wire [WIDTH-1:0] wire_d49_81;
	wire [WIDTH-1:0] wire_d49_82;
	wire [WIDTH-1:0] wire_d49_83;
	wire [WIDTH-1:0] wire_d49_84;
	wire [WIDTH-1:0] wire_d49_85;
	wire [WIDTH-1:0] wire_d49_86;
	wire [WIDTH-1:0] wire_d49_87;
	wire [WIDTH-1:0] wire_d49_88;
	wire [WIDTH-1:0] wire_d49_89;
	wire [WIDTH-1:0] wire_d49_90;
	wire [WIDTH-1:0] wire_d49_91;
	wire [WIDTH-1:0] wire_d49_92;
	wire [WIDTH-1:0] wire_d49_93;
	wire [WIDTH-1:0] wire_d49_94;
	wire [WIDTH-1:0] wire_d49_95;
	wire [WIDTH-1:0] wire_d49_96;
	wire [WIDTH-1:0] wire_d49_97;
	wire [WIDTH-1:0] wire_d49_98;
	wire [WIDTH-1:0] wire_d49_99;
	wire [WIDTH-1:0] wire_d49_100;
	wire [WIDTH-1:0] wire_d49_101;
	wire [WIDTH-1:0] wire_d49_102;
	wire [WIDTH-1:0] wire_d49_103;
	wire [WIDTH-1:0] wire_d49_104;
	wire [WIDTH-1:0] wire_d49_105;
	wire [WIDTH-1:0] wire_d49_106;
	wire [WIDTH-1:0] wire_d49_107;
	wire [WIDTH-1:0] wire_d49_108;
	wire [WIDTH-1:0] wire_d49_109;
	wire [WIDTH-1:0] wire_d49_110;
	wire [WIDTH-1:0] wire_d49_111;
	wire [WIDTH-1:0] wire_d49_112;
	wire [WIDTH-1:0] wire_d49_113;
	wire [WIDTH-1:0] wire_d49_114;
	wire [WIDTH-1:0] wire_d49_115;
	wire [WIDTH-1:0] wire_d49_116;
	wire [WIDTH-1:0] wire_d49_117;
	wire [WIDTH-1:0] wire_d49_118;
	wire [WIDTH-1:0] wire_d50_0;
	wire [WIDTH-1:0] wire_d50_1;
	wire [WIDTH-1:0] wire_d50_2;
	wire [WIDTH-1:0] wire_d50_3;
	wire [WIDTH-1:0] wire_d50_4;
	wire [WIDTH-1:0] wire_d50_5;
	wire [WIDTH-1:0] wire_d50_6;
	wire [WIDTH-1:0] wire_d50_7;
	wire [WIDTH-1:0] wire_d50_8;
	wire [WIDTH-1:0] wire_d50_9;
	wire [WIDTH-1:0] wire_d50_10;
	wire [WIDTH-1:0] wire_d50_11;
	wire [WIDTH-1:0] wire_d50_12;
	wire [WIDTH-1:0] wire_d50_13;
	wire [WIDTH-1:0] wire_d50_14;
	wire [WIDTH-1:0] wire_d50_15;
	wire [WIDTH-1:0] wire_d50_16;
	wire [WIDTH-1:0] wire_d50_17;
	wire [WIDTH-1:0] wire_d50_18;
	wire [WIDTH-1:0] wire_d50_19;
	wire [WIDTH-1:0] wire_d50_20;
	wire [WIDTH-1:0] wire_d50_21;
	wire [WIDTH-1:0] wire_d50_22;
	wire [WIDTH-1:0] wire_d50_23;
	wire [WIDTH-1:0] wire_d50_24;
	wire [WIDTH-1:0] wire_d50_25;
	wire [WIDTH-1:0] wire_d50_26;
	wire [WIDTH-1:0] wire_d50_27;
	wire [WIDTH-1:0] wire_d50_28;
	wire [WIDTH-1:0] wire_d50_29;
	wire [WIDTH-1:0] wire_d50_30;
	wire [WIDTH-1:0] wire_d50_31;
	wire [WIDTH-1:0] wire_d50_32;
	wire [WIDTH-1:0] wire_d50_33;
	wire [WIDTH-1:0] wire_d50_34;
	wire [WIDTH-1:0] wire_d50_35;
	wire [WIDTH-1:0] wire_d50_36;
	wire [WIDTH-1:0] wire_d50_37;
	wire [WIDTH-1:0] wire_d50_38;
	wire [WIDTH-1:0] wire_d50_39;
	wire [WIDTH-1:0] wire_d50_40;
	wire [WIDTH-1:0] wire_d50_41;
	wire [WIDTH-1:0] wire_d50_42;
	wire [WIDTH-1:0] wire_d50_43;
	wire [WIDTH-1:0] wire_d50_44;
	wire [WIDTH-1:0] wire_d50_45;
	wire [WIDTH-1:0] wire_d50_46;
	wire [WIDTH-1:0] wire_d50_47;
	wire [WIDTH-1:0] wire_d50_48;
	wire [WIDTH-1:0] wire_d50_49;
	wire [WIDTH-1:0] wire_d50_50;
	wire [WIDTH-1:0] wire_d50_51;
	wire [WIDTH-1:0] wire_d50_52;
	wire [WIDTH-1:0] wire_d50_53;
	wire [WIDTH-1:0] wire_d50_54;
	wire [WIDTH-1:0] wire_d50_55;
	wire [WIDTH-1:0] wire_d50_56;
	wire [WIDTH-1:0] wire_d50_57;
	wire [WIDTH-1:0] wire_d50_58;
	wire [WIDTH-1:0] wire_d50_59;
	wire [WIDTH-1:0] wire_d50_60;
	wire [WIDTH-1:0] wire_d50_61;
	wire [WIDTH-1:0] wire_d50_62;
	wire [WIDTH-1:0] wire_d50_63;
	wire [WIDTH-1:0] wire_d50_64;
	wire [WIDTH-1:0] wire_d50_65;
	wire [WIDTH-1:0] wire_d50_66;
	wire [WIDTH-1:0] wire_d50_67;
	wire [WIDTH-1:0] wire_d50_68;
	wire [WIDTH-1:0] wire_d50_69;
	wire [WIDTH-1:0] wire_d50_70;
	wire [WIDTH-1:0] wire_d50_71;
	wire [WIDTH-1:0] wire_d50_72;
	wire [WIDTH-1:0] wire_d50_73;
	wire [WIDTH-1:0] wire_d50_74;
	wire [WIDTH-1:0] wire_d50_75;
	wire [WIDTH-1:0] wire_d50_76;
	wire [WIDTH-1:0] wire_d50_77;
	wire [WIDTH-1:0] wire_d50_78;
	wire [WIDTH-1:0] wire_d50_79;
	wire [WIDTH-1:0] wire_d50_80;
	wire [WIDTH-1:0] wire_d50_81;
	wire [WIDTH-1:0] wire_d50_82;
	wire [WIDTH-1:0] wire_d50_83;
	wire [WIDTH-1:0] wire_d50_84;
	wire [WIDTH-1:0] wire_d50_85;
	wire [WIDTH-1:0] wire_d50_86;
	wire [WIDTH-1:0] wire_d50_87;
	wire [WIDTH-1:0] wire_d50_88;
	wire [WIDTH-1:0] wire_d50_89;
	wire [WIDTH-1:0] wire_d50_90;
	wire [WIDTH-1:0] wire_d50_91;
	wire [WIDTH-1:0] wire_d50_92;
	wire [WIDTH-1:0] wire_d50_93;
	wire [WIDTH-1:0] wire_d50_94;
	wire [WIDTH-1:0] wire_d50_95;
	wire [WIDTH-1:0] wire_d50_96;
	wire [WIDTH-1:0] wire_d50_97;
	wire [WIDTH-1:0] wire_d50_98;
	wire [WIDTH-1:0] wire_d50_99;
	wire [WIDTH-1:0] wire_d50_100;
	wire [WIDTH-1:0] wire_d50_101;
	wire [WIDTH-1:0] wire_d50_102;
	wire [WIDTH-1:0] wire_d50_103;
	wire [WIDTH-1:0] wire_d50_104;
	wire [WIDTH-1:0] wire_d50_105;
	wire [WIDTH-1:0] wire_d50_106;
	wire [WIDTH-1:0] wire_d50_107;
	wire [WIDTH-1:0] wire_d50_108;
	wire [WIDTH-1:0] wire_d50_109;
	wire [WIDTH-1:0] wire_d50_110;
	wire [WIDTH-1:0] wire_d50_111;
	wire [WIDTH-1:0] wire_d50_112;
	wire [WIDTH-1:0] wire_d50_113;
	wire [WIDTH-1:0] wire_d50_114;
	wire [WIDTH-1:0] wire_d50_115;
	wire [WIDTH-1:0] wire_d50_116;
	wire [WIDTH-1:0] wire_d50_117;
	wire [WIDTH-1:0] wire_d50_118;
	wire [WIDTH-1:0] wire_d51_0;
	wire [WIDTH-1:0] wire_d51_1;
	wire [WIDTH-1:0] wire_d51_2;
	wire [WIDTH-1:0] wire_d51_3;
	wire [WIDTH-1:0] wire_d51_4;
	wire [WIDTH-1:0] wire_d51_5;
	wire [WIDTH-1:0] wire_d51_6;
	wire [WIDTH-1:0] wire_d51_7;
	wire [WIDTH-1:0] wire_d51_8;
	wire [WIDTH-1:0] wire_d51_9;
	wire [WIDTH-1:0] wire_d51_10;
	wire [WIDTH-1:0] wire_d51_11;
	wire [WIDTH-1:0] wire_d51_12;
	wire [WIDTH-1:0] wire_d51_13;
	wire [WIDTH-1:0] wire_d51_14;
	wire [WIDTH-1:0] wire_d51_15;
	wire [WIDTH-1:0] wire_d51_16;
	wire [WIDTH-1:0] wire_d51_17;
	wire [WIDTH-1:0] wire_d51_18;
	wire [WIDTH-1:0] wire_d51_19;
	wire [WIDTH-1:0] wire_d51_20;
	wire [WIDTH-1:0] wire_d51_21;
	wire [WIDTH-1:0] wire_d51_22;
	wire [WIDTH-1:0] wire_d51_23;
	wire [WIDTH-1:0] wire_d51_24;
	wire [WIDTH-1:0] wire_d51_25;
	wire [WIDTH-1:0] wire_d51_26;
	wire [WIDTH-1:0] wire_d51_27;
	wire [WIDTH-1:0] wire_d51_28;
	wire [WIDTH-1:0] wire_d51_29;
	wire [WIDTH-1:0] wire_d51_30;
	wire [WIDTH-1:0] wire_d51_31;
	wire [WIDTH-1:0] wire_d51_32;
	wire [WIDTH-1:0] wire_d51_33;
	wire [WIDTH-1:0] wire_d51_34;
	wire [WIDTH-1:0] wire_d51_35;
	wire [WIDTH-1:0] wire_d51_36;
	wire [WIDTH-1:0] wire_d51_37;
	wire [WIDTH-1:0] wire_d51_38;
	wire [WIDTH-1:0] wire_d51_39;
	wire [WIDTH-1:0] wire_d51_40;
	wire [WIDTH-1:0] wire_d51_41;
	wire [WIDTH-1:0] wire_d51_42;
	wire [WIDTH-1:0] wire_d51_43;
	wire [WIDTH-1:0] wire_d51_44;
	wire [WIDTH-1:0] wire_d51_45;
	wire [WIDTH-1:0] wire_d51_46;
	wire [WIDTH-1:0] wire_d51_47;
	wire [WIDTH-1:0] wire_d51_48;
	wire [WIDTH-1:0] wire_d51_49;
	wire [WIDTH-1:0] wire_d51_50;
	wire [WIDTH-1:0] wire_d51_51;
	wire [WIDTH-1:0] wire_d51_52;
	wire [WIDTH-1:0] wire_d51_53;
	wire [WIDTH-1:0] wire_d51_54;
	wire [WIDTH-1:0] wire_d51_55;
	wire [WIDTH-1:0] wire_d51_56;
	wire [WIDTH-1:0] wire_d51_57;
	wire [WIDTH-1:0] wire_d51_58;
	wire [WIDTH-1:0] wire_d51_59;
	wire [WIDTH-1:0] wire_d51_60;
	wire [WIDTH-1:0] wire_d51_61;
	wire [WIDTH-1:0] wire_d51_62;
	wire [WIDTH-1:0] wire_d51_63;
	wire [WIDTH-1:0] wire_d51_64;
	wire [WIDTH-1:0] wire_d51_65;
	wire [WIDTH-1:0] wire_d51_66;
	wire [WIDTH-1:0] wire_d51_67;
	wire [WIDTH-1:0] wire_d51_68;
	wire [WIDTH-1:0] wire_d51_69;
	wire [WIDTH-1:0] wire_d51_70;
	wire [WIDTH-1:0] wire_d51_71;
	wire [WIDTH-1:0] wire_d51_72;
	wire [WIDTH-1:0] wire_d51_73;
	wire [WIDTH-1:0] wire_d51_74;
	wire [WIDTH-1:0] wire_d51_75;
	wire [WIDTH-1:0] wire_d51_76;
	wire [WIDTH-1:0] wire_d51_77;
	wire [WIDTH-1:0] wire_d51_78;
	wire [WIDTH-1:0] wire_d51_79;
	wire [WIDTH-1:0] wire_d51_80;
	wire [WIDTH-1:0] wire_d51_81;
	wire [WIDTH-1:0] wire_d51_82;
	wire [WIDTH-1:0] wire_d51_83;
	wire [WIDTH-1:0] wire_d51_84;
	wire [WIDTH-1:0] wire_d51_85;
	wire [WIDTH-1:0] wire_d51_86;
	wire [WIDTH-1:0] wire_d51_87;
	wire [WIDTH-1:0] wire_d51_88;
	wire [WIDTH-1:0] wire_d51_89;
	wire [WIDTH-1:0] wire_d51_90;
	wire [WIDTH-1:0] wire_d51_91;
	wire [WIDTH-1:0] wire_d51_92;
	wire [WIDTH-1:0] wire_d51_93;
	wire [WIDTH-1:0] wire_d51_94;
	wire [WIDTH-1:0] wire_d51_95;
	wire [WIDTH-1:0] wire_d51_96;
	wire [WIDTH-1:0] wire_d51_97;
	wire [WIDTH-1:0] wire_d51_98;
	wire [WIDTH-1:0] wire_d51_99;
	wire [WIDTH-1:0] wire_d51_100;
	wire [WIDTH-1:0] wire_d51_101;
	wire [WIDTH-1:0] wire_d51_102;
	wire [WIDTH-1:0] wire_d51_103;
	wire [WIDTH-1:0] wire_d51_104;
	wire [WIDTH-1:0] wire_d51_105;
	wire [WIDTH-1:0] wire_d51_106;
	wire [WIDTH-1:0] wire_d51_107;
	wire [WIDTH-1:0] wire_d51_108;
	wire [WIDTH-1:0] wire_d51_109;
	wire [WIDTH-1:0] wire_d51_110;
	wire [WIDTH-1:0] wire_d51_111;
	wire [WIDTH-1:0] wire_d51_112;
	wire [WIDTH-1:0] wire_d51_113;
	wire [WIDTH-1:0] wire_d51_114;
	wire [WIDTH-1:0] wire_d51_115;
	wire [WIDTH-1:0] wire_d51_116;
	wire [WIDTH-1:0] wire_d51_117;
	wire [WIDTH-1:0] wire_d51_118;
	wire [WIDTH-1:0] wire_d52_0;
	wire [WIDTH-1:0] wire_d52_1;
	wire [WIDTH-1:0] wire_d52_2;
	wire [WIDTH-1:0] wire_d52_3;
	wire [WIDTH-1:0] wire_d52_4;
	wire [WIDTH-1:0] wire_d52_5;
	wire [WIDTH-1:0] wire_d52_6;
	wire [WIDTH-1:0] wire_d52_7;
	wire [WIDTH-1:0] wire_d52_8;
	wire [WIDTH-1:0] wire_d52_9;
	wire [WIDTH-1:0] wire_d52_10;
	wire [WIDTH-1:0] wire_d52_11;
	wire [WIDTH-1:0] wire_d52_12;
	wire [WIDTH-1:0] wire_d52_13;
	wire [WIDTH-1:0] wire_d52_14;
	wire [WIDTH-1:0] wire_d52_15;
	wire [WIDTH-1:0] wire_d52_16;
	wire [WIDTH-1:0] wire_d52_17;
	wire [WIDTH-1:0] wire_d52_18;
	wire [WIDTH-1:0] wire_d52_19;
	wire [WIDTH-1:0] wire_d52_20;
	wire [WIDTH-1:0] wire_d52_21;
	wire [WIDTH-1:0] wire_d52_22;
	wire [WIDTH-1:0] wire_d52_23;
	wire [WIDTH-1:0] wire_d52_24;
	wire [WIDTH-1:0] wire_d52_25;
	wire [WIDTH-1:0] wire_d52_26;
	wire [WIDTH-1:0] wire_d52_27;
	wire [WIDTH-1:0] wire_d52_28;
	wire [WIDTH-1:0] wire_d52_29;
	wire [WIDTH-1:0] wire_d52_30;
	wire [WIDTH-1:0] wire_d52_31;
	wire [WIDTH-1:0] wire_d52_32;
	wire [WIDTH-1:0] wire_d52_33;
	wire [WIDTH-1:0] wire_d52_34;
	wire [WIDTH-1:0] wire_d52_35;
	wire [WIDTH-1:0] wire_d52_36;
	wire [WIDTH-1:0] wire_d52_37;
	wire [WIDTH-1:0] wire_d52_38;
	wire [WIDTH-1:0] wire_d52_39;
	wire [WIDTH-1:0] wire_d52_40;
	wire [WIDTH-1:0] wire_d52_41;
	wire [WIDTH-1:0] wire_d52_42;
	wire [WIDTH-1:0] wire_d52_43;
	wire [WIDTH-1:0] wire_d52_44;
	wire [WIDTH-1:0] wire_d52_45;
	wire [WIDTH-1:0] wire_d52_46;
	wire [WIDTH-1:0] wire_d52_47;
	wire [WIDTH-1:0] wire_d52_48;
	wire [WIDTH-1:0] wire_d52_49;
	wire [WIDTH-1:0] wire_d52_50;
	wire [WIDTH-1:0] wire_d52_51;
	wire [WIDTH-1:0] wire_d52_52;
	wire [WIDTH-1:0] wire_d52_53;
	wire [WIDTH-1:0] wire_d52_54;
	wire [WIDTH-1:0] wire_d52_55;
	wire [WIDTH-1:0] wire_d52_56;
	wire [WIDTH-1:0] wire_d52_57;
	wire [WIDTH-1:0] wire_d52_58;
	wire [WIDTH-1:0] wire_d52_59;
	wire [WIDTH-1:0] wire_d52_60;
	wire [WIDTH-1:0] wire_d52_61;
	wire [WIDTH-1:0] wire_d52_62;
	wire [WIDTH-1:0] wire_d52_63;
	wire [WIDTH-1:0] wire_d52_64;
	wire [WIDTH-1:0] wire_d52_65;
	wire [WIDTH-1:0] wire_d52_66;
	wire [WIDTH-1:0] wire_d52_67;
	wire [WIDTH-1:0] wire_d52_68;
	wire [WIDTH-1:0] wire_d52_69;
	wire [WIDTH-1:0] wire_d52_70;
	wire [WIDTH-1:0] wire_d52_71;
	wire [WIDTH-1:0] wire_d52_72;
	wire [WIDTH-1:0] wire_d52_73;
	wire [WIDTH-1:0] wire_d52_74;
	wire [WIDTH-1:0] wire_d52_75;
	wire [WIDTH-1:0] wire_d52_76;
	wire [WIDTH-1:0] wire_d52_77;
	wire [WIDTH-1:0] wire_d52_78;
	wire [WIDTH-1:0] wire_d52_79;
	wire [WIDTH-1:0] wire_d52_80;
	wire [WIDTH-1:0] wire_d52_81;
	wire [WIDTH-1:0] wire_d52_82;
	wire [WIDTH-1:0] wire_d52_83;
	wire [WIDTH-1:0] wire_d52_84;
	wire [WIDTH-1:0] wire_d52_85;
	wire [WIDTH-1:0] wire_d52_86;
	wire [WIDTH-1:0] wire_d52_87;
	wire [WIDTH-1:0] wire_d52_88;
	wire [WIDTH-1:0] wire_d52_89;
	wire [WIDTH-1:0] wire_d52_90;
	wire [WIDTH-1:0] wire_d52_91;
	wire [WIDTH-1:0] wire_d52_92;
	wire [WIDTH-1:0] wire_d52_93;
	wire [WIDTH-1:0] wire_d52_94;
	wire [WIDTH-1:0] wire_d52_95;
	wire [WIDTH-1:0] wire_d52_96;
	wire [WIDTH-1:0] wire_d52_97;
	wire [WIDTH-1:0] wire_d52_98;
	wire [WIDTH-1:0] wire_d52_99;
	wire [WIDTH-1:0] wire_d52_100;
	wire [WIDTH-1:0] wire_d52_101;
	wire [WIDTH-1:0] wire_d52_102;
	wire [WIDTH-1:0] wire_d52_103;
	wire [WIDTH-1:0] wire_d52_104;
	wire [WIDTH-1:0] wire_d52_105;
	wire [WIDTH-1:0] wire_d52_106;
	wire [WIDTH-1:0] wire_d52_107;
	wire [WIDTH-1:0] wire_d52_108;
	wire [WIDTH-1:0] wire_d52_109;
	wire [WIDTH-1:0] wire_d52_110;
	wire [WIDTH-1:0] wire_d52_111;
	wire [WIDTH-1:0] wire_d52_112;
	wire [WIDTH-1:0] wire_d52_113;
	wire [WIDTH-1:0] wire_d52_114;
	wire [WIDTH-1:0] wire_d52_115;
	wire [WIDTH-1:0] wire_d52_116;
	wire [WIDTH-1:0] wire_d52_117;
	wire [WIDTH-1:0] wire_d52_118;
	wire [WIDTH-1:0] wire_d53_0;
	wire [WIDTH-1:0] wire_d53_1;
	wire [WIDTH-1:0] wire_d53_2;
	wire [WIDTH-1:0] wire_d53_3;
	wire [WIDTH-1:0] wire_d53_4;
	wire [WIDTH-1:0] wire_d53_5;
	wire [WIDTH-1:0] wire_d53_6;
	wire [WIDTH-1:0] wire_d53_7;
	wire [WIDTH-1:0] wire_d53_8;
	wire [WIDTH-1:0] wire_d53_9;
	wire [WIDTH-1:0] wire_d53_10;
	wire [WIDTH-1:0] wire_d53_11;
	wire [WIDTH-1:0] wire_d53_12;
	wire [WIDTH-1:0] wire_d53_13;
	wire [WIDTH-1:0] wire_d53_14;
	wire [WIDTH-1:0] wire_d53_15;
	wire [WIDTH-1:0] wire_d53_16;
	wire [WIDTH-1:0] wire_d53_17;
	wire [WIDTH-1:0] wire_d53_18;
	wire [WIDTH-1:0] wire_d53_19;
	wire [WIDTH-1:0] wire_d53_20;
	wire [WIDTH-1:0] wire_d53_21;
	wire [WIDTH-1:0] wire_d53_22;
	wire [WIDTH-1:0] wire_d53_23;
	wire [WIDTH-1:0] wire_d53_24;
	wire [WIDTH-1:0] wire_d53_25;
	wire [WIDTH-1:0] wire_d53_26;
	wire [WIDTH-1:0] wire_d53_27;
	wire [WIDTH-1:0] wire_d53_28;
	wire [WIDTH-1:0] wire_d53_29;
	wire [WIDTH-1:0] wire_d53_30;
	wire [WIDTH-1:0] wire_d53_31;
	wire [WIDTH-1:0] wire_d53_32;
	wire [WIDTH-1:0] wire_d53_33;
	wire [WIDTH-1:0] wire_d53_34;
	wire [WIDTH-1:0] wire_d53_35;
	wire [WIDTH-1:0] wire_d53_36;
	wire [WIDTH-1:0] wire_d53_37;
	wire [WIDTH-1:0] wire_d53_38;
	wire [WIDTH-1:0] wire_d53_39;
	wire [WIDTH-1:0] wire_d53_40;
	wire [WIDTH-1:0] wire_d53_41;
	wire [WIDTH-1:0] wire_d53_42;
	wire [WIDTH-1:0] wire_d53_43;
	wire [WIDTH-1:0] wire_d53_44;
	wire [WIDTH-1:0] wire_d53_45;
	wire [WIDTH-1:0] wire_d53_46;
	wire [WIDTH-1:0] wire_d53_47;
	wire [WIDTH-1:0] wire_d53_48;
	wire [WIDTH-1:0] wire_d53_49;
	wire [WIDTH-1:0] wire_d53_50;
	wire [WIDTH-1:0] wire_d53_51;
	wire [WIDTH-1:0] wire_d53_52;
	wire [WIDTH-1:0] wire_d53_53;
	wire [WIDTH-1:0] wire_d53_54;
	wire [WIDTH-1:0] wire_d53_55;
	wire [WIDTH-1:0] wire_d53_56;
	wire [WIDTH-1:0] wire_d53_57;
	wire [WIDTH-1:0] wire_d53_58;
	wire [WIDTH-1:0] wire_d53_59;
	wire [WIDTH-1:0] wire_d53_60;
	wire [WIDTH-1:0] wire_d53_61;
	wire [WIDTH-1:0] wire_d53_62;
	wire [WIDTH-1:0] wire_d53_63;
	wire [WIDTH-1:0] wire_d53_64;
	wire [WIDTH-1:0] wire_d53_65;
	wire [WIDTH-1:0] wire_d53_66;
	wire [WIDTH-1:0] wire_d53_67;
	wire [WIDTH-1:0] wire_d53_68;
	wire [WIDTH-1:0] wire_d53_69;
	wire [WIDTH-1:0] wire_d53_70;
	wire [WIDTH-1:0] wire_d53_71;
	wire [WIDTH-1:0] wire_d53_72;
	wire [WIDTH-1:0] wire_d53_73;
	wire [WIDTH-1:0] wire_d53_74;
	wire [WIDTH-1:0] wire_d53_75;
	wire [WIDTH-1:0] wire_d53_76;
	wire [WIDTH-1:0] wire_d53_77;
	wire [WIDTH-1:0] wire_d53_78;
	wire [WIDTH-1:0] wire_d53_79;
	wire [WIDTH-1:0] wire_d53_80;
	wire [WIDTH-1:0] wire_d53_81;
	wire [WIDTH-1:0] wire_d53_82;
	wire [WIDTH-1:0] wire_d53_83;
	wire [WIDTH-1:0] wire_d53_84;
	wire [WIDTH-1:0] wire_d53_85;
	wire [WIDTH-1:0] wire_d53_86;
	wire [WIDTH-1:0] wire_d53_87;
	wire [WIDTH-1:0] wire_d53_88;
	wire [WIDTH-1:0] wire_d53_89;
	wire [WIDTH-1:0] wire_d53_90;
	wire [WIDTH-1:0] wire_d53_91;
	wire [WIDTH-1:0] wire_d53_92;
	wire [WIDTH-1:0] wire_d53_93;
	wire [WIDTH-1:0] wire_d53_94;
	wire [WIDTH-1:0] wire_d53_95;
	wire [WIDTH-1:0] wire_d53_96;
	wire [WIDTH-1:0] wire_d53_97;
	wire [WIDTH-1:0] wire_d53_98;
	wire [WIDTH-1:0] wire_d53_99;
	wire [WIDTH-1:0] wire_d53_100;
	wire [WIDTH-1:0] wire_d53_101;
	wire [WIDTH-1:0] wire_d53_102;
	wire [WIDTH-1:0] wire_d53_103;
	wire [WIDTH-1:0] wire_d53_104;
	wire [WIDTH-1:0] wire_d53_105;
	wire [WIDTH-1:0] wire_d53_106;
	wire [WIDTH-1:0] wire_d53_107;
	wire [WIDTH-1:0] wire_d53_108;
	wire [WIDTH-1:0] wire_d53_109;
	wire [WIDTH-1:0] wire_d53_110;
	wire [WIDTH-1:0] wire_d53_111;
	wire [WIDTH-1:0] wire_d53_112;
	wire [WIDTH-1:0] wire_d53_113;
	wire [WIDTH-1:0] wire_d53_114;
	wire [WIDTH-1:0] wire_d53_115;
	wire [WIDTH-1:0] wire_d53_116;
	wire [WIDTH-1:0] wire_d53_117;
	wire [WIDTH-1:0] wire_d53_118;
	wire [WIDTH-1:0] wire_d54_0;
	wire [WIDTH-1:0] wire_d54_1;
	wire [WIDTH-1:0] wire_d54_2;
	wire [WIDTH-1:0] wire_d54_3;
	wire [WIDTH-1:0] wire_d54_4;
	wire [WIDTH-1:0] wire_d54_5;
	wire [WIDTH-1:0] wire_d54_6;
	wire [WIDTH-1:0] wire_d54_7;
	wire [WIDTH-1:0] wire_d54_8;
	wire [WIDTH-1:0] wire_d54_9;
	wire [WIDTH-1:0] wire_d54_10;
	wire [WIDTH-1:0] wire_d54_11;
	wire [WIDTH-1:0] wire_d54_12;
	wire [WIDTH-1:0] wire_d54_13;
	wire [WIDTH-1:0] wire_d54_14;
	wire [WIDTH-1:0] wire_d54_15;
	wire [WIDTH-1:0] wire_d54_16;
	wire [WIDTH-1:0] wire_d54_17;
	wire [WIDTH-1:0] wire_d54_18;
	wire [WIDTH-1:0] wire_d54_19;
	wire [WIDTH-1:0] wire_d54_20;
	wire [WIDTH-1:0] wire_d54_21;
	wire [WIDTH-1:0] wire_d54_22;
	wire [WIDTH-1:0] wire_d54_23;
	wire [WIDTH-1:0] wire_d54_24;
	wire [WIDTH-1:0] wire_d54_25;
	wire [WIDTH-1:0] wire_d54_26;
	wire [WIDTH-1:0] wire_d54_27;
	wire [WIDTH-1:0] wire_d54_28;
	wire [WIDTH-1:0] wire_d54_29;
	wire [WIDTH-1:0] wire_d54_30;
	wire [WIDTH-1:0] wire_d54_31;
	wire [WIDTH-1:0] wire_d54_32;
	wire [WIDTH-1:0] wire_d54_33;
	wire [WIDTH-1:0] wire_d54_34;
	wire [WIDTH-1:0] wire_d54_35;
	wire [WIDTH-1:0] wire_d54_36;
	wire [WIDTH-1:0] wire_d54_37;
	wire [WIDTH-1:0] wire_d54_38;
	wire [WIDTH-1:0] wire_d54_39;
	wire [WIDTH-1:0] wire_d54_40;
	wire [WIDTH-1:0] wire_d54_41;
	wire [WIDTH-1:0] wire_d54_42;
	wire [WIDTH-1:0] wire_d54_43;
	wire [WIDTH-1:0] wire_d54_44;
	wire [WIDTH-1:0] wire_d54_45;
	wire [WIDTH-1:0] wire_d54_46;
	wire [WIDTH-1:0] wire_d54_47;
	wire [WIDTH-1:0] wire_d54_48;
	wire [WIDTH-1:0] wire_d54_49;
	wire [WIDTH-1:0] wire_d54_50;
	wire [WIDTH-1:0] wire_d54_51;
	wire [WIDTH-1:0] wire_d54_52;
	wire [WIDTH-1:0] wire_d54_53;
	wire [WIDTH-1:0] wire_d54_54;
	wire [WIDTH-1:0] wire_d54_55;
	wire [WIDTH-1:0] wire_d54_56;
	wire [WIDTH-1:0] wire_d54_57;
	wire [WIDTH-1:0] wire_d54_58;
	wire [WIDTH-1:0] wire_d54_59;
	wire [WIDTH-1:0] wire_d54_60;
	wire [WIDTH-1:0] wire_d54_61;
	wire [WIDTH-1:0] wire_d54_62;
	wire [WIDTH-1:0] wire_d54_63;
	wire [WIDTH-1:0] wire_d54_64;
	wire [WIDTH-1:0] wire_d54_65;
	wire [WIDTH-1:0] wire_d54_66;
	wire [WIDTH-1:0] wire_d54_67;
	wire [WIDTH-1:0] wire_d54_68;
	wire [WIDTH-1:0] wire_d54_69;
	wire [WIDTH-1:0] wire_d54_70;
	wire [WIDTH-1:0] wire_d54_71;
	wire [WIDTH-1:0] wire_d54_72;
	wire [WIDTH-1:0] wire_d54_73;
	wire [WIDTH-1:0] wire_d54_74;
	wire [WIDTH-1:0] wire_d54_75;
	wire [WIDTH-1:0] wire_d54_76;
	wire [WIDTH-1:0] wire_d54_77;
	wire [WIDTH-1:0] wire_d54_78;
	wire [WIDTH-1:0] wire_d54_79;
	wire [WIDTH-1:0] wire_d54_80;
	wire [WIDTH-1:0] wire_d54_81;
	wire [WIDTH-1:0] wire_d54_82;
	wire [WIDTH-1:0] wire_d54_83;
	wire [WIDTH-1:0] wire_d54_84;
	wire [WIDTH-1:0] wire_d54_85;
	wire [WIDTH-1:0] wire_d54_86;
	wire [WIDTH-1:0] wire_d54_87;
	wire [WIDTH-1:0] wire_d54_88;
	wire [WIDTH-1:0] wire_d54_89;
	wire [WIDTH-1:0] wire_d54_90;
	wire [WIDTH-1:0] wire_d54_91;
	wire [WIDTH-1:0] wire_d54_92;
	wire [WIDTH-1:0] wire_d54_93;
	wire [WIDTH-1:0] wire_d54_94;
	wire [WIDTH-1:0] wire_d54_95;
	wire [WIDTH-1:0] wire_d54_96;
	wire [WIDTH-1:0] wire_d54_97;
	wire [WIDTH-1:0] wire_d54_98;
	wire [WIDTH-1:0] wire_d54_99;
	wire [WIDTH-1:0] wire_d54_100;
	wire [WIDTH-1:0] wire_d54_101;
	wire [WIDTH-1:0] wire_d54_102;
	wire [WIDTH-1:0] wire_d54_103;
	wire [WIDTH-1:0] wire_d54_104;
	wire [WIDTH-1:0] wire_d54_105;
	wire [WIDTH-1:0] wire_d54_106;
	wire [WIDTH-1:0] wire_d54_107;
	wire [WIDTH-1:0] wire_d54_108;
	wire [WIDTH-1:0] wire_d54_109;
	wire [WIDTH-1:0] wire_d54_110;
	wire [WIDTH-1:0] wire_d54_111;
	wire [WIDTH-1:0] wire_d54_112;
	wire [WIDTH-1:0] wire_d54_113;
	wire [WIDTH-1:0] wire_d54_114;
	wire [WIDTH-1:0] wire_d54_115;
	wire [WIDTH-1:0] wire_d54_116;
	wire [WIDTH-1:0] wire_d54_117;
	wire [WIDTH-1:0] wire_d54_118;
	wire [WIDTH-1:0] wire_d55_0;
	wire [WIDTH-1:0] wire_d55_1;
	wire [WIDTH-1:0] wire_d55_2;
	wire [WIDTH-1:0] wire_d55_3;
	wire [WIDTH-1:0] wire_d55_4;
	wire [WIDTH-1:0] wire_d55_5;
	wire [WIDTH-1:0] wire_d55_6;
	wire [WIDTH-1:0] wire_d55_7;
	wire [WIDTH-1:0] wire_d55_8;
	wire [WIDTH-1:0] wire_d55_9;
	wire [WIDTH-1:0] wire_d55_10;
	wire [WIDTH-1:0] wire_d55_11;
	wire [WIDTH-1:0] wire_d55_12;
	wire [WIDTH-1:0] wire_d55_13;
	wire [WIDTH-1:0] wire_d55_14;
	wire [WIDTH-1:0] wire_d55_15;
	wire [WIDTH-1:0] wire_d55_16;
	wire [WIDTH-1:0] wire_d55_17;
	wire [WIDTH-1:0] wire_d55_18;
	wire [WIDTH-1:0] wire_d55_19;
	wire [WIDTH-1:0] wire_d55_20;
	wire [WIDTH-1:0] wire_d55_21;
	wire [WIDTH-1:0] wire_d55_22;
	wire [WIDTH-1:0] wire_d55_23;
	wire [WIDTH-1:0] wire_d55_24;
	wire [WIDTH-1:0] wire_d55_25;
	wire [WIDTH-1:0] wire_d55_26;
	wire [WIDTH-1:0] wire_d55_27;
	wire [WIDTH-1:0] wire_d55_28;
	wire [WIDTH-1:0] wire_d55_29;
	wire [WIDTH-1:0] wire_d55_30;
	wire [WIDTH-1:0] wire_d55_31;
	wire [WIDTH-1:0] wire_d55_32;
	wire [WIDTH-1:0] wire_d55_33;
	wire [WIDTH-1:0] wire_d55_34;
	wire [WIDTH-1:0] wire_d55_35;
	wire [WIDTH-1:0] wire_d55_36;
	wire [WIDTH-1:0] wire_d55_37;
	wire [WIDTH-1:0] wire_d55_38;
	wire [WIDTH-1:0] wire_d55_39;
	wire [WIDTH-1:0] wire_d55_40;
	wire [WIDTH-1:0] wire_d55_41;
	wire [WIDTH-1:0] wire_d55_42;
	wire [WIDTH-1:0] wire_d55_43;
	wire [WIDTH-1:0] wire_d55_44;
	wire [WIDTH-1:0] wire_d55_45;
	wire [WIDTH-1:0] wire_d55_46;
	wire [WIDTH-1:0] wire_d55_47;
	wire [WIDTH-1:0] wire_d55_48;
	wire [WIDTH-1:0] wire_d55_49;
	wire [WIDTH-1:0] wire_d55_50;
	wire [WIDTH-1:0] wire_d55_51;
	wire [WIDTH-1:0] wire_d55_52;
	wire [WIDTH-1:0] wire_d55_53;
	wire [WIDTH-1:0] wire_d55_54;
	wire [WIDTH-1:0] wire_d55_55;
	wire [WIDTH-1:0] wire_d55_56;
	wire [WIDTH-1:0] wire_d55_57;
	wire [WIDTH-1:0] wire_d55_58;
	wire [WIDTH-1:0] wire_d55_59;
	wire [WIDTH-1:0] wire_d55_60;
	wire [WIDTH-1:0] wire_d55_61;
	wire [WIDTH-1:0] wire_d55_62;
	wire [WIDTH-1:0] wire_d55_63;
	wire [WIDTH-1:0] wire_d55_64;
	wire [WIDTH-1:0] wire_d55_65;
	wire [WIDTH-1:0] wire_d55_66;
	wire [WIDTH-1:0] wire_d55_67;
	wire [WIDTH-1:0] wire_d55_68;
	wire [WIDTH-1:0] wire_d55_69;
	wire [WIDTH-1:0] wire_d55_70;
	wire [WIDTH-1:0] wire_d55_71;
	wire [WIDTH-1:0] wire_d55_72;
	wire [WIDTH-1:0] wire_d55_73;
	wire [WIDTH-1:0] wire_d55_74;
	wire [WIDTH-1:0] wire_d55_75;
	wire [WIDTH-1:0] wire_d55_76;
	wire [WIDTH-1:0] wire_d55_77;
	wire [WIDTH-1:0] wire_d55_78;
	wire [WIDTH-1:0] wire_d55_79;
	wire [WIDTH-1:0] wire_d55_80;
	wire [WIDTH-1:0] wire_d55_81;
	wire [WIDTH-1:0] wire_d55_82;
	wire [WIDTH-1:0] wire_d55_83;
	wire [WIDTH-1:0] wire_d55_84;
	wire [WIDTH-1:0] wire_d55_85;
	wire [WIDTH-1:0] wire_d55_86;
	wire [WIDTH-1:0] wire_d55_87;
	wire [WIDTH-1:0] wire_d55_88;
	wire [WIDTH-1:0] wire_d55_89;
	wire [WIDTH-1:0] wire_d55_90;
	wire [WIDTH-1:0] wire_d55_91;
	wire [WIDTH-1:0] wire_d55_92;
	wire [WIDTH-1:0] wire_d55_93;
	wire [WIDTH-1:0] wire_d55_94;
	wire [WIDTH-1:0] wire_d55_95;
	wire [WIDTH-1:0] wire_d55_96;
	wire [WIDTH-1:0] wire_d55_97;
	wire [WIDTH-1:0] wire_d55_98;
	wire [WIDTH-1:0] wire_d55_99;
	wire [WIDTH-1:0] wire_d55_100;
	wire [WIDTH-1:0] wire_d55_101;
	wire [WIDTH-1:0] wire_d55_102;
	wire [WIDTH-1:0] wire_d55_103;
	wire [WIDTH-1:0] wire_d55_104;
	wire [WIDTH-1:0] wire_d55_105;
	wire [WIDTH-1:0] wire_d55_106;
	wire [WIDTH-1:0] wire_d55_107;
	wire [WIDTH-1:0] wire_d55_108;
	wire [WIDTH-1:0] wire_d55_109;
	wire [WIDTH-1:0] wire_d55_110;
	wire [WIDTH-1:0] wire_d55_111;
	wire [WIDTH-1:0] wire_d55_112;
	wire [WIDTH-1:0] wire_d55_113;
	wire [WIDTH-1:0] wire_d55_114;
	wire [WIDTH-1:0] wire_d55_115;
	wire [WIDTH-1:0] wire_d55_116;
	wire [WIDTH-1:0] wire_d55_117;
	wire [WIDTH-1:0] wire_d55_118;
	wire [WIDTH-1:0] wire_d56_0;
	wire [WIDTH-1:0] wire_d56_1;
	wire [WIDTH-1:0] wire_d56_2;
	wire [WIDTH-1:0] wire_d56_3;
	wire [WIDTH-1:0] wire_d56_4;
	wire [WIDTH-1:0] wire_d56_5;
	wire [WIDTH-1:0] wire_d56_6;
	wire [WIDTH-1:0] wire_d56_7;
	wire [WIDTH-1:0] wire_d56_8;
	wire [WIDTH-1:0] wire_d56_9;
	wire [WIDTH-1:0] wire_d56_10;
	wire [WIDTH-1:0] wire_d56_11;
	wire [WIDTH-1:0] wire_d56_12;
	wire [WIDTH-1:0] wire_d56_13;
	wire [WIDTH-1:0] wire_d56_14;
	wire [WIDTH-1:0] wire_d56_15;
	wire [WIDTH-1:0] wire_d56_16;
	wire [WIDTH-1:0] wire_d56_17;
	wire [WIDTH-1:0] wire_d56_18;
	wire [WIDTH-1:0] wire_d56_19;
	wire [WIDTH-1:0] wire_d56_20;
	wire [WIDTH-1:0] wire_d56_21;
	wire [WIDTH-1:0] wire_d56_22;
	wire [WIDTH-1:0] wire_d56_23;
	wire [WIDTH-1:0] wire_d56_24;
	wire [WIDTH-1:0] wire_d56_25;
	wire [WIDTH-1:0] wire_d56_26;
	wire [WIDTH-1:0] wire_d56_27;
	wire [WIDTH-1:0] wire_d56_28;
	wire [WIDTH-1:0] wire_d56_29;
	wire [WIDTH-1:0] wire_d56_30;
	wire [WIDTH-1:0] wire_d56_31;
	wire [WIDTH-1:0] wire_d56_32;
	wire [WIDTH-1:0] wire_d56_33;
	wire [WIDTH-1:0] wire_d56_34;
	wire [WIDTH-1:0] wire_d56_35;
	wire [WIDTH-1:0] wire_d56_36;
	wire [WIDTH-1:0] wire_d56_37;
	wire [WIDTH-1:0] wire_d56_38;
	wire [WIDTH-1:0] wire_d56_39;
	wire [WIDTH-1:0] wire_d56_40;
	wire [WIDTH-1:0] wire_d56_41;
	wire [WIDTH-1:0] wire_d56_42;
	wire [WIDTH-1:0] wire_d56_43;
	wire [WIDTH-1:0] wire_d56_44;
	wire [WIDTH-1:0] wire_d56_45;
	wire [WIDTH-1:0] wire_d56_46;
	wire [WIDTH-1:0] wire_d56_47;
	wire [WIDTH-1:0] wire_d56_48;
	wire [WIDTH-1:0] wire_d56_49;
	wire [WIDTH-1:0] wire_d56_50;
	wire [WIDTH-1:0] wire_d56_51;
	wire [WIDTH-1:0] wire_d56_52;
	wire [WIDTH-1:0] wire_d56_53;
	wire [WIDTH-1:0] wire_d56_54;
	wire [WIDTH-1:0] wire_d56_55;
	wire [WIDTH-1:0] wire_d56_56;
	wire [WIDTH-1:0] wire_d56_57;
	wire [WIDTH-1:0] wire_d56_58;
	wire [WIDTH-1:0] wire_d56_59;
	wire [WIDTH-1:0] wire_d56_60;
	wire [WIDTH-1:0] wire_d56_61;
	wire [WIDTH-1:0] wire_d56_62;
	wire [WIDTH-1:0] wire_d56_63;
	wire [WIDTH-1:0] wire_d56_64;
	wire [WIDTH-1:0] wire_d56_65;
	wire [WIDTH-1:0] wire_d56_66;
	wire [WIDTH-1:0] wire_d56_67;
	wire [WIDTH-1:0] wire_d56_68;
	wire [WIDTH-1:0] wire_d56_69;
	wire [WIDTH-1:0] wire_d56_70;
	wire [WIDTH-1:0] wire_d56_71;
	wire [WIDTH-1:0] wire_d56_72;
	wire [WIDTH-1:0] wire_d56_73;
	wire [WIDTH-1:0] wire_d56_74;
	wire [WIDTH-1:0] wire_d56_75;
	wire [WIDTH-1:0] wire_d56_76;
	wire [WIDTH-1:0] wire_d56_77;
	wire [WIDTH-1:0] wire_d56_78;
	wire [WIDTH-1:0] wire_d56_79;
	wire [WIDTH-1:0] wire_d56_80;
	wire [WIDTH-1:0] wire_d56_81;
	wire [WIDTH-1:0] wire_d56_82;
	wire [WIDTH-1:0] wire_d56_83;
	wire [WIDTH-1:0] wire_d56_84;
	wire [WIDTH-1:0] wire_d56_85;
	wire [WIDTH-1:0] wire_d56_86;
	wire [WIDTH-1:0] wire_d56_87;
	wire [WIDTH-1:0] wire_d56_88;
	wire [WIDTH-1:0] wire_d56_89;
	wire [WIDTH-1:0] wire_d56_90;
	wire [WIDTH-1:0] wire_d56_91;
	wire [WIDTH-1:0] wire_d56_92;
	wire [WIDTH-1:0] wire_d56_93;
	wire [WIDTH-1:0] wire_d56_94;
	wire [WIDTH-1:0] wire_d56_95;
	wire [WIDTH-1:0] wire_d56_96;
	wire [WIDTH-1:0] wire_d56_97;
	wire [WIDTH-1:0] wire_d56_98;
	wire [WIDTH-1:0] wire_d56_99;
	wire [WIDTH-1:0] wire_d56_100;
	wire [WIDTH-1:0] wire_d56_101;
	wire [WIDTH-1:0] wire_d56_102;
	wire [WIDTH-1:0] wire_d56_103;
	wire [WIDTH-1:0] wire_d56_104;
	wire [WIDTH-1:0] wire_d56_105;
	wire [WIDTH-1:0] wire_d56_106;
	wire [WIDTH-1:0] wire_d56_107;
	wire [WIDTH-1:0] wire_d56_108;
	wire [WIDTH-1:0] wire_d56_109;
	wire [WIDTH-1:0] wire_d56_110;
	wire [WIDTH-1:0] wire_d56_111;
	wire [WIDTH-1:0] wire_d56_112;
	wire [WIDTH-1:0] wire_d56_113;
	wire [WIDTH-1:0] wire_d56_114;
	wire [WIDTH-1:0] wire_d56_115;
	wire [WIDTH-1:0] wire_d56_116;
	wire [WIDTH-1:0] wire_d56_117;
	wire [WIDTH-1:0] wire_d56_118;
	wire [WIDTH-1:0] wire_d57_0;
	wire [WIDTH-1:0] wire_d57_1;
	wire [WIDTH-1:0] wire_d57_2;
	wire [WIDTH-1:0] wire_d57_3;
	wire [WIDTH-1:0] wire_d57_4;
	wire [WIDTH-1:0] wire_d57_5;
	wire [WIDTH-1:0] wire_d57_6;
	wire [WIDTH-1:0] wire_d57_7;
	wire [WIDTH-1:0] wire_d57_8;
	wire [WIDTH-1:0] wire_d57_9;
	wire [WIDTH-1:0] wire_d57_10;
	wire [WIDTH-1:0] wire_d57_11;
	wire [WIDTH-1:0] wire_d57_12;
	wire [WIDTH-1:0] wire_d57_13;
	wire [WIDTH-1:0] wire_d57_14;
	wire [WIDTH-1:0] wire_d57_15;
	wire [WIDTH-1:0] wire_d57_16;
	wire [WIDTH-1:0] wire_d57_17;
	wire [WIDTH-1:0] wire_d57_18;
	wire [WIDTH-1:0] wire_d57_19;
	wire [WIDTH-1:0] wire_d57_20;
	wire [WIDTH-1:0] wire_d57_21;
	wire [WIDTH-1:0] wire_d57_22;
	wire [WIDTH-1:0] wire_d57_23;
	wire [WIDTH-1:0] wire_d57_24;
	wire [WIDTH-1:0] wire_d57_25;
	wire [WIDTH-1:0] wire_d57_26;
	wire [WIDTH-1:0] wire_d57_27;
	wire [WIDTH-1:0] wire_d57_28;
	wire [WIDTH-1:0] wire_d57_29;
	wire [WIDTH-1:0] wire_d57_30;
	wire [WIDTH-1:0] wire_d57_31;
	wire [WIDTH-1:0] wire_d57_32;
	wire [WIDTH-1:0] wire_d57_33;
	wire [WIDTH-1:0] wire_d57_34;
	wire [WIDTH-1:0] wire_d57_35;
	wire [WIDTH-1:0] wire_d57_36;
	wire [WIDTH-1:0] wire_d57_37;
	wire [WIDTH-1:0] wire_d57_38;
	wire [WIDTH-1:0] wire_d57_39;
	wire [WIDTH-1:0] wire_d57_40;
	wire [WIDTH-1:0] wire_d57_41;
	wire [WIDTH-1:0] wire_d57_42;
	wire [WIDTH-1:0] wire_d57_43;
	wire [WIDTH-1:0] wire_d57_44;
	wire [WIDTH-1:0] wire_d57_45;
	wire [WIDTH-1:0] wire_d57_46;
	wire [WIDTH-1:0] wire_d57_47;
	wire [WIDTH-1:0] wire_d57_48;
	wire [WIDTH-1:0] wire_d57_49;
	wire [WIDTH-1:0] wire_d57_50;
	wire [WIDTH-1:0] wire_d57_51;
	wire [WIDTH-1:0] wire_d57_52;
	wire [WIDTH-1:0] wire_d57_53;
	wire [WIDTH-1:0] wire_d57_54;
	wire [WIDTH-1:0] wire_d57_55;
	wire [WIDTH-1:0] wire_d57_56;
	wire [WIDTH-1:0] wire_d57_57;
	wire [WIDTH-1:0] wire_d57_58;
	wire [WIDTH-1:0] wire_d57_59;
	wire [WIDTH-1:0] wire_d57_60;
	wire [WIDTH-1:0] wire_d57_61;
	wire [WIDTH-1:0] wire_d57_62;
	wire [WIDTH-1:0] wire_d57_63;
	wire [WIDTH-1:0] wire_d57_64;
	wire [WIDTH-1:0] wire_d57_65;
	wire [WIDTH-1:0] wire_d57_66;
	wire [WIDTH-1:0] wire_d57_67;
	wire [WIDTH-1:0] wire_d57_68;
	wire [WIDTH-1:0] wire_d57_69;
	wire [WIDTH-1:0] wire_d57_70;
	wire [WIDTH-1:0] wire_d57_71;
	wire [WIDTH-1:0] wire_d57_72;
	wire [WIDTH-1:0] wire_d57_73;
	wire [WIDTH-1:0] wire_d57_74;
	wire [WIDTH-1:0] wire_d57_75;
	wire [WIDTH-1:0] wire_d57_76;
	wire [WIDTH-1:0] wire_d57_77;
	wire [WIDTH-1:0] wire_d57_78;
	wire [WIDTH-1:0] wire_d57_79;
	wire [WIDTH-1:0] wire_d57_80;
	wire [WIDTH-1:0] wire_d57_81;
	wire [WIDTH-1:0] wire_d57_82;
	wire [WIDTH-1:0] wire_d57_83;
	wire [WIDTH-1:0] wire_d57_84;
	wire [WIDTH-1:0] wire_d57_85;
	wire [WIDTH-1:0] wire_d57_86;
	wire [WIDTH-1:0] wire_d57_87;
	wire [WIDTH-1:0] wire_d57_88;
	wire [WIDTH-1:0] wire_d57_89;
	wire [WIDTH-1:0] wire_d57_90;
	wire [WIDTH-1:0] wire_d57_91;
	wire [WIDTH-1:0] wire_d57_92;
	wire [WIDTH-1:0] wire_d57_93;
	wire [WIDTH-1:0] wire_d57_94;
	wire [WIDTH-1:0] wire_d57_95;
	wire [WIDTH-1:0] wire_d57_96;
	wire [WIDTH-1:0] wire_d57_97;
	wire [WIDTH-1:0] wire_d57_98;
	wire [WIDTH-1:0] wire_d57_99;
	wire [WIDTH-1:0] wire_d57_100;
	wire [WIDTH-1:0] wire_d57_101;
	wire [WIDTH-1:0] wire_d57_102;
	wire [WIDTH-1:0] wire_d57_103;
	wire [WIDTH-1:0] wire_d57_104;
	wire [WIDTH-1:0] wire_d57_105;
	wire [WIDTH-1:0] wire_d57_106;
	wire [WIDTH-1:0] wire_d57_107;
	wire [WIDTH-1:0] wire_d57_108;
	wire [WIDTH-1:0] wire_d57_109;
	wire [WIDTH-1:0] wire_d57_110;
	wire [WIDTH-1:0] wire_d57_111;
	wire [WIDTH-1:0] wire_d57_112;
	wire [WIDTH-1:0] wire_d57_113;
	wire [WIDTH-1:0] wire_d57_114;
	wire [WIDTH-1:0] wire_d57_115;
	wire [WIDTH-1:0] wire_d57_116;
	wire [WIDTH-1:0] wire_d57_117;
	wire [WIDTH-1:0] wire_d57_118;
	wire [WIDTH-1:0] wire_d58_0;
	wire [WIDTH-1:0] wire_d58_1;
	wire [WIDTH-1:0] wire_d58_2;
	wire [WIDTH-1:0] wire_d58_3;
	wire [WIDTH-1:0] wire_d58_4;
	wire [WIDTH-1:0] wire_d58_5;
	wire [WIDTH-1:0] wire_d58_6;
	wire [WIDTH-1:0] wire_d58_7;
	wire [WIDTH-1:0] wire_d58_8;
	wire [WIDTH-1:0] wire_d58_9;
	wire [WIDTH-1:0] wire_d58_10;
	wire [WIDTH-1:0] wire_d58_11;
	wire [WIDTH-1:0] wire_d58_12;
	wire [WIDTH-1:0] wire_d58_13;
	wire [WIDTH-1:0] wire_d58_14;
	wire [WIDTH-1:0] wire_d58_15;
	wire [WIDTH-1:0] wire_d58_16;
	wire [WIDTH-1:0] wire_d58_17;
	wire [WIDTH-1:0] wire_d58_18;
	wire [WIDTH-1:0] wire_d58_19;
	wire [WIDTH-1:0] wire_d58_20;
	wire [WIDTH-1:0] wire_d58_21;
	wire [WIDTH-1:0] wire_d58_22;
	wire [WIDTH-1:0] wire_d58_23;
	wire [WIDTH-1:0] wire_d58_24;
	wire [WIDTH-1:0] wire_d58_25;
	wire [WIDTH-1:0] wire_d58_26;
	wire [WIDTH-1:0] wire_d58_27;
	wire [WIDTH-1:0] wire_d58_28;
	wire [WIDTH-1:0] wire_d58_29;
	wire [WIDTH-1:0] wire_d58_30;
	wire [WIDTH-1:0] wire_d58_31;
	wire [WIDTH-1:0] wire_d58_32;
	wire [WIDTH-1:0] wire_d58_33;
	wire [WIDTH-1:0] wire_d58_34;
	wire [WIDTH-1:0] wire_d58_35;
	wire [WIDTH-1:0] wire_d58_36;
	wire [WIDTH-1:0] wire_d58_37;
	wire [WIDTH-1:0] wire_d58_38;
	wire [WIDTH-1:0] wire_d58_39;
	wire [WIDTH-1:0] wire_d58_40;
	wire [WIDTH-1:0] wire_d58_41;
	wire [WIDTH-1:0] wire_d58_42;
	wire [WIDTH-1:0] wire_d58_43;
	wire [WIDTH-1:0] wire_d58_44;
	wire [WIDTH-1:0] wire_d58_45;
	wire [WIDTH-1:0] wire_d58_46;
	wire [WIDTH-1:0] wire_d58_47;
	wire [WIDTH-1:0] wire_d58_48;
	wire [WIDTH-1:0] wire_d58_49;
	wire [WIDTH-1:0] wire_d58_50;
	wire [WIDTH-1:0] wire_d58_51;
	wire [WIDTH-1:0] wire_d58_52;
	wire [WIDTH-1:0] wire_d58_53;
	wire [WIDTH-1:0] wire_d58_54;
	wire [WIDTH-1:0] wire_d58_55;
	wire [WIDTH-1:0] wire_d58_56;
	wire [WIDTH-1:0] wire_d58_57;
	wire [WIDTH-1:0] wire_d58_58;
	wire [WIDTH-1:0] wire_d58_59;
	wire [WIDTH-1:0] wire_d58_60;
	wire [WIDTH-1:0] wire_d58_61;
	wire [WIDTH-1:0] wire_d58_62;
	wire [WIDTH-1:0] wire_d58_63;
	wire [WIDTH-1:0] wire_d58_64;
	wire [WIDTH-1:0] wire_d58_65;
	wire [WIDTH-1:0] wire_d58_66;
	wire [WIDTH-1:0] wire_d58_67;
	wire [WIDTH-1:0] wire_d58_68;
	wire [WIDTH-1:0] wire_d58_69;
	wire [WIDTH-1:0] wire_d58_70;
	wire [WIDTH-1:0] wire_d58_71;
	wire [WIDTH-1:0] wire_d58_72;
	wire [WIDTH-1:0] wire_d58_73;
	wire [WIDTH-1:0] wire_d58_74;
	wire [WIDTH-1:0] wire_d58_75;
	wire [WIDTH-1:0] wire_d58_76;
	wire [WIDTH-1:0] wire_d58_77;
	wire [WIDTH-1:0] wire_d58_78;
	wire [WIDTH-1:0] wire_d58_79;
	wire [WIDTH-1:0] wire_d58_80;
	wire [WIDTH-1:0] wire_d58_81;
	wire [WIDTH-1:0] wire_d58_82;
	wire [WIDTH-1:0] wire_d58_83;
	wire [WIDTH-1:0] wire_d58_84;
	wire [WIDTH-1:0] wire_d58_85;
	wire [WIDTH-1:0] wire_d58_86;
	wire [WIDTH-1:0] wire_d58_87;
	wire [WIDTH-1:0] wire_d58_88;
	wire [WIDTH-1:0] wire_d58_89;
	wire [WIDTH-1:0] wire_d58_90;
	wire [WIDTH-1:0] wire_d58_91;
	wire [WIDTH-1:0] wire_d58_92;
	wire [WIDTH-1:0] wire_d58_93;
	wire [WIDTH-1:0] wire_d58_94;
	wire [WIDTH-1:0] wire_d58_95;
	wire [WIDTH-1:0] wire_d58_96;
	wire [WIDTH-1:0] wire_d58_97;
	wire [WIDTH-1:0] wire_d58_98;
	wire [WIDTH-1:0] wire_d58_99;
	wire [WIDTH-1:0] wire_d58_100;
	wire [WIDTH-1:0] wire_d58_101;
	wire [WIDTH-1:0] wire_d58_102;
	wire [WIDTH-1:0] wire_d58_103;
	wire [WIDTH-1:0] wire_d58_104;
	wire [WIDTH-1:0] wire_d58_105;
	wire [WIDTH-1:0] wire_d58_106;
	wire [WIDTH-1:0] wire_d58_107;
	wire [WIDTH-1:0] wire_d58_108;
	wire [WIDTH-1:0] wire_d58_109;
	wire [WIDTH-1:0] wire_d58_110;
	wire [WIDTH-1:0] wire_d58_111;
	wire [WIDTH-1:0] wire_d58_112;
	wire [WIDTH-1:0] wire_d58_113;
	wire [WIDTH-1:0] wire_d58_114;
	wire [WIDTH-1:0] wire_d58_115;
	wire [WIDTH-1:0] wire_d58_116;
	wire [WIDTH-1:0] wire_d58_117;
	wire [WIDTH-1:0] wire_d58_118;
	wire [WIDTH-1:0] wire_d59_0;
	wire [WIDTH-1:0] wire_d59_1;
	wire [WIDTH-1:0] wire_d59_2;
	wire [WIDTH-1:0] wire_d59_3;
	wire [WIDTH-1:0] wire_d59_4;
	wire [WIDTH-1:0] wire_d59_5;
	wire [WIDTH-1:0] wire_d59_6;
	wire [WIDTH-1:0] wire_d59_7;
	wire [WIDTH-1:0] wire_d59_8;
	wire [WIDTH-1:0] wire_d59_9;
	wire [WIDTH-1:0] wire_d59_10;
	wire [WIDTH-1:0] wire_d59_11;
	wire [WIDTH-1:0] wire_d59_12;
	wire [WIDTH-1:0] wire_d59_13;
	wire [WIDTH-1:0] wire_d59_14;
	wire [WIDTH-1:0] wire_d59_15;
	wire [WIDTH-1:0] wire_d59_16;
	wire [WIDTH-1:0] wire_d59_17;
	wire [WIDTH-1:0] wire_d59_18;
	wire [WIDTH-1:0] wire_d59_19;
	wire [WIDTH-1:0] wire_d59_20;
	wire [WIDTH-1:0] wire_d59_21;
	wire [WIDTH-1:0] wire_d59_22;
	wire [WIDTH-1:0] wire_d59_23;
	wire [WIDTH-1:0] wire_d59_24;
	wire [WIDTH-1:0] wire_d59_25;
	wire [WIDTH-1:0] wire_d59_26;
	wire [WIDTH-1:0] wire_d59_27;
	wire [WIDTH-1:0] wire_d59_28;
	wire [WIDTH-1:0] wire_d59_29;
	wire [WIDTH-1:0] wire_d59_30;
	wire [WIDTH-1:0] wire_d59_31;
	wire [WIDTH-1:0] wire_d59_32;
	wire [WIDTH-1:0] wire_d59_33;
	wire [WIDTH-1:0] wire_d59_34;
	wire [WIDTH-1:0] wire_d59_35;
	wire [WIDTH-1:0] wire_d59_36;
	wire [WIDTH-1:0] wire_d59_37;
	wire [WIDTH-1:0] wire_d59_38;
	wire [WIDTH-1:0] wire_d59_39;
	wire [WIDTH-1:0] wire_d59_40;
	wire [WIDTH-1:0] wire_d59_41;
	wire [WIDTH-1:0] wire_d59_42;
	wire [WIDTH-1:0] wire_d59_43;
	wire [WIDTH-1:0] wire_d59_44;
	wire [WIDTH-1:0] wire_d59_45;
	wire [WIDTH-1:0] wire_d59_46;
	wire [WIDTH-1:0] wire_d59_47;
	wire [WIDTH-1:0] wire_d59_48;
	wire [WIDTH-1:0] wire_d59_49;
	wire [WIDTH-1:0] wire_d59_50;
	wire [WIDTH-1:0] wire_d59_51;
	wire [WIDTH-1:0] wire_d59_52;
	wire [WIDTH-1:0] wire_d59_53;
	wire [WIDTH-1:0] wire_d59_54;
	wire [WIDTH-1:0] wire_d59_55;
	wire [WIDTH-1:0] wire_d59_56;
	wire [WIDTH-1:0] wire_d59_57;
	wire [WIDTH-1:0] wire_d59_58;
	wire [WIDTH-1:0] wire_d59_59;
	wire [WIDTH-1:0] wire_d59_60;
	wire [WIDTH-1:0] wire_d59_61;
	wire [WIDTH-1:0] wire_d59_62;
	wire [WIDTH-1:0] wire_d59_63;
	wire [WIDTH-1:0] wire_d59_64;
	wire [WIDTH-1:0] wire_d59_65;
	wire [WIDTH-1:0] wire_d59_66;
	wire [WIDTH-1:0] wire_d59_67;
	wire [WIDTH-1:0] wire_d59_68;
	wire [WIDTH-1:0] wire_d59_69;
	wire [WIDTH-1:0] wire_d59_70;
	wire [WIDTH-1:0] wire_d59_71;
	wire [WIDTH-1:0] wire_d59_72;
	wire [WIDTH-1:0] wire_d59_73;
	wire [WIDTH-1:0] wire_d59_74;
	wire [WIDTH-1:0] wire_d59_75;
	wire [WIDTH-1:0] wire_d59_76;
	wire [WIDTH-1:0] wire_d59_77;
	wire [WIDTH-1:0] wire_d59_78;
	wire [WIDTH-1:0] wire_d59_79;
	wire [WIDTH-1:0] wire_d59_80;
	wire [WIDTH-1:0] wire_d59_81;
	wire [WIDTH-1:0] wire_d59_82;
	wire [WIDTH-1:0] wire_d59_83;
	wire [WIDTH-1:0] wire_d59_84;
	wire [WIDTH-1:0] wire_d59_85;
	wire [WIDTH-1:0] wire_d59_86;
	wire [WIDTH-1:0] wire_d59_87;
	wire [WIDTH-1:0] wire_d59_88;
	wire [WIDTH-1:0] wire_d59_89;
	wire [WIDTH-1:0] wire_d59_90;
	wire [WIDTH-1:0] wire_d59_91;
	wire [WIDTH-1:0] wire_d59_92;
	wire [WIDTH-1:0] wire_d59_93;
	wire [WIDTH-1:0] wire_d59_94;
	wire [WIDTH-1:0] wire_d59_95;
	wire [WIDTH-1:0] wire_d59_96;
	wire [WIDTH-1:0] wire_d59_97;
	wire [WIDTH-1:0] wire_d59_98;
	wire [WIDTH-1:0] wire_d59_99;
	wire [WIDTH-1:0] wire_d59_100;
	wire [WIDTH-1:0] wire_d59_101;
	wire [WIDTH-1:0] wire_d59_102;
	wire [WIDTH-1:0] wire_d59_103;
	wire [WIDTH-1:0] wire_d59_104;
	wire [WIDTH-1:0] wire_d59_105;
	wire [WIDTH-1:0] wire_d59_106;
	wire [WIDTH-1:0] wire_d59_107;
	wire [WIDTH-1:0] wire_d59_108;
	wire [WIDTH-1:0] wire_d59_109;
	wire [WIDTH-1:0] wire_d59_110;
	wire [WIDTH-1:0] wire_d59_111;
	wire [WIDTH-1:0] wire_d59_112;
	wire [WIDTH-1:0] wire_d59_113;
	wire [WIDTH-1:0] wire_d59_114;
	wire [WIDTH-1:0] wire_d59_115;
	wire [WIDTH-1:0] wire_d59_116;
	wire [WIDTH-1:0] wire_d59_117;
	wire [WIDTH-1:0] wire_d59_118;
	wire [WIDTH-1:0] wire_d60_0;
	wire [WIDTH-1:0] wire_d60_1;
	wire [WIDTH-1:0] wire_d60_2;
	wire [WIDTH-1:0] wire_d60_3;
	wire [WIDTH-1:0] wire_d60_4;
	wire [WIDTH-1:0] wire_d60_5;
	wire [WIDTH-1:0] wire_d60_6;
	wire [WIDTH-1:0] wire_d60_7;
	wire [WIDTH-1:0] wire_d60_8;
	wire [WIDTH-1:0] wire_d60_9;
	wire [WIDTH-1:0] wire_d60_10;
	wire [WIDTH-1:0] wire_d60_11;
	wire [WIDTH-1:0] wire_d60_12;
	wire [WIDTH-1:0] wire_d60_13;
	wire [WIDTH-1:0] wire_d60_14;
	wire [WIDTH-1:0] wire_d60_15;
	wire [WIDTH-1:0] wire_d60_16;
	wire [WIDTH-1:0] wire_d60_17;
	wire [WIDTH-1:0] wire_d60_18;
	wire [WIDTH-1:0] wire_d60_19;
	wire [WIDTH-1:0] wire_d60_20;
	wire [WIDTH-1:0] wire_d60_21;
	wire [WIDTH-1:0] wire_d60_22;
	wire [WIDTH-1:0] wire_d60_23;
	wire [WIDTH-1:0] wire_d60_24;
	wire [WIDTH-1:0] wire_d60_25;
	wire [WIDTH-1:0] wire_d60_26;
	wire [WIDTH-1:0] wire_d60_27;
	wire [WIDTH-1:0] wire_d60_28;
	wire [WIDTH-1:0] wire_d60_29;
	wire [WIDTH-1:0] wire_d60_30;
	wire [WIDTH-1:0] wire_d60_31;
	wire [WIDTH-1:0] wire_d60_32;
	wire [WIDTH-1:0] wire_d60_33;
	wire [WIDTH-1:0] wire_d60_34;
	wire [WIDTH-1:0] wire_d60_35;
	wire [WIDTH-1:0] wire_d60_36;
	wire [WIDTH-1:0] wire_d60_37;
	wire [WIDTH-1:0] wire_d60_38;
	wire [WIDTH-1:0] wire_d60_39;
	wire [WIDTH-1:0] wire_d60_40;
	wire [WIDTH-1:0] wire_d60_41;
	wire [WIDTH-1:0] wire_d60_42;
	wire [WIDTH-1:0] wire_d60_43;
	wire [WIDTH-1:0] wire_d60_44;
	wire [WIDTH-1:0] wire_d60_45;
	wire [WIDTH-1:0] wire_d60_46;
	wire [WIDTH-1:0] wire_d60_47;
	wire [WIDTH-1:0] wire_d60_48;
	wire [WIDTH-1:0] wire_d60_49;
	wire [WIDTH-1:0] wire_d60_50;
	wire [WIDTH-1:0] wire_d60_51;
	wire [WIDTH-1:0] wire_d60_52;
	wire [WIDTH-1:0] wire_d60_53;
	wire [WIDTH-1:0] wire_d60_54;
	wire [WIDTH-1:0] wire_d60_55;
	wire [WIDTH-1:0] wire_d60_56;
	wire [WIDTH-1:0] wire_d60_57;
	wire [WIDTH-1:0] wire_d60_58;
	wire [WIDTH-1:0] wire_d60_59;
	wire [WIDTH-1:0] wire_d60_60;
	wire [WIDTH-1:0] wire_d60_61;
	wire [WIDTH-1:0] wire_d60_62;
	wire [WIDTH-1:0] wire_d60_63;
	wire [WIDTH-1:0] wire_d60_64;
	wire [WIDTH-1:0] wire_d60_65;
	wire [WIDTH-1:0] wire_d60_66;
	wire [WIDTH-1:0] wire_d60_67;
	wire [WIDTH-1:0] wire_d60_68;
	wire [WIDTH-1:0] wire_d60_69;
	wire [WIDTH-1:0] wire_d60_70;
	wire [WIDTH-1:0] wire_d60_71;
	wire [WIDTH-1:0] wire_d60_72;
	wire [WIDTH-1:0] wire_d60_73;
	wire [WIDTH-1:0] wire_d60_74;
	wire [WIDTH-1:0] wire_d60_75;
	wire [WIDTH-1:0] wire_d60_76;
	wire [WIDTH-1:0] wire_d60_77;
	wire [WIDTH-1:0] wire_d60_78;
	wire [WIDTH-1:0] wire_d60_79;
	wire [WIDTH-1:0] wire_d60_80;
	wire [WIDTH-1:0] wire_d60_81;
	wire [WIDTH-1:0] wire_d60_82;
	wire [WIDTH-1:0] wire_d60_83;
	wire [WIDTH-1:0] wire_d60_84;
	wire [WIDTH-1:0] wire_d60_85;
	wire [WIDTH-1:0] wire_d60_86;
	wire [WIDTH-1:0] wire_d60_87;
	wire [WIDTH-1:0] wire_d60_88;
	wire [WIDTH-1:0] wire_d60_89;
	wire [WIDTH-1:0] wire_d60_90;
	wire [WIDTH-1:0] wire_d60_91;
	wire [WIDTH-1:0] wire_d60_92;
	wire [WIDTH-1:0] wire_d60_93;
	wire [WIDTH-1:0] wire_d60_94;
	wire [WIDTH-1:0] wire_d60_95;
	wire [WIDTH-1:0] wire_d60_96;
	wire [WIDTH-1:0] wire_d60_97;
	wire [WIDTH-1:0] wire_d60_98;
	wire [WIDTH-1:0] wire_d60_99;
	wire [WIDTH-1:0] wire_d60_100;
	wire [WIDTH-1:0] wire_d60_101;
	wire [WIDTH-1:0] wire_d60_102;
	wire [WIDTH-1:0] wire_d60_103;
	wire [WIDTH-1:0] wire_d60_104;
	wire [WIDTH-1:0] wire_d60_105;
	wire [WIDTH-1:0] wire_d60_106;
	wire [WIDTH-1:0] wire_d60_107;
	wire [WIDTH-1:0] wire_d60_108;
	wire [WIDTH-1:0] wire_d60_109;
	wire [WIDTH-1:0] wire_d60_110;
	wire [WIDTH-1:0] wire_d60_111;
	wire [WIDTH-1:0] wire_d60_112;
	wire [WIDTH-1:0] wire_d60_113;
	wire [WIDTH-1:0] wire_d60_114;
	wire [WIDTH-1:0] wire_d60_115;
	wire [WIDTH-1:0] wire_d60_116;
	wire [WIDTH-1:0] wire_d60_117;
	wire [WIDTH-1:0] wire_d60_118;
	wire [WIDTH-1:0] wire_d61_0;
	wire [WIDTH-1:0] wire_d61_1;
	wire [WIDTH-1:0] wire_d61_2;
	wire [WIDTH-1:0] wire_d61_3;
	wire [WIDTH-1:0] wire_d61_4;
	wire [WIDTH-1:0] wire_d61_5;
	wire [WIDTH-1:0] wire_d61_6;
	wire [WIDTH-1:0] wire_d61_7;
	wire [WIDTH-1:0] wire_d61_8;
	wire [WIDTH-1:0] wire_d61_9;
	wire [WIDTH-1:0] wire_d61_10;
	wire [WIDTH-1:0] wire_d61_11;
	wire [WIDTH-1:0] wire_d61_12;
	wire [WIDTH-1:0] wire_d61_13;
	wire [WIDTH-1:0] wire_d61_14;
	wire [WIDTH-1:0] wire_d61_15;
	wire [WIDTH-1:0] wire_d61_16;
	wire [WIDTH-1:0] wire_d61_17;
	wire [WIDTH-1:0] wire_d61_18;
	wire [WIDTH-1:0] wire_d61_19;
	wire [WIDTH-1:0] wire_d61_20;
	wire [WIDTH-1:0] wire_d61_21;
	wire [WIDTH-1:0] wire_d61_22;
	wire [WIDTH-1:0] wire_d61_23;
	wire [WIDTH-1:0] wire_d61_24;
	wire [WIDTH-1:0] wire_d61_25;
	wire [WIDTH-1:0] wire_d61_26;
	wire [WIDTH-1:0] wire_d61_27;
	wire [WIDTH-1:0] wire_d61_28;
	wire [WIDTH-1:0] wire_d61_29;
	wire [WIDTH-1:0] wire_d61_30;
	wire [WIDTH-1:0] wire_d61_31;
	wire [WIDTH-1:0] wire_d61_32;
	wire [WIDTH-1:0] wire_d61_33;
	wire [WIDTH-1:0] wire_d61_34;
	wire [WIDTH-1:0] wire_d61_35;
	wire [WIDTH-1:0] wire_d61_36;
	wire [WIDTH-1:0] wire_d61_37;
	wire [WIDTH-1:0] wire_d61_38;
	wire [WIDTH-1:0] wire_d61_39;
	wire [WIDTH-1:0] wire_d61_40;
	wire [WIDTH-1:0] wire_d61_41;
	wire [WIDTH-1:0] wire_d61_42;
	wire [WIDTH-1:0] wire_d61_43;
	wire [WIDTH-1:0] wire_d61_44;
	wire [WIDTH-1:0] wire_d61_45;
	wire [WIDTH-1:0] wire_d61_46;
	wire [WIDTH-1:0] wire_d61_47;
	wire [WIDTH-1:0] wire_d61_48;
	wire [WIDTH-1:0] wire_d61_49;
	wire [WIDTH-1:0] wire_d61_50;
	wire [WIDTH-1:0] wire_d61_51;
	wire [WIDTH-1:0] wire_d61_52;
	wire [WIDTH-1:0] wire_d61_53;
	wire [WIDTH-1:0] wire_d61_54;
	wire [WIDTH-1:0] wire_d61_55;
	wire [WIDTH-1:0] wire_d61_56;
	wire [WIDTH-1:0] wire_d61_57;
	wire [WIDTH-1:0] wire_d61_58;
	wire [WIDTH-1:0] wire_d61_59;
	wire [WIDTH-1:0] wire_d61_60;
	wire [WIDTH-1:0] wire_d61_61;
	wire [WIDTH-1:0] wire_d61_62;
	wire [WIDTH-1:0] wire_d61_63;
	wire [WIDTH-1:0] wire_d61_64;
	wire [WIDTH-1:0] wire_d61_65;
	wire [WIDTH-1:0] wire_d61_66;
	wire [WIDTH-1:0] wire_d61_67;
	wire [WIDTH-1:0] wire_d61_68;
	wire [WIDTH-1:0] wire_d61_69;
	wire [WIDTH-1:0] wire_d61_70;
	wire [WIDTH-1:0] wire_d61_71;
	wire [WIDTH-1:0] wire_d61_72;
	wire [WIDTH-1:0] wire_d61_73;
	wire [WIDTH-1:0] wire_d61_74;
	wire [WIDTH-1:0] wire_d61_75;
	wire [WIDTH-1:0] wire_d61_76;
	wire [WIDTH-1:0] wire_d61_77;
	wire [WIDTH-1:0] wire_d61_78;
	wire [WIDTH-1:0] wire_d61_79;
	wire [WIDTH-1:0] wire_d61_80;
	wire [WIDTH-1:0] wire_d61_81;
	wire [WIDTH-1:0] wire_d61_82;
	wire [WIDTH-1:0] wire_d61_83;
	wire [WIDTH-1:0] wire_d61_84;
	wire [WIDTH-1:0] wire_d61_85;
	wire [WIDTH-1:0] wire_d61_86;
	wire [WIDTH-1:0] wire_d61_87;
	wire [WIDTH-1:0] wire_d61_88;
	wire [WIDTH-1:0] wire_d61_89;
	wire [WIDTH-1:0] wire_d61_90;
	wire [WIDTH-1:0] wire_d61_91;
	wire [WIDTH-1:0] wire_d61_92;
	wire [WIDTH-1:0] wire_d61_93;
	wire [WIDTH-1:0] wire_d61_94;
	wire [WIDTH-1:0] wire_d61_95;
	wire [WIDTH-1:0] wire_d61_96;
	wire [WIDTH-1:0] wire_d61_97;
	wire [WIDTH-1:0] wire_d61_98;
	wire [WIDTH-1:0] wire_d61_99;
	wire [WIDTH-1:0] wire_d61_100;
	wire [WIDTH-1:0] wire_d61_101;
	wire [WIDTH-1:0] wire_d61_102;
	wire [WIDTH-1:0] wire_d61_103;
	wire [WIDTH-1:0] wire_d61_104;
	wire [WIDTH-1:0] wire_d61_105;
	wire [WIDTH-1:0] wire_d61_106;
	wire [WIDTH-1:0] wire_d61_107;
	wire [WIDTH-1:0] wire_d61_108;
	wire [WIDTH-1:0] wire_d61_109;
	wire [WIDTH-1:0] wire_d61_110;
	wire [WIDTH-1:0] wire_d61_111;
	wire [WIDTH-1:0] wire_d61_112;
	wire [WIDTH-1:0] wire_d61_113;
	wire [WIDTH-1:0] wire_d61_114;
	wire [WIDTH-1:0] wire_d61_115;
	wire [WIDTH-1:0] wire_d61_116;
	wire [WIDTH-1:0] wire_d61_117;
	wire [WIDTH-1:0] wire_d61_118;
	wire [WIDTH-1:0] wire_d62_0;
	wire [WIDTH-1:0] wire_d62_1;
	wire [WIDTH-1:0] wire_d62_2;
	wire [WIDTH-1:0] wire_d62_3;
	wire [WIDTH-1:0] wire_d62_4;
	wire [WIDTH-1:0] wire_d62_5;
	wire [WIDTH-1:0] wire_d62_6;
	wire [WIDTH-1:0] wire_d62_7;
	wire [WIDTH-1:0] wire_d62_8;
	wire [WIDTH-1:0] wire_d62_9;
	wire [WIDTH-1:0] wire_d62_10;
	wire [WIDTH-1:0] wire_d62_11;
	wire [WIDTH-1:0] wire_d62_12;
	wire [WIDTH-1:0] wire_d62_13;
	wire [WIDTH-1:0] wire_d62_14;
	wire [WIDTH-1:0] wire_d62_15;
	wire [WIDTH-1:0] wire_d62_16;
	wire [WIDTH-1:0] wire_d62_17;
	wire [WIDTH-1:0] wire_d62_18;
	wire [WIDTH-1:0] wire_d62_19;
	wire [WIDTH-1:0] wire_d62_20;
	wire [WIDTH-1:0] wire_d62_21;
	wire [WIDTH-1:0] wire_d62_22;
	wire [WIDTH-1:0] wire_d62_23;
	wire [WIDTH-1:0] wire_d62_24;
	wire [WIDTH-1:0] wire_d62_25;
	wire [WIDTH-1:0] wire_d62_26;
	wire [WIDTH-1:0] wire_d62_27;
	wire [WIDTH-1:0] wire_d62_28;
	wire [WIDTH-1:0] wire_d62_29;
	wire [WIDTH-1:0] wire_d62_30;
	wire [WIDTH-1:0] wire_d62_31;
	wire [WIDTH-1:0] wire_d62_32;
	wire [WIDTH-1:0] wire_d62_33;
	wire [WIDTH-1:0] wire_d62_34;
	wire [WIDTH-1:0] wire_d62_35;
	wire [WIDTH-1:0] wire_d62_36;
	wire [WIDTH-1:0] wire_d62_37;
	wire [WIDTH-1:0] wire_d62_38;
	wire [WIDTH-1:0] wire_d62_39;
	wire [WIDTH-1:0] wire_d62_40;
	wire [WIDTH-1:0] wire_d62_41;
	wire [WIDTH-1:0] wire_d62_42;
	wire [WIDTH-1:0] wire_d62_43;
	wire [WIDTH-1:0] wire_d62_44;
	wire [WIDTH-1:0] wire_d62_45;
	wire [WIDTH-1:0] wire_d62_46;
	wire [WIDTH-1:0] wire_d62_47;
	wire [WIDTH-1:0] wire_d62_48;
	wire [WIDTH-1:0] wire_d62_49;
	wire [WIDTH-1:0] wire_d62_50;
	wire [WIDTH-1:0] wire_d62_51;
	wire [WIDTH-1:0] wire_d62_52;
	wire [WIDTH-1:0] wire_d62_53;
	wire [WIDTH-1:0] wire_d62_54;
	wire [WIDTH-1:0] wire_d62_55;
	wire [WIDTH-1:0] wire_d62_56;
	wire [WIDTH-1:0] wire_d62_57;
	wire [WIDTH-1:0] wire_d62_58;
	wire [WIDTH-1:0] wire_d62_59;
	wire [WIDTH-1:0] wire_d62_60;
	wire [WIDTH-1:0] wire_d62_61;
	wire [WIDTH-1:0] wire_d62_62;
	wire [WIDTH-1:0] wire_d62_63;
	wire [WIDTH-1:0] wire_d62_64;
	wire [WIDTH-1:0] wire_d62_65;
	wire [WIDTH-1:0] wire_d62_66;
	wire [WIDTH-1:0] wire_d62_67;
	wire [WIDTH-1:0] wire_d62_68;
	wire [WIDTH-1:0] wire_d62_69;
	wire [WIDTH-1:0] wire_d62_70;
	wire [WIDTH-1:0] wire_d62_71;
	wire [WIDTH-1:0] wire_d62_72;
	wire [WIDTH-1:0] wire_d62_73;
	wire [WIDTH-1:0] wire_d62_74;
	wire [WIDTH-1:0] wire_d62_75;
	wire [WIDTH-1:0] wire_d62_76;
	wire [WIDTH-1:0] wire_d62_77;
	wire [WIDTH-1:0] wire_d62_78;
	wire [WIDTH-1:0] wire_d62_79;
	wire [WIDTH-1:0] wire_d62_80;
	wire [WIDTH-1:0] wire_d62_81;
	wire [WIDTH-1:0] wire_d62_82;
	wire [WIDTH-1:0] wire_d62_83;
	wire [WIDTH-1:0] wire_d62_84;
	wire [WIDTH-1:0] wire_d62_85;
	wire [WIDTH-1:0] wire_d62_86;
	wire [WIDTH-1:0] wire_d62_87;
	wire [WIDTH-1:0] wire_d62_88;
	wire [WIDTH-1:0] wire_d62_89;
	wire [WIDTH-1:0] wire_d62_90;
	wire [WIDTH-1:0] wire_d62_91;
	wire [WIDTH-1:0] wire_d62_92;
	wire [WIDTH-1:0] wire_d62_93;
	wire [WIDTH-1:0] wire_d62_94;
	wire [WIDTH-1:0] wire_d62_95;
	wire [WIDTH-1:0] wire_d62_96;
	wire [WIDTH-1:0] wire_d62_97;
	wire [WIDTH-1:0] wire_d62_98;
	wire [WIDTH-1:0] wire_d62_99;
	wire [WIDTH-1:0] wire_d62_100;
	wire [WIDTH-1:0] wire_d62_101;
	wire [WIDTH-1:0] wire_d62_102;
	wire [WIDTH-1:0] wire_d62_103;
	wire [WIDTH-1:0] wire_d62_104;
	wire [WIDTH-1:0] wire_d62_105;
	wire [WIDTH-1:0] wire_d62_106;
	wire [WIDTH-1:0] wire_d62_107;
	wire [WIDTH-1:0] wire_d62_108;
	wire [WIDTH-1:0] wire_d62_109;
	wire [WIDTH-1:0] wire_d62_110;
	wire [WIDTH-1:0] wire_d62_111;
	wire [WIDTH-1:0] wire_d62_112;
	wire [WIDTH-1:0] wire_d62_113;
	wire [WIDTH-1:0] wire_d62_114;
	wire [WIDTH-1:0] wire_d62_115;
	wire [WIDTH-1:0] wire_d62_116;
	wire [WIDTH-1:0] wire_d62_117;
	wire [WIDTH-1:0] wire_d62_118;
	wire [WIDTH-1:0] wire_d63_0;
	wire [WIDTH-1:0] wire_d63_1;
	wire [WIDTH-1:0] wire_d63_2;
	wire [WIDTH-1:0] wire_d63_3;
	wire [WIDTH-1:0] wire_d63_4;
	wire [WIDTH-1:0] wire_d63_5;
	wire [WIDTH-1:0] wire_d63_6;
	wire [WIDTH-1:0] wire_d63_7;
	wire [WIDTH-1:0] wire_d63_8;
	wire [WIDTH-1:0] wire_d63_9;
	wire [WIDTH-1:0] wire_d63_10;
	wire [WIDTH-1:0] wire_d63_11;
	wire [WIDTH-1:0] wire_d63_12;
	wire [WIDTH-1:0] wire_d63_13;
	wire [WIDTH-1:0] wire_d63_14;
	wire [WIDTH-1:0] wire_d63_15;
	wire [WIDTH-1:0] wire_d63_16;
	wire [WIDTH-1:0] wire_d63_17;
	wire [WIDTH-1:0] wire_d63_18;
	wire [WIDTH-1:0] wire_d63_19;
	wire [WIDTH-1:0] wire_d63_20;
	wire [WIDTH-1:0] wire_d63_21;
	wire [WIDTH-1:0] wire_d63_22;
	wire [WIDTH-1:0] wire_d63_23;
	wire [WIDTH-1:0] wire_d63_24;
	wire [WIDTH-1:0] wire_d63_25;
	wire [WIDTH-1:0] wire_d63_26;
	wire [WIDTH-1:0] wire_d63_27;
	wire [WIDTH-1:0] wire_d63_28;
	wire [WIDTH-1:0] wire_d63_29;
	wire [WIDTH-1:0] wire_d63_30;
	wire [WIDTH-1:0] wire_d63_31;
	wire [WIDTH-1:0] wire_d63_32;
	wire [WIDTH-1:0] wire_d63_33;
	wire [WIDTH-1:0] wire_d63_34;
	wire [WIDTH-1:0] wire_d63_35;
	wire [WIDTH-1:0] wire_d63_36;
	wire [WIDTH-1:0] wire_d63_37;
	wire [WIDTH-1:0] wire_d63_38;
	wire [WIDTH-1:0] wire_d63_39;
	wire [WIDTH-1:0] wire_d63_40;
	wire [WIDTH-1:0] wire_d63_41;
	wire [WIDTH-1:0] wire_d63_42;
	wire [WIDTH-1:0] wire_d63_43;
	wire [WIDTH-1:0] wire_d63_44;
	wire [WIDTH-1:0] wire_d63_45;
	wire [WIDTH-1:0] wire_d63_46;
	wire [WIDTH-1:0] wire_d63_47;
	wire [WIDTH-1:0] wire_d63_48;
	wire [WIDTH-1:0] wire_d63_49;
	wire [WIDTH-1:0] wire_d63_50;
	wire [WIDTH-1:0] wire_d63_51;
	wire [WIDTH-1:0] wire_d63_52;
	wire [WIDTH-1:0] wire_d63_53;
	wire [WIDTH-1:0] wire_d63_54;
	wire [WIDTH-1:0] wire_d63_55;
	wire [WIDTH-1:0] wire_d63_56;
	wire [WIDTH-1:0] wire_d63_57;
	wire [WIDTH-1:0] wire_d63_58;
	wire [WIDTH-1:0] wire_d63_59;
	wire [WIDTH-1:0] wire_d63_60;
	wire [WIDTH-1:0] wire_d63_61;
	wire [WIDTH-1:0] wire_d63_62;
	wire [WIDTH-1:0] wire_d63_63;
	wire [WIDTH-1:0] wire_d63_64;
	wire [WIDTH-1:0] wire_d63_65;
	wire [WIDTH-1:0] wire_d63_66;
	wire [WIDTH-1:0] wire_d63_67;
	wire [WIDTH-1:0] wire_d63_68;
	wire [WIDTH-1:0] wire_d63_69;
	wire [WIDTH-1:0] wire_d63_70;
	wire [WIDTH-1:0] wire_d63_71;
	wire [WIDTH-1:0] wire_d63_72;
	wire [WIDTH-1:0] wire_d63_73;
	wire [WIDTH-1:0] wire_d63_74;
	wire [WIDTH-1:0] wire_d63_75;
	wire [WIDTH-1:0] wire_d63_76;
	wire [WIDTH-1:0] wire_d63_77;
	wire [WIDTH-1:0] wire_d63_78;
	wire [WIDTH-1:0] wire_d63_79;
	wire [WIDTH-1:0] wire_d63_80;
	wire [WIDTH-1:0] wire_d63_81;
	wire [WIDTH-1:0] wire_d63_82;
	wire [WIDTH-1:0] wire_d63_83;
	wire [WIDTH-1:0] wire_d63_84;
	wire [WIDTH-1:0] wire_d63_85;
	wire [WIDTH-1:0] wire_d63_86;
	wire [WIDTH-1:0] wire_d63_87;
	wire [WIDTH-1:0] wire_d63_88;
	wire [WIDTH-1:0] wire_d63_89;
	wire [WIDTH-1:0] wire_d63_90;
	wire [WIDTH-1:0] wire_d63_91;
	wire [WIDTH-1:0] wire_d63_92;
	wire [WIDTH-1:0] wire_d63_93;
	wire [WIDTH-1:0] wire_d63_94;
	wire [WIDTH-1:0] wire_d63_95;
	wire [WIDTH-1:0] wire_d63_96;
	wire [WIDTH-1:0] wire_d63_97;
	wire [WIDTH-1:0] wire_d63_98;
	wire [WIDTH-1:0] wire_d63_99;
	wire [WIDTH-1:0] wire_d63_100;
	wire [WIDTH-1:0] wire_d63_101;
	wire [WIDTH-1:0] wire_d63_102;
	wire [WIDTH-1:0] wire_d63_103;
	wire [WIDTH-1:0] wire_d63_104;
	wire [WIDTH-1:0] wire_d63_105;
	wire [WIDTH-1:0] wire_d63_106;
	wire [WIDTH-1:0] wire_d63_107;
	wire [WIDTH-1:0] wire_d63_108;
	wire [WIDTH-1:0] wire_d63_109;
	wire [WIDTH-1:0] wire_d63_110;
	wire [WIDTH-1:0] wire_d63_111;
	wire [WIDTH-1:0] wire_d63_112;
	wire [WIDTH-1:0] wire_d63_113;
	wire [WIDTH-1:0] wire_d63_114;
	wire [WIDTH-1:0] wire_d63_115;
	wire [WIDTH-1:0] wire_d63_116;
	wire [WIDTH-1:0] wire_d63_117;
	wire [WIDTH-1:0] wire_d63_118;
	wire [WIDTH-1:0] wire_d64_0;
	wire [WIDTH-1:0] wire_d64_1;
	wire [WIDTH-1:0] wire_d64_2;
	wire [WIDTH-1:0] wire_d64_3;
	wire [WIDTH-1:0] wire_d64_4;
	wire [WIDTH-1:0] wire_d64_5;
	wire [WIDTH-1:0] wire_d64_6;
	wire [WIDTH-1:0] wire_d64_7;
	wire [WIDTH-1:0] wire_d64_8;
	wire [WIDTH-1:0] wire_d64_9;
	wire [WIDTH-1:0] wire_d64_10;
	wire [WIDTH-1:0] wire_d64_11;
	wire [WIDTH-1:0] wire_d64_12;
	wire [WIDTH-1:0] wire_d64_13;
	wire [WIDTH-1:0] wire_d64_14;
	wire [WIDTH-1:0] wire_d64_15;
	wire [WIDTH-1:0] wire_d64_16;
	wire [WIDTH-1:0] wire_d64_17;
	wire [WIDTH-1:0] wire_d64_18;
	wire [WIDTH-1:0] wire_d64_19;
	wire [WIDTH-1:0] wire_d64_20;
	wire [WIDTH-1:0] wire_d64_21;
	wire [WIDTH-1:0] wire_d64_22;
	wire [WIDTH-1:0] wire_d64_23;
	wire [WIDTH-1:0] wire_d64_24;
	wire [WIDTH-1:0] wire_d64_25;
	wire [WIDTH-1:0] wire_d64_26;
	wire [WIDTH-1:0] wire_d64_27;
	wire [WIDTH-1:0] wire_d64_28;
	wire [WIDTH-1:0] wire_d64_29;
	wire [WIDTH-1:0] wire_d64_30;
	wire [WIDTH-1:0] wire_d64_31;
	wire [WIDTH-1:0] wire_d64_32;
	wire [WIDTH-1:0] wire_d64_33;
	wire [WIDTH-1:0] wire_d64_34;
	wire [WIDTH-1:0] wire_d64_35;
	wire [WIDTH-1:0] wire_d64_36;
	wire [WIDTH-1:0] wire_d64_37;
	wire [WIDTH-1:0] wire_d64_38;
	wire [WIDTH-1:0] wire_d64_39;
	wire [WIDTH-1:0] wire_d64_40;
	wire [WIDTH-1:0] wire_d64_41;
	wire [WIDTH-1:0] wire_d64_42;
	wire [WIDTH-1:0] wire_d64_43;
	wire [WIDTH-1:0] wire_d64_44;
	wire [WIDTH-1:0] wire_d64_45;
	wire [WIDTH-1:0] wire_d64_46;
	wire [WIDTH-1:0] wire_d64_47;
	wire [WIDTH-1:0] wire_d64_48;
	wire [WIDTH-1:0] wire_d64_49;
	wire [WIDTH-1:0] wire_d64_50;
	wire [WIDTH-1:0] wire_d64_51;
	wire [WIDTH-1:0] wire_d64_52;
	wire [WIDTH-1:0] wire_d64_53;
	wire [WIDTH-1:0] wire_d64_54;
	wire [WIDTH-1:0] wire_d64_55;
	wire [WIDTH-1:0] wire_d64_56;
	wire [WIDTH-1:0] wire_d64_57;
	wire [WIDTH-1:0] wire_d64_58;
	wire [WIDTH-1:0] wire_d64_59;
	wire [WIDTH-1:0] wire_d64_60;
	wire [WIDTH-1:0] wire_d64_61;
	wire [WIDTH-1:0] wire_d64_62;
	wire [WIDTH-1:0] wire_d64_63;
	wire [WIDTH-1:0] wire_d64_64;
	wire [WIDTH-1:0] wire_d64_65;
	wire [WIDTH-1:0] wire_d64_66;
	wire [WIDTH-1:0] wire_d64_67;
	wire [WIDTH-1:0] wire_d64_68;
	wire [WIDTH-1:0] wire_d64_69;
	wire [WIDTH-1:0] wire_d64_70;
	wire [WIDTH-1:0] wire_d64_71;
	wire [WIDTH-1:0] wire_d64_72;
	wire [WIDTH-1:0] wire_d64_73;
	wire [WIDTH-1:0] wire_d64_74;
	wire [WIDTH-1:0] wire_d64_75;
	wire [WIDTH-1:0] wire_d64_76;
	wire [WIDTH-1:0] wire_d64_77;
	wire [WIDTH-1:0] wire_d64_78;
	wire [WIDTH-1:0] wire_d64_79;
	wire [WIDTH-1:0] wire_d64_80;
	wire [WIDTH-1:0] wire_d64_81;
	wire [WIDTH-1:0] wire_d64_82;
	wire [WIDTH-1:0] wire_d64_83;
	wire [WIDTH-1:0] wire_d64_84;
	wire [WIDTH-1:0] wire_d64_85;
	wire [WIDTH-1:0] wire_d64_86;
	wire [WIDTH-1:0] wire_d64_87;
	wire [WIDTH-1:0] wire_d64_88;
	wire [WIDTH-1:0] wire_d64_89;
	wire [WIDTH-1:0] wire_d64_90;
	wire [WIDTH-1:0] wire_d64_91;
	wire [WIDTH-1:0] wire_d64_92;
	wire [WIDTH-1:0] wire_d64_93;
	wire [WIDTH-1:0] wire_d64_94;
	wire [WIDTH-1:0] wire_d64_95;
	wire [WIDTH-1:0] wire_d64_96;
	wire [WIDTH-1:0] wire_d64_97;
	wire [WIDTH-1:0] wire_d64_98;
	wire [WIDTH-1:0] wire_d64_99;
	wire [WIDTH-1:0] wire_d64_100;
	wire [WIDTH-1:0] wire_d64_101;
	wire [WIDTH-1:0] wire_d64_102;
	wire [WIDTH-1:0] wire_d64_103;
	wire [WIDTH-1:0] wire_d64_104;
	wire [WIDTH-1:0] wire_d64_105;
	wire [WIDTH-1:0] wire_d64_106;
	wire [WIDTH-1:0] wire_d64_107;
	wire [WIDTH-1:0] wire_d64_108;
	wire [WIDTH-1:0] wire_d64_109;
	wire [WIDTH-1:0] wire_d64_110;
	wire [WIDTH-1:0] wire_d64_111;
	wire [WIDTH-1:0] wire_d64_112;
	wire [WIDTH-1:0] wire_d64_113;
	wire [WIDTH-1:0] wire_d64_114;
	wire [WIDTH-1:0] wire_d64_115;
	wire [WIDTH-1:0] wire_d64_116;
	wire [WIDTH-1:0] wire_d64_117;
	wire [WIDTH-1:0] wire_d64_118;
	wire [WIDTH-1:0] wire_d65_0;
	wire [WIDTH-1:0] wire_d65_1;
	wire [WIDTH-1:0] wire_d65_2;
	wire [WIDTH-1:0] wire_d65_3;
	wire [WIDTH-1:0] wire_d65_4;
	wire [WIDTH-1:0] wire_d65_5;
	wire [WIDTH-1:0] wire_d65_6;
	wire [WIDTH-1:0] wire_d65_7;
	wire [WIDTH-1:0] wire_d65_8;
	wire [WIDTH-1:0] wire_d65_9;
	wire [WIDTH-1:0] wire_d65_10;
	wire [WIDTH-1:0] wire_d65_11;
	wire [WIDTH-1:0] wire_d65_12;
	wire [WIDTH-1:0] wire_d65_13;
	wire [WIDTH-1:0] wire_d65_14;
	wire [WIDTH-1:0] wire_d65_15;
	wire [WIDTH-1:0] wire_d65_16;
	wire [WIDTH-1:0] wire_d65_17;
	wire [WIDTH-1:0] wire_d65_18;
	wire [WIDTH-1:0] wire_d65_19;
	wire [WIDTH-1:0] wire_d65_20;
	wire [WIDTH-1:0] wire_d65_21;
	wire [WIDTH-1:0] wire_d65_22;
	wire [WIDTH-1:0] wire_d65_23;
	wire [WIDTH-1:0] wire_d65_24;
	wire [WIDTH-1:0] wire_d65_25;
	wire [WIDTH-1:0] wire_d65_26;
	wire [WIDTH-1:0] wire_d65_27;
	wire [WIDTH-1:0] wire_d65_28;
	wire [WIDTH-1:0] wire_d65_29;
	wire [WIDTH-1:0] wire_d65_30;
	wire [WIDTH-1:0] wire_d65_31;
	wire [WIDTH-1:0] wire_d65_32;
	wire [WIDTH-1:0] wire_d65_33;
	wire [WIDTH-1:0] wire_d65_34;
	wire [WIDTH-1:0] wire_d65_35;
	wire [WIDTH-1:0] wire_d65_36;
	wire [WIDTH-1:0] wire_d65_37;
	wire [WIDTH-1:0] wire_d65_38;
	wire [WIDTH-1:0] wire_d65_39;
	wire [WIDTH-1:0] wire_d65_40;
	wire [WIDTH-1:0] wire_d65_41;
	wire [WIDTH-1:0] wire_d65_42;
	wire [WIDTH-1:0] wire_d65_43;
	wire [WIDTH-1:0] wire_d65_44;
	wire [WIDTH-1:0] wire_d65_45;
	wire [WIDTH-1:0] wire_d65_46;
	wire [WIDTH-1:0] wire_d65_47;
	wire [WIDTH-1:0] wire_d65_48;
	wire [WIDTH-1:0] wire_d65_49;
	wire [WIDTH-1:0] wire_d65_50;
	wire [WIDTH-1:0] wire_d65_51;
	wire [WIDTH-1:0] wire_d65_52;
	wire [WIDTH-1:0] wire_d65_53;
	wire [WIDTH-1:0] wire_d65_54;
	wire [WIDTH-1:0] wire_d65_55;
	wire [WIDTH-1:0] wire_d65_56;
	wire [WIDTH-1:0] wire_d65_57;
	wire [WIDTH-1:0] wire_d65_58;
	wire [WIDTH-1:0] wire_d65_59;
	wire [WIDTH-1:0] wire_d65_60;
	wire [WIDTH-1:0] wire_d65_61;
	wire [WIDTH-1:0] wire_d65_62;
	wire [WIDTH-1:0] wire_d65_63;
	wire [WIDTH-1:0] wire_d65_64;
	wire [WIDTH-1:0] wire_d65_65;
	wire [WIDTH-1:0] wire_d65_66;
	wire [WIDTH-1:0] wire_d65_67;
	wire [WIDTH-1:0] wire_d65_68;
	wire [WIDTH-1:0] wire_d65_69;
	wire [WIDTH-1:0] wire_d65_70;
	wire [WIDTH-1:0] wire_d65_71;
	wire [WIDTH-1:0] wire_d65_72;
	wire [WIDTH-1:0] wire_d65_73;
	wire [WIDTH-1:0] wire_d65_74;
	wire [WIDTH-1:0] wire_d65_75;
	wire [WIDTH-1:0] wire_d65_76;
	wire [WIDTH-1:0] wire_d65_77;
	wire [WIDTH-1:0] wire_d65_78;
	wire [WIDTH-1:0] wire_d65_79;
	wire [WIDTH-1:0] wire_d65_80;
	wire [WIDTH-1:0] wire_d65_81;
	wire [WIDTH-1:0] wire_d65_82;
	wire [WIDTH-1:0] wire_d65_83;
	wire [WIDTH-1:0] wire_d65_84;
	wire [WIDTH-1:0] wire_d65_85;
	wire [WIDTH-1:0] wire_d65_86;
	wire [WIDTH-1:0] wire_d65_87;
	wire [WIDTH-1:0] wire_d65_88;
	wire [WIDTH-1:0] wire_d65_89;
	wire [WIDTH-1:0] wire_d65_90;
	wire [WIDTH-1:0] wire_d65_91;
	wire [WIDTH-1:0] wire_d65_92;
	wire [WIDTH-1:0] wire_d65_93;
	wire [WIDTH-1:0] wire_d65_94;
	wire [WIDTH-1:0] wire_d65_95;
	wire [WIDTH-1:0] wire_d65_96;
	wire [WIDTH-1:0] wire_d65_97;
	wire [WIDTH-1:0] wire_d65_98;
	wire [WIDTH-1:0] wire_d65_99;
	wire [WIDTH-1:0] wire_d65_100;
	wire [WIDTH-1:0] wire_d65_101;
	wire [WIDTH-1:0] wire_d65_102;
	wire [WIDTH-1:0] wire_d65_103;
	wire [WIDTH-1:0] wire_d65_104;
	wire [WIDTH-1:0] wire_d65_105;
	wire [WIDTH-1:0] wire_d65_106;
	wire [WIDTH-1:0] wire_d65_107;
	wire [WIDTH-1:0] wire_d65_108;
	wire [WIDTH-1:0] wire_d65_109;
	wire [WIDTH-1:0] wire_d65_110;
	wire [WIDTH-1:0] wire_d65_111;
	wire [WIDTH-1:0] wire_d65_112;
	wire [WIDTH-1:0] wire_d65_113;
	wire [WIDTH-1:0] wire_d65_114;
	wire [WIDTH-1:0] wire_d65_115;
	wire [WIDTH-1:0] wire_d65_116;
	wire [WIDTH-1:0] wire_d65_117;
	wire [WIDTH-1:0] wire_d65_118;
	wire [WIDTH-1:0] wire_d66_0;
	wire [WIDTH-1:0] wire_d66_1;
	wire [WIDTH-1:0] wire_d66_2;
	wire [WIDTH-1:0] wire_d66_3;
	wire [WIDTH-1:0] wire_d66_4;
	wire [WIDTH-1:0] wire_d66_5;
	wire [WIDTH-1:0] wire_d66_6;
	wire [WIDTH-1:0] wire_d66_7;
	wire [WIDTH-1:0] wire_d66_8;
	wire [WIDTH-1:0] wire_d66_9;
	wire [WIDTH-1:0] wire_d66_10;
	wire [WIDTH-1:0] wire_d66_11;
	wire [WIDTH-1:0] wire_d66_12;
	wire [WIDTH-1:0] wire_d66_13;
	wire [WIDTH-1:0] wire_d66_14;
	wire [WIDTH-1:0] wire_d66_15;
	wire [WIDTH-1:0] wire_d66_16;
	wire [WIDTH-1:0] wire_d66_17;
	wire [WIDTH-1:0] wire_d66_18;
	wire [WIDTH-1:0] wire_d66_19;
	wire [WIDTH-1:0] wire_d66_20;
	wire [WIDTH-1:0] wire_d66_21;
	wire [WIDTH-1:0] wire_d66_22;
	wire [WIDTH-1:0] wire_d66_23;
	wire [WIDTH-1:0] wire_d66_24;
	wire [WIDTH-1:0] wire_d66_25;
	wire [WIDTH-1:0] wire_d66_26;
	wire [WIDTH-1:0] wire_d66_27;
	wire [WIDTH-1:0] wire_d66_28;
	wire [WIDTH-1:0] wire_d66_29;
	wire [WIDTH-1:0] wire_d66_30;
	wire [WIDTH-1:0] wire_d66_31;
	wire [WIDTH-1:0] wire_d66_32;
	wire [WIDTH-1:0] wire_d66_33;
	wire [WIDTH-1:0] wire_d66_34;
	wire [WIDTH-1:0] wire_d66_35;
	wire [WIDTH-1:0] wire_d66_36;
	wire [WIDTH-1:0] wire_d66_37;
	wire [WIDTH-1:0] wire_d66_38;
	wire [WIDTH-1:0] wire_d66_39;
	wire [WIDTH-1:0] wire_d66_40;
	wire [WIDTH-1:0] wire_d66_41;
	wire [WIDTH-1:0] wire_d66_42;
	wire [WIDTH-1:0] wire_d66_43;
	wire [WIDTH-1:0] wire_d66_44;
	wire [WIDTH-1:0] wire_d66_45;
	wire [WIDTH-1:0] wire_d66_46;
	wire [WIDTH-1:0] wire_d66_47;
	wire [WIDTH-1:0] wire_d66_48;
	wire [WIDTH-1:0] wire_d66_49;
	wire [WIDTH-1:0] wire_d66_50;
	wire [WIDTH-1:0] wire_d66_51;
	wire [WIDTH-1:0] wire_d66_52;
	wire [WIDTH-1:0] wire_d66_53;
	wire [WIDTH-1:0] wire_d66_54;
	wire [WIDTH-1:0] wire_d66_55;
	wire [WIDTH-1:0] wire_d66_56;
	wire [WIDTH-1:0] wire_d66_57;
	wire [WIDTH-1:0] wire_d66_58;
	wire [WIDTH-1:0] wire_d66_59;
	wire [WIDTH-1:0] wire_d66_60;
	wire [WIDTH-1:0] wire_d66_61;
	wire [WIDTH-1:0] wire_d66_62;
	wire [WIDTH-1:0] wire_d66_63;
	wire [WIDTH-1:0] wire_d66_64;
	wire [WIDTH-1:0] wire_d66_65;
	wire [WIDTH-1:0] wire_d66_66;
	wire [WIDTH-1:0] wire_d66_67;
	wire [WIDTH-1:0] wire_d66_68;
	wire [WIDTH-1:0] wire_d66_69;
	wire [WIDTH-1:0] wire_d66_70;
	wire [WIDTH-1:0] wire_d66_71;
	wire [WIDTH-1:0] wire_d66_72;
	wire [WIDTH-1:0] wire_d66_73;
	wire [WIDTH-1:0] wire_d66_74;
	wire [WIDTH-1:0] wire_d66_75;
	wire [WIDTH-1:0] wire_d66_76;
	wire [WIDTH-1:0] wire_d66_77;
	wire [WIDTH-1:0] wire_d66_78;
	wire [WIDTH-1:0] wire_d66_79;
	wire [WIDTH-1:0] wire_d66_80;
	wire [WIDTH-1:0] wire_d66_81;
	wire [WIDTH-1:0] wire_d66_82;
	wire [WIDTH-1:0] wire_d66_83;
	wire [WIDTH-1:0] wire_d66_84;
	wire [WIDTH-1:0] wire_d66_85;
	wire [WIDTH-1:0] wire_d66_86;
	wire [WIDTH-1:0] wire_d66_87;
	wire [WIDTH-1:0] wire_d66_88;
	wire [WIDTH-1:0] wire_d66_89;
	wire [WIDTH-1:0] wire_d66_90;
	wire [WIDTH-1:0] wire_d66_91;
	wire [WIDTH-1:0] wire_d66_92;
	wire [WIDTH-1:0] wire_d66_93;
	wire [WIDTH-1:0] wire_d66_94;
	wire [WIDTH-1:0] wire_d66_95;
	wire [WIDTH-1:0] wire_d66_96;
	wire [WIDTH-1:0] wire_d66_97;
	wire [WIDTH-1:0] wire_d66_98;
	wire [WIDTH-1:0] wire_d66_99;
	wire [WIDTH-1:0] wire_d66_100;
	wire [WIDTH-1:0] wire_d66_101;
	wire [WIDTH-1:0] wire_d66_102;
	wire [WIDTH-1:0] wire_d66_103;
	wire [WIDTH-1:0] wire_d66_104;
	wire [WIDTH-1:0] wire_d66_105;
	wire [WIDTH-1:0] wire_d66_106;
	wire [WIDTH-1:0] wire_d66_107;
	wire [WIDTH-1:0] wire_d66_108;
	wire [WIDTH-1:0] wire_d66_109;
	wire [WIDTH-1:0] wire_d66_110;
	wire [WIDTH-1:0] wire_d66_111;
	wire [WIDTH-1:0] wire_d66_112;
	wire [WIDTH-1:0] wire_d66_113;
	wire [WIDTH-1:0] wire_d66_114;
	wire [WIDTH-1:0] wire_d66_115;
	wire [WIDTH-1:0] wire_d66_116;
	wire [WIDTH-1:0] wire_d66_117;
	wire [WIDTH-1:0] wire_d66_118;
	wire [WIDTH-1:0] wire_d67_0;
	wire [WIDTH-1:0] wire_d67_1;
	wire [WIDTH-1:0] wire_d67_2;
	wire [WIDTH-1:0] wire_d67_3;
	wire [WIDTH-1:0] wire_d67_4;
	wire [WIDTH-1:0] wire_d67_5;
	wire [WIDTH-1:0] wire_d67_6;
	wire [WIDTH-1:0] wire_d67_7;
	wire [WIDTH-1:0] wire_d67_8;
	wire [WIDTH-1:0] wire_d67_9;
	wire [WIDTH-1:0] wire_d67_10;
	wire [WIDTH-1:0] wire_d67_11;
	wire [WIDTH-1:0] wire_d67_12;
	wire [WIDTH-1:0] wire_d67_13;
	wire [WIDTH-1:0] wire_d67_14;
	wire [WIDTH-1:0] wire_d67_15;
	wire [WIDTH-1:0] wire_d67_16;
	wire [WIDTH-1:0] wire_d67_17;
	wire [WIDTH-1:0] wire_d67_18;
	wire [WIDTH-1:0] wire_d67_19;
	wire [WIDTH-1:0] wire_d67_20;
	wire [WIDTH-1:0] wire_d67_21;
	wire [WIDTH-1:0] wire_d67_22;
	wire [WIDTH-1:0] wire_d67_23;
	wire [WIDTH-1:0] wire_d67_24;
	wire [WIDTH-1:0] wire_d67_25;
	wire [WIDTH-1:0] wire_d67_26;
	wire [WIDTH-1:0] wire_d67_27;
	wire [WIDTH-1:0] wire_d67_28;
	wire [WIDTH-1:0] wire_d67_29;
	wire [WIDTH-1:0] wire_d67_30;
	wire [WIDTH-1:0] wire_d67_31;
	wire [WIDTH-1:0] wire_d67_32;
	wire [WIDTH-1:0] wire_d67_33;
	wire [WIDTH-1:0] wire_d67_34;
	wire [WIDTH-1:0] wire_d67_35;
	wire [WIDTH-1:0] wire_d67_36;
	wire [WIDTH-1:0] wire_d67_37;
	wire [WIDTH-1:0] wire_d67_38;
	wire [WIDTH-1:0] wire_d67_39;
	wire [WIDTH-1:0] wire_d67_40;
	wire [WIDTH-1:0] wire_d67_41;
	wire [WIDTH-1:0] wire_d67_42;
	wire [WIDTH-1:0] wire_d67_43;
	wire [WIDTH-1:0] wire_d67_44;
	wire [WIDTH-1:0] wire_d67_45;
	wire [WIDTH-1:0] wire_d67_46;
	wire [WIDTH-1:0] wire_d67_47;
	wire [WIDTH-1:0] wire_d67_48;
	wire [WIDTH-1:0] wire_d67_49;
	wire [WIDTH-1:0] wire_d67_50;
	wire [WIDTH-1:0] wire_d67_51;
	wire [WIDTH-1:0] wire_d67_52;
	wire [WIDTH-1:0] wire_d67_53;
	wire [WIDTH-1:0] wire_d67_54;
	wire [WIDTH-1:0] wire_d67_55;
	wire [WIDTH-1:0] wire_d67_56;
	wire [WIDTH-1:0] wire_d67_57;
	wire [WIDTH-1:0] wire_d67_58;
	wire [WIDTH-1:0] wire_d67_59;
	wire [WIDTH-1:0] wire_d67_60;
	wire [WIDTH-1:0] wire_d67_61;
	wire [WIDTH-1:0] wire_d67_62;
	wire [WIDTH-1:0] wire_d67_63;
	wire [WIDTH-1:0] wire_d67_64;
	wire [WIDTH-1:0] wire_d67_65;
	wire [WIDTH-1:0] wire_d67_66;
	wire [WIDTH-1:0] wire_d67_67;
	wire [WIDTH-1:0] wire_d67_68;
	wire [WIDTH-1:0] wire_d67_69;
	wire [WIDTH-1:0] wire_d67_70;
	wire [WIDTH-1:0] wire_d67_71;
	wire [WIDTH-1:0] wire_d67_72;
	wire [WIDTH-1:0] wire_d67_73;
	wire [WIDTH-1:0] wire_d67_74;
	wire [WIDTH-1:0] wire_d67_75;
	wire [WIDTH-1:0] wire_d67_76;
	wire [WIDTH-1:0] wire_d67_77;
	wire [WIDTH-1:0] wire_d67_78;
	wire [WIDTH-1:0] wire_d67_79;
	wire [WIDTH-1:0] wire_d67_80;
	wire [WIDTH-1:0] wire_d67_81;
	wire [WIDTH-1:0] wire_d67_82;
	wire [WIDTH-1:0] wire_d67_83;
	wire [WIDTH-1:0] wire_d67_84;
	wire [WIDTH-1:0] wire_d67_85;
	wire [WIDTH-1:0] wire_d67_86;
	wire [WIDTH-1:0] wire_d67_87;
	wire [WIDTH-1:0] wire_d67_88;
	wire [WIDTH-1:0] wire_d67_89;
	wire [WIDTH-1:0] wire_d67_90;
	wire [WIDTH-1:0] wire_d67_91;
	wire [WIDTH-1:0] wire_d67_92;
	wire [WIDTH-1:0] wire_d67_93;
	wire [WIDTH-1:0] wire_d67_94;
	wire [WIDTH-1:0] wire_d67_95;
	wire [WIDTH-1:0] wire_d67_96;
	wire [WIDTH-1:0] wire_d67_97;
	wire [WIDTH-1:0] wire_d67_98;
	wire [WIDTH-1:0] wire_d67_99;
	wire [WIDTH-1:0] wire_d67_100;
	wire [WIDTH-1:0] wire_d67_101;
	wire [WIDTH-1:0] wire_d67_102;
	wire [WIDTH-1:0] wire_d67_103;
	wire [WIDTH-1:0] wire_d67_104;
	wire [WIDTH-1:0] wire_d67_105;
	wire [WIDTH-1:0] wire_d67_106;
	wire [WIDTH-1:0] wire_d67_107;
	wire [WIDTH-1:0] wire_d67_108;
	wire [WIDTH-1:0] wire_d67_109;
	wire [WIDTH-1:0] wire_d67_110;
	wire [WIDTH-1:0] wire_d67_111;
	wire [WIDTH-1:0] wire_d67_112;
	wire [WIDTH-1:0] wire_d67_113;
	wire [WIDTH-1:0] wire_d67_114;
	wire [WIDTH-1:0] wire_d67_115;
	wire [WIDTH-1:0] wire_d67_116;
	wire [WIDTH-1:0] wire_d67_117;
	wire [WIDTH-1:0] wire_d67_118;
	wire [WIDTH-1:0] wire_d68_0;
	wire [WIDTH-1:0] wire_d68_1;
	wire [WIDTH-1:0] wire_d68_2;
	wire [WIDTH-1:0] wire_d68_3;
	wire [WIDTH-1:0] wire_d68_4;
	wire [WIDTH-1:0] wire_d68_5;
	wire [WIDTH-1:0] wire_d68_6;
	wire [WIDTH-1:0] wire_d68_7;
	wire [WIDTH-1:0] wire_d68_8;
	wire [WIDTH-1:0] wire_d68_9;
	wire [WIDTH-1:0] wire_d68_10;
	wire [WIDTH-1:0] wire_d68_11;
	wire [WIDTH-1:0] wire_d68_12;
	wire [WIDTH-1:0] wire_d68_13;
	wire [WIDTH-1:0] wire_d68_14;
	wire [WIDTH-1:0] wire_d68_15;
	wire [WIDTH-1:0] wire_d68_16;
	wire [WIDTH-1:0] wire_d68_17;
	wire [WIDTH-1:0] wire_d68_18;
	wire [WIDTH-1:0] wire_d68_19;
	wire [WIDTH-1:0] wire_d68_20;
	wire [WIDTH-1:0] wire_d68_21;
	wire [WIDTH-1:0] wire_d68_22;
	wire [WIDTH-1:0] wire_d68_23;
	wire [WIDTH-1:0] wire_d68_24;
	wire [WIDTH-1:0] wire_d68_25;
	wire [WIDTH-1:0] wire_d68_26;
	wire [WIDTH-1:0] wire_d68_27;
	wire [WIDTH-1:0] wire_d68_28;
	wire [WIDTH-1:0] wire_d68_29;
	wire [WIDTH-1:0] wire_d68_30;
	wire [WIDTH-1:0] wire_d68_31;
	wire [WIDTH-1:0] wire_d68_32;
	wire [WIDTH-1:0] wire_d68_33;
	wire [WIDTH-1:0] wire_d68_34;
	wire [WIDTH-1:0] wire_d68_35;
	wire [WIDTH-1:0] wire_d68_36;
	wire [WIDTH-1:0] wire_d68_37;
	wire [WIDTH-1:0] wire_d68_38;
	wire [WIDTH-1:0] wire_d68_39;
	wire [WIDTH-1:0] wire_d68_40;
	wire [WIDTH-1:0] wire_d68_41;
	wire [WIDTH-1:0] wire_d68_42;
	wire [WIDTH-1:0] wire_d68_43;
	wire [WIDTH-1:0] wire_d68_44;
	wire [WIDTH-1:0] wire_d68_45;
	wire [WIDTH-1:0] wire_d68_46;
	wire [WIDTH-1:0] wire_d68_47;
	wire [WIDTH-1:0] wire_d68_48;
	wire [WIDTH-1:0] wire_d68_49;
	wire [WIDTH-1:0] wire_d68_50;
	wire [WIDTH-1:0] wire_d68_51;
	wire [WIDTH-1:0] wire_d68_52;
	wire [WIDTH-1:0] wire_d68_53;
	wire [WIDTH-1:0] wire_d68_54;
	wire [WIDTH-1:0] wire_d68_55;
	wire [WIDTH-1:0] wire_d68_56;
	wire [WIDTH-1:0] wire_d68_57;
	wire [WIDTH-1:0] wire_d68_58;
	wire [WIDTH-1:0] wire_d68_59;
	wire [WIDTH-1:0] wire_d68_60;
	wire [WIDTH-1:0] wire_d68_61;
	wire [WIDTH-1:0] wire_d68_62;
	wire [WIDTH-1:0] wire_d68_63;
	wire [WIDTH-1:0] wire_d68_64;
	wire [WIDTH-1:0] wire_d68_65;
	wire [WIDTH-1:0] wire_d68_66;
	wire [WIDTH-1:0] wire_d68_67;
	wire [WIDTH-1:0] wire_d68_68;
	wire [WIDTH-1:0] wire_d68_69;
	wire [WIDTH-1:0] wire_d68_70;
	wire [WIDTH-1:0] wire_d68_71;
	wire [WIDTH-1:0] wire_d68_72;
	wire [WIDTH-1:0] wire_d68_73;
	wire [WIDTH-1:0] wire_d68_74;
	wire [WIDTH-1:0] wire_d68_75;
	wire [WIDTH-1:0] wire_d68_76;
	wire [WIDTH-1:0] wire_d68_77;
	wire [WIDTH-1:0] wire_d68_78;
	wire [WIDTH-1:0] wire_d68_79;
	wire [WIDTH-1:0] wire_d68_80;
	wire [WIDTH-1:0] wire_d68_81;
	wire [WIDTH-1:0] wire_d68_82;
	wire [WIDTH-1:0] wire_d68_83;
	wire [WIDTH-1:0] wire_d68_84;
	wire [WIDTH-1:0] wire_d68_85;
	wire [WIDTH-1:0] wire_d68_86;
	wire [WIDTH-1:0] wire_d68_87;
	wire [WIDTH-1:0] wire_d68_88;
	wire [WIDTH-1:0] wire_d68_89;
	wire [WIDTH-1:0] wire_d68_90;
	wire [WIDTH-1:0] wire_d68_91;
	wire [WIDTH-1:0] wire_d68_92;
	wire [WIDTH-1:0] wire_d68_93;
	wire [WIDTH-1:0] wire_d68_94;
	wire [WIDTH-1:0] wire_d68_95;
	wire [WIDTH-1:0] wire_d68_96;
	wire [WIDTH-1:0] wire_d68_97;
	wire [WIDTH-1:0] wire_d68_98;
	wire [WIDTH-1:0] wire_d68_99;
	wire [WIDTH-1:0] wire_d68_100;
	wire [WIDTH-1:0] wire_d68_101;
	wire [WIDTH-1:0] wire_d68_102;
	wire [WIDTH-1:0] wire_d68_103;
	wire [WIDTH-1:0] wire_d68_104;
	wire [WIDTH-1:0] wire_d68_105;
	wire [WIDTH-1:0] wire_d68_106;
	wire [WIDTH-1:0] wire_d68_107;
	wire [WIDTH-1:0] wire_d68_108;
	wire [WIDTH-1:0] wire_d68_109;
	wire [WIDTH-1:0] wire_d68_110;
	wire [WIDTH-1:0] wire_d68_111;
	wire [WIDTH-1:0] wire_d68_112;
	wire [WIDTH-1:0] wire_d68_113;
	wire [WIDTH-1:0] wire_d68_114;
	wire [WIDTH-1:0] wire_d68_115;
	wire [WIDTH-1:0] wire_d68_116;
	wire [WIDTH-1:0] wire_d68_117;
	wire [WIDTH-1:0] wire_d68_118;
	wire [WIDTH-1:0] wire_d69_0;
	wire [WIDTH-1:0] wire_d69_1;
	wire [WIDTH-1:0] wire_d69_2;
	wire [WIDTH-1:0] wire_d69_3;
	wire [WIDTH-1:0] wire_d69_4;
	wire [WIDTH-1:0] wire_d69_5;
	wire [WIDTH-1:0] wire_d69_6;
	wire [WIDTH-1:0] wire_d69_7;
	wire [WIDTH-1:0] wire_d69_8;
	wire [WIDTH-1:0] wire_d69_9;
	wire [WIDTH-1:0] wire_d69_10;
	wire [WIDTH-1:0] wire_d69_11;
	wire [WIDTH-1:0] wire_d69_12;
	wire [WIDTH-1:0] wire_d69_13;
	wire [WIDTH-1:0] wire_d69_14;
	wire [WIDTH-1:0] wire_d69_15;
	wire [WIDTH-1:0] wire_d69_16;
	wire [WIDTH-1:0] wire_d69_17;
	wire [WIDTH-1:0] wire_d69_18;
	wire [WIDTH-1:0] wire_d69_19;
	wire [WIDTH-1:0] wire_d69_20;
	wire [WIDTH-1:0] wire_d69_21;
	wire [WIDTH-1:0] wire_d69_22;
	wire [WIDTH-1:0] wire_d69_23;
	wire [WIDTH-1:0] wire_d69_24;
	wire [WIDTH-1:0] wire_d69_25;
	wire [WIDTH-1:0] wire_d69_26;
	wire [WIDTH-1:0] wire_d69_27;
	wire [WIDTH-1:0] wire_d69_28;
	wire [WIDTH-1:0] wire_d69_29;
	wire [WIDTH-1:0] wire_d69_30;
	wire [WIDTH-1:0] wire_d69_31;
	wire [WIDTH-1:0] wire_d69_32;
	wire [WIDTH-1:0] wire_d69_33;
	wire [WIDTH-1:0] wire_d69_34;
	wire [WIDTH-1:0] wire_d69_35;
	wire [WIDTH-1:0] wire_d69_36;
	wire [WIDTH-1:0] wire_d69_37;
	wire [WIDTH-1:0] wire_d69_38;
	wire [WIDTH-1:0] wire_d69_39;
	wire [WIDTH-1:0] wire_d69_40;
	wire [WIDTH-1:0] wire_d69_41;
	wire [WIDTH-1:0] wire_d69_42;
	wire [WIDTH-1:0] wire_d69_43;
	wire [WIDTH-1:0] wire_d69_44;
	wire [WIDTH-1:0] wire_d69_45;
	wire [WIDTH-1:0] wire_d69_46;
	wire [WIDTH-1:0] wire_d69_47;
	wire [WIDTH-1:0] wire_d69_48;
	wire [WIDTH-1:0] wire_d69_49;
	wire [WIDTH-1:0] wire_d69_50;
	wire [WIDTH-1:0] wire_d69_51;
	wire [WIDTH-1:0] wire_d69_52;
	wire [WIDTH-1:0] wire_d69_53;
	wire [WIDTH-1:0] wire_d69_54;
	wire [WIDTH-1:0] wire_d69_55;
	wire [WIDTH-1:0] wire_d69_56;
	wire [WIDTH-1:0] wire_d69_57;
	wire [WIDTH-1:0] wire_d69_58;
	wire [WIDTH-1:0] wire_d69_59;
	wire [WIDTH-1:0] wire_d69_60;
	wire [WIDTH-1:0] wire_d69_61;
	wire [WIDTH-1:0] wire_d69_62;
	wire [WIDTH-1:0] wire_d69_63;
	wire [WIDTH-1:0] wire_d69_64;
	wire [WIDTH-1:0] wire_d69_65;
	wire [WIDTH-1:0] wire_d69_66;
	wire [WIDTH-1:0] wire_d69_67;
	wire [WIDTH-1:0] wire_d69_68;
	wire [WIDTH-1:0] wire_d69_69;
	wire [WIDTH-1:0] wire_d69_70;
	wire [WIDTH-1:0] wire_d69_71;
	wire [WIDTH-1:0] wire_d69_72;
	wire [WIDTH-1:0] wire_d69_73;
	wire [WIDTH-1:0] wire_d69_74;
	wire [WIDTH-1:0] wire_d69_75;
	wire [WIDTH-1:0] wire_d69_76;
	wire [WIDTH-1:0] wire_d69_77;
	wire [WIDTH-1:0] wire_d69_78;
	wire [WIDTH-1:0] wire_d69_79;
	wire [WIDTH-1:0] wire_d69_80;
	wire [WIDTH-1:0] wire_d69_81;
	wire [WIDTH-1:0] wire_d69_82;
	wire [WIDTH-1:0] wire_d69_83;
	wire [WIDTH-1:0] wire_d69_84;
	wire [WIDTH-1:0] wire_d69_85;
	wire [WIDTH-1:0] wire_d69_86;
	wire [WIDTH-1:0] wire_d69_87;
	wire [WIDTH-1:0] wire_d69_88;
	wire [WIDTH-1:0] wire_d69_89;
	wire [WIDTH-1:0] wire_d69_90;
	wire [WIDTH-1:0] wire_d69_91;
	wire [WIDTH-1:0] wire_d69_92;
	wire [WIDTH-1:0] wire_d69_93;
	wire [WIDTH-1:0] wire_d69_94;
	wire [WIDTH-1:0] wire_d69_95;
	wire [WIDTH-1:0] wire_d69_96;
	wire [WIDTH-1:0] wire_d69_97;
	wire [WIDTH-1:0] wire_d69_98;
	wire [WIDTH-1:0] wire_d69_99;
	wire [WIDTH-1:0] wire_d69_100;
	wire [WIDTH-1:0] wire_d69_101;
	wire [WIDTH-1:0] wire_d69_102;
	wire [WIDTH-1:0] wire_d69_103;
	wire [WIDTH-1:0] wire_d69_104;
	wire [WIDTH-1:0] wire_d69_105;
	wire [WIDTH-1:0] wire_d69_106;
	wire [WIDTH-1:0] wire_d69_107;
	wire [WIDTH-1:0] wire_d69_108;
	wire [WIDTH-1:0] wire_d69_109;
	wire [WIDTH-1:0] wire_d69_110;
	wire [WIDTH-1:0] wire_d69_111;
	wire [WIDTH-1:0] wire_d69_112;
	wire [WIDTH-1:0] wire_d69_113;
	wire [WIDTH-1:0] wire_d69_114;
	wire [WIDTH-1:0] wire_d69_115;
	wire [WIDTH-1:0] wire_d69_116;
	wire [WIDTH-1:0] wire_d69_117;
	wire [WIDTH-1:0] wire_d69_118;
	wire [WIDTH-1:0] wire_d70_0;
	wire [WIDTH-1:0] wire_d70_1;
	wire [WIDTH-1:0] wire_d70_2;
	wire [WIDTH-1:0] wire_d70_3;
	wire [WIDTH-1:0] wire_d70_4;
	wire [WIDTH-1:0] wire_d70_5;
	wire [WIDTH-1:0] wire_d70_6;
	wire [WIDTH-1:0] wire_d70_7;
	wire [WIDTH-1:0] wire_d70_8;
	wire [WIDTH-1:0] wire_d70_9;
	wire [WIDTH-1:0] wire_d70_10;
	wire [WIDTH-1:0] wire_d70_11;
	wire [WIDTH-1:0] wire_d70_12;
	wire [WIDTH-1:0] wire_d70_13;
	wire [WIDTH-1:0] wire_d70_14;
	wire [WIDTH-1:0] wire_d70_15;
	wire [WIDTH-1:0] wire_d70_16;
	wire [WIDTH-1:0] wire_d70_17;
	wire [WIDTH-1:0] wire_d70_18;
	wire [WIDTH-1:0] wire_d70_19;
	wire [WIDTH-1:0] wire_d70_20;
	wire [WIDTH-1:0] wire_d70_21;
	wire [WIDTH-1:0] wire_d70_22;
	wire [WIDTH-1:0] wire_d70_23;
	wire [WIDTH-1:0] wire_d70_24;
	wire [WIDTH-1:0] wire_d70_25;
	wire [WIDTH-1:0] wire_d70_26;
	wire [WIDTH-1:0] wire_d70_27;
	wire [WIDTH-1:0] wire_d70_28;
	wire [WIDTH-1:0] wire_d70_29;
	wire [WIDTH-1:0] wire_d70_30;
	wire [WIDTH-1:0] wire_d70_31;
	wire [WIDTH-1:0] wire_d70_32;
	wire [WIDTH-1:0] wire_d70_33;
	wire [WIDTH-1:0] wire_d70_34;
	wire [WIDTH-1:0] wire_d70_35;
	wire [WIDTH-1:0] wire_d70_36;
	wire [WIDTH-1:0] wire_d70_37;
	wire [WIDTH-1:0] wire_d70_38;
	wire [WIDTH-1:0] wire_d70_39;
	wire [WIDTH-1:0] wire_d70_40;
	wire [WIDTH-1:0] wire_d70_41;
	wire [WIDTH-1:0] wire_d70_42;
	wire [WIDTH-1:0] wire_d70_43;
	wire [WIDTH-1:0] wire_d70_44;
	wire [WIDTH-1:0] wire_d70_45;
	wire [WIDTH-1:0] wire_d70_46;
	wire [WIDTH-1:0] wire_d70_47;
	wire [WIDTH-1:0] wire_d70_48;
	wire [WIDTH-1:0] wire_d70_49;
	wire [WIDTH-1:0] wire_d70_50;
	wire [WIDTH-1:0] wire_d70_51;
	wire [WIDTH-1:0] wire_d70_52;
	wire [WIDTH-1:0] wire_d70_53;
	wire [WIDTH-1:0] wire_d70_54;
	wire [WIDTH-1:0] wire_d70_55;
	wire [WIDTH-1:0] wire_d70_56;
	wire [WIDTH-1:0] wire_d70_57;
	wire [WIDTH-1:0] wire_d70_58;
	wire [WIDTH-1:0] wire_d70_59;
	wire [WIDTH-1:0] wire_d70_60;
	wire [WIDTH-1:0] wire_d70_61;
	wire [WIDTH-1:0] wire_d70_62;
	wire [WIDTH-1:0] wire_d70_63;
	wire [WIDTH-1:0] wire_d70_64;
	wire [WIDTH-1:0] wire_d70_65;
	wire [WIDTH-1:0] wire_d70_66;
	wire [WIDTH-1:0] wire_d70_67;
	wire [WIDTH-1:0] wire_d70_68;
	wire [WIDTH-1:0] wire_d70_69;
	wire [WIDTH-1:0] wire_d70_70;
	wire [WIDTH-1:0] wire_d70_71;
	wire [WIDTH-1:0] wire_d70_72;
	wire [WIDTH-1:0] wire_d70_73;
	wire [WIDTH-1:0] wire_d70_74;
	wire [WIDTH-1:0] wire_d70_75;
	wire [WIDTH-1:0] wire_d70_76;
	wire [WIDTH-1:0] wire_d70_77;
	wire [WIDTH-1:0] wire_d70_78;
	wire [WIDTH-1:0] wire_d70_79;
	wire [WIDTH-1:0] wire_d70_80;
	wire [WIDTH-1:0] wire_d70_81;
	wire [WIDTH-1:0] wire_d70_82;
	wire [WIDTH-1:0] wire_d70_83;
	wire [WIDTH-1:0] wire_d70_84;
	wire [WIDTH-1:0] wire_d70_85;
	wire [WIDTH-1:0] wire_d70_86;
	wire [WIDTH-1:0] wire_d70_87;
	wire [WIDTH-1:0] wire_d70_88;
	wire [WIDTH-1:0] wire_d70_89;
	wire [WIDTH-1:0] wire_d70_90;
	wire [WIDTH-1:0] wire_d70_91;
	wire [WIDTH-1:0] wire_d70_92;
	wire [WIDTH-1:0] wire_d70_93;
	wire [WIDTH-1:0] wire_d70_94;
	wire [WIDTH-1:0] wire_d70_95;
	wire [WIDTH-1:0] wire_d70_96;
	wire [WIDTH-1:0] wire_d70_97;
	wire [WIDTH-1:0] wire_d70_98;
	wire [WIDTH-1:0] wire_d70_99;
	wire [WIDTH-1:0] wire_d70_100;
	wire [WIDTH-1:0] wire_d70_101;
	wire [WIDTH-1:0] wire_d70_102;
	wire [WIDTH-1:0] wire_d70_103;
	wire [WIDTH-1:0] wire_d70_104;
	wire [WIDTH-1:0] wire_d70_105;
	wire [WIDTH-1:0] wire_d70_106;
	wire [WIDTH-1:0] wire_d70_107;
	wire [WIDTH-1:0] wire_d70_108;
	wire [WIDTH-1:0] wire_d70_109;
	wire [WIDTH-1:0] wire_d70_110;
	wire [WIDTH-1:0] wire_d70_111;
	wire [WIDTH-1:0] wire_d70_112;
	wire [WIDTH-1:0] wire_d70_113;
	wire [WIDTH-1:0] wire_d70_114;
	wire [WIDTH-1:0] wire_d70_115;
	wire [WIDTH-1:0] wire_d70_116;
	wire [WIDTH-1:0] wire_d70_117;
	wire [WIDTH-1:0] wire_d70_118;
	wire [WIDTH-1:0] wire_d71_0;
	wire [WIDTH-1:0] wire_d71_1;
	wire [WIDTH-1:0] wire_d71_2;
	wire [WIDTH-1:0] wire_d71_3;
	wire [WIDTH-1:0] wire_d71_4;
	wire [WIDTH-1:0] wire_d71_5;
	wire [WIDTH-1:0] wire_d71_6;
	wire [WIDTH-1:0] wire_d71_7;
	wire [WIDTH-1:0] wire_d71_8;
	wire [WIDTH-1:0] wire_d71_9;
	wire [WIDTH-1:0] wire_d71_10;
	wire [WIDTH-1:0] wire_d71_11;
	wire [WIDTH-1:0] wire_d71_12;
	wire [WIDTH-1:0] wire_d71_13;
	wire [WIDTH-1:0] wire_d71_14;
	wire [WIDTH-1:0] wire_d71_15;
	wire [WIDTH-1:0] wire_d71_16;
	wire [WIDTH-1:0] wire_d71_17;
	wire [WIDTH-1:0] wire_d71_18;
	wire [WIDTH-1:0] wire_d71_19;
	wire [WIDTH-1:0] wire_d71_20;
	wire [WIDTH-1:0] wire_d71_21;
	wire [WIDTH-1:0] wire_d71_22;
	wire [WIDTH-1:0] wire_d71_23;
	wire [WIDTH-1:0] wire_d71_24;
	wire [WIDTH-1:0] wire_d71_25;
	wire [WIDTH-1:0] wire_d71_26;
	wire [WIDTH-1:0] wire_d71_27;
	wire [WIDTH-1:0] wire_d71_28;
	wire [WIDTH-1:0] wire_d71_29;
	wire [WIDTH-1:0] wire_d71_30;
	wire [WIDTH-1:0] wire_d71_31;
	wire [WIDTH-1:0] wire_d71_32;
	wire [WIDTH-1:0] wire_d71_33;
	wire [WIDTH-1:0] wire_d71_34;
	wire [WIDTH-1:0] wire_d71_35;
	wire [WIDTH-1:0] wire_d71_36;
	wire [WIDTH-1:0] wire_d71_37;
	wire [WIDTH-1:0] wire_d71_38;
	wire [WIDTH-1:0] wire_d71_39;
	wire [WIDTH-1:0] wire_d71_40;
	wire [WIDTH-1:0] wire_d71_41;
	wire [WIDTH-1:0] wire_d71_42;
	wire [WIDTH-1:0] wire_d71_43;
	wire [WIDTH-1:0] wire_d71_44;
	wire [WIDTH-1:0] wire_d71_45;
	wire [WIDTH-1:0] wire_d71_46;
	wire [WIDTH-1:0] wire_d71_47;
	wire [WIDTH-1:0] wire_d71_48;
	wire [WIDTH-1:0] wire_d71_49;
	wire [WIDTH-1:0] wire_d71_50;
	wire [WIDTH-1:0] wire_d71_51;
	wire [WIDTH-1:0] wire_d71_52;
	wire [WIDTH-1:0] wire_d71_53;
	wire [WIDTH-1:0] wire_d71_54;
	wire [WIDTH-1:0] wire_d71_55;
	wire [WIDTH-1:0] wire_d71_56;
	wire [WIDTH-1:0] wire_d71_57;
	wire [WIDTH-1:0] wire_d71_58;
	wire [WIDTH-1:0] wire_d71_59;
	wire [WIDTH-1:0] wire_d71_60;
	wire [WIDTH-1:0] wire_d71_61;
	wire [WIDTH-1:0] wire_d71_62;
	wire [WIDTH-1:0] wire_d71_63;
	wire [WIDTH-1:0] wire_d71_64;
	wire [WIDTH-1:0] wire_d71_65;
	wire [WIDTH-1:0] wire_d71_66;
	wire [WIDTH-1:0] wire_d71_67;
	wire [WIDTH-1:0] wire_d71_68;
	wire [WIDTH-1:0] wire_d71_69;
	wire [WIDTH-1:0] wire_d71_70;
	wire [WIDTH-1:0] wire_d71_71;
	wire [WIDTH-1:0] wire_d71_72;
	wire [WIDTH-1:0] wire_d71_73;
	wire [WIDTH-1:0] wire_d71_74;
	wire [WIDTH-1:0] wire_d71_75;
	wire [WIDTH-1:0] wire_d71_76;
	wire [WIDTH-1:0] wire_d71_77;
	wire [WIDTH-1:0] wire_d71_78;
	wire [WIDTH-1:0] wire_d71_79;
	wire [WIDTH-1:0] wire_d71_80;
	wire [WIDTH-1:0] wire_d71_81;
	wire [WIDTH-1:0] wire_d71_82;
	wire [WIDTH-1:0] wire_d71_83;
	wire [WIDTH-1:0] wire_d71_84;
	wire [WIDTH-1:0] wire_d71_85;
	wire [WIDTH-1:0] wire_d71_86;
	wire [WIDTH-1:0] wire_d71_87;
	wire [WIDTH-1:0] wire_d71_88;
	wire [WIDTH-1:0] wire_d71_89;
	wire [WIDTH-1:0] wire_d71_90;
	wire [WIDTH-1:0] wire_d71_91;
	wire [WIDTH-1:0] wire_d71_92;
	wire [WIDTH-1:0] wire_d71_93;
	wire [WIDTH-1:0] wire_d71_94;
	wire [WIDTH-1:0] wire_d71_95;
	wire [WIDTH-1:0] wire_d71_96;
	wire [WIDTH-1:0] wire_d71_97;
	wire [WIDTH-1:0] wire_d71_98;
	wire [WIDTH-1:0] wire_d71_99;
	wire [WIDTH-1:0] wire_d71_100;
	wire [WIDTH-1:0] wire_d71_101;
	wire [WIDTH-1:0] wire_d71_102;
	wire [WIDTH-1:0] wire_d71_103;
	wire [WIDTH-1:0] wire_d71_104;
	wire [WIDTH-1:0] wire_d71_105;
	wire [WIDTH-1:0] wire_d71_106;
	wire [WIDTH-1:0] wire_d71_107;
	wire [WIDTH-1:0] wire_d71_108;
	wire [WIDTH-1:0] wire_d71_109;
	wire [WIDTH-1:0] wire_d71_110;
	wire [WIDTH-1:0] wire_d71_111;
	wire [WIDTH-1:0] wire_d71_112;
	wire [WIDTH-1:0] wire_d71_113;
	wire [WIDTH-1:0] wire_d71_114;
	wire [WIDTH-1:0] wire_d71_115;
	wire [WIDTH-1:0] wire_d71_116;
	wire [WIDTH-1:0] wire_d71_117;
	wire [WIDTH-1:0] wire_d71_118;
	wire [WIDTH-1:0] wire_d72_0;
	wire [WIDTH-1:0] wire_d72_1;
	wire [WIDTH-1:0] wire_d72_2;
	wire [WIDTH-1:0] wire_d72_3;
	wire [WIDTH-1:0] wire_d72_4;
	wire [WIDTH-1:0] wire_d72_5;
	wire [WIDTH-1:0] wire_d72_6;
	wire [WIDTH-1:0] wire_d72_7;
	wire [WIDTH-1:0] wire_d72_8;
	wire [WIDTH-1:0] wire_d72_9;
	wire [WIDTH-1:0] wire_d72_10;
	wire [WIDTH-1:0] wire_d72_11;
	wire [WIDTH-1:0] wire_d72_12;
	wire [WIDTH-1:0] wire_d72_13;
	wire [WIDTH-1:0] wire_d72_14;
	wire [WIDTH-1:0] wire_d72_15;
	wire [WIDTH-1:0] wire_d72_16;
	wire [WIDTH-1:0] wire_d72_17;
	wire [WIDTH-1:0] wire_d72_18;
	wire [WIDTH-1:0] wire_d72_19;
	wire [WIDTH-1:0] wire_d72_20;
	wire [WIDTH-1:0] wire_d72_21;
	wire [WIDTH-1:0] wire_d72_22;
	wire [WIDTH-1:0] wire_d72_23;
	wire [WIDTH-1:0] wire_d72_24;
	wire [WIDTH-1:0] wire_d72_25;
	wire [WIDTH-1:0] wire_d72_26;
	wire [WIDTH-1:0] wire_d72_27;
	wire [WIDTH-1:0] wire_d72_28;
	wire [WIDTH-1:0] wire_d72_29;
	wire [WIDTH-1:0] wire_d72_30;
	wire [WIDTH-1:0] wire_d72_31;
	wire [WIDTH-1:0] wire_d72_32;
	wire [WIDTH-1:0] wire_d72_33;
	wire [WIDTH-1:0] wire_d72_34;
	wire [WIDTH-1:0] wire_d72_35;
	wire [WIDTH-1:0] wire_d72_36;
	wire [WIDTH-1:0] wire_d72_37;
	wire [WIDTH-1:0] wire_d72_38;
	wire [WIDTH-1:0] wire_d72_39;
	wire [WIDTH-1:0] wire_d72_40;
	wire [WIDTH-1:0] wire_d72_41;
	wire [WIDTH-1:0] wire_d72_42;
	wire [WIDTH-1:0] wire_d72_43;
	wire [WIDTH-1:0] wire_d72_44;
	wire [WIDTH-1:0] wire_d72_45;
	wire [WIDTH-1:0] wire_d72_46;
	wire [WIDTH-1:0] wire_d72_47;
	wire [WIDTH-1:0] wire_d72_48;
	wire [WIDTH-1:0] wire_d72_49;
	wire [WIDTH-1:0] wire_d72_50;
	wire [WIDTH-1:0] wire_d72_51;
	wire [WIDTH-1:0] wire_d72_52;
	wire [WIDTH-1:0] wire_d72_53;
	wire [WIDTH-1:0] wire_d72_54;
	wire [WIDTH-1:0] wire_d72_55;
	wire [WIDTH-1:0] wire_d72_56;
	wire [WIDTH-1:0] wire_d72_57;
	wire [WIDTH-1:0] wire_d72_58;
	wire [WIDTH-1:0] wire_d72_59;
	wire [WIDTH-1:0] wire_d72_60;
	wire [WIDTH-1:0] wire_d72_61;
	wire [WIDTH-1:0] wire_d72_62;
	wire [WIDTH-1:0] wire_d72_63;
	wire [WIDTH-1:0] wire_d72_64;
	wire [WIDTH-1:0] wire_d72_65;
	wire [WIDTH-1:0] wire_d72_66;
	wire [WIDTH-1:0] wire_d72_67;
	wire [WIDTH-1:0] wire_d72_68;
	wire [WIDTH-1:0] wire_d72_69;
	wire [WIDTH-1:0] wire_d72_70;
	wire [WIDTH-1:0] wire_d72_71;
	wire [WIDTH-1:0] wire_d72_72;
	wire [WIDTH-1:0] wire_d72_73;
	wire [WIDTH-1:0] wire_d72_74;
	wire [WIDTH-1:0] wire_d72_75;
	wire [WIDTH-1:0] wire_d72_76;
	wire [WIDTH-1:0] wire_d72_77;
	wire [WIDTH-1:0] wire_d72_78;
	wire [WIDTH-1:0] wire_d72_79;
	wire [WIDTH-1:0] wire_d72_80;
	wire [WIDTH-1:0] wire_d72_81;
	wire [WIDTH-1:0] wire_d72_82;
	wire [WIDTH-1:0] wire_d72_83;
	wire [WIDTH-1:0] wire_d72_84;
	wire [WIDTH-1:0] wire_d72_85;
	wire [WIDTH-1:0] wire_d72_86;
	wire [WIDTH-1:0] wire_d72_87;
	wire [WIDTH-1:0] wire_d72_88;
	wire [WIDTH-1:0] wire_d72_89;
	wire [WIDTH-1:0] wire_d72_90;
	wire [WIDTH-1:0] wire_d72_91;
	wire [WIDTH-1:0] wire_d72_92;
	wire [WIDTH-1:0] wire_d72_93;
	wire [WIDTH-1:0] wire_d72_94;
	wire [WIDTH-1:0] wire_d72_95;
	wire [WIDTH-1:0] wire_d72_96;
	wire [WIDTH-1:0] wire_d72_97;
	wire [WIDTH-1:0] wire_d72_98;
	wire [WIDTH-1:0] wire_d72_99;
	wire [WIDTH-1:0] wire_d72_100;
	wire [WIDTH-1:0] wire_d72_101;
	wire [WIDTH-1:0] wire_d72_102;
	wire [WIDTH-1:0] wire_d72_103;
	wire [WIDTH-1:0] wire_d72_104;
	wire [WIDTH-1:0] wire_d72_105;
	wire [WIDTH-1:0] wire_d72_106;
	wire [WIDTH-1:0] wire_d72_107;
	wire [WIDTH-1:0] wire_d72_108;
	wire [WIDTH-1:0] wire_d72_109;
	wire [WIDTH-1:0] wire_d72_110;
	wire [WIDTH-1:0] wire_d72_111;
	wire [WIDTH-1:0] wire_d72_112;
	wire [WIDTH-1:0] wire_d72_113;
	wire [WIDTH-1:0] wire_d72_114;
	wire [WIDTH-1:0] wire_d72_115;
	wire [WIDTH-1:0] wire_d72_116;
	wire [WIDTH-1:0] wire_d72_117;
	wire [WIDTH-1:0] wire_d72_118;
	wire [WIDTH-1:0] wire_d73_0;
	wire [WIDTH-1:0] wire_d73_1;
	wire [WIDTH-1:0] wire_d73_2;
	wire [WIDTH-1:0] wire_d73_3;
	wire [WIDTH-1:0] wire_d73_4;
	wire [WIDTH-1:0] wire_d73_5;
	wire [WIDTH-1:0] wire_d73_6;
	wire [WIDTH-1:0] wire_d73_7;
	wire [WIDTH-1:0] wire_d73_8;
	wire [WIDTH-1:0] wire_d73_9;
	wire [WIDTH-1:0] wire_d73_10;
	wire [WIDTH-1:0] wire_d73_11;
	wire [WIDTH-1:0] wire_d73_12;
	wire [WIDTH-1:0] wire_d73_13;
	wire [WIDTH-1:0] wire_d73_14;
	wire [WIDTH-1:0] wire_d73_15;
	wire [WIDTH-1:0] wire_d73_16;
	wire [WIDTH-1:0] wire_d73_17;
	wire [WIDTH-1:0] wire_d73_18;
	wire [WIDTH-1:0] wire_d73_19;
	wire [WIDTH-1:0] wire_d73_20;
	wire [WIDTH-1:0] wire_d73_21;
	wire [WIDTH-1:0] wire_d73_22;
	wire [WIDTH-1:0] wire_d73_23;
	wire [WIDTH-1:0] wire_d73_24;
	wire [WIDTH-1:0] wire_d73_25;
	wire [WIDTH-1:0] wire_d73_26;
	wire [WIDTH-1:0] wire_d73_27;
	wire [WIDTH-1:0] wire_d73_28;
	wire [WIDTH-1:0] wire_d73_29;
	wire [WIDTH-1:0] wire_d73_30;
	wire [WIDTH-1:0] wire_d73_31;
	wire [WIDTH-1:0] wire_d73_32;
	wire [WIDTH-1:0] wire_d73_33;
	wire [WIDTH-1:0] wire_d73_34;
	wire [WIDTH-1:0] wire_d73_35;
	wire [WIDTH-1:0] wire_d73_36;
	wire [WIDTH-1:0] wire_d73_37;
	wire [WIDTH-1:0] wire_d73_38;
	wire [WIDTH-1:0] wire_d73_39;
	wire [WIDTH-1:0] wire_d73_40;
	wire [WIDTH-1:0] wire_d73_41;
	wire [WIDTH-1:0] wire_d73_42;
	wire [WIDTH-1:0] wire_d73_43;
	wire [WIDTH-1:0] wire_d73_44;
	wire [WIDTH-1:0] wire_d73_45;
	wire [WIDTH-1:0] wire_d73_46;
	wire [WIDTH-1:0] wire_d73_47;
	wire [WIDTH-1:0] wire_d73_48;
	wire [WIDTH-1:0] wire_d73_49;
	wire [WIDTH-1:0] wire_d73_50;
	wire [WIDTH-1:0] wire_d73_51;
	wire [WIDTH-1:0] wire_d73_52;
	wire [WIDTH-1:0] wire_d73_53;
	wire [WIDTH-1:0] wire_d73_54;
	wire [WIDTH-1:0] wire_d73_55;
	wire [WIDTH-1:0] wire_d73_56;
	wire [WIDTH-1:0] wire_d73_57;
	wire [WIDTH-1:0] wire_d73_58;
	wire [WIDTH-1:0] wire_d73_59;
	wire [WIDTH-1:0] wire_d73_60;
	wire [WIDTH-1:0] wire_d73_61;
	wire [WIDTH-1:0] wire_d73_62;
	wire [WIDTH-1:0] wire_d73_63;
	wire [WIDTH-1:0] wire_d73_64;
	wire [WIDTH-1:0] wire_d73_65;
	wire [WIDTH-1:0] wire_d73_66;
	wire [WIDTH-1:0] wire_d73_67;
	wire [WIDTH-1:0] wire_d73_68;
	wire [WIDTH-1:0] wire_d73_69;
	wire [WIDTH-1:0] wire_d73_70;
	wire [WIDTH-1:0] wire_d73_71;
	wire [WIDTH-1:0] wire_d73_72;
	wire [WIDTH-1:0] wire_d73_73;
	wire [WIDTH-1:0] wire_d73_74;
	wire [WIDTH-1:0] wire_d73_75;
	wire [WIDTH-1:0] wire_d73_76;
	wire [WIDTH-1:0] wire_d73_77;
	wire [WIDTH-1:0] wire_d73_78;
	wire [WIDTH-1:0] wire_d73_79;
	wire [WIDTH-1:0] wire_d73_80;
	wire [WIDTH-1:0] wire_d73_81;
	wire [WIDTH-1:0] wire_d73_82;
	wire [WIDTH-1:0] wire_d73_83;
	wire [WIDTH-1:0] wire_d73_84;
	wire [WIDTH-1:0] wire_d73_85;
	wire [WIDTH-1:0] wire_d73_86;
	wire [WIDTH-1:0] wire_d73_87;
	wire [WIDTH-1:0] wire_d73_88;
	wire [WIDTH-1:0] wire_d73_89;
	wire [WIDTH-1:0] wire_d73_90;
	wire [WIDTH-1:0] wire_d73_91;
	wire [WIDTH-1:0] wire_d73_92;
	wire [WIDTH-1:0] wire_d73_93;
	wire [WIDTH-1:0] wire_d73_94;
	wire [WIDTH-1:0] wire_d73_95;
	wire [WIDTH-1:0] wire_d73_96;
	wire [WIDTH-1:0] wire_d73_97;
	wire [WIDTH-1:0] wire_d73_98;
	wire [WIDTH-1:0] wire_d73_99;
	wire [WIDTH-1:0] wire_d73_100;
	wire [WIDTH-1:0] wire_d73_101;
	wire [WIDTH-1:0] wire_d73_102;
	wire [WIDTH-1:0] wire_d73_103;
	wire [WIDTH-1:0] wire_d73_104;
	wire [WIDTH-1:0] wire_d73_105;
	wire [WIDTH-1:0] wire_d73_106;
	wire [WIDTH-1:0] wire_d73_107;
	wire [WIDTH-1:0] wire_d73_108;
	wire [WIDTH-1:0] wire_d73_109;
	wire [WIDTH-1:0] wire_d73_110;
	wire [WIDTH-1:0] wire_d73_111;
	wire [WIDTH-1:0] wire_d73_112;
	wire [WIDTH-1:0] wire_d73_113;
	wire [WIDTH-1:0] wire_d73_114;
	wire [WIDTH-1:0] wire_d73_115;
	wire [WIDTH-1:0] wire_d73_116;
	wire [WIDTH-1:0] wire_d73_117;
	wire [WIDTH-1:0] wire_d73_118;
	wire [WIDTH-1:0] wire_d74_0;
	wire [WIDTH-1:0] wire_d74_1;
	wire [WIDTH-1:0] wire_d74_2;
	wire [WIDTH-1:0] wire_d74_3;
	wire [WIDTH-1:0] wire_d74_4;
	wire [WIDTH-1:0] wire_d74_5;
	wire [WIDTH-1:0] wire_d74_6;
	wire [WIDTH-1:0] wire_d74_7;
	wire [WIDTH-1:0] wire_d74_8;
	wire [WIDTH-1:0] wire_d74_9;
	wire [WIDTH-1:0] wire_d74_10;
	wire [WIDTH-1:0] wire_d74_11;
	wire [WIDTH-1:0] wire_d74_12;
	wire [WIDTH-1:0] wire_d74_13;
	wire [WIDTH-1:0] wire_d74_14;
	wire [WIDTH-1:0] wire_d74_15;
	wire [WIDTH-1:0] wire_d74_16;
	wire [WIDTH-1:0] wire_d74_17;
	wire [WIDTH-1:0] wire_d74_18;
	wire [WIDTH-1:0] wire_d74_19;
	wire [WIDTH-1:0] wire_d74_20;
	wire [WIDTH-1:0] wire_d74_21;
	wire [WIDTH-1:0] wire_d74_22;
	wire [WIDTH-1:0] wire_d74_23;
	wire [WIDTH-1:0] wire_d74_24;
	wire [WIDTH-1:0] wire_d74_25;
	wire [WIDTH-1:0] wire_d74_26;
	wire [WIDTH-1:0] wire_d74_27;
	wire [WIDTH-1:0] wire_d74_28;
	wire [WIDTH-1:0] wire_d74_29;
	wire [WIDTH-1:0] wire_d74_30;
	wire [WIDTH-1:0] wire_d74_31;
	wire [WIDTH-1:0] wire_d74_32;
	wire [WIDTH-1:0] wire_d74_33;
	wire [WIDTH-1:0] wire_d74_34;
	wire [WIDTH-1:0] wire_d74_35;
	wire [WIDTH-1:0] wire_d74_36;
	wire [WIDTH-1:0] wire_d74_37;
	wire [WIDTH-1:0] wire_d74_38;
	wire [WIDTH-1:0] wire_d74_39;
	wire [WIDTH-1:0] wire_d74_40;
	wire [WIDTH-1:0] wire_d74_41;
	wire [WIDTH-1:0] wire_d74_42;
	wire [WIDTH-1:0] wire_d74_43;
	wire [WIDTH-1:0] wire_d74_44;
	wire [WIDTH-1:0] wire_d74_45;
	wire [WIDTH-1:0] wire_d74_46;
	wire [WIDTH-1:0] wire_d74_47;
	wire [WIDTH-1:0] wire_d74_48;
	wire [WIDTH-1:0] wire_d74_49;
	wire [WIDTH-1:0] wire_d74_50;
	wire [WIDTH-1:0] wire_d74_51;
	wire [WIDTH-1:0] wire_d74_52;
	wire [WIDTH-1:0] wire_d74_53;
	wire [WIDTH-1:0] wire_d74_54;
	wire [WIDTH-1:0] wire_d74_55;
	wire [WIDTH-1:0] wire_d74_56;
	wire [WIDTH-1:0] wire_d74_57;
	wire [WIDTH-1:0] wire_d74_58;
	wire [WIDTH-1:0] wire_d74_59;
	wire [WIDTH-1:0] wire_d74_60;
	wire [WIDTH-1:0] wire_d74_61;
	wire [WIDTH-1:0] wire_d74_62;
	wire [WIDTH-1:0] wire_d74_63;
	wire [WIDTH-1:0] wire_d74_64;
	wire [WIDTH-1:0] wire_d74_65;
	wire [WIDTH-1:0] wire_d74_66;
	wire [WIDTH-1:0] wire_d74_67;
	wire [WIDTH-1:0] wire_d74_68;
	wire [WIDTH-1:0] wire_d74_69;
	wire [WIDTH-1:0] wire_d74_70;
	wire [WIDTH-1:0] wire_d74_71;
	wire [WIDTH-1:0] wire_d74_72;
	wire [WIDTH-1:0] wire_d74_73;
	wire [WIDTH-1:0] wire_d74_74;
	wire [WIDTH-1:0] wire_d74_75;
	wire [WIDTH-1:0] wire_d74_76;
	wire [WIDTH-1:0] wire_d74_77;
	wire [WIDTH-1:0] wire_d74_78;
	wire [WIDTH-1:0] wire_d74_79;
	wire [WIDTH-1:0] wire_d74_80;
	wire [WIDTH-1:0] wire_d74_81;
	wire [WIDTH-1:0] wire_d74_82;
	wire [WIDTH-1:0] wire_d74_83;
	wire [WIDTH-1:0] wire_d74_84;
	wire [WIDTH-1:0] wire_d74_85;
	wire [WIDTH-1:0] wire_d74_86;
	wire [WIDTH-1:0] wire_d74_87;
	wire [WIDTH-1:0] wire_d74_88;
	wire [WIDTH-1:0] wire_d74_89;
	wire [WIDTH-1:0] wire_d74_90;
	wire [WIDTH-1:0] wire_d74_91;
	wire [WIDTH-1:0] wire_d74_92;
	wire [WIDTH-1:0] wire_d74_93;
	wire [WIDTH-1:0] wire_d74_94;
	wire [WIDTH-1:0] wire_d74_95;
	wire [WIDTH-1:0] wire_d74_96;
	wire [WIDTH-1:0] wire_d74_97;
	wire [WIDTH-1:0] wire_d74_98;
	wire [WIDTH-1:0] wire_d74_99;
	wire [WIDTH-1:0] wire_d74_100;
	wire [WIDTH-1:0] wire_d74_101;
	wire [WIDTH-1:0] wire_d74_102;
	wire [WIDTH-1:0] wire_d74_103;
	wire [WIDTH-1:0] wire_d74_104;
	wire [WIDTH-1:0] wire_d74_105;
	wire [WIDTH-1:0] wire_d74_106;
	wire [WIDTH-1:0] wire_d74_107;
	wire [WIDTH-1:0] wire_d74_108;
	wire [WIDTH-1:0] wire_d74_109;
	wire [WIDTH-1:0] wire_d74_110;
	wire [WIDTH-1:0] wire_d74_111;
	wire [WIDTH-1:0] wire_d74_112;
	wire [WIDTH-1:0] wire_d74_113;
	wire [WIDTH-1:0] wire_d74_114;
	wire [WIDTH-1:0] wire_d74_115;
	wire [WIDTH-1:0] wire_d74_116;
	wire [WIDTH-1:0] wire_d74_117;
	wire [WIDTH-1:0] wire_d74_118;
	wire [WIDTH-1:0] wire_d75_0;
	wire [WIDTH-1:0] wire_d75_1;
	wire [WIDTH-1:0] wire_d75_2;
	wire [WIDTH-1:0] wire_d75_3;
	wire [WIDTH-1:0] wire_d75_4;
	wire [WIDTH-1:0] wire_d75_5;
	wire [WIDTH-1:0] wire_d75_6;
	wire [WIDTH-1:0] wire_d75_7;
	wire [WIDTH-1:0] wire_d75_8;
	wire [WIDTH-1:0] wire_d75_9;
	wire [WIDTH-1:0] wire_d75_10;
	wire [WIDTH-1:0] wire_d75_11;
	wire [WIDTH-1:0] wire_d75_12;
	wire [WIDTH-1:0] wire_d75_13;
	wire [WIDTH-1:0] wire_d75_14;
	wire [WIDTH-1:0] wire_d75_15;
	wire [WIDTH-1:0] wire_d75_16;
	wire [WIDTH-1:0] wire_d75_17;
	wire [WIDTH-1:0] wire_d75_18;
	wire [WIDTH-1:0] wire_d75_19;
	wire [WIDTH-1:0] wire_d75_20;
	wire [WIDTH-1:0] wire_d75_21;
	wire [WIDTH-1:0] wire_d75_22;
	wire [WIDTH-1:0] wire_d75_23;
	wire [WIDTH-1:0] wire_d75_24;
	wire [WIDTH-1:0] wire_d75_25;
	wire [WIDTH-1:0] wire_d75_26;
	wire [WIDTH-1:0] wire_d75_27;
	wire [WIDTH-1:0] wire_d75_28;
	wire [WIDTH-1:0] wire_d75_29;
	wire [WIDTH-1:0] wire_d75_30;
	wire [WIDTH-1:0] wire_d75_31;
	wire [WIDTH-1:0] wire_d75_32;
	wire [WIDTH-1:0] wire_d75_33;
	wire [WIDTH-1:0] wire_d75_34;
	wire [WIDTH-1:0] wire_d75_35;
	wire [WIDTH-1:0] wire_d75_36;
	wire [WIDTH-1:0] wire_d75_37;
	wire [WIDTH-1:0] wire_d75_38;
	wire [WIDTH-1:0] wire_d75_39;
	wire [WIDTH-1:0] wire_d75_40;
	wire [WIDTH-1:0] wire_d75_41;
	wire [WIDTH-1:0] wire_d75_42;
	wire [WIDTH-1:0] wire_d75_43;
	wire [WIDTH-1:0] wire_d75_44;
	wire [WIDTH-1:0] wire_d75_45;
	wire [WIDTH-1:0] wire_d75_46;
	wire [WIDTH-1:0] wire_d75_47;
	wire [WIDTH-1:0] wire_d75_48;
	wire [WIDTH-1:0] wire_d75_49;
	wire [WIDTH-1:0] wire_d75_50;
	wire [WIDTH-1:0] wire_d75_51;
	wire [WIDTH-1:0] wire_d75_52;
	wire [WIDTH-1:0] wire_d75_53;
	wire [WIDTH-1:0] wire_d75_54;
	wire [WIDTH-1:0] wire_d75_55;
	wire [WIDTH-1:0] wire_d75_56;
	wire [WIDTH-1:0] wire_d75_57;
	wire [WIDTH-1:0] wire_d75_58;
	wire [WIDTH-1:0] wire_d75_59;
	wire [WIDTH-1:0] wire_d75_60;
	wire [WIDTH-1:0] wire_d75_61;
	wire [WIDTH-1:0] wire_d75_62;
	wire [WIDTH-1:0] wire_d75_63;
	wire [WIDTH-1:0] wire_d75_64;
	wire [WIDTH-1:0] wire_d75_65;
	wire [WIDTH-1:0] wire_d75_66;
	wire [WIDTH-1:0] wire_d75_67;
	wire [WIDTH-1:0] wire_d75_68;
	wire [WIDTH-1:0] wire_d75_69;
	wire [WIDTH-1:0] wire_d75_70;
	wire [WIDTH-1:0] wire_d75_71;
	wire [WIDTH-1:0] wire_d75_72;
	wire [WIDTH-1:0] wire_d75_73;
	wire [WIDTH-1:0] wire_d75_74;
	wire [WIDTH-1:0] wire_d75_75;
	wire [WIDTH-1:0] wire_d75_76;
	wire [WIDTH-1:0] wire_d75_77;
	wire [WIDTH-1:0] wire_d75_78;
	wire [WIDTH-1:0] wire_d75_79;
	wire [WIDTH-1:0] wire_d75_80;
	wire [WIDTH-1:0] wire_d75_81;
	wire [WIDTH-1:0] wire_d75_82;
	wire [WIDTH-1:0] wire_d75_83;
	wire [WIDTH-1:0] wire_d75_84;
	wire [WIDTH-1:0] wire_d75_85;
	wire [WIDTH-1:0] wire_d75_86;
	wire [WIDTH-1:0] wire_d75_87;
	wire [WIDTH-1:0] wire_d75_88;
	wire [WIDTH-1:0] wire_d75_89;
	wire [WIDTH-1:0] wire_d75_90;
	wire [WIDTH-1:0] wire_d75_91;
	wire [WIDTH-1:0] wire_d75_92;
	wire [WIDTH-1:0] wire_d75_93;
	wire [WIDTH-1:0] wire_d75_94;
	wire [WIDTH-1:0] wire_d75_95;
	wire [WIDTH-1:0] wire_d75_96;
	wire [WIDTH-1:0] wire_d75_97;
	wire [WIDTH-1:0] wire_d75_98;
	wire [WIDTH-1:0] wire_d75_99;
	wire [WIDTH-1:0] wire_d75_100;
	wire [WIDTH-1:0] wire_d75_101;
	wire [WIDTH-1:0] wire_d75_102;
	wire [WIDTH-1:0] wire_d75_103;
	wire [WIDTH-1:0] wire_d75_104;
	wire [WIDTH-1:0] wire_d75_105;
	wire [WIDTH-1:0] wire_d75_106;
	wire [WIDTH-1:0] wire_d75_107;
	wire [WIDTH-1:0] wire_d75_108;
	wire [WIDTH-1:0] wire_d75_109;
	wire [WIDTH-1:0] wire_d75_110;
	wire [WIDTH-1:0] wire_d75_111;
	wire [WIDTH-1:0] wire_d75_112;
	wire [WIDTH-1:0] wire_d75_113;
	wire [WIDTH-1:0] wire_d75_114;
	wire [WIDTH-1:0] wire_d75_115;
	wire [WIDTH-1:0] wire_d75_116;
	wire [WIDTH-1:0] wire_d75_117;
	wire [WIDTH-1:0] wire_d75_118;
	wire [WIDTH-1:0] wire_d76_0;
	wire [WIDTH-1:0] wire_d76_1;
	wire [WIDTH-1:0] wire_d76_2;
	wire [WIDTH-1:0] wire_d76_3;
	wire [WIDTH-1:0] wire_d76_4;
	wire [WIDTH-1:0] wire_d76_5;
	wire [WIDTH-1:0] wire_d76_6;
	wire [WIDTH-1:0] wire_d76_7;
	wire [WIDTH-1:0] wire_d76_8;
	wire [WIDTH-1:0] wire_d76_9;
	wire [WIDTH-1:0] wire_d76_10;
	wire [WIDTH-1:0] wire_d76_11;
	wire [WIDTH-1:0] wire_d76_12;
	wire [WIDTH-1:0] wire_d76_13;
	wire [WIDTH-1:0] wire_d76_14;
	wire [WIDTH-1:0] wire_d76_15;
	wire [WIDTH-1:0] wire_d76_16;
	wire [WIDTH-1:0] wire_d76_17;
	wire [WIDTH-1:0] wire_d76_18;
	wire [WIDTH-1:0] wire_d76_19;
	wire [WIDTH-1:0] wire_d76_20;
	wire [WIDTH-1:0] wire_d76_21;
	wire [WIDTH-1:0] wire_d76_22;
	wire [WIDTH-1:0] wire_d76_23;
	wire [WIDTH-1:0] wire_d76_24;
	wire [WIDTH-1:0] wire_d76_25;
	wire [WIDTH-1:0] wire_d76_26;
	wire [WIDTH-1:0] wire_d76_27;
	wire [WIDTH-1:0] wire_d76_28;
	wire [WIDTH-1:0] wire_d76_29;
	wire [WIDTH-1:0] wire_d76_30;
	wire [WIDTH-1:0] wire_d76_31;
	wire [WIDTH-1:0] wire_d76_32;
	wire [WIDTH-1:0] wire_d76_33;
	wire [WIDTH-1:0] wire_d76_34;
	wire [WIDTH-1:0] wire_d76_35;
	wire [WIDTH-1:0] wire_d76_36;
	wire [WIDTH-1:0] wire_d76_37;
	wire [WIDTH-1:0] wire_d76_38;
	wire [WIDTH-1:0] wire_d76_39;
	wire [WIDTH-1:0] wire_d76_40;
	wire [WIDTH-1:0] wire_d76_41;
	wire [WIDTH-1:0] wire_d76_42;
	wire [WIDTH-1:0] wire_d76_43;
	wire [WIDTH-1:0] wire_d76_44;
	wire [WIDTH-1:0] wire_d76_45;
	wire [WIDTH-1:0] wire_d76_46;
	wire [WIDTH-1:0] wire_d76_47;
	wire [WIDTH-1:0] wire_d76_48;
	wire [WIDTH-1:0] wire_d76_49;
	wire [WIDTH-1:0] wire_d76_50;
	wire [WIDTH-1:0] wire_d76_51;
	wire [WIDTH-1:0] wire_d76_52;
	wire [WIDTH-1:0] wire_d76_53;
	wire [WIDTH-1:0] wire_d76_54;
	wire [WIDTH-1:0] wire_d76_55;
	wire [WIDTH-1:0] wire_d76_56;
	wire [WIDTH-1:0] wire_d76_57;
	wire [WIDTH-1:0] wire_d76_58;
	wire [WIDTH-1:0] wire_d76_59;
	wire [WIDTH-1:0] wire_d76_60;
	wire [WIDTH-1:0] wire_d76_61;
	wire [WIDTH-1:0] wire_d76_62;
	wire [WIDTH-1:0] wire_d76_63;
	wire [WIDTH-1:0] wire_d76_64;
	wire [WIDTH-1:0] wire_d76_65;
	wire [WIDTH-1:0] wire_d76_66;
	wire [WIDTH-1:0] wire_d76_67;
	wire [WIDTH-1:0] wire_d76_68;
	wire [WIDTH-1:0] wire_d76_69;
	wire [WIDTH-1:0] wire_d76_70;
	wire [WIDTH-1:0] wire_d76_71;
	wire [WIDTH-1:0] wire_d76_72;
	wire [WIDTH-1:0] wire_d76_73;
	wire [WIDTH-1:0] wire_d76_74;
	wire [WIDTH-1:0] wire_d76_75;
	wire [WIDTH-1:0] wire_d76_76;
	wire [WIDTH-1:0] wire_d76_77;
	wire [WIDTH-1:0] wire_d76_78;
	wire [WIDTH-1:0] wire_d76_79;
	wire [WIDTH-1:0] wire_d76_80;
	wire [WIDTH-1:0] wire_d76_81;
	wire [WIDTH-1:0] wire_d76_82;
	wire [WIDTH-1:0] wire_d76_83;
	wire [WIDTH-1:0] wire_d76_84;
	wire [WIDTH-1:0] wire_d76_85;
	wire [WIDTH-1:0] wire_d76_86;
	wire [WIDTH-1:0] wire_d76_87;
	wire [WIDTH-1:0] wire_d76_88;
	wire [WIDTH-1:0] wire_d76_89;
	wire [WIDTH-1:0] wire_d76_90;
	wire [WIDTH-1:0] wire_d76_91;
	wire [WIDTH-1:0] wire_d76_92;
	wire [WIDTH-1:0] wire_d76_93;
	wire [WIDTH-1:0] wire_d76_94;
	wire [WIDTH-1:0] wire_d76_95;
	wire [WIDTH-1:0] wire_d76_96;
	wire [WIDTH-1:0] wire_d76_97;
	wire [WIDTH-1:0] wire_d76_98;
	wire [WIDTH-1:0] wire_d76_99;
	wire [WIDTH-1:0] wire_d76_100;
	wire [WIDTH-1:0] wire_d76_101;
	wire [WIDTH-1:0] wire_d76_102;
	wire [WIDTH-1:0] wire_d76_103;
	wire [WIDTH-1:0] wire_d76_104;
	wire [WIDTH-1:0] wire_d76_105;
	wire [WIDTH-1:0] wire_d76_106;
	wire [WIDTH-1:0] wire_d76_107;
	wire [WIDTH-1:0] wire_d76_108;
	wire [WIDTH-1:0] wire_d76_109;
	wire [WIDTH-1:0] wire_d76_110;
	wire [WIDTH-1:0] wire_d76_111;
	wire [WIDTH-1:0] wire_d76_112;
	wire [WIDTH-1:0] wire_d76_113;
	wire [WIDTH-1:0] wire_d76_114;
	wire [WIDTH-1:0] wire_d76_115;
	wire [WIDTH-1:0] wire_d76_116;
	wire [WIDTH-1:0] wire_d76_117;
	wire [WIDTH-1:0] wire_d76_118;
	wire [WIDTH-1:0] wire_d77_0;
	wire [WIDTH-1:0] wire_d77_1;
	wire [WIDTH-1:0] wire_d77_2;
	wire [WIDTH-1:0] wire_d77_3;
	wire [WIDTH-1:0] wire_d77_4;
	wire [WIDTH-1:0] wire_d77_5;
	wire [WIDTH-1:0] wire_d77_6;
	wire [WIDTH-1:0] wire_d77_7;
	wire [WIDTH-1:0] wire_d77_8;
	wire [WIDTH-1:0] wire_d77_9;
	wire [WIDTH-1:0] wire_d77_10;
	wire [WIDTH-1:0] wire_d77_11;
	wire [WIDTH-1:0] wire_d77_12;
	wire [WIDTH-1:0] wire_d77_13;
	wire [WIDTH-1:0] wire_d77_14;
	wire [WIDTH-1:0] wire_d77_15;
	wire [WIDTH-1:0] wire_d77_16;
	wire [WIDTH-1:0] wire_d77_17;
	wire [WIDTH-1:0] wire_d77_18;
	wire [WIDTH-1:0] wire_d77_19;
	wire [WIDTH-1:0] wire_d77_20;
	wire [WIDTH-1:0] wire_d77_21;
	wire [WIDTH-1:0] wire_d77_22;
	wire [WIDTH-1:0] wire_d77_23;
	wire [WIDTH-1:0] wire_d77_24;
	wire [WIDTH-1:0] wire_d77_25;
	wire [WIDTH-1:0] wire_d77_26;
	wire [WIDTH-1:0] wire_d77_27;
	wire [WIDTH-1:0] wire_d77_28;
	wire [WIDTH-1:0] wire_d77_29;
	wire [WIDTH-1:0] wire_d77_30;
	wire [WIDTH-1:0] wire_d77_31;
	wire [WIDTH-1:0] wire_d77_32;
	wire [WIDTH-1:0] wire_d77_33;
	wire [WIDTH-1:0] wire_d77_34;
	wire [WIDTH-1:0] wire_d77_35;
	wire [WIDTH-1:0] wire_d77_36;
	wire [WIDTH-1:0] wire_d77_37;
	wire [WIDTH-1:0] wire_d77_38;
	wire [WIDTH-1:0] wire_d77_39;
	wire [WIDTH-1:0] wire_d77_40;
	wire [WIDTH-1:0] wire_d77_41;
	wire [WIDTH-1:0] wire_d77_42;
	wire [WIDTH-1:0] wire_d77_43;
	wire [WIDTH-1:0] wire_d77_44;
	wire [WIDTH-1:0] wire_d77_45;
	wire [WIDTH-1:0] wire_d77_46;
	wire [WIDTH-1:0] wire_d77_47;
	wire [WIDTH-1:0] wire_d77_48;
	wire [WIDTH-1:0] wire_d77_49;
	wire [WIDTH-1:0] wire_d77_50;
	wire [WIDTH-1:0] wire_d77_51;
	wire [WIDTH-1:0] wire_d77_52;
	wire [WIDTH-1:0] wire_d77_53;
	wire [WIDTH-1:0] wire_d77_54;
	wire [WIDTH-1:0] wire_d77_55;
	wire [WIDTH-1:0] wire_d77_56;
	wire [WIDTH-1:0] wire_d77_57;
	wire [WIDTH-1:0] wire_d77_58;
	wire [WIDTH-1:0] wire_d77_59;
	wire [WIDTH-1:0] wire_d77_60;
	wire [WIDTH-1:0] wire_d77_61;
	wire [WIDTH-1:0] wire_d77_62;
	wire [WIDTH-1:0] wire_d77_63;
	wire [WIDTH-1:0] wire_d77_64;
	wire [WIDTH-1:0] wire_d77_65;
	wire [WIDTH-1:0] wire_d77_66;
	wire [WIDTH-1:0] wire_d77_67;
	wire [WIDTH-1:0] wire_d77_68;
	wire [WIDTH-1:0] wire_d77_69;
	wire [WIDTH-1:0] wire_d77_70;
	wire [WIDTH-1:0] wire_d77_71;
	wire [WIDTH-1:0] wire_d77_72;
	wire [WIDTH-1:0] wire_d77_73;
	wire [WIDTH-1:0] wire_d77_74;
	wire [WIDTH-1:0] wire_d77_75;
	wire [WIDTH-1:0] wire_d77_76;
	wire [WIDTH-1:0] wire_d77_77;
	wire [WIDTH-1:0] wire_d77_78;
	wire [WIDTH-1:0] wire_d77_79;
	wire [WIDTH-1:0] wire_d77_80;
	wire [WIDTH-1:0] wire_d77_81;
	wire [WIDTH-1:0] wire_d77_82;
	wire [WIDTH-1:0] wire_d77_83;
	wire [WIDTH-1:0] wire_d77_84;
	wire [WIDTH-1:0] wire_d77_85;
	wire [WIDTH-1:0] wire_d77_86;
	wire [WIDTH-1:0] wire_d77_87;
	wire [WIDTH-1:0] wire_d77_88;
	wire [WIDTH-1:0] wire_d77_89;
	wire [WIDTH-1:0] wire_d77_90;
	wire [WIDTH-1:0] wire_d77_91;
	wire [WIDTH-1:0] wire_d77_92;
	wire [WIDTH-1:0] wire_d77_93;
	wire [WIDTH-1:0] wire_d77_94;
	wire [WIDTH-1:0] wire_d77_95;
	wire [WIDTH-1:0] wire_d77_96;
	wire [WIDTH-1:0] wire_d77_97;
	wire [WIDTH-1:0] wire_d77_98;
	wire [WIDTH-1:0] wire_d77_99;
	wire [WIDTH-1:0] wire_d77_100;
	wire [WIDTH-1:0] wire_d77_101;
	wire [WIDTH-1:0] wire_d77_102;
	wire [WIDTH-1:0] wire_d77_103;
	wire [WIDTH-1:0] wire_d77_104;
	wire [WIDTH-1:0] wire_d77_105;
	wire [WIDTH-1:0] wire_d77_106;
	wire [WIDTH-1:0] wire_d77_107;
	wire [WIDTH-1:0] wire_d77_108;
	wire [WIDTH-1:0] wire_d77_109;
	wire [WIDTH-1:0] wire_d77_110;
	wire [WIDTH-1:0] wire_d77_111;
	wire [WIDTH-1:0] wire_d77_112;
	wire [WIDTH-1:0] wire_d77_113;
	wire [WIDTH-1:0] wire_d77_114;
	wire [WIDTH-1:0] wire_d77_115;
	wire [WIDTH-1:0] wire_d77_116;
	wire [WIDTH-1:0] wire_d77_117;
	wire [WIDTH-1:0] wire_d77_118;
	wire [WIDTH-1:0] wire_d78_0;
	wire [WIDTH-1:0] wire_d78_1;
	wire [WIDTH-1:0] wire_d78_2;
	wire [WIDTH-1:0] wire_d78_3;
	wire [WIDTH-1:0] wire_d78_4;
	wire [WIDTH-1:0] wire_d78_5;
	wire [WIDTH-1:0] wire_d78_6;
	wire [WIDTH-1:0] wire_d78_7;
	wire [WIDTH-1:0] wire_d78_8;
	wire [WIDTH-1:0] wire_d78_9;
	wire [WIDTH-1:0] wire_d78_10;
	wire [WIDTH-1:0] wire_d78_11;
	wire [WIDTH-1:0] wire_d78_12;
	wire [WIDTH-1:0] wire_d78_13;
	wire [WIDTH-1:0] wire_d78_14;
	wire [WIDTH-1:0] wire_d78_15;
	wire [WIDTH-1:0] wire_d78_16;
	wire [WIDTH-1:0] wire_d78_17;
	wire [WIDTH-1:0] wire_d78_18;
	wire [WIDTH-1:0] wire_d78_19;
	wire [WIDTH-1:0] wire_d78_20;
	wire [WIDTH-1:0] wire_d78_21;
	wire [WIDTH-1:0] wire_d78_22;
	wire [WIDTH-1:0] wire_d78_23;
	wire [WIDTH-1:0] wire_d78_24;
	wire [WIDTH-1:0] wire_d78_25;
	wire [WIDTH-1:0] wire_d78_26;
	wire [WIDTH-1:0] wire_d78_27;
	wire [WIDTH-1:0] wire_d78_28;
	wire [WIDTH-1:0] wire_d78_29;
	wire [WIDTH-1:0] wire_d78_30;
	wire [WIDTH-1:0] wire_d78_31;
	wire [WIDTH-1:0] wire_d78_32;
	wire [WIDTH-1:0] wire_d78_33;
	wire [WIDTH-1:0] wire_d78_34;
	wire [WIDTH-1:0] wire_d78_35;
	wire [WIDTH-1:0] wire_d78_36;
	wire [WIDTH-1:0] wire_d78_37;
	wire [WIDTH-1:0] wire_d78_38;
	wire [WIDTH-1:0] wire_d78_39;
	wire [WIDTH-1:0] wire_d78_40;
	wire [WIDTH-1:0] wire_d78_41;
	wire [WIDTH-1:0] wire_d78_42;
	wire [WIDTH-1:0] wire_d78_43;
	wire [WIDTH-1:0] wire_d78_44;
	wire [WIDTH-1:0] wire_d78_45;
	wire [WIDTH-1:0] wire_d78_46;
	wire [WIDTH-1:0] wire_d78_47;
	wire [WIDTH-1:0] wire_d78_48;
	wire [WIDTH-1:0] wire_d78_49;
	wire [WIDTH-1:0] wire_d78_50;
	wire [WIDTH-1:0] wire_d78_51;
	wire [WIDTH-1:0] wire_d78_52;
	wire [WIDTH-1:0] wire_d78_53;
	wire [WIDTH-1:0] wire_d78_54;
	wire [WIDTH-1:0] wire_d78_55;
	wire [WIDTH-1:0] wire_d78_56;
	wire [WIDTH-1:0] wire_d78_57;
	wire [WIDTH-1:0] wire_d78_58;
	wire [WIDTH-1:0] wire_d78_59;
	wire [WIDTH-1:0] wire_d78_60;
	wire [WIDTH-1:0] wire_d78_61;
	wire [WIDTH-1:0] wire_d78_62;
	wire [WIDTH-1:0] wire_d78_63;
	wire [WIDTH-1:0] wire_d78_64;
	wire [WIDTH-1:0] wire_d78_65;
	wire [WIDTH-1:0] wire_d78_66;
	wire [WIDTH-1:0] wire_d78_67;
	wire [WIDTH-1:0] wire_d78_68;
	wire [WIDTH-1:0] wire_d78_69;
	wire [WIDTH-1:0] wire_d78_70;
	wire [WIDTH-1:0] wire_d78_71;
	wire [WIDTH-1:0] wire_d78_72;
	wire [WIDTH-1:0] wire_d78_73;
	wire [WIDTH-1:0] wire_d78_74;
	wire [WIDTH-1:0] wire_d78_75;
	wire [WIDTH-1:0] wire_d78_76;
	wire [WIDTH-1:0] wire_d78_77;
	wire [WIDTH-1:0] wire_d78_78;
	wire [WIDTH-1:0] wire_d78_79;
	wire [WIDTH-1:0] wire_d78_80;
	wire [WIDTH-1:0] wire_d78_81;
	wire [WIDTH-1:0] wire_d78_82;
	wire [WIDTH-1:0] wire_d78_83;
	wire [WIDTH-1:0] wire_d78_84;
	wire [WIDTH-1:0] wire_d78_85;
	wire [WIDTH-1:0] wire_d78_86;
	wire [WIDTH-1:0] wire_d78_87;
	wire [WIDTH-1:0] wire_d78_88;
	wire [WIDTH-1:0] wire_d78_89;
	wire [WIDTH-1:0] wire_d78_90;
	wire [WIDTH-1:0] wire_d78_91;
	wire [WIDTH-1:0] wire_d78_92;
	wire [WIDTH-1:0] wire_d78_93;
	wire [WIDTH-1:0] wire_d78_94;
	wire [WIDTH-1:0] wire_d78_95;
	wire [WIDTH-1:0] wire_d78_96;
	wire [WIDTH-1:0] wire_d78_97;
	wire [WIDTH-1:0] wire_d78_98;
	wire [WIDTH-1:0] wire_d78_99;
	wire [WIDTH-1:0] wire_d78_100;
	wire [WIDTH-1:0] wire_d78_101;
	wire [WIDTH-1:0] wire_d78_102;
	wire [WIDTH-1:0] wire_d78_103;
	wire [WIDTH-1:0] wire_d78_104;
	wire [WIDTH-1:0] wire_d78_105;
	wire [WIDTH-1:0] wire_d78_106;
	wire [WIDTH-1:0] wire_d78_107;
	wire [WIDTH-1:0] wire_d78_108;
	wire [WIDTH-1:0] wire_d78_109;
	wire [WIDTH-1:0] wire_d78_110;
	wire [WIDTH-1:0] wire_d78_111;
	wire [WIDTH-1:0] wire_d78_112;
	wire [WIDTH-1:0] wire_d78_113;
	wire [WIDTH-1:0] wire_d78_114;
	wire [WIDTH-1:0] wire_d78_115;
	wire [WIDTH-1:0] wire_d78_116;
	wire [WIDTH-1:0] wire_d78_117;
	wire [WIDTH-1:0] wire_d78_118;
	wire [WIDTH-1:0] wire_d79_0;
	wire [WIDTH-1:0] wire_d79_1;
	wire [WIDTH-1:0] wire_d79_2;
	wire [WIDTH-1:0] wire_d79_3;
	wire [WIDTH-1:0] wire_d79_4;
	wire [WIDTH-1:0] wire_d79_5;
	wire [WIDTH-1:0] wire_d79_6;
	wire [WIDTH-1:0] wire_d79_7;
	wire [WIDTH-1:0] wire_d79_8;
	wire [WIDTH-1:0] wire_d79_9;
	wire [WIDTH-1:0] wire_d79_10;
	wire [WIDTH-1:0] wire_d79_11;
	wire [WIDTH-1:0] wire_d79_12;
	wire [WIDTH-1:0] wire_d79_13;
	wire [WIDTH-1:0] wire_d79_14;
	wire [WIDTH-1:0] wire_d79_15;
	wire [WIDTH-1:0] wire_d79_16;
	wire [WIDTH-1:0] wire_d79_17;
	wire [WIDTH-1:0] wire_d79_18;
	wire [WIDTH-1:0] wire_d79_19;
	wire [WIDTH-1:0] wire_d79_20;
	wire [WIDTH-1:0] wire_d79_21;
	wire [WIDTH-1:0] wire_d79_22;
	wire [WIDTH-1:0] wire_d79_23;
	wire [WIDTH-1:0] wire_d79_24;
	wire [WIDTH-1:0] wire_d79_25;
	wire [WIDTH-1:0] wire_d79_26;
	wire [WIDTH-1:0] wire_d79_27;
	wire [WIDTH-1:0] wire_d79_28;
	wire [WIDTH-1:0] wire_d79_29;
	wire [WIDTH-1:0] wire_d79_30;
	wire [WIDTH-1:0] wire_d79_31;
	wire [WIDTH-1:0] wire_d79_32;
	wire [WIDTH-1:0] wire_d79_33;
	wire [WIDTH-1:0] wire_d79_34;
	wire [WIDTH-1:0] wire_d79_35;
	wire [WIDTH-1:0] wire_d79_36;
	wire [WIDTH-1:0] wire_d79_37;
	wire [WIDTH-1:0] wire_d79_38;
	wire [WIDTH-1:0] wire_d79_39;
	wire [WIDTH-1:0] wire_d79_40;
	wire [WIDTH-1:0] wire_d79_41;
	wire [WIDTH-1:0] wire_d79_42;
	wire [WIDTH-1:0] wire_d79_43;
	wire [WIDTH-1:0] wire_d79_44;
	wire [WIDTH-1:0] wire_d79_45;
	wire [WIDTH-1:0] wire_d79_46;
	wire [WIDTH-1:0] wire_d79_47;
	wire [WIDTH-1:0] wire_d79_48;
	wire [WIDTH-1:0] wire_d79_49;
	wire [WIDTH-1:0] wire_d79_50;
	wire [WIDTH-1:0] wire_d79_51;
	wire [WIDTH-1:0] wire_d79_52;
	wire [WIDTH-1:0] wire_d79_53;
	wire [WIDTH-1:0] wire_d79_54;
	wire [WIDTH-1:0] wire_d79_55;
	wire [WIDTH-1:0] wire_d79_56;
	wire [WIDTH-1:0] wire_d79_57;
	wire [WIDTH-1:0] wire_d79_58;
	wire [WIDTH-1:0] wire_d79_59;
	wire [WIDTH-1:0] wire_d79_60;
	wire [WIDTH-1:0] wire_d79_61;
	wire [WIDTH-1:0] wire_d79_62;
	wire [WIDTH-1:0] wire_d79_63;
	wire [WIDTH-1:0] wire_d79_64;
	wire [WIDTH-1:0] wire_d79_65;
	wire [WIDTH-1:0] wire_d79_66;
	wire [WIDTH-1:0] wire_d79_67;
	wire [WIDTH-1:0] wire_d79_68;
	wire [WIDTH-1:0] wire_d79_69;
	wire [WIDTH-1:0] wire_d79_70;
	wire [WIDTH-1:0] wire_d79_71;
	wire [WIDTH-1:0] wire_d79_72;
	wire [WIDTH-1:0] wire_d79_73;
	wire [WIDTH-1:0] wire_d79_74;
	wire [WIDTH-1:0] wire_d79_75;
	wire [WIDTH-1:0] wire_d79_76;
	wire [WIDTH-1:0] wire_d79_77;
	wire [WIDTH-1:0] wire_d79_78;
	wire [WIDTH-1:0] wire_d79_79;
	wire [WIDTH-1:0] wire_d79_80;
	wire [WIDTH-1:0] wire_d79_81;
	wire [WIDTH-1:0] wire_d79_82;
	wire [WIDTH-1:0] wire_d79_83;
	wire [WIDTH-1:0] wire_d79_84;
	wire [WIDTH-1:0] wire_d79_85;
	wire [WIDTH-1:0] wire_d79_86;
	wire [WIDTH-1:0] wire_d79_87;
	wire [WIDTH-1:0] wire_d79_88;
	wire [WIDTH-1:0] wire_d79_89;
	wire [WIDTH-1:0] wire_d79_90;
	wire [WIDTH-1:0] wire_d79_91;
	wire [WIDTH-1:0] wire_d79_92;
	wire [WIDTH-1:0] wire_d79_93;
	wire [WIDTH-1:0] wire_d79_94;
	wire [WIDTH-1:0] wire_d79_95;
	wire [WIDTH-1:0] wire_d79_96;
	wire [WIDTH-1:0] wire_d79_97;
	wire [WIDTH-1:0] wire_d79_98;
	wire [WIDTH-1:0] wire_d79_99;
	wire [WIDTH-1:0] wire_d79_100;
	wire [WIDTH-1:0] wire_d79_101;
	wire [WIDTH-1:0] wire_d79_102;
	wire [WIDTH-1:0] wire_d79_103;
	wire [WIDTH-1:0] wire_d79_104;
	wire [WIDTH-1:0] wire_d79_105;
	wire [WIDTH-1:0] wire_d79_106;
	wire [WIDTH-1:0] wire_d79_107;
	wire [WIDTH-1:0] wire_d79_108;
	wire [WIDTH-1:0] wire_d79_109;
	wire [WIDTH-1:0] wire_d79_110;
	wire [WIDTH-1:0] wire_d79_111;
	wire [WIDTH-1:0] wire_d79_112;
	wire [WIDTH-1:0] wire_d79_113;
	wire [WIDTH-1:0] wire_d79_114;
	wire [WIDTH-1:0] wire_d79_115;
	wire [WIDTH-1:0] wire_d79_116;
	wire [WIDTH-1:0] wire_d79_117;
	wire [WIDTH-1:0] wire_d79_118;
	wire [WIDTH-1:0] wire_d80_0;
	wire [WIDTH-1:0] wire_d80_1;
	wire [WIDTH-1:0] wire_d80_2;
	wire [WIDTH-1:0] wire_d80_3;
	wire [WIDTH-1:0] wire_d80_4;
	wire [WIDTH-1:0] wire_d80_5;
	wire [WIDTH-1:0] wire_d80_6;
	wire [WIDTH-1:0] wire_d80_7;
	wire [WIDTH-1:0] wire_d80_8;
	wire [WIDTH-1:0] wire_d80_9;
	wire [WIDTH-1:0] wire_d80_10;
	wire [WIDTH-1:0] wire_d80_11;
	wire [WIDTH-1:0] wire_d80_12;
	wire [WIDTH-1:0] wire_d80_13;
	wire [WIDTH-1:0] wire_d80_14;
	wire [WIDTH-1:0] wire_d80_15;
	wire [WIDTH-1:0] wire_d80_16;
	wire [WIDTH-1:0] wire_d80_17;
	wire [WIDTH-1:0] wire_d80_18;
	wire [WIDTH-1:0] wire_d80_19;
	wire [WIDTH-1:0] wire_d80_20;
	wire [WIDTH-1:0] wire_d80_21;
	wire [WIDTH-1:0] wire_d80_22;
	wire [WIDTH-1:0] wire_d80_23;
	wire [WIDTH-1:0] wire_d80_24;
	wire [WIDTH-1:0] wire_d80_25;
	wire [WIDTH-1:0] wire_d80_26;
	wire [WIDTH-1:0] wire_d80_27;
	wire [WIDTH-1:0] wire_d80_28;
	wire [WIDTH-1:0] wire_d80_29;
	wire [WIDTH-1:0] wire_d80_30;
	wire [WIDTH-1:0] wire_d80_31;
	wire [WIDTH-1:0] wire_d80_32;
	wire [WIDTH-1:0] wire_d80_33;
	wire [WIDTH-1:0] wire_d80_34;
	wire [WIDTH-1:0] wire_d80_35;
	wire [WIDTH-1:0] wire_d80_36;
	wire [WIDTH-1:0] wire_d80_37;
	wire [WIDTH-1:0] wire_d80_38;
	wire [WIDTH-1:0] wire_d80_39;
	wire [WIDTH-1:0] wire_d80_40;
	wire [WIDTH-1:0] wire_d80_41;
	wire [WIDTH-1:0] wire_d80_42;
	wire [WIDTH-1:0] wire_d80_43;
	wire [WIDTH-1:0] wire_d80_44;
	wire [WIDTH-1:0] wire_d80_45;
	wire [WIDTH-1:0] wire_d80_46;
	wire [WIDTH-1:0] wire_d80_47;
	wire [WIDTH-1:0] wire_d80_48;
	wire [WIDTH-1:0] wire_d80_49;
	wire [WIDTH-1:0] wire_d80_50;
	wire [WIDTH-1:0] wire_d80_51;
	wire [WIDTH-1:0] wire_d80_52;
	wire [WIDTH-1:0] wire_d80_53;
	wire [WIDTH-1:0] wire_d80_54;
	wire [WIDTH-1:0] wire_d80_55;
	wire [WIDTH-1:0] wire_d80_56;
	wire [WIDTH-1:0] wire_d80_57;
	wire [WIDTH-1:0] wire_d80_58;
	wire [WIDTH-1:0] wire_d80_59;
	wire [WIDTH-1:0] wire_d80_60;
	wire [WIDTH-1:0] wire_d80_61;
	wire [WIDTH-1:0] wire_d80_62;
	wire [WIDTH-1:0] wire_d80_63;
	wire [WIDTH-1:0] wire_d80_64;
	wire [WIDTH-1:0] wire_d80_65;
	wire [WIDTH-1:0] wire_d80_66;
	wire [WIDTH-1:0] wire_d80_67;
	wire [WIDTH-1:0] wire_d80_68;
	wire [WIDTH-1:0] wire_d80_69;
	wire [WIDTH-1:0] wire_d80_70;
	wire [WIDTH-1:0] wire_d80_71;
	wire [WIDTH-1:0] wire_d80_72;
	wire [WIDTH-1:0] wire_d80_73;
	wire [WIDTH-1:0] wire_d80_74;
	wire [WIDTH-1:0] wire_d80_75;
	wire [WIDTH-1:0] wire_d80_76;
	wire [WIDTH-1:0] wire_d80_77;
	wire [WIDTH-1:0] wire_d80_78;
	wire [WIDTH-1:0] wire_d80_79;
	wire [WIDTH-1:0] wire_d80_80;
	wire [WIDTH-1:0] wire_d80_81;
	wire [WIDTH-1:0] wire_d80_82;
	wire [WIDTH-1:0] wire_d80_83;
	wire [WIDTH-1:0] wire_d80_84;
	wire [WIDTH-1:0] wire_d80_85;
	wire [WIDTH-1:0] wire_d80_86;
	wire [WIDTH-1:0] wire_d80_87;
	wire [WIDTH-1:0] wire_d80_88;
	wire [WIDTH-1:0] wire_d80_89;
	wire [WIDTH-1:0] wire_d80_90;
	wire [WIDTH-1:0] wire_d80_91;
	wire [WIDTH-1:0] wire_d80_92;
	wire [WIDTH-1:0] wire_d80_93;
	wire [WIDTH-1:0] wire_d80_94;
	wire [WIDTH-1:0] wire_d80_95;
	wire [WIDTH-1:0] wire_d80_96;
	wire [WIDTH-1:0] wire_d80_97;
	wire [WIDTH-1:0] wire_d80_98;
	wire [WIDTH-1:0] wire_d80_99;
	wire [WIDTH-1:0] wire_d80_100;
	wire [WIDTH-1:0] wire_d80_101;
	wire [WIDTH-1:0] wire_d80_102;
	wire [WIDTH-1:0] wire_d80_103;
	wire [WIDTH-1:0] wire_d80_104;
	wire [WIDTH-1:0] wire_d80_105;
	wire [WIDTH-1:0] wire_d80_106;
	wire [WIDTH-1:0] wire_d80_107;
	wire [WIDTH-1:0] wire_d80_108;
	wire [WIDTH-1:0] wire_d80_109;
	wire [WIDTH-1:0] wire_d80_110;
	wire [WIDTH-1:0] wire_d80_111;
	wire [WIDTH-1:0] wire_d80_112;
	wire [WIDTH-1:0] wire_d80_113;
	wire [WIDTH-1:0] wire_d80_114;
	wire [WIDTH-1:0] wire_d80_115;
	wire [WIDTH-1:0] wire_d80_116;
	wire [WIDTH-1:0] wire_d80_117;
	wire [WIDTH-1:0] wire_d80_118;
	wire [WIDTH-1:0] wire_d81_0;
	wire [WIDTH-1:0] wire_d81_1;
	wire [WIDTH-1:0] wire_d81_2;
	wire [WIDTH-1:0] wire_d81_3;
	wire [WIDTH-1:0] wire_d81_4;
	wire [WIDTH-1:0] wire_d81_5;
	wire [WIDTH-1:0] wire_d81_6;
	wire [WIDTH-1:0] wire_d81_7;
	wire [WIDTH-1:0] wire_d81_8;
	wire [WIDTH-1:0] wire_d81_9;
	wire [WIDTH-1:0] wire_d81_10;
	wire [WIDTH-1:0] wire_d81_11;
	wire [WIDTH-1:0] wire_d81_12;
	wire [WIDTH-1:0] wire_d81_13;
	wire [WIDTH-1:0] wire_d81_14;
	wire [WIDTH-1:0] wire_d81_15;
	wire [WIDTH-1:0] wire_d81_16;
	wire [WIDTH-1:0] wire_d81_17;
	wire [WIDTH-1:0] wire_d81_18;
	wire [WIDTH-1:0] wire_d81_19;
	wire [WIDTH-1:0] wire_d81_20;
	wire [WIDTH-1:0] wire_d81_21;
	wire [WIDTH-1:0] wire_d81_22;
	wire [WIDTH-1:0] wire_d81_23;
	wire [WIDTH-1:0] wire_d81_24;
	wire [WIDTH-1:0] wire_d81_25;
	wire [WIDTH-1:0] wire_d81_26;
	wire [WIDTH-1:0] wire_d81_27;
	wire [WIDTH-1:0] wire_d81_28;
	wire [WIDTH-1:0] wire_d81_29;
	wire [WIDTH-1:0] wire_d81_30;
	wire [WIDTH-1:0] wire_d81_31;
	wire [WIDTH-1:0] wire_d81_32;
	wire [WIDTH-1:0] wire_d81_33;
	wire [WIDTH-1:0] wire_d81_34;
	wire [WIDTH-1:0] wire_d81_35;
	wire [WIDTH-1:0] wire_d81_36;
	wire [WIDTH-1:0] wire_d81_37;
	wire [WIDTH-1:0] wire_d81_38;
	wire [WIDTH-1:0] wire_d81_39;
	wire [WIDTH-1:0] wire_d81_40;
	wire [WIDTH-1:0] wire_d81_41;
	wire [WIDTH-1:0] wire_d81_42;
	wire [WIDTH-1:0] wire_d81_43;
	wire [WIDTH-1:0] wire_d81_44;
	wire [WIDTH-1:0] wire_d81_45;
	wire [WIDTH-1:0] wire_d81_46;
	wire [WIDTH-1:0] wire_d81_47;
	wire [WIDTH-1:0] wire_d81_48;
	wire [WIDTH-1:0] wire_d81_49;
	wire [WIDTH-1:0] wire_d81_50;
	wire [WIDTH-1:0] wire_d81_51;
	wire [WIDTH-1:0] wire_d81_52;
	wire [WIDTH-1:0] wire_d81_53;
	wire [WIDTH-1:0] wire_d81_54;
	wire [WIDTH-1:0] wire_d81_55;
	wire [WIDTH-1:0] wire_d81_56;
	wire [WIDTH-1:0] wire_d81_57;
	wire [WIDTH-1:0] wire_d81_58;
	wire [WIDTH-1:0] wire_d81_59;
	wire [WIDTH-1:0] wire_d81_60;
	wire [WIDTH-1:0] wire_d81_61;
	wire [WIDTH-1:0] wire_d81_62;
	wire [WIDTH-1:0] wire_d81_63;
	wire [WIDTH-1:0] wire_d81_64;
	wire [WIDTH-1:0] wire_d81_65;
	wire [WIDTH-1:0] wire_d81_66;
	wire [WIDTH-1:0] wire_d81_67;
	wire [WIDTH-1:0] wire_d81_68;
	wire [WIDTH-1:0] wire_d81_69;
	wire [WIDTH-1:0] wire_d81_70;
	wire [WIDTH-1:0] wire_d81_71;
	wire [WIDTH-1:0] wire_d81_72;
	wire [WIDTH-1:0] wire_d81_73;
	wire [WIDTH-1:0] wire_d81_74;
	wire [WIDTH-1:0] wire_d81_75;
	wire [WIDTH-1:0] wire_d81_76;
	wire [WIDTH-1:0] wire_d81_77;
	wire [WIDTH-1:0] wire_d81_78;
	wire [WIDTH-1:0] wire_d81_79;
	wire [WIDTH-1:0] wire_d81_80;
	wire [WIDTH-1:0] wire_d81_81;
	wire [WIDTH-1:0] wire_d81_82;
	wire [WIDTH-1:0] wire_d81_83;
	wire [WIDTH-1:0] wire_d81_84;
	wire [WIDTH-1:0] wire_d81_85;
	wire [WIDTH-1:0] wire_d81_86;
	wire [WIDTH-1:0] wire_d81_87;
	wire [WIDTH-1:0] wire_d81_88;
	wire [WIDTH-1:0] wire_d81_89;
	wire [WIDTH-1:0] wire_d81_90;
	wire [WIDTH-1:0] wire_d81_91;
	wire [WIDTH-1:0] wire_d81_92;
	wire [WIDTH-1:0] wire_d81_93;
	wire [WIDTH-1:0] wire_d81_94;
	wire [WIDTH-1:0] wire_d81_95;
	wire [WIDTH-1:0] wire_d81_96;
	wire [WIDTH-1:0] wire_d81_97;
	wire [WIDTH-1:0] wire_d81_98;
	wire [WIDTH-1:0] wire_d81_99;
	wire [WIDTH-1:0] wire_d81_100;
	wire [WIDTH-1:0] wire_d81_101;
	wire [WIDTH-1:0] wire_d81_102;
	wire [WIDTH-1:0] wire_d81_103;
	wire [WIDTH-1:0] wire_d81_104;
	wire [WIDTH-1:0] wire_d81_105;
	wire [WIDTH-1:0] wire_d81_106;
	wire [WIDTH-1:0] wire_d81_107;
	wire [WIDTH-1:0] wire_d81_108;
	wire [WIDTH-1:0] wire_d81_109;
	wire [WIDTH-1:0] wire_d81_110;
	wire [WIDTH-1:0] wire_d81_111;
	wire [WIDTH-1:0] wire_d81_112;
	wire [WIDTH-1:0] wire_d81_113;
	wire [WIDTH-1:0] wire_d81_114;
	wire [WIDTH-1:0] wire_d81_115;
	wire [WIDTH-1:0] wire_d81_116;
	wire [WIDTH-1:0] wire_d81_117;
	wire [WIDTH-1:0] wire_d81_118;
	wire [WIDTH-1:0] wire_d82_0;
	wire [WIDTH-1:0] wire_d82_1;
	wire [WIDTH-1:0] wire_d82_2;
	wire [WIDTH-1:0] wire_d82_3;
	wire [WIDTH-1:0] wire_d82_4;
	wire [WIDTH-1:0] wire_d82_5;
	wire [WIDTH-1:0] wire_d82_6;
	wire [WIDTH-1:0] wire_d82_7;
	wire [WIDTH-1:0] wire_d82_8;
	wire [WIDTH-1:0] wire_d82_9;
	wire [WIDTH-1:0] wire_d82_10;
	wire [WIDTH-1:0] wire_d82_11;
	wire [WIDTH-1:0] wire_d82_12;
	wire [WIDTH-1:0] wire_d82_13;
	wire [WIDTH-1:0] wire_d82_14;
	wire [WIDTH-1:0] wire_d82_15;
	wire [WIDTH-1:0] wire_d82_16;
	wire [WIDTH-1:0] wire_d82_17;
	wire [WIDTH-1:0] wire_d82_18;
	wire [WIDTH-1:0] wire_d82_19;
	wire [WIDTH-1:0] wire_d82_20;
	wire [WIDTH-1:0] wire_d82_21;
	wire [WIDTH-1:0] wire_d82_22;
	wire [WIDTH-1:0] wire_d82_23;
	wire [WIDTH-1:0] wire_d82_24;
	wire [WIDTH-1:0] wire_d82_25;
	wire [WIDTH-1:0] wire_d82_26;
	wire [WIDTH-1:0] wire_d82_27;
	wire [WIDTH-1:0] wire_d82_28;
	wire [WIDTH-1:0] wire_d82_29;
	wire [WIDTH-1:0] wire_d82_30;
	wire [WIDTH-1:0] wire_d82_31;
	wire [WIDTH-1:0] wire_d82_32;
	wire [WIDTH-1:0] wire_d82_33;
	wire [WIDTH-1:0] wire_d82_34;
	wire [WIDTH-1:0] wire_d82_35;
	wire [WIDTH-1:0] wire_d82_36;
	wire [WIDTH-1:0] wire_d82_37;
	wire [WIDTH-1:0] wire_d82_38;
	wire [WIDTH-1:0] wire_d82_39;
	wire [WIDTH-1:0] wire_d82_40;
	wire [WIDTH-1:0] wire_d82_41;
	wire [WIDTH-1:0] wire_d82_42;
	wire [WIDTH-1:0] wire_d82_43;
	wire [WIDTH-1:0] wire_d82_44;
	wire [WIDTH-1:0] wire_d82_45;
	wire [WIDTH-1:0] wire_d82_46;
	wire [WIDTH-1:0] wire_d82_47;
	wire [WIDTH-1:0] wire_d82_48;
	wire [WIDTH-1:0] wire_d82_49;
	wire [WIDTH-1:0] wire_d82_50;
	wire [WIDTH-1:0] wire_d82_51;
	wire [WIDTH-1:0] wire_d82_52;
	wire [WIDTH-1:0] wire_d82_53;
	wire [WIDTH-1:0] wire_d82_54;
	wire [WIDTH-1:0] wire_d82_55;
	wire [WIDTH-1:0] wire_d82_56;
	wire [WIDTH-1:0] wire_d82_57;
	wire [WIDTH-1:0] wire_d82_58;
	wire [WIDTH-1:0] wire_d82_59;
	wire [WIDTH-1:0] wire_d82_60;
	wire [WIDTH-1:0] wire_d82_61;
	wire [WIDTH-1:0] wire_d82_62;
	wire [WIDTH-1:0] wire_d82_63;
	wire [WIDTH-1:0] wire_d82_64;
	wire [WIDTH-1:0] wire_d82_65;
	wire [WIDTH-1:0] wire_d82_66;
	wire [WIDTH-1:0] wire_d82_67;
	wire [WIDTH-1:0] wire_d82_68;
	wire [WIDTH-1:0] wire_d82_69;
	wire [WIDTH-1:0] wire_d82_70;
	wire [WIDTH-1:0] wire_d82_71;
	wire [WIDTH-1:0] wire_d82_72;
	wire [WIDTH-1:0] wire_d82_73;
	wire [WIDTH-1:0] wire_d82_74;
	wire [WIDTH-1:0] wire_d82_75;
	wire [WIDTH-1:0] wire_d82_76;
	wire [WIDTH-1:0] wire_d82_77;
	wire [WIDTH-1:0] wire_d82_78;
	wire [WIDTH-1:0] wire_d82_79;
	wire [WIDTH-1:0] wire_d82_80;
	wire [WIDTH-1:0] wire_d82_81;
	wire [WIDTH-1:0] wire_d82_82;
	wire [WIDTH-1:0] wire_d82_83;
	wire [WIDTH-1:0] wire_d82_84;
	wire [WIDTH-1:0] wire_d82_85;
	wire [WIDTH-1:0] wire_d82_86;
	wire [WIDTH-1:0] wire_d82_87;
	wire [WIDTH-1:0] wire_d82_88;
	wire [WIDTH-1:0] wire_d82_89;
	wire [WIDTH-1:0] wire_d82_90;
	wire [WIDTH-1:0] wire_d82_91;
	wire [WIDTH-1:0] wire_d82_92;
	wire [WIDTH-1:0] wire_d82_93;
	wire [WIDTH-1:0] wire_d82_94;
	wire [WIDTH-1:0] wire_d82_95;
	wire [WIDTH-1:0] wire_d82_96;
	wire [WIDTH-1:0] wire_d82_97;
	wire [WIDTH-1:0] wire_d82_98;
	wire [WIDTH-1:0] wire_d82_99;
	wire [WIDTH-1:0] wire_d82_100;
	wire [WIDTH-1:0] wire_d82_101;
	wire [WIDTH-1:0] wire_d82_102;
	wire [WIDTH-1:0] wire_d82_103;
	wire [WIDTH-1:0] wire_d82_104;
	wire [WIDTH-1:0] wire_d82_105;
	wire [WIDTH-1:0] wire_d82_106;
	wire [WIDTH-1:0] wire_d82_107;
	wire [WIDTH-1:0] wire_d82_108;
	wire [WIDTH-1:0] wire_d82_109;
	wire [WIDTH-1:0] wire_d82_110;
	wire [WIDTH-1:0] wire_d82_111;
	wire [WIDTH-1:0] wire_d82_112;
	wire [WIDTH-1:0] wire_d82_113;
	wire [WIDTH-1:0] wire_d82_114;
	wire [WIDTH-1:0] wire_d82_115;
	wire [WIDTH-1:0] wire_d82_116;
	wire [WIDTH-1:0] wire_d82_117;
	wire [WIDTH-1:0] wire_d82_118;
	wire [WIDTH-1:0] wire_d83_0;
	wire [WIDTH-1:0] wire_d83_1;
	wire [WIDTH-1:0] wire_d83_2;
	wire [WIDTH-1:0] wire_d83_3;
	wire [WIDTH-1:0] wire_d83_4;
	wire [WIDTH-1:0] wire_d83_5;
	wire [WIDTH-1:0] wire_d83_6;
	wire [WIDTH-1:0] wire_d83_7;
	wire [WIDTH-1:0] wire_d83_8;
	wire [WIDTH-1:0] wire_d83_9;
	wire [WIDTH-1:0] wire_d83_10;
	wire [WIDTH-1:0] wire_d83_11;
	wire [WIDTH-1:0] wire_d83_12;
	wire [WIDTH-1:0] wire_d83_13;
	wire [WIDTH-1:0] wire_d83_14;
	wire [WIDTH-1:0] wire_d83_15;
	wire [WIDTH-1:0] wire_d83_16;
	wire [WIDTH-1:0] wire_d83_17;
	wire [WIDTH-1:0] wire_d83_18;
	wire [WIDTH-1:0] wire_d83_19;
	wire [WIDTH-1:0] wire_d83_20;
	wire [WIDTH-1:0] wire_d83_21;
	wire [WIDTH-1:0] wire_d83_22;
	wire [WIDTH-1:0] wire_d83_23;
	wire [WIDTH-1:0] wire_d83_24;
	wire [WIDTH-1:0] wire_d83_25;
	wire [WIDTH-1:0] wire_d83_26;
	wire [WIDTH-1:0] wire_d83_27;
	wire [WIDTH-1:0] wire_d83_28;
	wire [WIDTH-1:0] wire_d83_29;
	wire [WIDTH-1:0] wire_d83_30;
	wire [WIDTH-1:0] wire_d83_31;
	wire [WIDTH-1:0] wire_d83_32;
	wire [WIDTH-1:0] wire_d83_33;
	wire [WIDTH-1:0] wire_d83_34;
	wire [WIDTH-1:0] wire_d83_35;
	wire [WIDTH-1:0] wire_d83_36;
	wire [WIDTH-1:0] wire_d83_37;
	wire [WIDTH-1:0] wire_d83_38;
	wire [WIDTH-1:0] wire_d83_39;
	wire [WIDTH-1:0] wire_d83_40;
	wire [WIDTH-1:0] wire_d83_41;
	wire [WIDTH-1:0] wire_d83_42;
	wire [WIDTH-1:0] wire_d83_43;
	wire [WIDTH-1:0] wire_d83_44;
	wire [WIDTH-1:0] wire_d83_45;
	wire [WIDTH-1:0] wire_d83_46;
	wire [WIDTH-1:0] wire_d83_47;
	wire [WIDTH-1:0] wire_d83_48;
	wire [WIDTH-1:0] wire_d83_49;
	wire [WIDTH-1:0] wire_d83_50;
	wire [WIDTH-1:0] wire_d83_51;
	wire [WIDTH-1:0] wire_d83_52;
	wire [WIDTH-1:0] wire_d83_53;
	wire [WIDTH-1:0] wire_d83_54;
	wire [WIDTH-1:0] wire_d83_55;
	wire [WIDTH-1:0] wire_d83_56;
	wire [WIDTH-1:0] wire_d83_57;
	wire [WIDTH-1:0] wire_d83_58;
	wire [WIDTH-1:0] wire_d83_59;
	wire [WIDTH-1:0] wire_d83_60;
	wire [WIDTH-1:0] wire_d83_61;
	wire [WIDTH-1:0] wire_d83_62;
	wire [WIDTH-1:0] wire_d83_63;
	wire [WIDTH-1:0] wire_d83_64;
	wire [WIDTH-1:0] wire_d83_65;
	wire [WIDTH-1:0] wire_d83_66;
	wire [WIDTH-1:0] wire_d83_67;
	wire [WIDTH-1:0] wire_d83_68;
	wire [WIDTH-1:0] wire_d83_69;
	wire [WIDTH-1:0] wire_d83_70;
	wire [WIDTH-1:0] wire_d83_71;
	wire [WIDTH-1:0] wire_d83_72;
	wire [WIDTH-1:0] wire_d83_73;
	wire [WIDTH-1:0] wire_d83_74;
	wire [WIDTH-1:0] wire_d83_75;
	wire [WIDTH-1:0] wire_d83_76;
	wire [WIDTH-1:0] wire_d83_77;
	wire [WIDTH-1:0] wire_d83_78;
	wire [WIDTH-1:0] wire_d83_79;
	wire [WIDTH-1:0] wire_d83_80;
	wire [WIDTH-1:0] wire_d83_81;
	wire [WIDTH-1:0] wire_d83_82;
	wire [WIDTH-1:0] wire_d83_83;
	wire [WIDTH-1:0] wire_d83_84;
	wire [WIDTH-1:0] wire_d83_85;
	wire [WIDTH-1:0] wire_d83_86;
	wire [WIDTH-1:0] wire_d83_87;
	wire [WIDTH-1:0] wire_d83_88;
	wire [WIDTH-1:0] wire_d83_89;
	wire [WIDTH-1:0] wire_d83_90;
	wire [WIDTH-1:0] wire_d83_91;
	wire [WIDTH-1:0] wire_d83_92;
	wire [WIDTH-1:0] wire_d83_93;
	wire [WIDTH-1:0] wire_d83_94;
	wire [WIDTH-1:0] wire_d83_95;
	wire [WIDTH-1:0] wire_d83_96;
	wire [WIDTH-1:0] wire_d83_97;
	wire [WIDTH-1:0] wire_d83_98;
	wire [WIDTH-1:0] wire_d83_99;
	wire [WIDTH-1:0] wire_d83_100;
	wire [WIDTH-1:0] wire_d83_101;
	wire [WIDTH-1:0] wire_d83_102;
	wire [WIDTH-1:0] wire_d83_103;
	wire [WIDTH-1:0] wire_d83_104;
	wire [WIDTH-1:0] wire_d83_105;
	wire [WIDTH-1:0] wire_d83_106;
	wire [WIDTH-1:0] wire_d83_107;
	wire [WIDTH-1:0] wire_d83_108;
	wire [WIDTH-1:0] wire_d83_109;
	wire [WIDTH-1:0] wire_d83_110;
	wire [WIDTH-1:0] wire_d83_111;
	wire [WIDTH-1:0] wire_d83_112;
	wire [WIDTH-1:0] wire_d83_113;
	wire [WIDTH-1:0] wire_d83_114;
	wire [WIDTH-1:0] wire_d83_115;
	wire [WIDTH-1:0] wire_d83_116;
	wire [WIDTH-1:0] wire_d83_117;
	wire [WIDTH-1:0] wire_d83_118;
	wire [WIDTH-1:0] wire_d84_0;
	wire [WIDTH-1:0] wire_d84_1;
	wire [WIDTH-1:0] wire_d84_2;
	wire [WIDTH-1:0] wire_d84_3;
	wire [WIDTH-1:0] wire_d84_4;
	wire [WIDTH-1:0] wire_d84_5;
	wire [WIDTH-1:0] wire_d84_6;
	wire [WIDTH-1:0] wire_d84_7;
	wire [WIDTH-1:0] wire_d84_8;
	wire [WIDTH-1:0] wire_d84_9;
	wire [WIDTH-1:0] wire_d84_10;
	wire [WIDTH-1:0] wire_d84_11;
	wire [WIDTH-1:0] wire_d84_12;
	wire [WIDTH-1:0] wire_d84_13;
	wire [WIDTH-1:0] wire_d84_14;
	wire [WIDTH-1:0] wire_d84_15;
	wire [WIDTH-1:0] wire_d84_16;
	wire [WIDTH-1:0] wire_d84_17;
	wire [WIDTH-1:0] wire_d84_18;
	wire [WIDTH-1:0] wire_d84_19;
	wire [WIDTH-1:0] wire_d84_20;
	wire [WIDTH-1:0] wire_d84_21;
	wire [WIDTH-1:0] wire_d84_22;
	wire [WIDTH-1:0] wire_d84_23;
	wire [WIDTH-1:0] wire_d84_24;
	wire [WIDTH-1:0] wire_d84_25;
	wire [WIDTH-1:0] wire_d84_26;
	wire [WIDTH-1:0] wire_d84_27;
	wire [WIDTH-1:0] wire_d84_28;
	wire [WIDTH-1:0] wire_d84_29;
	wire [WIDTH-1:0] wire_d84_30;
	wire [WIDTH-1:0] wire_d84_31;
	wire [WIDTH-1:0] wire_d84_32;
	wire [WIDTH-1:0] wire_d84_33;
	wire [WIDTH-1:0] wire_d84_34;
	wire [WIDTH-1:0] wire_d84_35;
	wire [WIDTH-1:0] wire_d84_36;
	wire [WIDTH-1:0] wire_d84_37;
	wire [WIDTH-1:0] wire_d84_38;
	wire [WIDTH-1:0] wire_d84_39;
	wire [WIDTH-1:0] wire_d84_40;
	wire [WIDTH-1:0] wire_d84_41;
	wire [WIDTH-1:0] wire_d84_42;
	wire [WIDTH-1:0] wire_d84_43;
	wire [WIDTH-1:0] wire_d84_44;
	wire [WIDTH-1:0] wire_d84_45;
	wire [WIDTH-1:0] wire_d84_46;
	wire [WIDTH-1:0] wire_d84_47;
	wire [WIDTH-1:0] wire_d84_48;
	wire [WIDTH-1:0] wire_d84_49;
	wire [WIDTH-1:0] wire_d84_50;
	wire [WIDTH-1:0] wire_d84_51;
	wire [WIDTH-1:0] wire_d84_52;
	wire [WIDTH-1:0] wire_d84_53;
	wire [WIDTH-1:0] wire_d84_54;
	wire [WIDTH-1:0] wire_d84_55;
	wire [WIDTH-1:0] wire_d84_56;
	wire [WIDTH-1:0] wire_d84_57;
	wire [WIDTH-1:0] wire_d84_58;
	wire [WIDTH-1:0] wire_d84_59;
	wire [WIDTH-1:0] wire_d84_60;
	wire [WIDTH-1:0] wire_d84_61;
	wire [WIDTH-1:0] wire_d84_62;
	wire [WIDTH-1:0] wire_d84_63;
	wire [WIDTH-1:0] wire_d84_64;
	wire [WIDTH-1:0] wire_d84_65;
	wire [WIDTH-1:0] wire_d84_66;
	wire [WIDTH-1:0] wire_d84_67;
	wire [WIDTH-1:0] wire_d84_68;
	wire [WIDTH-1:0] wire_d84_69;
	wire [WIDTH-1:0] wire_d84_70;
	wire [WIDTH-1:0] wire_d84_71;
	wire [WIDTH-1:0] wire_d84_72;
	wire [WIDTH-1:0] wire_d84_73;
	wire [WIDTH-1:0] wire_d84_74;
	wire [WIDTH-1:0] wire_d84_75;
	wire [WIDTH-1:0] wire_d84_76;
	wire [WIDTH-1:0] wire_d84_77;
	wire [WIDTH-1:0] wire_d84_78;
	wire [WIDTH-1:0] wire_d84_79;
	wire [WIDTH-1:0] wire_d84_80;
	wire [WIDTH-1:0] wire_d84_81;
	wire [WIDTH-1:0] wire_d84_82;
	wire [WIDTH-1:0] wire_d84_83;
	wire [WIDTH-1:0] wire_d84_84;
	wire [WIDTH-1:0] wire_d84_85;
	wire [WIDTH-1:0] wire_d84_86;
	wire [WIDTH-1:0] wire_d84_87;
	wire [WIDTH-1:0] wire_d84_88;
	wire [WIDTH-1:0] wire_d84_89;
	wire [WIDTH-1:0] wire_d84_90;
	wire [WIDTH-1:0] wire_d84_91;
	wire [WIDTH-1:0] wire_d84_92;
	wire [WIDTH-1:0] wire_d84_93;
	wire [WIDTH-1:0] wire_d84_94;
	wire [WIDTH-1:0] wire_d84_95;
	wire [WIDTH-1:0] wire_d84_96;
	wire [WIDTH-1:0] wire_d84_97;
	wire [WIDTH-1:0] wire_d84_98;
	wire [WIDTH-1:0] wire_d84_99;
	wire [WIDTH-1:0] wire_d84_100;
	wire [WIDTH-1:0] wire_d84_101;
	wire [WIDTH-1:0] wire_d84_102;
	wire [WIDTH-1:0] wire_d84_103;
	wire [WIDTH-1:0] wire_d84_104;
	wire [WIDTH-1:0] wire_d84_105;
	wire [WIDTH-1:0] wire_d84_106;
	wire [WIDTH-1:0] wire_d84_107;
	wire [WIDTH-1:0] wire_d84_108;
	wire [WIDTH-1:0] wire_d84_109;
	wire [WIDTH-1:0] wire_d84_110;
	wire [WIDTH-1:0] wire_d84_111;
	wire [WIDTH-1:0] wire_d84_112;
	wire [WIDTH-1:0] wire_d84_113;
	wire [WIDTH-1:0] wire_d84_114;
	wire [WIDTH-1:0] wire_d84_115;
	wire [WIDTH-1:0] wire_d84_116;
	wire [WIDTH-1:0] wire_d84_117;
	wire [WIDTH-1:0] wire_d84_118;
	wire [WIDTH-1:0] wire_d85_0;
	wire [WIDTH-1:0] wire_d85_1;
	wire [WIDTH-1:0] wire_d85_2;
	wire [WIDTH-1:0] wire_d85_3;
	wire [WIDTH-1:0] wire_d85_4;
	wire [WIDTH-1:0] wire_d85_5;
	wire [WIDTH-1:0] wire_d85_6;
	wire [WIDTH-1:0] wire_d85_7;
	wire [WIDTH-1:0] wire_d85_8;
	wire [WIDTH-1:0] wire_d85_9;
	wire [WIDTH-1:0] wire_d85_10;
	wire [WIDTH-1:0] wire_d85_11;
	wire [WIDTH-1:0] wire_d85_12;
	wire [WIDTH-1:0] wire_d85_13;
	wire [WIDTH-1:0] wire_d85_14;
	wire [WIDTH-1:0] wire_d85_15;
	wire [WIDTH-1:0] wire_d85_16;
	wire [WIDTH-1:0] wire_d85_17;
	wire [WIDTH-1:0] wire_d85_18;
	wire [WIDTH-1:0] wire_d85_19;
	wire [WIDTH-1:0] wire_d85_20;
	wire [WIDTH-1:0] wire_d85_21;
	wire [WIDTH-1:0] wire_d85_22;
	wire [WIDTH-1:0] wire_d85_23;
	wire [WIDTH-1:0] wire_d85_24;
	wire [WIDTH-1:0] wire_d85_25;
	wire [WIDTH-1:0] wire_d85_26;
	wire [WIDTH-1:0] wire_d85_27;
	wire [WIDTH-1:0] wire_d85_28;
	wire [WIDTH-1:0] wire_d85_29;
	wire [WIDTH-1:0] wire_d85_30;
	wire [WIDTH-1:0] wire_d85_31;
	wire [WIDTH-1:0] wire_d85_32;
	wire [WIDTH-1:0] wire_d85_33;
	wire [WIDTH-1:0] wire_d85_34;
	wire [WIDTH-1:0] wire_d85_35;
	wire [WIDTH-1:0] wire_d85_36;
	wire [WIDTH-1:0] wire_d85_37;
	wire [WIDTH-1:0] wire_d85_38;
	wire [WIDTH-1:0] wire_d85_39;
	wire [WIDTH-1:0] wire_d85_40;
	wire [WIDTH-1:0] wire_d85_41;
	wire [WIDTH-1:0] wire_d85_42;
	wire [WIDTH-1:0] wire_d85_43;
	wire [WIDTH-1:0] wire_d85_44;
	wire [WIDTH-1:0] wire_d85_45;
	wire [WIDTH-1:0] wire_d85_46;
	wire [WIDTH-1:0] wire_d85_47;
	wire [WIDTH-1:0] wire_d85_48;
	wire [WIDTH-1:0] wire_d85_49;
	wire [WIDTH-1:0] wire_d85_50;
	wire [WIDTH-1:0] wire_d85_51;
	wire [WIDTH-1:0] wire_d85_52;
	wire [WIDTH-1:0] wire_d85_53;
	wire [WIDTH-1:0] wire_d85_54;
	wire [WIDTH-1:0] wire_d85_55;
	wire [WIDTH-1:0] wire_d85_56;
	wire [WIDTH-1:0] wire_d85_57;
	wire [WIDTH-1:0] wire_d85_58;
	wire [WIDTH-1:0] wire_d85_59;
	wire [WIDTH-1:0] wire_d85_60;
	wire [WIDTH-1:0] wire_d85_61;
	wire [WIDTH-1:0] wire_d85_62;
	wire [WIDTH-1:0] wire_d85_63;
	wire [WIDTH-1:0] wire_d85_64;
	wire [WIDTH-1:0] wire_d85_65;
	wire [WIDTH-1:0] wire_d85_66;
	wire [WIDTH-1:0] wire_d85_67;
	wire [WIDTH-1:0] wire_d85_68;
	wire [WIDTH-1:0] wire_d85_69;
	wire [WIDTH-1:0] wire_d85_70;
	wire [WIDTH-1:0] wire_d85_71;
	wire [WIDTH-1:0] wire_d85_72;
	wire [WIDTH-1:0] wire_d85_73;
	wire [WIDTH-1:0] wire_d85_74;
	wire [WIDTH-1:0] wire_d85_75;
	wire [WIDTH-1:0] wire_d85_76;
	wire [WIDTH-1:0] wire_d85_77;
	wire [WIDTH-1:0] wire_d85_78;
	wire [WIDTH-1:0] wire_d85_79;
	wire [WIDTH-1:0] wire_d85_80;
	wire [WIDTH-1:0] wire_d85_81;
	wire [WIDTH-1:0] wire_d85_82;
	wire [WIDTH-1:0] wire_d85_83;
	wire [WIDTH-1:0] wire_d85_84;
	wire [WIDTH-1:0] wire_d85_85;
	wire [WIDTH-1:0] wire_d85_86;
	wire [WIDTH-1:0] wire_d85_87;
	wire [WIDTH-1:0] wire_d85_88;
	wire [WIDTH-1:0] wire_d85_89;
	wire [WIDTH-1:0] wire_d85_90;
	wire [WIDTH-1:0] wire_d85_91;
	wire [WIDTH-1:0] wire_d85_92;
	wire [WIDTH-1:0] wire_d85_93;
	wire [WIDTH-1:0] wire_d85_94;
	wire [WIDTH-1:0] wire_d85_95;
	wire [WIDTH-1:0] wire_d85_96;
	wire [WIDTH-1:0] wire_d85_97;
	wire [WIDTH-1:0] wire_d85_98;
	wire [WIDTH-1:0] wire_d85_99;
	wire [WIDTH-1:0] wire_d85_100;
	wire [WIDTH-1:0] wire_d85_101;
	wire [WIDTH-1:0] wire_d85_102;
	wire [WIDTH-1:0] wire_d85_103;
	wire [WIDTH-1:0] wire_d85_104;
	wire [WIDTH-1:0] wire_d85_105;
	wire [WIDTH-1:0] wire_d85_106;
	wire [WIDTH-1:0] wire_d85_107;
	wire [WIDTH-1:0] wire_d85_108;
	wire [WIDTH-1:0] wire_d85_109;
	wire [WIDTH-1:0] wire_d85_110;
	wire [WIDTH-1:0] wire_d85_111;
	wire [WIDTH-1:0] wire_d85_112;
	wire [WIDTH-1:0] wire_d85_113;
	wire [WIDTH-1:0] wire_d85_114;
	wire [WIDTH-1:0] wire_d85_115;
	wire [WIDTH-1:0] wire_d85_116;
	wire [WIDTH-1:0] wire_d85_117;
	wire [WIDTH-1:0] wire_d85_118;
	wire [WIDTH-1:0] wire_d86_0;
	wire [WIDTH-1:0] wire_d86_1;
	wire [WIDTH-1:0] wire_d86_2;
	wire [WIDTH-1:0] wire_d86_3;
	wire [WIDTH-1:0] wire_d86_4;
	wire [WIDTH-1:0] wire_d86_5;
	wire [WIDTH-1:0] wire_d86_6;
	wire [WIDTH-1:0] wire_d86_7;
	wire [WIDTH-1:0] wire_d86_8;
	wire [WIDTH-1:0] wire_d86_9;
	wire [WIDTH-1:0] wire_d86_10;
	wire [WIDTH-1:0] wire_d86_11;
	wire [WIDTH-1:0] wire_d86_12;
	wire [WIDTH-1:0] wire_d86_13;
	wire [WIDTH-1:0] wire_d86_14;
	wire [WIDTH-1:0] wire_d86_15;
	wire [WIDTH-1:0] wire_d86_16;
	wire [WIDTH-1:0] wire_d86_17;
	wire [WIDTH-1:0] wire_d86_18;
	wire [WIDTH-1:0] wire_d86_19;
	wire [WIDTH-1:0] wire_d86_20;
	wire [WIDTH-1:0] wire_d86_21;
	wire [WIDTH-1:0] wire_d86_22;
	wire [WIDTH-1:0] wire_d86_23;
	wire [WIDTH-1:0] wire_d86_24;
	wire [WIDTH-1:0] wire_d86_25;
	wire [WIDTH-1:0] wire_d86_26;
	wire [WIDTH-1:0] wire_d86_27;
	wire [WIDTH-1:0] wire_d86_28;
	wire [WIDTH-1:0] wire_d86_29;
	wire [WIDTH-1:0] wire_d86_30;
	wire [WIDTH-1:0] wire_d86_31;
	wire [WIDTH-1:0] wire_d86_32;
	wire [WIDTH-1:0] wire_d86_33;
	wire [WIDTH-1:0] wire_d86_34;
	wire [WIDTH-1:0] wire_d86_35;
	wire [WIDTH-1:0] wire_d86_36;
	wire [WIDTH-1:0] wire_d86_37;
	wire [WIDTH-1:0] wire_d86_38;
	wire [WIDTH-1:0] wire_d86_39;
	wire [WIDTH-1:0] wire_d86_40;
	wire [WIDTH-1:0] wire_d86_41;
	wire [WIDTH-1:0] wire_d86_42;
	wire [WIDTH-1:0] wire_d86_43;
	wire [WIDTH-1:0] wire_d86_44;
	wire [WIDTH-1:0] wire_d86_45;
	wire [WIDTH-1:0] wire_d86_46;
	wire [WIDTH-1:0] wire_d86_47;
	wire [WIDTH-1:0] wire_d86_48;
	wire [WIDTH-1:0] wire_d86_49;
	wire [WIDTH-1:0] wire_d86_50;
	wire [WIDTH-1:0] wire_d86_51;
	wire [WIDTH-1:0] wire_d86_52;
	wire [WIDTH-1:0] wire_d86_53;
	wire [WIDTH-1:0] wire_d86_54;
	wire [WIDTH-1:0] wire_d86_55;
	wire [WIDTH-1:0] wire_d86_56;
	wire [WIDTH-1:0] wire_d86_57;
	wire [WIDTH-1:0] wire_d86_58;
	wire [WIDTH-1:0] wire_d86_59;
	wire [WIDTH-1:0] wire_d86_60;
	wire [WIDTH-1:0] wire_d86_61;
	wire [WIDTH-1:0] wire_d86_62;
	wire [WIDTH-1:0] wire_d86_63;
	wire [WIDTH-1:0] wire_d86_64;
	wire [WIDTH-1:0] wire_d86_65;
	wire [WIDTH-1:0] wire_d86_66;
	wire [WIDTH-1:0] wire_d86_67;
	wire [WIDTH-1:0] wire_d86_68;
	wire [WIDTH-1:0] wire_d86_69;
	wire [WIDTH-1:0] wire_d86_70;
	wire [WIDTH-1:0] wire_d86_71;
	wire [WIDTH-1:0] wire_d86_72;
	wire [WIDTH-1:0] wire_d86_73;
	wire [WIDTH-1:0] wire_d86_74;
	wire [WIDTH-1:0] wire_d86_75;
	wire [WIDTH-1:0] wire_d86_76;
	wire [WIDTH-1:0] wire_d86_77;
	wire [WIDTH-1:0] wire_d86_78;
	wire [WIDTH-1:0] wire_d86_79;
	wire [WIDTH-1:0] wire_d86_80;
	wire [WIDTH-1:0] wire_d86_81;
	wire [WIDTH-1:0] wire_d86_82;
	wire [WIDTH-1:0] wire_d86_83;
	wire [WIDTH-1:0] wire_d86_84;
	wire [WIDTH-1:0] wire_d86_85;
	wire [WIDTH-1:0] wire_d86_86;
	wire [WIDTH-1:0] wire_d86_87;
	wire [WIDTH-1:0] wire_d86_88;
	wire [WIDTH-1:0] wire_d86_89;
	wire [WIDTH-1:0] wire_d86_90;
	wire [WIDTH-1:0] wire_d86_91;
	wire [WIDTH-1:0] wire_d86_92;
	wire [WIDTH-1:0] wire_d86_93;
	wire [WIDTH-1:0] wire_d86_94;
	wire [WIDTH-1:0] wire_d86_95;
	wire [WIDTH-1:0] wire_d86_96;
	wire [WIDTH-1:0] wire_d86_97;
	wire [WIDTH-1:0] wire_d86_98;
	wire [WIDTH-1:0] wire_d86_99;
	wire [WIDTH-1:0] wire_d86_100;
	wire [WIDTH-1:0] wire_d86_101;
	wire [WIDTH-1:0] wire_d86_102;
	wire [WIDTH-1:0] wire_d86_103;
	wire [WIDTH-1:0] wire_d86_104;
	wire [WIDTH-1:0] wire_d86_105;
	wire [WIDTH-1:0] wire_d86_106;
	wire [WIDTH-1:0] wire_d86_107;
	wire [WIDTH-1:0] wire_d86_108;
	wire [WIDTH-1:0] wire_d86_109;
	wire [WIDTH-1:0] wire_d86_110;
	wire [WIDTH-1:0] wire_d86_111;
	wire [WIDTH-1:0] wire_d86_112;
	wire [WIDTH-1:0] wire_d86_113;
	wire [WIDTH-1:0] wire_d86_114;
	wire [WIDTH-1:0] wire_d86_115;
	wire [WIDTH-1:0] wire_d86_116;
	wire [WIDTH-1:0] wire_d86_117;
	wire [WIDTH-1:0] wire_d86_118;
	wire [WIDTH-1:0] wire_d87_0;
	wire [WIDTH-1:0] wire_d87_1;
	wire [WIDTH-1:0] wire_d87_2;
	wire [WIDTH-1:0] wire_d87_3;
	wire [WIDTH-1:0] wire_d87_4;
	wire [WIDTH-1:0] wire_d87_5;
	wire [WIDTH-1:0] wire_d87_6;
	wire [WIDTH-1:0] wire_d87_7;
	wire [WIDTH-1:0] wire_d87_8;
	wire [WIDTH-1:0] wire_d87_9;
	wire [WIDTH-1:0] wire_d87_10;
	wire [WIDTH-1:0] wire_d87_11;
	wire [WIDTH-1:0] wire_d87_12;
	wire [WIDTH-1:0] wire_d87_13;
	wire [WIDTH-1:0] wire_d87_14;
	wire [WIDTH-1:0] wire_d87_15;
	wire [WIDTH-1:0] wire_d87_16;
	wire [WIDTH-1:0] wire_d87_17;
	wire [WIDTH-1:0] wire_d87_18;
	wire [WIDTH-1:0] wire_d87_19;
	wire [WIDTH-1:0] wire_d87_20;
	wire [WIDTH-1:0] wire_d87_21;
	wire [WIDTH-1:0] wire_d87_22;
	wire [WIDTH-1:0] wire_d87_23;
	wire [WIDTH-1:0] wire_d87_24;
	wire [WIDTH-1:0] wire_d87_25;
	wire [WIDTH-1:0] wire_d87_26;
	wire [WIDTH-1:0] wire_d87_27;
	wire [WIDTH-1:0] wire_d87_28;
	wire [WIDTH-1:0] wire_d87_29;
	wire [WIDTH-1:0] wire_d87_30;
	wire [WIDTH-1:0] wire_d87_31;
	wire [WIDTH-1:0] wire_d87_32;
	wire [WIDTH-1:0] wire_d87_33;
	wire [WIDTH-1:0] wire_d87_34;
	wire [WIDTH-1:0] wire_d87_35;
	wire [WIDTH-1:0] wire_d87_36;
	wire [WIDTH-1:0] wire_d87_37;
	wire [WIDTH-1:0] wire_d87_38;
	wire [WIDTH-1:0] wire_d87_39;
	wire [WIDTH-1:0] wire_d87_40;
	wire [WIDTH-1:0] wire_d87_41;
	wire [WIDTH-1:0] wire_d87_42;
	wire [WIDTH-1:0] wire_d87_43;
	wire [WIDTH-1:0] wire_d87_44;
	wire [WIDTH-1:0] wire_d87_45;
	wire [WIDTH-1:0] wire_d87_46;
	wire [WIDTH-1:0] wire_d87_47;
	wire [WIDTH-1:0] wire_d87_48;
	wire [WIDTH-1:0] wire_d87_49;
	wire [WIDTH-1:0] wire_d87_50;
	wire [WIDTH-1:0] wire_d87_51;
	wire [WIDTH-1:0] wire_d87_52;
	wire [WIDTH-1:0] wire_d87_53;
	wire [WIDTH-1:0] wire_d87_54;
	wire [WIDTH-1:0] wire_d87_55;
	wire [WIDTH-1:0] wire_d87_56;
	wire [WIDTH-1:0] wire_d87_57;
	wire [WIDTH-1:0] wire_d87_58;
	wire [WIDTH-1:0] wire_d87_59;
	wire [WIDTH-1:0] wire_d87_60;
	wire [WIDTH-1:0] wire_d87_61;
	wire [WIDTH-1:0] wire_d87_62;
	wire [WIDTH-1:0] wire_d87_63;
	wire [WIDTH-1:0] wire_d87_64;
	wire [WIDTH-1:0] wire_d87_65;
	wire [WIDTH-1:0] wire_d87_66;
	wire [WIDTH-1:0] wire_d87_67;
	wire [WIDTH-1:0] wire_d87_68;
	wire [WIDTH-1:0] wire_d87_69;
	wire [WIDTH-1:0] wire_d87_70;
	wire [WIDTH-1:0] wire_d87_71;
	wire [WIDTH-1:0] wire_d87_72;
	wire [WIDTH-1:0] wire_d87_73;
	wire [WIDTH-1:0] wire_d87_74;
	wire [WIDTH-1:0] wire_d87_75;
	wire [WIDTH-1:0] wire_d87_76;
	wire [WIDTH-1:0] wire_d87_77;
	wire [WIDTH-1:0] wire_d87_78;
	wire [WIDTH-1:0] wire_d87_79;
	wire [WIDTH-1:0] wire_d87_80;
	wire [WIDTH-1:0] wire_d87_81;
	wire [WIDTH-1:0] wire_d87_82;
	wire [WIDTH-1:0] wire_d87_83;
	wire [WIDTH-1:0] wire_d87_84;
	wire [WIDTH-1:0] wire_d87_85;
	wire [WIDTH-1:0] wire_d87_86;
	wire [WIDTH-1:0] wire_d87_87;
	wire [WIDTH-1:0] wire_d87_88;
	wire [WIDTH-1:0] wire_d87_89;
	wire [WIDTH-1:0] wire_d87_90;
	wire [WIDTH-1:0] wire_d87_91;
	wire [WIDTH-1:0] wire_d87_92;
	wire [WIDTH-1:0] wire_d87_93;
	wire [WIDTH-1:0] wire_d87_94;
	wire [WIDTH-1:0] wire_d87_95;
	wire [WIDTH-1:0] wire_d87_96;
	wire [WIDTH-1:0] wire_d87_97;
	wire [WIDTH-1:0] wire_d87_98;
	wire [WIDTH-1:0] wire_d87_99;
	wire [WIDTH-1:0] wire_d87_100;
	wire [WIDTH-1:0] wire_d87_101;
	wire [WIDTH-1:0] wire_d87_102;
	wire [WIDTH-1:0] wire_d87_103;
	wire [WIDTH-1:0] wire_d87_104;
	wire [WIDTH-1:0] wire_d87_105;
	wire [WIDTH-1:0] wire_d87_106;
	wire [WIDTH-1:0] wire_d87_107;
	wire [WIDTH-1:0] wire_d87_108;
	wire [WIDTH-1:0] wire_d87_109;
	wire [WIDTH-1:0] wire_d87_110;
	wire [WIDTH-1:0] wire_d87_111;
	wire [WIDTH-1:0] wire_d87_112;
	wire [WIDTH-1:0] wire_d87_113;
	wire [WIDTH-1:0] wire_d87_114;
	wire [WIDTH-1:0] wire_d87_115;
	wire [WIDTH-1:0] wire_d87_116;
	wire [WIDTH-1:0] wire_d87_117;
	wire [WIDTH-1:0] wire_d87_118;
	wire [WIDTH-1:0] wire_d88_0;
	wire [WIDTH-1:0] wire_d88_1;
	wire [WIDTH-1:0] wire_d88_2;
	wire [WIDTH-1:0] wire_d88_3;
	wire [WIDTH-1:0] wire_d88_4;
	wire [WIDTH-1:0] wire_d88_5;
	wire [WIDTH-1:0] wire_d88_6;
	wire [WIDTH-1:0] wire_d88_7;
	wire [WIDTH-1:0] wire_d88_8;
	wire [WIDTH-1:0] wire_d88_9;
	wire [WIDTH-1:0] wire_d88_10;
	wire [WIDTH-1:0] wire_d88_11;
	wire [WIDTH-1:0] wire_d88_12;
	wire [WIDTH-1:0] wire_d88_13;
	wire [WIDTH-1:0] wire_d88_14;
	wire [WIDTH-1:0] wire_d88_15;
	wire [WIDTH-1:0] wire_d88_16;
	wire [WIDTH-1:0] wire_d88_17;
	wire [WIDTH-1:0] wire_d88_18;
	wire [WIDTH-1:0] wire_d88_19;
	wire [WIDTH-1:0] wire_d88_20;
	wire [WIDTH-1:0] wire_d88_21;
	wire [WIDTH-1:0] wire_d88_22;
	wire [WIDTH-1:0] wire_d88_23;
	wire [WIDTH-1:0] wire_d88_24;
	wire [WIDTH-1:0] wire_d88_25;
	wire [WIDTH-1:0] wire_d88_26;
	wire [WIDTH-1:0] wire_d88_27;
	wire [WIDTH-1:0] wire_d88_28;
	wire [WIDTH-1:0] wire_d88_29;
	wire [WIDTH-1:0] wire_d88_30;
	wire [WIDTH-1:0] wire_d88_31;
	wire [WIDTH-1:0] wire_d88_32;
	wire [WIDTH-1:0] wire_d88_33;
	wire [WIDTH-1:0] wire_d88_34;
	wire [WIDTH-1:0] wire_d88_35;
	wire [WIDTH-1:0] wire_d88_36;
	wire [WIDTH-1:0] wire_d88_37;
	wire [WIDTH-1:0] wire_d88_38;
	wire [WIDTH-1:0] wire_d88_39;
	wire [WIDTH-1:0] wire_d88_40;
	wire [WIDTH-1:0] wire_d88_41;
	wire [WIDTH-1:0] wire_d88_42;
	wire [WIDTH-1:0] wire_d88_43;
	wire [WIDTH-1:0] wire_d88_44;
	wire [WIDTH-1:0] wire_d88_45;
	wire [WIDTH-1:0] wire_d88_46;
	wire [WIDTH-1:0] wire_d88_47;
	wire [WIDTH-1:0] wire_d88_48;
	wire [WIDTH-1:0] wire_d88_49;
	wire [WIDTH-1:0] wire_d88_50;
	wire [WIDTH-1:0] wire_d88_51;
	wire [WIDTH-1:0] wire_d88_52;
	wire [WIDTH-1:0] wire_d88_53;
	wire [WIDTH-1:0] wire_d88_54;
	wire [WIDTH-1:0] wire_d88_55;
	wire [WIDTH-1:0] wire_d88_56;
	wire [WIDTH-1:0] wire_d88_57;
	wire [WIDTH-1:0] wire_d88_58;
	wire [WIDTH-1:0] wire_d88_59;
	wire [WIDTH-1:0] wire_d88_60;
	wire [WIDTH-1:0] wire_d88_61;
	wire [WIDTH-1:0] wire_d88_62;
	wire [WIDTH-1:0] wire_d88_63;
	wire [WIDTH-1:0] wire_d88_64;
	wire [WIDTH-1:0] wire_d88_65;
	wire [WIDTH-1:0] wire_d88_66;
	wire [WIDTH-1:0] wire_d88_67;
	wire [WIDTH-1:0] wire_d88_68;
	wire [WIDTH-1:0] wire_d88_69;
	wire [WIDTH-1:0] wire_d88_70;
	wire [WIDTH-1:0] wire_d88_71;
	wire [WIDTH-1:0] wire_d88_72;
	wire [WIDTH-1:0] wire_d88_73;
	wire [WIDTH-1:0] wire_d88_74;
	wire [WIDTH-1:0] wire_d88_75;
	wire [WIDTH-1:0] wire_d88_76;
	wire [WIDTH-1:0] wire_d88_77;
	wire [WIDTH-1:0] wire_d88_78;
	wire [WIDTH-1:0] wire_d88_79;
	wire [WIDTH-1:0] wire_d88_80;
	wire [WIDTH-1:0] wire_d88_81;
	wire [WIDTH-1:0] wire_d88_82;
	wire [WIDTH-1:0] wire_d88_83;
	wire [WIDTH-1:0] wire_d88_84;
	wire [WIDTH-1:0] wire_d88_85;
	wire [WIDTH-1:0] wire_d88_86;
	wire [WIDTH-1:0] wire_d88_87;
	wire [WIDTH-1:0] wire_d88_88;
	wire [WIDTH-1:0] wire_d88_89;
	wire [WIDTH-1:0] wire_d88_90;
	wire [WIDTH-1:0] wire_d88_91;
	wire [WIDTH-1:0] wire_d88_92;
	wire [WIDTH-1:0] wire_d88_93;
	wire [WIDTH-1:0] wire_d88_94;
	wire [WIDTH-1:0] wire_d88_95;
	wire [WIDTH-1:0] wire_d88_96;
	wire [WIDTH-1:0] wire_d88_97;
	wire [WIDTH-1:0] wire_d88_98;
	wire [WIDTH-1:0] wire_d88_99;
	wire [WIDTH-1:0] wire_d88_100;
	wire [WIDTH-1:0] wire_d88_101;
	wire [WIDTH-1:0] wire_d88_102;
	wire [WIDTH-1:0] wire_d88_103;
	wire [WIDTH-1:0] wire_d88_104;
	wire [WIDTH-1:0] wire_d88_105;
	wire [WIDTH-1:0] wire_d88_106;
	wire [WIDTH-1:0] wire_d88_107;
	wire [WIDTH-1:0] wire_d88_108;
	wire [WIDTH-1:0] wire_d88_109;
	wire [WIDTH-1:0] wire_d88_110;
	wire [WIDTH-1:0] wire_d88_111;
	wire [WIDTH-1:0] wire_d88_112;
	wire [WIDTH-1:0] wire_d88_113;
	wire [WIDTH-1:0] wire_d88_114;
	wire [WIDTH-1:0] wire_d88_115;
	wire [WIDTH-1:0] wire_d88_116;
	wire [WIDTH-1:0] wire_d88_117;
	wire [WIDTH-1:0] wire_d88_118;
	wire [WIDTH-1:0] wire_d89_0;
	wire [WIDTH-1:0] wire_d89_1;
	wire [WIDTH-1:0] wire_d89_2;
	wire [WIDTH-1:0] wire_d89_3;
	wire [WIDTH-1:0] wire_d89_4;
	wire [WIDTH-1:0] wire_d89_5;
	wire [WIDTH-1:0] wire_d89_6;
	wire [WIDTH-1:0] wire_d89_7;
	wire [WIDTH-1:0] wire_d89_8;
	wire [WIDTH-1:0] wire_d89_9;
	wire [WIDTH-1:0] wire_d89_10;
	wire [WIDTH-1:0] wire_d89_11;
	wire [WIDTH-1:0] wire_d89_12;
	wire [WIDTH-1:0] wire_d89_13;
	wire [WIDTH-1:0] wire_d89_14;
	wire [WIDTH-1:0] wire_d89_15;
	wire [WIDTH-1:0] wire_d89_16;
	wire [WIDTH-1:0] wire_d89_17;
	wire [WIDTH-1:0] wire_d89_18;
	wire [WIDTH-1:0] wire_d89_19;
	wire [WIDTH-1:0] wire_d89_20;
	wire [WIDTH-1:0] wire_d89_21;
	wire [WIDTH-1:0] wire_d89_22;
	wire [WIDTH-1:0] wire_d89_23;
	wire [WIDTH-1:0] wire_d89_24;
	wire [WIDTH-1:0] wire_d89_25;
	wire [WIDTH-1:0] wire_d89_26;
	wire [WIDTH-1:0] wire_d89_27;
	wire [WIDTH-1:0] wire_d89_28;
	wire [WIDTH-1:0] wire_d89_29;
	wire [WIDTH-1:0] wire_d89_30;
	wire [WIDTH-1:0] wire_d89_31;
	wire [WIDTH-1:0] wire_d89_32;
	wire [WIDTH-1:0] wire_d89_33;
	wire [WIDTH-1:0] wire_d89_34;
	wire [WIDTH-1:0] wire_d89_35;
	wire [WIDTH-1:0] wire_d89_36;
	wire [WIDTH-1:0] wire_d89_37;
	wire [WIDTH-1:0] wire_d89_38;
	wire [WIDTH-1:0] wire_d89_39;
	wire [WIDTH-1:0] wire_d89_40;
	wire [WIDTH-1:0] wire_d89_41;
	wire [WIDTH-1:0] wire_d89_42;
	wire [WIDTH-1:0] wire_d89_43;
	wire [WIDTH-1:0] wire_d89_44;
	wire [WIDTH-1:0] wire_d89_45;
	wire [WIDTH-1:0] wire_d89_46;
	wire [WIDTH-1:0] wire_d89_47;
	wire [WIDTH-1:0] wire_d89_48;
	wire [WIDTH-1:0] wire_d89_49;
	wire [WIDTH-1:0] wire_d89_50;
	wire [WIDTH-1:0] wire_d89_51;
	wire [WIDTH-1:0] wire_d89_52;
	wire [WIDTH-1:0] wire_d89_53;
	wire [WIDTH-1:0] wire_d89_54;
	wire [WIDTH-1:0] wire_d89_55;
	wire [WIDTH-1:0] wire_d89_56;
	wire [WIDTH-1:0] wire_d89_57;
	wire [WIDTH-1:0] wire_d89_58;
	wire [WIDTH-1:0] wire_d89_59;
	wire [WIDTH-1:0] wire_d89_60;
	wire [WIDTH-1:0] wire_d89_61;
	wire [WIDTH-1:0] wire_d89_62;
	wire [WIDTH-1:0] wire_d89_63;
	wire [WIDTH-1:0] wire_d89_64;
	wire [WIDTH-1:0] wire_d89_65;
	wire [WIDTH-1:0] wire_d89_66;
	wire [WIDTH-1:0] wire_d89_67;
	wire [WIDTH-1:0] wire_d89_68;
	wire [WIDTH-1:0] wire_d89_69;
	wire [WIDTH-1:0] wire_d89_70;
	wire [WIDTH-1:0] wire_d89_71;
	wire [WIDTH-1:0] wire_d89_72;
	wire [WIDTH-1:0] wire_d89_73;
	wire [WIDTH-1:0] wire_d89_74;
	wire [WIDTH-1:0] wire_d89_75;
	wire [WIDTH-1:0] wire_d89_76;
	wire [WIDTH-1:0] wire_d89_77;
	wire [WIDTH-1:0] wire_d89_78;
	wire [WIDTH-1:0] wire_d89_79;
	wire [WIDTH-1:0] wire_d89_80;
	wire [WIDTH-1:0] wire_d89_81;
	wire [WIDTH-1:0] wire_d89_82;
	wire [WIDTH-1:0] wire_d89_83;
	wire [WIDTH-1:0] wire_d89_84;
	wire [WIDTH-1:0] wire_d89_85;
	wire [WIDTH-1:0] wire_d89_86;
	wire [WIDTH-1:0] wire_d89_87;
	wire [WIDTH-1:0] wire_d89_88;
	wire [WIDTH-1:0] wire_d89_89;
	wire [WIDTH-1:0] wire_d89_90;
	wire [WIDTH-1:0] wire_d89_91;
	wire [WIDTH-1:0] wire_d89_92;
	wire [WIDTH-1:0] wire_d89_93;
	wire [WIDTH-1:0] wire_d89_94;
	wire [WIDTH-1:0] wire_d89_95;
	wire [WIDTH-1:0] wire_d89_96;
	wire [WIDTH-1:0] wire_d89_97;
	wire [WIDTH-1:0] wire_d89_98;
	wire [WIDTH-1:0] wire_d89_99;
	wire [WIDTH-1:0] wire_d89_100;
	wire [WIDTH-1:0] wire_d89_101;
	wire [WIDTH-1:0] wire_d89_102;
	wire [WIDTH-1:0] wire_d89_103;
	wire [WIDTH-1:0] wire_d89_104;
	wire [WIDTH-1:0] wire_d89_105;
	wire [WIDTH-1:0] wire_d89_106;
	wire [WIDTH-1:0] wire_d89_107;
	wire [WIDTH-1:0] wire_d89_108;
	wire [WIDTH-1:0] wire_d89_109;
	wire [WIDTH-1:0] wire_d89_110;
	wire [WIDTH-1:0] wire_d89_111;
	wire [WIDTH-1:0] wire_d89_112;
	wire [WIDTH-1:0] wire_d89_113;
	wire [WIDTH-1:0] wire_d89_114;
	wire [WIDTH-1:0] wire_d89_115;
	wire [WIDTH-1:0] wire_d89_116;
	wire [WIDTH-1:0] wire_d89_117;
	wire [WIDTH-1:0] wire_d89_118;
	wire [WIDTH-1:0] wire_d90_0;
	wire [WIDTH-1:0] wire_d90_1;
	wire [WIDTH-1:0] wire_d90_2;
	wire [WIDTH-1:0] wire_d90_3;
	wire [WIDTH-1:0] wire_d90_4;
	wire [WIDTH-1:0] wire_d90_5;
	wire [WIDTH-1:0] wire_d90_6;
	wire [WIDTH-1:0] wire_d90_7;
	wire [WIDTH-1:0] wire_d90_8;
	wire [WIDTH-1:0] wire_d90_9;
	wire [WIDTH-1:0] wire_d90_10;
	wire [WIDTH-1:0] wire_d90_11;
	wire [WIDTH-1:0] wire_d90_12;
	wire [WIDTH-1:0] wire_d90_13;
	wire [WIDTH-1:0] wire_d90_14;
	wire [WIDTH-1:0] wire_d90_15;
	wire [WIDTH-1:0] wire_d90_16;
	wire [WIDTH-1:0] wire_d90_17;
	wire [WIDTH-1:0] wire_d90_18;
	wire [WIDTH-1:0] wire_d90_19;
	wire [WIDTH-1:0] wire_d90_20;
	wire [WIDTH-1:0] wire_d90_21;
	wire [WIDTH-1:0] wire_d90_22;
	wire [WIDTH-1:0] wire_d90_23;
	wire [WIDTH-1:0] wire_d90_24;
	wire [WIDTH-1:0] wire_d90_25;
	wire [WIDTH-1:0] wire_d90_26;
	wire [WIDTH-1:0] wire_d90_27;
	wire [WIDTH-1:0] wire_d90_28;
	wire [WIDTH-1:0] wire_d90_29;
	wire [WIDTH-1:0] wire_d90_30;
	wire [WIDTH-1:0] wire_d90_31;
	wire [WIDTH-1:0] wire_d90_32;
	wire [WIDTH-1:0] wire_d90_33;
	wire [WIDTH-1:0] wire_d90_34;
	wire [WIDTH-1:0] wire_d90_35;
	wire [WIDTH-1:0] wire_d90_36;
	wire [WIDTH-1:0] wire_d90_37;
	wire [WIDTH-1:0] wire_d90_38;
	wire [WIDTH-1:0] wire_d90_39;
	wire [WIDTH-1:0] wire_d90_40;
	wire [WIDTH-1:0] wire_d90_41;
	wire [WIDTH-1:0] wire_d90_42;
	wire [WIDTH-1:0] wire_d90_43;
	wire [WIDTH-1:0] wire_d90_44;
	wire [WIDTH-1:0] wire_d90_45;
	wire [WIDTH-1:0] wire_d90_46;
	wire [WIDTH-1:0] wire_d90_47;
	wire [WIDTH-1:0] wire_d90_48;
	wire [WIDTH-1:0] wire_d90_49;
	wire [WIDTH-1:0] wire_d90_50;
	wire [WIDTH-1:0] wire_d90_51;
	wire [WIDTH-1:0] wire_d90_52;
	wire [WIDTH-1:0] wire_d90_53;
	wire [WIDTH-1:0] wire_d90_54;
	wire [WIDTH-1:0] wire_d90_55;
	wire [WIDTH-1:0] wire_d90_56;
	wire [WIDTH-1:0] wire_d90_57;
	wire [WIDTH-1:0] wire_d90_58;
	wire [WIDTH-1:0] wire_d90_59;
	wire [WIDTH-1:0] wire_d90_60;
	wire [WIDTH-1:0] wire_d90_61;
	wire [WIDTH-1:0] wire_d90_62;
	wire [WIDTH-1:0] wire_d90_63;
	wire [WIDTH-1:0] wire_d90_64;
	wire [WIDTH-1:0] wire_d90_65;
	wire [WIDTH-1:0] wire_d90_66;
	wire [WIDTH-1:0] wire_d90_67;
	wire [WIDTH-1:0] wire_d90_68;
	wire [WIDTH-1:0] wire_d90_69;
	wire [WIDTH-1:0] wire_d90_70;
	wire [WIDTH-1:0] wire_d90_71;
	wire [WIDTH-1:0] wire_d90_72;
	wire [WIDTH-1:0] wire_d90_73;
	wire [WIDTH-1:0] wire_d90_74;
	wire [WIDTH-1:0] wire_d90_75;
	wire [WIDTH-1:0] wire_d90_76;
	wire [WIDTH-1:0] wire_d90_77;
	wire [WIDTH-1:0] wire_d90_78;
	wire [WIDTH-1:0] wire_d90_79;
	wire [WIDTH-1:0] wire_d90_80;
	wire [WIDTH-1:0] wire_d90_81;
	wire [WIDTH-1:0] wire_d90_82;
	wire [WIDTH-1:0] wire_d90_83;
	wire [WIDTH-1:0] wire_d90_84;
	wire [WIDTH-1:0] wire_d90_85;
	wire [WIDTH-1:0] wire_d90_86;
	wire [WIDTH-1:0] wire_d90_87;
	wire [WIDTH-1:0] wire_d90_88;
	wire [WIDTH-1:0] wire_d90_89;
	wire [WIDTH-1:0] wire_d90_90;
	wire [WIDTH-1:0] wire_d90_91;
	wire [WIDTH-1:0] wire_d90_92;
	wire [WIDTH-1:0] wire_d90_93;
	wire [WIDTH-1:0] wire_d90_94;
	wire [WIDTH-1:0] wire_d90_95;
	wire [WIDTH-1:0] wire_d90_96;
	wire [WIDTH-1:0] wire_d90_97;
	wire [WIDTH-1:0] wire_d90_98;
	wire [WIDTH-1:0] wire_d90_99;
	wire [WIDTH-1:0] wire_d90_100;
	wire [WIDTH-1:0] wire_d90_101;
	wire [WIDTH-1:0] wire_d90_102;
	wire [WIDTH-1:0] wire_d90_103;
	wire [WIDTH-1:0] wire_d90_104;
	wire [WIDTH-1:0] wire_d90_105;
	wire [WIDTH-1:0] wire_d90_106;
	wire [WIDTH-1:0] wire_d90_107;
	wire [WIDTH-1:0] wire_d90_108;
	wire [WIDTH-1:0] wire_d90_109;
	wire [WIDTH-1:0] wire_d90_110;
	wire [WIDTH-1:0] wire_d90_111;
	wire [WIDTH-1:0] wire_d90_112;
	wire [WIDTH-1:0] wire_d90_113;
	wire [WIDTH-1:0] wire_d90_114;
	wire [WIDTH-1:0] wire_d90_115;
	wire [WIDTH-1:0] wire_d90_116;
	wire [WIDTH-1:0] wire_d90_117;
	wire [WIDTH-1:0] wire_d90_118;
	wire [WIDTH-1:0] wire_d91_0;
	wire [WIDTH-1:0] wire_d91_1;
	wire [WIDTH-1:0] wire_d91_2;
	wire [WIDTH-1:0] wire_d91_3;
	wire [WIDTH-1:0] wire_d91_4;
	wire [WIDTH-1:0] wire_d91_5;
	wire [WIDTH-1:0] wire_d91_6;
	wire [WIDTH-1:0] wire_d91_7;
	wire [WIDTH-1:0] wire_d91_8;
	wire [WIDTH-1:0] wire_d91_9;
	wire [WIDTH-1:0] wire_d91_10;
	wire [WIDTH-1:0] wire_d91_11;
	wire [WIDTH-1:0] wire_d91_12;
	wire [WIDTH-1:0] wire_d91_13;
	wire [WIDTH-1:0] wire_d91_14;
	wire [WIDTH-1:0] wire_d91_15;
	wire [WIDTH-1:0] wire_d91_16;
	wire [WIDTH-1:0] wire_d91_17;
	wire [WIDTH-1:0] wire_d91_18;
	wire [WIDTH-1:0] wire_d91_19;
	wire [WIDTH-1:0] wire_d91_20;
	wire [WIDTH-1:0] wire_d91_21;
	wire [WIDTH-1:0] wire_d91_22;
	wire [WIDTH-1:0] wire_d91_23;
	wire [WIDTH-1:0] wire_d91_24;
	wire [WIDTH-1:0] wire_d91_25;
	wire [WIDTH-1:0] wire_d91_26;
	wire [WIDTH-1:0] wire_d91_27;
	wire [WIDTH-1:0] wire_d91_28;
	wire [WIDTH-1:0] wire_d91_29;
	wire [WIDTH-1:0] wire_d91_30;
	wire [WIDTH-1:0] wire_d91_31;
	wire [WIDTH-1:0] wire_d91_32;
	wire [WIDTH-1:0] wire_d91_33;
	wire [WIDTH-1:0] wire_d91_34;
	wire [WIDTH-1:0] wire_d91_35;
	wire [WIDTH-1:0] wire_d91_36;
	wire [WIDTH-1:0] wire_d91_37;
	wire [WIDTH-1:0] wire_d91_38;
	wire [WIDTH-1:0] wire_d91_39;
	wire [WIDTH-1:0] wire_d91_40;
	wire [WIDTH-1:0] wire_d91_41;
	wire [WIDTH-1:0] wire_d91_42;
	wire [WIDTH-1:0] wire_d91_43;
	wire [WIDTH-1:0] wire_d91_44;
	wire [WIDTH-1:0] wire_d91_45;
	wire [WIDTH-1:0] wire_d91_46;
	wire [WIDTH-1:0] wire_d91_47;
	wire [WIDTH-1:0] wire_d91_48;
	wire [WIDTH-1:0] wire_d91_49;
	wire [WIDTH-1:0] wire_d91_50;
	wire [WIDTH-1:0] wire_d91_51;
	wire [WIDTH-1:0] wire_d91_52;
	wire [WIDTH-1:0] wire_d91_53;
	wire [WIDTH-1:0] wire_d91_54;
	wire [WIDTH-1:0] wire_d91_55;
	wire [WIDTH-1:0] wire_d91_56;
	wire [WIDTH-1:0] wire_d91_57;
	wire [WIDTH-1:0] wire_d91_58;
	wire [WIDTH-1:0] wire_d91_59;
	wire [WIDTH-1:0] wire_d91_60;
	wire [WIDTH-1:0] wire_d91_61;
	wire [WIDTH-1:0] wire_d91_62;
	wire [WIDTH-1:0] wire_d91_63;
	wire [WIDTH-1:0] wire_d91_64;
	wire [WIDTH-1:0] wire_d91_65;
	wire [WIDTH-1:0] wire_d91_66;
	wire [WIDTH-1:0] wire_d91_67;
	wire [WIDTH-1:0] wire_d91_68;
	wire [WIDTH-1:0] wire_d91_69;
	wire [WIDTH-1:0] wire_d91_70;
	wire [WIDTH-1:0] wire_d91_71;
	wire [WIDTH-1:0] wire_d91_72;
	wire [WIDTH-1:0] wire_d91_73;
	wire [WIDTH-1:0] wire_d91_74;
	wire [WIDTH-1:0] wire_d91_75;
	wire [WIDTH-1:0] wire_d91_76;
	wire [WIDTH-1:0] wire_d91_77;
	wire [WIDTH-1:0] wire_d91_78;
	wire [WIDTH-1:0] wire_d91_79;
	wire [WIDTH-1:0] wire_d91_80;
	wire [WIDTH-1:0] wire_d91_81;
	wire [WIDTH-1:0] wire_d91_82;
	wire [WIDTH-1:0] wire_d91_83;
	wire [WIDTH-1:0] wire_d91_84;
	wire [WIDTH-1:0] wire_d91_85;
	wire [WIDTH-1:0] wire_d91_86;
	wire [WIDTH-1:0] wire_d91_87;
	wire [WIDTH-1:0] wire_d91_88;
	wire [WIDTH-1:0] wire_d91_89;
	wire [WIDTH-1:0] wire_d91_90;
	wire [WIDTH-1:0] wire_d91_91;
	wire [WIDTH-1:0] wire_d91_92;
	wire [WIDTH-1:0] wire_d91_93;
	wire [WIDTH-1:0] wire_d91_94;
	wire [WIDTH-1:0] wire_d91_95;
	wire [WIDTH-1:0] wire_d91_96;
	wire [WIDTH-1:0] wire_d91_97;
	wire [WIDTH-1:0] wire_d91_98;
	wire [WIDTH-1:0] wire_d91_99;
	wire [WIDTH-1:0] wire_d91_100;
	wire [WIDTH-1:0] wire_d91_101;
	wire [WIDTH-1:0] wire_d91_102;
	wire [WIDTH-1:0] wire_d91_103;
	wire [WIDTH-1:0] wire_d91_104;
	wire [WIDTH-1:0] wire_d91_105;
	wire [WIDTH-1:0] wire_d91_106;
	wire [WIDTH-1:0] wire_d91_107;
	wire [WIDTH-1:0] wire_d91_108;
	wire [WIDTH-1:0] wire_d91_109;
	wire [WIDTH-1:0] wire_d91_110;
	wire [WIDTH-1:0] wire_d91_111;
	wire [WIDTH-1:0] wire_d91_112;
	wire [WIDTH-1:0] wire_d91_113;
	wire [WIDTH-1:0] wire_d91_114;
	wire [WIDTH-1:0] wire_d91_115;
	wire [WIDTH-1:0] wire_d91_116;
	wire [WIDTH-1:0] wire_d91_117;
	wire [WIDTH-1:0] wire_d91_118;
	wire [WIDTH-1:0] wire_d92_0;
	wire [WIDTH-1:0] wire_d92_1;
	wire [WIDTH-1:0] wire_d92_2;
	wire [WIDTH-1:0] wire_d92_3;
	wire [WIDTH-1:0] wire_d92_4;
	wire [WIDTH-1:0] wire_d92_5;
	wire [WIDTH-1:0] wire_d92_6;
	wire [WIDTH-1:0] wire_d92_7;
	wire [WIDTH-1:0] wire_d92_8;
	wire [WIDTH-1:0] wire_d92_9;
	wire [WIDTH-1:0] wire_d92_10;
	wire [WIDTH-1:0] wire_d92_11;
	wire [WIDTH-1:0] wire_d92_12;
	wire [WIDTH-1:0] wire_d92_13;
	wire [WIDTH-1:0] wire_d92_14;
	wire [WIDTH-1:0] wire_d92_15;
	wire [WIDTH-1:0] wire_d92_16;
	wire [WIDTH-1:0] wire_d92_17;
	wire [WIDTH-1:0] wire_d92_18;
	wire [WIDTH-1:0] wire_d92_19;
	wire [WIDTH-1:0] wire_d92_20;
	wire [WIDTH-1:0] wire_d92_21;
	wire [WIDTH-1:0] wire_d92_22;
	wire [WIDTH-1:0] wire_d92_23;
	wire [WIDTH-1:0] wire_d92_24;
	wire [WIDTH-1:0] wire_d92_25;
	wire [WIDTH-1:0] wire_d92_26;
	wire [WIDTH-1:0] wire_d92_27;
	wire [WIDTH-1:0] wire_d92_28;
	wire [WIDTH-1:0] wire_d92_29;
	wire [WIDTH-1:0] wire_d92_30;
	wire [WIDTH-1:0] wire_d92_31;
	wire [WIDTH-1:0] wire_d92_32;
	wire [WIDTH-1:0] wire_d92_33;
	wire [WIDTH-1:0] wire_d92_34;
	wire [WIDTH-1:0] wire_d92_35;
	wire [WIDTH-1:0] wire_d92_36;
	wire [WIDTH-1:0] wire_d92_37;
	wire [WIDTH-1:0] wire_d92_38;
	wire [WIDTH-1:0] wire_d92_39;
	wire [WIDTH-1:0] wire_d92_40;
	wire [WIDTH-1:0] wire_d92_41;
	wire [WIDTH-1:0] wire_d92_42;
	wire [WIDTH-1:0] wire_d92_43;
	wire [WIDTH-1:0] wire_d92_44;
	wire [WIDTH-1:0] wire_d92_45;
	wire [WIDTH-1:0] wire_d92_46;
	wire [WIDTH-1:0] wire_d92_47;
	wire [WIDTH-1:0] wire_d92_48;
	wire [WIDTH-1:0] wire_d92_49;
	wire [WIDTH-1:0] wire_d92_50;
	wire [WIDTH-1:0] wire_d92_51;
	wire [WIDTH-1:0] wire_d92_52;
	wire [WIDTH-1:0] wire_d92_53;
	wire [WIDTH-1:0] wire_d92_54;
	wire [WIDTH-1:0] wire_d92_55;
	wire [WIDTH-1:0] wire_d92_56;
	wire [WIDTH-1:0] wire_d92_57;
	wire [WIDTH-1:0] wire_d92_58;
	wire [WIDTH-1:0] wire_d92_59;
	wire [WIDTH-1:0] wire_d92_60;
	wire [WIDTH-1:0] wire_d92_61;
	wire [WIDTH-1:0] wire_d92_62;
	wire [WIDTH-1:0] wire_d92_63;
	wire [WIDTH-1:0] wire_d92_64;
	wire [WIDTH-1:0] wire_d92_65;
	wire [WIDTH-1:0] wire_d92_66;
	wire [WIDTH-1:0] wire_d92_67;
	wire [WIDTH-1:0] wire_d92_68;
	wire [WIDTH-1:0] wire_d92_69;
	wire [WIDTH-1:0] wire_d92_70;
	wire [WIDTH-1:0] wire_d92_71;
	wire [WIDTH-1:0] wire_d92_72;
	wire [WIDTH-1:0] wire_d92_73;
	wire [WIDTH-1:0] wire_d92_74;
	wire [WIDTH-1:0] wire_d92_75;
	wire [WIDTH-1:0] wire_d92_76;
	wire [WIDTH-1:0] wire_d92_77;
	wire [WIDTH-1:0] wire_d92_78;
	wire [WIDTH-1:0] wire_d92_79;
	wire [WIDTH-1:0] wire_d92_80;
	wire [WIDTH-1:0] wire_d92_81;
	wire [WIDTH-1:0] wire_d92_82;
	wire [WIDTH-1:0] wire_d92_83;
	wire [WIDTH-1:0] wire_d92_84;
	wire [WIDTH-1:0] wire_d92_85;
	wire [WIDTH-1:0] wire_d92_86;
	wire [WIDTH-1:0] wire_d92_87;
	wire [WIDTH-1:0] wire_d92_88;
	wire [WIDTH-1:0] wire_d92_89;
	wire [WIDTH-1:0] wire_d92_90;
	wire [WIDTH-1:0] wire_d92_91;
	wire [WIDTH-1:0] wire_d92_92;
	wire [WIDTH-1:0] wire_d92_93;
	wire [WIDTH-1:0] wire_d92_94;
	wire [WIDTH-1:0] wire_d92_95;
	wire [WIDTH-1:0] wire_d92_96;
	wire [WIDTH-1:0] wire_d92_97;
	wire [WIDTH-1:0] wire_d92_98;
	wire [WIDTH-1:0] wire_d92_99;
	wire [WIDTH-1:0] wire_d92_100;
	wire [WIDTH-1:0] wire_d92_101;
	wire [WIDTH-1:0] wire_d92_102;
	wire [WIDTH-1:0] wire_d92_103;
	wire [WIDTH-1:0] wire_d92_104;
	wire [WIDTH-1:0] wire_d92_105;
	wire [WIDTH-1:0] wire_d92_106;
	wire [WIDTH-1:0] wire_d92_107;
	wire [WIDTH-1:0] wire_d92_108;
	wire [WIDTH-1:0] wire_d92_109;
	wire [WIDTH-1:0] wire_d92_110;
	wire [WIDTH-1:0] wire_d92_111;
	wire [WIDTH-1:0] wire_d92_112;
	wire [WIDTH-1:0] wire_d92_113;
	wire [WIDTH-1:0] wire_d92_114;
	wire [WIDTH-1:0] wire_d92_115;
	wire [WIDTH-1:0] wire_d92_116;
	wire [WIDTH-1:0] wire_d92_117;
	wire [WIDTH-1:0] wire_d92_118;
	wire [WIDTH-1:0] wire_d93_0;
	wire [WIDTH-1:0] wire_d93_1;
	wire [WIDTH-1:0] wire_d93_2;
	wire [WIDTH-1:0] wire_d93_3;
	wire [WIDTH-1:0] wire_d93_4;
	wire [WIDTH-1:0] wire_d93_5;
	wire [WIDTH-1:0] wire_d93_6;
	wire [WIDTH-1:0] wire_d93_7;
	wire [WIDTH-1:0] wire_d93_8;
	wire [WIDTH-1:0] wire_d93_9;
	wire [WIDTH-1:0] wire_d93_10;
	wire [WIDTH-1:0] wire_d93_11;
	wire [WIDTH-1:0] wire_d93_12;
	wire [WIDTH-1:0] wire_d93_13;
	wire [WIDTH-1:0] wire_d93_14;
	wire [WIDTH-1:0] wire_d93_15;
	wire [WIDTH-1:0] wire_d93_16;
	wire [WIDTH-1:0] wire_d93_17;
	wire [WIDTH-1:0] wire_d93_18;
	wire [WIDTH-1:0] wire_d93_19;
	wire [WIDTH-1:0] wire_d93_20;
	wire [WIDTH-1:0] wire_d93_21;
	wire [WIDTH-1:0] wire_d93_22;
	wire [WIDTH-1:0] wire_d93_23;
	wire [WIDTH-1:0] wire_d93_24;
	wire [WIDTH-1:0] wire_d93_25;
	wire [WIDTH-1:0] wire_d93_26;
	wire [WIDTH-1:0] wire_d93_27;
	wire [WIDTH-1:0] wire_d93_28;
	wire [WIDTH-1:0] wire_d93_29;
	wire [WIDTH-1:0] wire_d93_30;
	wire [WIDTH-1:0] wire_d93_31;
	wire [WIDTH-1:0] wire_d93_32;
	wire [WIDTH-1:0] wire_d93_33;
	wire [WIDTH-1:0] wire_d93_34;
	wire [WIDTH-1:0] wire_d93_35;
	wire [WIDTH-1:0] wire_d93_36;
	wire [WIDTH-1:0] wire_d93_37;
	wire [WIDTH-1:0] wire_d93_38;
	wire [WIDTH-1:0] wire_d93_39;
	wire [WIDTH-1:0] wire_d93_40;
	wire [WIDTH-1:0] wire_d93_41;
	wire [WIDTH-1:0] wire_d93_42;
	wire [WIDTH-1:0] wire_d93_43;
	wire [WIDTH-1:0] wire_d93_44;
	wire [WIDTH-1:0] wire_d93_45;
	wire [WIDTH-1:0] wire_d93_46;
	wire [WIDTH-1:0] wire_d93_47;
	wire [WIDTH-1:0] wire_d93_48;
	wire [WIDTH-1:0] wire_d93_49;
	wire [WIDTH-1:0] wire_d93_50;
	wire [WIDTH-1:0] wire_d93_51;
	wire [WIDTH-1:0] wire_d93_52;
	wire [WIDTH-1:0] wire_d93_53;
	wire [WIDTH-1:0] wire_d93_54;
	wire [WIDTH-1:0] wire_d93_55;
	wire [WIDTH-1:0] wire_d93_56;
	wire [WIDTH-1:0] wire_d93_57;
	wire [WIDTH-1:0] wire_d93_58;
	wire [WIDTH-1:0] wire_d93_59;
	wire [WIDTH-1:0] wire_d93_60;
	wire [WIDTH-1:0] wire_d93_61;
	wire [WIDTH-1:0] wire_d93_62;
	wire [WIDTH-1:0] wire_d93_63;
	wire [WIDTH-1:0] wire_d93_64;
	wire [WIDTH-1:0] wire_d93_65;
	wire [WIDTH-1:0] wire_d93_66;
	wire [WIDTH-1:0] wire_d93_67;
	wire [WIDTH-1:0] wire_d93_68;
	wire [WIDTH-1:0] wire_d93_69;
	wire [WIDTH-1:0] wire_d93_70;
	wire [WIDTH-1:0] wire_d93_71;
	wire [WIDTH-1:0] wire_d93_72;
	wire [WIDTH-1:0] wire_d93_73;
	wire [WIDTH-1:0] wire_d93_74;
	wire [WIDTH-1:0] wire_d93_75;
	wire [WIDTH-1:0] wire_d93_76;
	wire [WIDTH-1:0] wire_d93_77;
	wire [WIDTH-1:0] wire_d93_78;
	wire [WIDTH-1:0] wire_d93_79;
	wire [WIDTH-1:0] wire_d93_80;
	wire [WIDTH-1:0] wire_d93_81;
	wire [WIDTH-1:0] wire_d93_82;
	wire [WIDTH-1:0] wire_d93_83;
	wire [WIDTH-1:0] wire_d93_84;
	wire [WIDTH-1:0] wire_d93_85;
	wire [WIDTH-1:0] wire_d93_86;
	wire [WIDTH-1:0] wire_d93_87;
	wire [WIDTH-1:0] wire_d93_88;
	wire [WIDTH-1:0] wire_d93_89;
	wire [WIDTH-1:0] wire_d93_90;
	wire [WIDTH-1:0] wire_d93_91;
	wire [WIDTH-1:0] wire_d93_92;
	wire [WIDTH-1:0] wire_d93_93;
	wire [WIDTH-1:0] wire_d93_94;
	wire [WIDTH-1:0] wire_d93_95;
	wire [WIDTH-1:0] wire_d93_96;
	wire [WIDTH-1:0] wire_d93_97;
	wire [WIDTH-1:0] wire_d93_98;
	wire [WIDTH-1:0] wire_d93_99;
	wire [WIDTH-1:0] wire_d93_100;
	wire [WIDTH-1:0] wire_d93_101;
	wire [WIDTH-1:0] wire_d93_102;
	wire [WIDTH-1:0] wire_d93_103;
	wire [WIDTH-1:0] wire_d93_104;
	wire [WIDTH-1:0] wire_d93_105;
	wire [WIDTH-1:0] wire_d93_106;
	wire [WIDTH-1:0] wire_d93_107;
	wire [WIDTH-1:0] wire_d93_108;
	wire [WIDTH-1:0] wire_d93_109;
	wire [WIDTH-1:0] wire_d93_110;
	wire [WIDTH-1:0] wire_d93_111;
	wire [WIDTH-1:0] wire_d93_112;
	wire [WIDTH-1:0] wire_d93_113;
	wire [WIDTH-1:0] wire_d93_114;
	wire [WIDTH-1:0] wire_d93_115;
	wire [WIDTH-1:0] wire_d93_116;
	wire [WIDTH-1:0] wire_d93_117;
	wire [WIDTH-1:0] wire_d93_118;
	wire [WIDTH-1:0] wire_d94_0;
	wire [WIDTH-1:0] wire_d94_1;
	wire [WIDTH-1:0] wire_d94_2;
	wire [WIDTH-1:0] wire_d94_3;
	wire [WIDTH-1:0] wire_d94_4;
	wire [WIDTH-1:0] wire_d94_5;
	wire [WIDTH-1:0] wire_d94_6;
	wire [WIDTH-1:0] wire_d94_7;
	wire [WIDTH-1:0] wire_d94_8;
	wire [WIDTH-1:0] wire_d94_9;
	wire [WIDTH-1:0] wire_d94_10;
	wire [WIDTH-1:0] wire_d94_11;
	wire [WIDTH-1:0] wire_d94_12;
	wire [WIDTH-1:0] wire_d94_13;
	wire [WIDTH-1:0] wire_d94_14;
	wire [WIDTH-1:0] wire_d94_15;
	wire [WIDTH-1:0] wire_d94_16;
	wire [WIDTH-1:0] wire_d94_17;
	wire [WIDTH-1:0] wire_d94_18;
	wire [WIDTH-1:0] wire_d94_19;
	wire [WIDTH-1:0] wire_d94_20;
	wire [WIDTH-1:0] wire_d94_21;
	wire [WIDTH-1:0] wire_d94_22;
	wire [WIDTH-1:0] wire_d94_23;
	wire [WIDTH-1:0] wire_d94_24;
	wire [WIDTH-1:0] wire_d94_25;
	wire [WIDTH-1:0] wire_d94_26;
	wire [WIDTH-1:0] wire_d94_27;
	wire [WIDTH-1:0] wire_d94_28;
	wire [WIDTH-1:0] wire_d94_29;
	wire [WIDTH-1:0] wire_d94_30;
	wire [WIDTH-1:0] wire_d94_31;
	wire [WIDTH-1:0] wire_d94_32;
	wire [WIDTH-1:0] wire_d94_33;
	wire [WIDTH-1:0] wire_d94_34;
	wire [WIDTH-1:0] wire_d94_35;
	wire [WIDTH-1:0] wire_d94_36;
	wire [WIDTH-1:0] wire_d94_37;
	wire [WIDTH-1:0] wire_d94_38;
	wire [WIDTH-1:0] wire_d94_39;
	wire [WIDTH-1:0] wire_d94_40;
	wire [WIDTH-1:0] wire_d94_41;
	wire [WIDTH-1:0] wire_d94_42;
	wire [WIDTH-1:0] wire_d94_43;
	wire [WIDTH-1:0] wire_d94_44;
	wire [WIDTH-1:0] wire_d94_45;
	wire [WIDTH-1:0] wire_d94_46;
	wire [WIDTH-1:0] wire_d94_47;
	wire [WIDTH-1:0] wire_d94_48;
	wire [WIDTH-1:0] wire_d94_49;
	wire [WIDTH-1:0] wire_d94_50;
	wire [WIDTH-1:0] wire_d94_51;
	wire [WIDTH-1:0] wire_d94_52;
	wire [WIDTH-1:0] wire_d94_53;
	wire [WIDTH-1:0] wire_d94_54;
	wire [WIDTH-1:0] wire_d94_55;
	wire [WIDTH-1:0] wire_d94_56;
	wire [WIDTH-1:0] wire_d94_57;
	wire [WIDTH-1:0] wire_d94_58;
	wire [WIDTH-1:0] wire_d94_59;
	wire [WIDTH-1:0] wire_d94_60;
	wire [WIDTH-1:0] wire_d94_61;
	wire [WIDTH-1:0] wire_d94_62;
	wire [WIDTH-1:0] wire_d94_63;
	wire [WIDTH-1:0] wire_d94_64;
	wire [WIDTH-1:0] wire_d94_65;
	wire [WIDTH-1:0] wire_d94_66;
	wire [WIDTH-1:0] wire_d94_67;
	wire [WIDTH-1:0] wire_d94_68;
	wire [WIDTH-1:0] wire_d94_69;
	wire [WIDTH-1:0] wire_d94_70;
	wire [WIDTH-1:0] wire_d94_71;
	wire [WIDTH-1:0] wire_d94_72;
	wire [WIDTH-1:0] wire_d94_73;
	wire [WIDTH-1:0] wire_d94_74;
	wire [WIDTH-1:0] wire_d94_75;
	wire [WIDTH-1:0] wire_d94_76;
	wire [WIDTH-1:0] wire_d94_77;
	wire [WIDTH-1:0] wire_d94_78;
	wire [WIDTH-1:0] wire_d94_79;
	wire [WIDTH-1:0] wire_d94_80;
	wire [WIDTH-1:0] wire_d94_81;
	wire [WIDTH-1:0] wire_d94_82;
	wire [WIDTH-1:0] wire_d94_83;
	wire [WIDTH-1:0] wire_d94_84;
	wire [WIDTH-1:0] wire_d94_85;
	wire [WIDTH-1:0] wire_d94_86;
	wire [WIDTH-1:0] wire_d94_87;
	wire [WIDTH-1:0] wire_d94_88;
	wire [WIDTH-1:0] wire_d94_89;
	wire [WIDTH-1:0] wire_d94_90;
	wire [WIDTH-1:0] wire_d94_91;
	wire [WIDTH-1:0] wire_d94_92;
	wire [WIDTH-1:0] wire_d94_93;
	wire [WIDTH-1:0] wire_d94_94;
	wire [WIDTH-1:0] wire_d94_95;
	wire [WIDTH-1:0] wire_d94_96;
	wire [WIDTH-1:0] wire_d94_97;
	wire [WIDTH-1:0] wire_d94_98;
	wire [WIDTH-1:0] wire_d94_99;
	wire [WIDTH-1:0] wire_d94_100;
	wire [WIDTH-1:0] wire_d94_101;
	wire [WIDTH-1:0] wire_d94_102;
	wire [WIDTH-1:0] wire_d94_103;
	wire [WIDTH-1:0] wire_d94_104;
	wire [WIDTH-1:0] wire_d94_105;
	wire [WIDTH-1:0] wire_d94_106;
	wire [WIDTH-1:0] wire_d94_107;
	wire [WIDTH-1:0] wire_d94_108;
	wire [WIDTH-1:0] wire_d94_109;
	wire [WIDTH-1:0] wire_d94_110;
	wire [WIDTH-1:0] wire_d94_111;
	wire [WIDTH-1:0] wire_d94_112;
	wire [WIDTH-1:0] wire_d94_113;
	wire [WIDTH-1:0] wire_d94_114;
	wire [WIDTH-1:0] wire_d94_115;
	wire [WIDTH-1:0] wire_d94_116;
	wire [WIDTH-1:0] wire_d94_117;
	wire [WIDTH-1:0] wire_d94_118;
	wire [WIDTH-1:0] wire_d95_0;
	wire [WIDTH-1:0] wire_d95_1;
	wire [WIDTH-1:0] wire_d95_2;
	wire [WIDTH-1:0] wire_d95_3;
	wire [WIDTH-1:0] wire_d95_4;
	wire [WIDTH-1:0] wire_d95_5;
	wire [WIDTH-1:0] wire_d95_6;
	wire [WIDTH-1:0] wire_d95_7;
	wire [WIDTH-1:0] wire_d95_8;
	wire [WIDTH-1:0] wire_d95_9;
	wire [WIDTH-1:0] wire_d95_10;
	wire [WIDTH-1:0] wire_d95_11;
	wire [WIDTH-1:0] wire_d95_12;
	wire [WIDTH-1:0] wire_d95_13;
	wire [WIDTH-1:0] wire_d95_14;
	wire [WIDTH-1:0] wire_d95_15;
	wire [WIDTH-1:0] wire_d95_16;
	wire [WIDTH-1:0] wire_d95_17;
	wire [WIDTH-1:0] wire_d95_18;
	wire [WIDTH-1:0] wire_d95_19;
	wire [WIDTH-1:0] wire_d95_20;
	wire [WIDTH-1:0] wire_d95_21;
	wire [WIDTH-1:0] wire_d95_22;
	wire [WIDTH-1:0] wire_d95_23;
	wire [WIDTH-1:0] wire_d95_24;
	wire [WIDTH-1:0] wire_d95_25;
	wire [WIDTH-1:0] wire_d95_26;
	wire [WIDTH-1:0] wire_d95_27;
	wire [WIDTH-1:0] wire_d95_28;
	wire [WIDTH-1:0] wire_d95_29;
	wire [WIDTH-1:0] wire_d95_30;
	wire [WIDTH-1:0] wire_d95_31;
	wire [WIDTH-1:0] wire_d95_32;
	wire [WIDTH-1:0] wire_d95_33;
	wire [WIDTH-1:0] wire_d95_34;
	wire [WIDTH-1:0] wire_d95_35;
	wire [WIDTH-1:0] wire_d95_36;
	wire [WIDTH-1:0] wire_d95_37;
	wire [WIDTH-1:0] wire_d95_38;
	wire [WIDTH-1:0] wire_d95_39;
	wire [WIDTH-1:0] wire_d95_40;
	wire [WIDTH-1:0] wire_d95_41;
	wire [WIDTH-1:0] wire_d95_42;
	wire [WIDTH-1:0] wire_d95_43;
	wire [WIDTH-1:0] wire_d95_44;
	wire [WIDTH-1:0] wire_d95_45;
	wire [WIDTH-1:0] wire_d95_46;
	wire [WIDTH-1:0] wire_d95_47;
	wire [WIDTH-1:0] wire_d95_48;
	wire [WIDTH-1:0] wire_d95_49;
	wire [WIDTH-1:0] wire_d95_50;
	wire [WIDTH-1:0] wire_d95_51;
	wire [WIDTH-1:0] wire_d95_52;
	wire [WIDTH-1:0] wire_d95_53;
	wire [WIDTH-1:0] wire_d95_54;
	wire [WIDTH-1:0] wire_d95_55;
	wire [WIDTH-1:0] wire_d95_56;
	wire [WIDTH-1:0] wire_d95_57;
	wire [WIDTH-1:0] wire_d95_58;
	wire [WIDTH-1:0] wire_d95_59;
	wire [WIDTH-1:0] wire_d95_60;
	wire [WIDTH-1:0] wire_d95_61;
	wire [WIDTH-1:0] wire_d95_62;
	wire [WIDTH-1:0] wire_d95_63;
	wire [WIDTH-1:0] wire_d95_64;
	wire [WIDTH-1:0] wire_d95_65;
	wire [WIDTH-1:0] wire_d95_66;
	wire [WIDTH-1:0] wire_d95_67;
	wire [WIDTH-1:0] wire_d95_68;
	wire [WIDTH-1:0] wire_d95_69;
	wire [WIDTH-1:0] wire_d95_70;
	wire [WIDTH-1:0] wire_d95_71;
	wire [WIDTH-1:0] wire_d95_72;
	wire [WIDTH-1:0] wire_d95_73;
	wire [WIDTH-1:0] wire_d95_74;
	wire [WIDTH-1:0] wire_d95_75;
	wire [WIDTH-1:0] wire_d95_76;
	wire [WIDTH-1:0] wire_d95_77;
	wire [WIDTH-1:0] wire_d95_78;
	wire [WIDTH-1:0] wire_d95_79;
	wire [WIDTH-1:0] wire_d95_80;
	wire [WIDTH-1:0] wire_d95_81;
	wire [WIDTH-1:0] wire_d95_82;
	wire [WIDTH-1:0] wire_d95_83;
	wire [WIDTH-1:0] wire_d95_84;
	wire [WIDTH-1:0] wire_d95_85;
	wire [WIDTH-1:0] wire_d95_86;
	wire [WIDTH-1:0] wire_d95_87;
	wire [WIDTH-1:0] wire_d95_88;
	wire [WIDTH-1:0] wire_d95_89;
	wire [WIDTH-1:0] wire_d95_90;
	wire [WIDTH-1:0] wire_d95_91;
	wire [WIDTH-1:0] wire_d95_92;
	wire [WIDTH-1:0] wire_d95_93;
	wire [WIDTH-1:0] wire_d95_94;
	wire [WIDTH-1:0] wire_d95_95;
	wire [WIDTH-1:0] wire_d95_96;
	wire [WIDTH-1:0] wire_d95_97;
	wire [WIDTH-1:0] wire_d95_98;
	wire [WIDTH-1:0] wire_d95_99;
	wire [WIDTH-1:0] wire_d95_100;
	wire [WIDTH-1:0] wire_d95_101;
	wire [WIDTH-1:0] wire_d95_102;
	wire [WIDTH-1:0] wire_d95_103;
	wire [WIDTH-1:0] wire_d95_104;
	wire [WIDTH-1:0] wire_d95_105;
	wire [WIDTH-1:0] wire_d95_106;
	wire [WIDTH-1:0] wire_d95_107;
	wire [WIDTH-1:0] wire_d95_108;
	wire [WIDTH-1:0] wire_d95_109;
	wire [WIDTH-1:0] wire_d95_110;
	wire [WIDTH-1:0] wire_d95_111;
	wire [WIDTH-1:0] wire_d95_112;
	wire [WIDTH-1:0] wire_d95_113;
	wire [WIDTH-1:0] wire_d95_114;
	wire [WIDTH-1:0] wire_d95_115;
	wire [WIDTH-1:0] wire_d95_116;
	wire [WIDTH-1:0] wire_d95_117;
	wire [WIDTH-1:0] wire_d95_118;
	wire [WIDTH-1:0] wire_d96_0;
	wire [WIDTH-1:0] wire_d96_1;
	wire [WIDTH-1:0] wire_d96_2;
	wire [WIDTH-1:0] wire_d96_3;
	wire [WIDTH-1:0] wire_d96_4;
	wire [WIDTH-1:0] wire_d96_5;
	wire [WIDTH-1:0] wire_d96_6;
	wire [WIDTH-1:0] wire_d96_7;
	wire [WIDTH-1:0] wire_d96_8;
	wire [WIDTH-1:0] wire_d96_9;
	wire [WIDTH-1:0] wire_d96_10;
	wire [WIDTH-1:0] wire_d96_11;
	wire [WIDTH-1:0] wire_d96_12;
	wire [WIDTH-1:0] wire_d96_13;
	wire [WIDTH-1:0] wire_d96_14;
	wire [WIDTH-1:0] wire_d96_15;
	wire [WIDTH-1:0] wire_d96_16;
	wire [WIDTH-1:0] wire_d96_17;
	wire [WIDTH-1:0] wire_d96_18;
	wire [WIDTH-1:0] wire_d96_19;
	wire [WIDTH-1:0] wire_d96_20;
	wire [WIDTH-1:0] wire_d96_21;
	wire [WIDTH-1:0] wire_d96_22;
	wire [WIDTH-1:0] wire_d96_23;
	wire [WIDTH-1:0] wire_d96_24;
	wire [WIDTH-1:0] wire_d96_25;
	wire [WIDTH-1:0] wire_d96_26;
	wire [WIDTH-1:0] wire_d96_27;
	wire [WIDTH-1:0] wire_d96_28;
	wire [WIDTH-1:0] wire_d96_29;
	wire [WIDTH-1:0] wire_d96_30;
	wire [WIDTH-1:0] wire_d96_31;
	wire [WIDTH-1:0] wire_d96_32;
	wire [WIDTH-1:0] wire_d96_33;
	wire [WIDTH-1:0] wire_d96_34;
	wire [WIDTH-1:0] wire_d96_35;
	wire [WIDTH-1:0] wire_d96_36;
	wire [WIDTH-1:0] wire_d96_37;
	wire [WIDTH-1:0] wire_d96_38;
	wire [WIDTH-1:0] wire_d96_39;
	wire [WIDTH-1:0] wire_d96_40;
	wire [WIDTH-1:0] wire_d96_41;
	wire [WIDTH-1:0] wire_d96_42;
	wire [WIDTH-1:0] wire_d96_43;
	wire [WIDTH-1:0] wire_d96_44;
	wire [WIDTH-1:0] wire_d96_45;
	wire [WIDTH-1:0] wire_d96_46;
	wire [WIDTH-1:0] wire_d96_47;
	wire [WIDTH-1:0] wire_d96_48;
	wire [WIDTH-1:0] wire_d96_49;
	wire [WIDTH-1:0] wire_d96_50;
	wire [WIDTH-1:0] wire_d96_51;
	wire [WIDTH-1:0] wire_d96_52;
	wire [WIDTH-1:0] wire_d96_53;
	wire [WIDTH-1:0] wire_d96_54;
	wire [WIDTH-1:0] wire_d96_55;
	wire [WIDTH-1:0] wire_d96_56;
	wire [WIDTH-1:0] wire_d96_57;
	wire [WIDTH-1:0] wire_d96_58;
	wire [WIDTH-1:0] wire_d96_59;
	wire [WIDTH-1:0] wire_d96_60;
	wire [WIDTH-1:0] wire_d96_61;
	wire [WIDTH-1:0] wire_d96_62;
	wire [WIDTH-1:0] wire_d96_63;
	wire [WIDTH-1:0] wire_d96_64;
	wire [WIDTH-1:0] wire_d96_65;
	wire [WIDTH-1:0] wire_d96_66;
	wire [WIDTH-1:0] wire_d96_67;
	wire [WIDTH-1:0] wire_d96_68;
	wire [WIDTH-1:0] wire_d96_69;
	wire [WIDTH-1:0] wire_d96_70;
	wire [WIDTH-1:0] wire_d96_71;
	wire [WIDTH-1:0] wire_d96_72;
	wire [WIDTH-1:0] wire_d96_73;
	wire [WIDTH-1:0] wire_d96_74;
	wire [WIDTH-1:0] wire_d96_75;
	wire [WIDTH-1:0] wire_d96_76;
	wire [WIDTH-1:0] wire_d96_77;
	wire [WIDTH-1:0] wire_d96_78;
	wire [WIDTH-1:0] wire_d96_79;
	wire [WIDTH-1:0] wire_d96_80;
	wire [WIDTH-1:0] wire_d96_81;
	wire [WIDTH-1:0] wire_d96_82;
	wire [WIDTH-1:0] wire_d96_83;
	wire [WIDTH-1:0] wire_d96_84;
	wire [WIDTH-1:0] wire_d96_85;
	wire [WIDTH-1:0] wire_d96_86;
	wire [WIDTH-1:0] wire_d96_87;
	wire [WIDTH-1:0] wire_d96_88;
	wire [WIDTH-1:0] wire_d96_89;
	wire [WIDTH-1:0] wire_d96_90;
	wire [WIDTH-1:0] wire_d96_91;
	wire [WIDTH-1:0] wire_d96_92;
	wire [WIDTH-1:0] wire_d96_93;
	wire [WIDTH-1:0] wire_d96_94;
	wire [WIDTH-1:0] wire_d96_95;
	wire [WIDTH-1:0] wire_d96_96;
	wire [WIDTH-1:0] wire_d96_97;
	wire [WIDTH-1:0] wire_d96_98;
	wire [WIDTH-1:0] wire_d96_99;
	wire [WIDTH-1:0] wire_d96_100;
	wire [WIDTH-1:0] wire_d96_101;
	wire [WIDTH-1:0] wire_d96_102;
	wire [WIDTH-1:0] wire_d96_103;
	wire [WIDTH-1:0] wire_d96_104;
	wire [WIDTH-1:0] wire_d96_105;
	wire [WIDTH-1:0] wire_d96_106;
	wire [WIDTH-1:0] wire_d96_107;
	wire [WIDTH-1:0] wire_d96_108;
	wire [WIDTH-1:0] wire_d96_109;
	wire [WIDTH-1:0] wire_d96_110;
	wire [WIDTH-1:0] wire_d96_111;
	wire [WIDTH-1:0] wire_d96_112;
	wire [WIDTH-1:0] wire_d96_113;
	wire [WIDTH-1:0] wire_d96_114;
	wire [WIDTH-1:0] wire_d96_115;
	wire [WIDTH-1:0] wire_d96_116;
	wire [WIDTH-1:0] wire_d96_117;
	wire [WIDTH-1:0] wire_d96_118;
	wire [WIDTH-1:0] wire_d97_0;
	wire [WIDTH-1:0] wire_d97_1;
	wire [WIDTH-1:0] wire_d97_2;
	wire [WIDTH-1:0] wire_d97_3;
	wire [WIDTH-1:0] wire_d97_4;
	wire [WIDTH-1:0] wire_d97_5;
	wire [WIDTH-1:0] wire_d97_6;
	wire [WIDTH-1:0] wire_d97_7;
	wire [WIDTH-1:0] wire_d97_8;
	wire [WIDTH-1:0] wire_d97_9;
	wire [WIDTH-1:0] wire_d97_10;
	wire [WIDTH-1:0] wire_d97_11;
	wire [WIDTH-1:0] wire_d97_12;
	wire [WIDTH-1:0] wire_d97_13;
	wire [WIDTH-1:0] wire_d97_14;
	wire [WIDTH-1:0] wire_d97_15;
	wire [WIDTH-1:0] wire_d97_16;
	wire [WIDTH-1:0] wire_d97_17;
	wire [WIDTH-1:0] wire_d97_18;
	wire [WIDTH-1:0] wire_d97_19;
	wire [WIDTH-1:0] wire_d97_20;
	wire [WIDTH-1:0] wire_d97_21;
	wire [WIDTH-1:0] wire_d97_22;
	wire [WIDTH-1:0] wire_d97_23;
	wire [WIDTH-1:0] wire_d97_24;
	wire [WIDTH-1:0] wire_d97_25;
	wire [WIDTH-1:0] wire_d97_26;
	wire [WIDTH-1:0] wire_d97_27;
	wire [WIDTH-1:0] wire_d97_28;
	wire [WIDTH-1:0] wire_d97_29;
	wire [WIDTH-1:0] wire_d97_30;
	wire [WIDTH-1:0] wire_d97_31;
	wire [WIDTH-1:0] wire_d97_32;
	wire [WIDTH-1:0] wire_d97_33;
	wire [WIDTH-1:0] wire_d97_34;
	wire [WIDTH-1:0] wire_d97_35;
	wire [WIDTH-1:0] wire_d97_36;
	wire [WIDTH-1:0] wire_d97_37;
	wire [WIDTH-1:0] wire_d97_38;
	wire [WIDTH-1:0] wire_d97_39;
	wire [WIDTH-1:0] wire_d97_40;
	wire [WIDTH-1:0] wire_d97_41;
	wire [WIDTH-1:0] wire_d97_42;
	wire [WIDTH-1:0] wire_d97_43;
	wire [WIDTH-1:0] wire_d97_44;
	wire [WIDTH-1:0] wire_d97_45;
	wire [WIDTH-1:0] wire_d97_46;
	wire [WIDTH-1:0] wire_d97_47;
	wire [WIDTH-1:0] wire_d97_48;
	wire [WIDTH-1:0] wire_d97_49;
	wire [WIDTH-1:0] wire_d97_50;
	wire [WIDTH-1:0] wire_d97_51;
	wire [WIDTH-1:0] wire_d97_52;
	wire [WIDTH-1:0] wire_d97_53;
	wire [WIDTH-1:0] wire_d97_54;
	wire [WIDTH-1:0] wire_d97_55;
	wire [WIDTH-1:0] wire_d97_56;
	wire [WIDTH-1:0] wire_d97_57;
	wire [WIDTH-1:0] wire_d97_58;
	wire [WIDTH-1:0] wire_d97_59;
	wire [WIDTH-1:0] wire_d97_60;
	wire [WIDTH-1:0] wire_d97_61;
	wire [WIDTH-1:0] wire_d97_62;
	wire [WIDTH-1:0] wire_d97_63;
	wire [WIDTH-1:0] wire_d97_64;
	wire [WIDTH-1:0] wire_d97_65;
	wire [WIDTH-1:0] wire_d97_66;
	wire [WIDTH-1:0] wire_d97_67;
	wire [WIDTH-1:0] wire_d97_68;
	wire [WIDTH-1:0] wire_d97_69;
	wire [WIDTH-1:0] wire_d97_70;
	wire [WIDTH-1:0] wire_d97_71;
	wire [WIDTH-1:0] wire_d97_72;
	wire [WIDTH-1:0] wire_d97_73;
	wire [WIDTH-1:0] wire_d97_74;
	wire [WIDTH-1:0] wire_d97_75;
	wire [WIDTH-1:0] wire_d97_76;
	wire [WIDTH-1:0] wire_d97_77;
	wire [WIDTH-1:0] wire_d97_78;
	wire [WIDTH-1:0] wire_d97_79;
	wire [WIDTH-1:0] wire_d97_80;
	wire [WIDTH-1:0] wire_d97_81;
	wire [WIDTH-1:0] wire_d97_82;
	wire [WIDTH-1:0] wire_d97_83;
	wire [WIDTH-1:0] wire_d97_84;
	wire [WIDTH-1:0] wire_d97_85;
	wire [WIDTH-1:0] wire_d97_86;
	wire [WIDTH-1:0] wire_d97_87;
	wire [WIDTH-1:0] wire_d97_88;
	wire [WIDTH-1:0] wire_d97_89;
	wire [WIDTH-1:0] wire_d97_90;
	wire [WIDTH-1:0] wire_d97_91;
	wire [WIDTH-1:0] wire_d97_92;
	wire [WIDTH-1:0] wire_d97_93;
	wire [WIDTH-1:0] wire_d97_94;
	wire [WIDTH-1:0] wire_d97_95;
	wire [WIDTH-1:0] wire_d97_96;
	wire [WIDTH-1:0] wire_d97_97;
	wire [WIDTH-1:0] wire_d97_98;
	wire [WIDTH-1:0] wire_d97_99;
	wire [WIDTH-1:0] wire_d97_100;
	wire [WIDTH-1:0] wire_d97_101;
	wire [WIDTH-1:0] wire_d97_102;
	wire [WIDTH-1:0] wire_d97_103;
	wire [WIDTH-1:0] wire_d97_104;
	wire [WIDTH-1:0] wire_d97_105;
	wire [WIDTH-1:0] wire_d97_106;
	wire [WIDTH-1:0] wire_d97_107;
	wire [WIDTH-1:0] wire_d97_108;
	wire [WIDTH-1:0] wire_d97_109;
	wire [WIDTH-1:0] wire_d97_110;
	wire [WIDTH-1:0] wire_d97_111;
	wire [WIDTH-1:0] wire_d97_112;
	wire [WIDTH-1:0] wire_d97_113;
	wire [WIDTH-1:0] wire_d97_114;
	wire [WIDTH-1:0] wire_d97_115;
	wire [WIDTH-1:0] wire_d97_116;
	wire [WIDTH-1:0] wire_d97_117;
	wire [WIDTH-1:0] wire_d97_118;
	wire [WIDTH-1:0] wire_d98_0;
	wire [WIDTH-1:0] wire_d98_1;
	wire [WIDTH-1:0] wire_d98_2;
	wire [WIDTH-1:0] wire_d98_3;
	wire [WIDTH-1:0] wire_d98_4;
	wire [WIDTH-1:0] wire_d98_5;
	wire [WIDTH-1:0] wire_d98_6;
	wire [WIDTH-1:0] wire_d98_7;
	wire [WIDTH-1:0] wire_d98_8;
	wire [WIDTH-1:0] wire_d98_9;
	wire [WIDTH-1:0] wire_d98_10;
	wire [WIDTH-1:0] wire_d98_11;
	wire [WIDTH-1:0] wire_d98_12;
	wire [WIDTH-1:0] wire_d98_13;
	wire [WIDTH-1:0] wire_d98_14;
	wire [WIDTH-1:0] wire_d98_15;
	wire [WIDTH-1:0] wire_d98_16;
	wire [WIDTH-1:0] wire_d98_17;
	wire [WIDTH-1:0] wire_d98_18;
	wire [WIDTH-1:0] wire_d98_19;
	wire [WIDTH-1:0] wire_d98_20;
	wire [WIDTH-1:0] wire_d98_21;
	wire [WIDTH-1:0] wire_d98_22;
	wire [WIDTH-1:0] wire_d98_23;
	wire [WIDTH-1:0] wire_d98_24;
	wire [WIDTH-1:0] wire_d98_25;
	wire [WIDTH-1:0] wire_d98_26;
	wire [WIDTH-1:0] wire_d98_27;
	wire [WIDTH-1:0] wire_d98_28;
	wire [WIDTH-1:0] wire_d98_29;
	wire [WIDTH-1:0] wire_d98_30;
	wire [WIDTH-1:0] wire_d98_31;
	wire [WIDTH-1:0] wire_d98_32;
	wire [WIDTH-1:0] wire_d98_33;
	wire [WIDTH-1:0] wire_d98_34;
	wire [WIDTH-1:0] wire_d98_35;
	wire [WIDTH-1:0] wire_d98_36;
	wire [WIDTH-1:0] wire_d98_37;
	wire [WIDTH-1:0] wire_d98_38;
	wire [WIDTH-1:0] wire_d98_39;
	wire [WIDTH-1:0] wire_d98_40;
	wire [WIDTH-1:0] wire_d98_41;
	wire [WIDTH-1:0] wire_d98_42;
	wire [WIDTH-1:0] wire_d98_43;
	wire [WIDTH-1:0] wire_d98_44;
	wire [WIDTH-1:0] wire_d98_45;
	wire [WIDTH-1:0] wire_d98_46;
	wire [WIDTH-1:0] wire_d98_47;
	wire [WIDTH-1:0] wire_d98_48;
	wire [WIDTH-1:0] wire_d98_49;
	wire [WIDTH-1:0] wire_d98_50;
	wire [WIDTH-1:0] wire_d98_51;
	wire [WIDTH-1:0] wire_d98_52;
	wire [WIDTH-1:0] wire_d98_53;
	wire [WIDTH-1:0] wire_d98_54;
	wire [WIDTH-1:0] wire_d98_55;
	wire [WIDTH-1:0] wire_d98_56;
	wire [WIDTH-1:0] wire_d98_57;
	wire [WIDTH-1:0] wire_d98_58;
	wire [WIDTH-1:0] wire_d98_59;
	wire [WIDTH-1:0] wire_d98_60;
	wire [WIDTH-1:0] wire_d98_61;
	wire [WIDTH-1:0] wire_d98_62;
	wire [WIDTH-1:0] wire_d98_63;
	wire [WIDTH-1:0] wire_d98_64;
	wire [WIDTH-1:0] wire_d98_65;
	wire [WIDTH-1:0] wire_d98_66;
	wire [WIDTH-1:0] wire_d98_67;
	wire [WIDTH-1:0] wire_d98_68;
	wire [WIDTH-1:0] wire_d98_69;
	wire [WIDTH-1:0] wire_d98_70;
	wire [WIDTH-1:0] wire_d98_71;
	wire [WIDTH-1:0] wire_d98_72;
	wire [WIDTH-1:0] wire_d98_73;
	wire [WIDTH-1:0] wire_d98_74;
	wire [WIDTH-1:0] wire_d98_75;
	wire [WIDTH-1:0] wire_d98_76;
	wire [WIDTH-1:0] wire_d98_77;
	wire [WIDTH-1:0] wire_d98_78;
	wire [WIDTH-1:0] wire_d98_79;
	wire [WIDTH-1:0] wire_d98_80;
	wire [WIDTH-1:0] wire_d98_81;
	wire [WIDTH-1:0] wire_d98_82;
	wire [WIDTH-1:0] wire_d98_83;
	wire [WIDTH-1:0] wire_d98_84;
	wire [WIDTH-1:0] wire_d98_85;
	wire [WIDTH-1:0] wire_d98_86;
	wire [WIDTH-1:0] wire_d98_87;
	wire [WIDTH-1:0] wire_d98_88;
	wire [WIDTH-1:0] wire_d98_89;
	wire [WIDTH-1:0] wire_d98_90;
	wire [WIDTH-1:0] wire_d98_91;
	wire [WIDTH-1:0] wire_d98_92;
	wire [WIDTH-1:0] wire_d98_93;
	wire [WIDTH-1:0] wire_d98_94;
	wire [WIDTH-1:0] wire_d98_95;
	wire [WIDTH-1:0] wire_d98_96;
	wire [WIDTH-1:0] wire_d98_97;
	wire [WIDTH-1:0] wire_d98_98;
	wire [WIDTH-1:0] wire_d98_99;
	wire [WIDTH-1:0] wire_d98_100;
	wire [WIDTH-1:0] wire_d98_101;
	wire [WIDTH-1:0] wire_d98_102;
	wire [WIDTH-1:0] wire_d98_103;
	wire [WIDTH-1:0] wire_d98_104;
	wire [WIDTH-1:0] wire_d98_105;
	wire [WIDTH-1:0] wire_d98_106;
	wire [WIDTH-1:0] wire_d98_107;
	wire [WIDTH-1:0] wire_d98_108;
	wire [WIDTH-1:0] wire_d98_109;
	wire [WIDTH-1:0] wire_d98_110;
	wire [WIDTH-1:0] wire_d98_111;
	wire [WIDTH-1:0] wire_d98_112;
	wire [WIDTH-1:0] wire_d98_113;
	wire [WIDTH-1:0] wire_d98_114;
	wire [WIDTH-1:0] wire_d98_115;
	wire [WIDTH-1:0] wire_d98_116;
	wire [WIDTH-1:0] wire_d98_117;
	wire [WIDTH-1:0] wire_d98_118;
	wire [WIDTH-1:0] wire_d99_0;
	wire [WIDTH-1:0] wire_d99_1;
	wire [WIDTH-1:0] wire_d99_2;
	wire [WIDTH-1:0] wire_d99_3;
	wire [WIDTH-1:0] wire_d99_4;
	wire [WIDTH-1:0] wire_d99_5;
	wire [WIDTH-1:0] wire_d99_6;
	wire [WIDTH-1:0] wire_d99_7;
	wire [WIDTH-1:0] wire_d99_8;
	wire [WIDTH-1:0] wire_d99_9;
	wire [WIDTH-1:0] wire_d99_10;
	wire [WIDTH-1:0] wire_d99_11;
	wire [WIDTH-1:0] wire_d99_12;
	wire [WIDTH-1:0] wire_d99_13;
	wire [WIDTH-1:0] wire_d99_14;
	wire [WIDTH-1:0] wire_d99_15;
	wire [WIDTH-1:0] wire_d99_16;
	wire [WIDTH-1:0] wire_d99_17;
	wire [WIDTH-1:0] wire_d99_18;
	wire [WIDTH-1:0] wire_d99_19;
	wire [WIDTH-1:0] wire_d99_20;
	wire [WIDTH-1:0] wire_d99_21;
	wire [WIDTH-1:0] wire_d99_22;
	wire [WIDTH-1:0] wire_d99_23;
	wire [WIDTH-1:0] wire_d99_24;
	wire [WIDTH-1:0] wire_d99_25;
	wire [WIDTH-1:0] wire_d99_26;
	wire [WIDTH-1:0] wire_d99_27;
	wire [WIDTH-1:0] wire_d99_28;
	wire [WIDTH-1:0] wire_d99_29;
	wire [WIDTH-1:0] wire_d99_30;
	wire [WIDTH-1:0] wire_d99_31;
	wire [WIDTH-1:0] wire_d99_32;
	wire [WIDTH-1:0] wire_d99_33;
	wire [WIDTH-1:0] wire_d99_34;
	wire [WIDTH-1:0] wire_d99_35;
	wire [WIDTH-1:0] wire_d99_36;
	wire [WIDTH-1:0] wire_d99_37;
	wire [WIDTH-1:0] wire_d99_38;
	wire [WIDTH-1:0] wire_d99_39;
	wire [WIDTH-1:0] wire_d99_40;
	wire [WIDTH-1:0] wire_d99_41;
	wire [WIDTH-1:0] wire_d99_42;
	wire [WIDTH-1:0] wire_d99_43;
	wire [WIDTH-1:0] wire_d99_44;
	wire [WIDTH-1:0] wire_d99_45;
	wire [WIDTH-1:0] wire_d99_46;
	wire [WIDTH-1:0] wire_d99_47;
	wire [WIDTH-1:0] wire_d99_48;
	wire [WIDTH-1:0] wire_d99_49;
	wire [WIDTH-1:0] wire_d99_50;
	wire [WIDTH-1:0] wire_d99_51;
	wire [WIDTH-1:0] wire_d99_52;
	wire [WIDTH-1:0] wire_d99_53;
	wire [WIDTH-1:0] wire_d99_54;
	wire [WIDTH-1:0] wire_d99_55;
	wire [WIDTH-1:0] wire_d99_56;
	wire [WIDTH-1:0] wire_d99_57;
	wire [WIDTH-1:0] wire_d99_58;
	wire [WIDTH-1:0] wire_d99_59;
	wire [WIDTH-1:0] wire_d99_60;
	wire [WIDTH-1:0] wire_d99_61;
	wire [WIDTH-1:0] wire_d99_62;
	wire [WIDTH-1:0] wire_d99_63;
	wire [WIDTH-1:0] wire_d99_64;
	wire [WIDTH-1:0] wire_d99_65;
	wire [WIDTH-1:0] wire_d99_66;
	wire [WIDTH-1:0] wire_d99_67;
	wire [WIDTH-1:0] wire_d99_68;
	wire [WIDTH-1:0] wire_d99_69;
	wire [WIDTH-1:0] wire_d99_70;
	wire [WIDTH-1:0] wire_d99_71;
	wire [WIDTH-1:0] wire_d99_72;
	wire [WIDTH-1:0] wire_d99_73;
	wire [WIDTH-1:0] wire_d99_74;
	wire [WIDTH-1:0] wire_d99_75;
	wire [WIDTH-1:0] wire_d99_76;
	wire [WIDTH-1:0] wire_d99_77;
	wire [WIDTH-1:0] wire_d99_78;
	wire [WIDTH-1:0] wire_d99_79;
	wire [WIDTH-1:0] wire_d99_80;
	wire [WIDTH-1:0] wire_d99_81;
	wire [WIDTH-1:0] wire_d99_82;
	wire [WIDTH-1:0] wire_d99_83;
	wire [WIDTH-1:0] wire_d99_84;
	wire [WIDTH-1:0] wire_d99_85;
	wire [WIDTH-1:0] wire_d99_86;
	wire [WIDTH-1:0] wire_d99_87;
	wire [WIDTH-1:0] wire_d99_88;
	wire [WIDTH-1:0] wire_d99_89;
	wire [WIDTH-1:0] wire_d99_90;
	wire [WIDTH-1:0] wire_d99_91;
	wire [WIDTH-1:0] wire_d99_92;
	wire [WIDTH-1:0] wire_d99_93;
	wire [WIDTH-1:0] wire_d99_94;
	wire [WIDTH-1:0] wire_d99_95;
	wire [WIDTH-1:0] wire_d99_96;
	wire [WIDTH-1:0] wire_d99_97;
	wire [WIDTH-1:0] wire_d99_98;
	wire [WIDTH-1:0] wire_d99_99;
	wire [WIDTH-1:0] wire_d99_100;
	wire [WIDTH-1:0] wire_d99_101;
	wire [WIDTH-1:0] wire_d99_102;
	wire [WIDTH-1:0] wire_d99_103;
	wire [WIDTH-1:0] wire_d99_104;
	wire [WIDTH-1:0] wire_d99_105;
	wire [WIDTH-1:0] wire_d99_106;
	wire [WIDTH-1:0] wire_d99_107;
	wire [WIDTH-1:0] wire_d99_108;
	wire [WIDTH-1:0] wire_d99_109;
	wire [WIDTH-1:0] wire_d99_110;
	wire [WIDTH-1:0] wire_d99_111;
	wire [WIDTH-1:0] wire_d99_112;
	wire [WIDTH-1:0] wire_d99_113;
	wire [WIDTH-1:0] wire_d99_114;
	wire [WIDTH-1:0] wire_d99_115;
	wire [WIDTH-1:0] wire_d99_116;
	wire [WIDTH-1:0] wire_d99_117;
	wire [WIDTH-1:0] wire_d99_118;

	invertion #(.WIDTH(WIDTH)) invertion_instance100(.data_in(d_in0),.data_out(wire_d0_0),.clk(clk),.rst(rst));            //channel 1
	register #(.WIDTH(WIDTH)) register_instance101(.data_in(wire_d0_0),.data_out(wire_d0_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance102(.data_in(wire_d0_1),.data_out(wire_d0_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance103(.data_in(wire_d0_2),.data_out(wire_d0_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance104(.data_in(wire_d0_3),.data_out(wire_d0_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance105(.data_in(wire_d0_4),.data_out(wire_d0_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance106(.data_in(wire_d0_5),.data_out(wire_d0_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance107(.data_in(wire_d0_6),.data_out(wire_d0_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance108(.data_in(wire_d0_7),.data_out(wire_d0_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance109(.data_in(wire_d0_8),.data_out(wire_d0_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1010(.data_in(wire_d0_9),.data_out(wire_d0_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1011(.data_in(wire_d0_10),.data_out(wire_d0_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1012(.data_in(wire_d0_11),.data_out(wire_d0_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1013(.data_in(wire_d0_12),.data_out(wire_d0_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1014(.data_in(wire_d0_13),.data_out(wire_d0_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1015(.data_in(wire_d0_14),.data_out(wire_d0_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1016(.data_in(wire_d0_15),.data_out(wire_d0_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1017(.data_in(wire_d0_16),.data_out(wire_d0_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1018(.data_in(wire_d0_17),.data_out(wire_d0_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1019(.data_in(wire_d0_18),.data_out(wire_d0_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1020(.data_in(wire_d0_19),.data_out(wire_d0_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1021(.data_in(wire_d0_20),.data_out(wire_d0_21),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1022(.data_in(wire_d0_21),.data_out(wire_d0_22),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1023(.data_in(wire_d0_22),.data_out(wire_d0_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1024(.data_in(wire_d0_23),.data_out(wire_d0_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1025(.data_in(wire_d0_24),.data_out(wire_d0_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1026(.data_in(wire_d0_25),.data_out(wire_d0_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1027(.data_in(wire_d0_26),.data_out(wire_d0_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1028(.data_in(wire_d0_27),.data_out(wire_d0_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1029(.data_in(wire_d0_28),.data_out(wire_d0_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1030(.data_in(wire_d0_29),.data_out(wire_d0_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1031(.data_in(wire_d0_30),.data_out(wire_d0_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1032(.data_in(wire_d0_31),.data_out(wire_d0_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1033(.data_in(wire_d0_32),.data_out(wire_d0_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1034(.data_in(wire_d0_33),.data_out(wire_d0_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1035(.data_in(wire_d0_34),.data_out(wire_d0_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1036(.data_in(wire_d0_35),.data_out(wire_d0_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1037(.data_in(wire_d0_36),.data_out(wire_d0_37),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1038(.data_in(wire_d0_37),.data_out(wire_d0_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1039(.data_in(wire_d0_38),.data_out(wire_d0_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1040(.data_in(wire_d0_39),.data_out(wire_d0_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1041(.data_in(wire_d0_40),.data_out(wire_d0_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1042(.data_in(wire_d0_41),.data_out(wire_d0_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1043(.data_in(wire_d0_42),.data_out(wire_d0_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1044(.data_in(wire_d0_43),.data_out(wire_d0_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1045(.data_in(wire_d0_44),.data_out(wire_d0_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1046(.data_in(wire_d0_45),.data_out(wire_d0_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1047(.data_in(wire_d0_46),.data_out(wire_d0_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1048(.data_in(wire_d0_47),.data_out(wire_d0_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1049(.data_in(wire_d0_48),.data_out(wire_d0_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1050(.data_in(wire_d0_49),.data_out(wire_d0_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1051(.data_in(wire_d0_50),.data_out(wire_d0_51),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1052(.data_in(wire_d0_51),.data_out(wire_d0_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1053(.data_in(wire_d0_52),.data_out(wire_d0_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1054(.data_in(wire_d0_53),.data_out(wire_d0_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1055(.data_in(wire_d0_54),.data_out(wire_d0_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1056(.data_in(wire_d0_55),.data_out(wire_d0_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1057(.data_in(wire_d0_56),.data_out(wire_d0_57),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1058(.data_in(wire_d0_57),.data_out(wire_d0_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1059(.data_in(wire_d0_58),.data_out(wire_d0_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1060(.data_in(wire_d0_59),.data_out(wire_d0_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1061(.data_in(wire_d0_60),.data_out(wire_d0_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1062(.data_in(wire_d0_61),.data_out(wire_d0_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1063(.data_in(wire_d0_62),.data_out(wire_d0_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1064(.data_in(wire_d0_63),.data_out(wire_d0_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1065(.data_in(wire_d0_64),.data_out(wire_d0_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1066(.data_in(wire_d0_65),.data_out(wire_d0_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1067(.data_in(wire_d0_66),.data_out(wire_d0_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1068(.data_in(wire_d0_67),.data_out(wire_d0_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1069(.data_in(wire_d0_68),.data_out(wire_d0_69),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1070(.data_in(wire_d0_69),.data_out(wire_d0_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1071(.data_in(wire_d0_70),.data_out(wire_d0_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1072(.data_in(wire_d0_71),.data_out(wire_d0_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1073(.data_in(wire_d0_72),.data_out(wire_d0_73),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1074(.data_in(wire_d0_73),.data_out(wire_d0_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1075(.data_in(wire_d0_74),.data_out(wire_d0_75),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1076(.data_in(wire_d0_75),.data_out(wire_d0_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1077(.data_in(wire_d0_76),.data_out(wire_d0_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1078(.data_in(wire_d0_77),.data_out(wire_d0_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1079(.data_in(wire_d0_78),.data_out(wire_d0_79),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1080(.data_in(wire_d0_79),.data_out(wire_d0_80),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1081(.data_in(wire_d0_80),.data_out(wire_d0_81),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1082(.data_in(wire_d0_81),.data_out(wire_d0_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1083(.data_in(wire_d0_82),.data_out(wire_d0_83),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1084(.data_in(wire_d0_83),.data_out(wire_d0_84),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1085(.data_in(wire_d0_84),.data_out(wire_d0_85),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1086(.data_in(wire_d0_85),.data_out(wire_d0_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1087(.data_in(wire_d0_86),.data_out(wire_d0_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1088(.data_in(wire_d0_87),.data_out(wire_d0_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1089(.data_in(wire_d0_88),.data_out(wire_d0_89),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1090(.data_in(wire_d0_89),.data_out(wire_d0_90),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1091(.data_in(wire_d0_90),.data_out(wire_d0_91),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1092(.data_in(wire_d0_91),.data_out(wire_d0_92),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1093(.data_in(wire_d0_92),.data_out(wire_d0_93),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1094(.data_in(wire_d0_93),.data_out(wire_d0_94),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1095(.data_in(wire_d0_94),.data_out(wire_d0_95),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1096(.data_in(wire_d0_95),.data_out(wire_d0_96),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1097(.data_in(wire_d0_96),.data_out(wire_d0_97),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1098(.data_in(wire_d0_97),.data_out(wire_d0_98),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1099(.data_in(wire_d0_98),.data_out(wire_d0_99),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance10100(.data_in(wire_d0_99),.data_out(wire_d0_100),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10101(.data_in(wire_d0_100),.data_out(wire_d0_101),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance10102(.data_in(wire_d0_101),.data_out(wire_d0_102),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10103(.data_in(wire_d0_102),.data_out(wire_d0_103),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance10104(.data_in(wire_d0_103),.data_out(wire_d0_104),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance10105(.data_in(wire_d0_104),.data_out(wire_d0_105),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance10106(.data_in(wire_d0_105),.data_out(wire_d0_106),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10107(.data_in(wire_d0_106),.data_out(wire_d0_107),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance10108(.data_in(wire_d0_107),.data_out(wire_d0_108),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance10109(.data_in(wire_d0_108),.data_out(wire_d0_109),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance10110(.data_in(wire_d0_109),.data_out(wire_d0_110),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance10111(.data_in(wire_d0_110),.data_out(wire_d0_111),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10112(.data_in(wire_d0_111),.data_out(wire_d0_112),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance10113(.data_in(wire_d0_112),.data_out(wire_d0_113),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10114(.data_in(wire_d0_113),.data_out(wire_d0_114),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance10115(.data_in(wire_d0_114),.data_out(wire_d0_115),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10116(.data_in(wire_d0_115),.data_out(wire_d0_116),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10117(.data_in(wire_d0_116),.data_out(wire_d0_117),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance10118(.data_in(wire_d0_117),.data_out(wire_d0_118),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance10119(.data_in(wire_d0_118),.data_out(d_out0),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance210(.data_in(d_in1),.data_out(wire_d1_0),.clk(clk),.rst(rst));            //channel 2
	register #(.WIDTH(WIDTH)) register_instance211(.data_in(wire_d1_0),.data_out(wire_d1_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212(.data_in(wire_d1_1),.data_out(wire_d1_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance213(.data_in(wire_d1_2),.data_out(wire_d1_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance214(.data_in(wire_d1_3),.data_out(wire_d1_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance215(.data_in(wire_d1_4),.data_out(wire_d1_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance216(.data_in(wire_d1_5),.data_out(wire_d1_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance217(.data_in(wire_d1_6),.data_out(wire_d1_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance218(.data_in(wire_d1_7),.data_out(wire_d1_8),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance219(.data_in(wire_d1_8),.data_out(wire_d1_9),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2110(.data_in(wire_d1_9),.data_out(wire_d1_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2111(.data_in(wire_d1_10),.data_out(wire_d1_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2112(.data_in(wire_d1_11),.data_out(wire_d1_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2113(.data_in(wire_d1_12),.data_out(wire_d1_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2114(.data_in(wire_d1_13),.data_out(wire_d1_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2115(.data_in(wire_d1_14),.data_out(wire_d1_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2116(.data_in(wire_d1_15),.data_out(wire_d1_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2117(.data_in(wire_d1_16),.data_out(wire_d1_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2118(.data_in(wire_d1_17),.data_out(wire_d1_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2119(.data_in(wire_d1_18),.data_out(wire_d1_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2120(.data_in(wire_d1_19),.data_out(wire_d1_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2121(.data_in(wire_d1_20),.data_out(wire_d1_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2122(.data_in(wire_d1_21),.data_out(wire_d1_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2123(.data_in(wire_d1_22),.data_out(wire_d1_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2124(.data_in(wire_d1_23),.data_out(wire_d1_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2125(.data_in(wire_d1_24),.data_out(wire_d1_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2126(.data_in(wire_d1_25),.data_out(wire_d1_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2127(.data_in(wire_d1_26),.data_out(wire_d1_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2128(.data_in(wire_d1_27),.data_out(wire_d1_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2129(.data_in(wire_d1_28),.data_out(wire_d1_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2130(.data_in(wire_d1_29),.data_out(wire_d1_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2131(.data_in(wire_d1_30),.data_out(wire_d1_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2132(.data_in(wire_d1_31),.data_out(wire_d1_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2133(.data_in(wire_d1_32),.data_out(wire_d1_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2134(.data_in(wire_d1_33),.data_out(wire_d1_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2135(.data_in(wire_d1_34),.data_out(wire_d1_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2136(.data_in(wire_d1_35),.data_out(wire_d1_36),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2137(.data_in(wire_d1_36),.data_out(wire_d1_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2138(.data_in(wire_d1_37),.data_out(wire_d1_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2139(.data_in(wire_d1_38),.data_out(wire_d1_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2140(.data_in(wire_d1_39),.data_out(wire_d1_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2141(.data_in(wire_d1_40),.data_out(wire_d1_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2142(.data_in(wire_d1_41),.data_out(wire_d1_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2143(.data_in(wire_d1_42),.data_out(wire_d1_43),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2144(.data_in(wire_d1_43),.data_out(wire_d1_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2145(.data_in(wire_d1_44),.data_out(wire_d1_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2146(.data_in(wire_d1_45),.data_out(wire_d1_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2147(.data_in(wire_d1_46),.data_out(wire_d1_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2148(.data_in(wire_d1_47),.data_out(wire_d1_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2149(.data_in(wire_d1_48),.data_out(wire_d1_49),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2150(.data_in(wire_d1_49),.data_out(wire_d1_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2151(.data_in(wire_d1_50),.data_out(wire_d1_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2152(.data_in(wire_d1_51),.data_out(wire_d1_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2153(.data_in(wire_d1_52),.data_out(wire_d1_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2154(.data_in(wire_d1_53),.data_out(wire_d1_54),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2155(.data_in(wire_d1_54),.data_out(wire_d1_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2156(.data_in(wire_d1_55),.data_out(wire_d1_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2157(.data_in(wire_d1_56),.data_out(wire_d1_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2158(.data_in(wire_d1_57),.data_out(wire_d1_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2159(.data_in(wire_d1_58),.data_out(wire_d1_59),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2160(.data_in(wire_d1_59),.data_out(wire_d1_60),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2161(.data_in(wire_d1_60),.data_out(wire_d1_61),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2162(.data_in(wire_d1_61),.data_out(wire_d1_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2163(.data_in(wire_d1_62),.data_out(wire_d1_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2164(.data_in(wire_d1_63),.data_out(wire_d1_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2165(.data_in(wire_d1_64),.data_out(wire_d1_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2166(.data_in(wire_d1_65),.data_out(wire_d1_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2167(.data_in(wire_d1_66),.data_out(wire_d1_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2168(.data_in(wire_d1_67),.data_out(wire_d1_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2169(.data_in(wire_d1_68),.data_out(wire_d1_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2170(.data_in(wire_d1_69),.data_out(wire_d1_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2171(.data_in(wire_d1_70),.data_out(wire_d1_71),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2172(.data_in(wire_d1_71),.data_out(wire_d1_72),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2173(.data_in(wire_d1_72),.data_out(wire_d1_73),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2174(.data_in(wire_d1_73),.data_out(wire_d1_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2175(.data_in(wire_d1_74),.data_out(wire_d1_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2176(.data_in(wire_d1_75),.data_out(wire_d1_76),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2177(.data_in(wire_d1_76),.data_out(wire_d1_77),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2178(.data_in(wire_d1_77),.data_out(wire_d1_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2179(.data_in(wire_d1_78),.data_out(wire_d1_79),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2180(.data_in(wire_d1_79),.data_out(wire_d1_80),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2181(.data_in(wire_d1_80),.data_out(wire_d1_81),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2182(.data_in(wire_d1_81),.data_out(wire_d1_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2183(.data_in(wire_d1_82),.data_out(wire_d1_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2184(.data_in(wire_d1_83),.data_out(wire_d1_84),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2185(.data_in(wire_d1_84),.data_out(wire_d1_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2186(.data_in(wire_d1_85),.data_out(wire_d1_86),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2187(.data_in(wire_d1_86),.data_out(wire_d1_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2188(.data_in(wire_d1_87),.data_out(wire_d1_88),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2189(.data_in(wire_d1_88),.data_out(wire_d1_89),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2190(.data_in(wire_d1_89),.data_out(wire_d1_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2191(.data_in(wire_d1_90),.data_out(wire_d1_91),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2192(.data_in(wire_d1_91),.data_out(wire_d1_92),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2193(.data_in(wire_d1_92),.data_out(wire_d1_93),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2194(.data_in(wire_d1_93),.data_out(wire_d1_94),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2195(.data_in(wire_d1_94),.data_out(wire_d1_95),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2196(.data_in(wire_d1_95),.data_out(wire_d1_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2197(.data_in(wire_d1_96),.data_out(wire_d1_97),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2198(.data_in(wire_d1_97),.data_out(wire_d1_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2199(.data_in(wire_d1_98),.data_out(wire_d1_99),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance21100(.data_in(wire_d1_99),.data_out(wire_d1_100),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance21101(.data_in(wire_d1_100),.data_out(wire_d1_101),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance21102(.data_in(wire_d1_101),.data_out(wire_d1_102),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance21103(.data_in(wire_d1_102),.data_out(wire_d1_103),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance21104(.data_in(wire_d1_103),.data_out(wire_d1_104),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance21105(.data_in(wire_d1_104),.data_out(wire_d1_105),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance21106(.data_in(wire_d1_105),.data_out(wire_d1_106),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance21107(.data_in(wire_d1_106),.data_out(wire_d1_107),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance21108(.data_in(wire_d1_107),.data_out(wire_d1_108),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance21109(.data_in(wire_d1_108),.data_out(wire_d1_109),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance21110(.data_in(wire_d1_109),.data_out(wire_d1_110),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance21111(.data_in(wire_d1_110),.data_out(wire_d1_111),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance21112(.data_in(wire_d1_111),.data_out(wire_d1_112),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance21113(.data_in(wire_d1_112),.data_out(wire_d1_113),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance21114(.data_in(wire_d1_113),.data_out(wire_d1_114),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21115(.data_in(wire_d1_114),.data_out(wire_d1_115),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance21116(.data_in(wire_d1_115),.data_out(wire_d1_116),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance21117(.data_in(wire_d1_116),.data_out(wire_d1_117),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance21118(.data_in(wire_d1_117),.data_out(wire_d1_118),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance21119(.data_in(wire_d1_118),.data_out(d_out1),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance320(.data_in(d_in2),.data_out(wire_d2_0),.clk(clk),.rst(rst));            //channel 3
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance321(.data_in(wire_d2_0),.data_out(wire_d2_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance322(.data_in(wire_d2_1),.data_out(wire_d2_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323(.data_in(wire_d2_2),.data_out(wire_d2_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance324(.data_in(wire_d2_3),.data_out(wire_d2_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance325(.data_in(wire_d2_4),.data_out(wire_d2_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance326(.data_in(wire_d2_5),.data_out(wire_d2_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance327(.data_in(wire_d2_6),.data_out(wire_d2_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance328(.data_in(wire_d2_7),.data_out(wire_d2_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance329(.data_in(wire_d2_8),.data_out(wire_d2_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3210(.data_in(wire_d2_9),.data_out(wire_d2_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3211(.data_in(wire_d2_10),.data_out(wire_d2_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3212(.data_in(wire_d2_11),.data_out(wire_d2_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3213(.data_in(wire_d2_12),.data_out(wire_d2_13),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3214(.data_in(wire_d2_13),.data_out(wire_d2_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3215(.data_in(wire_d2_14),.data_out(wire_d2_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3216(.data_in(wire_d2_15),.data_out(wire_d2_16),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3217(.data_in(wire_d2_16),.data_out(wire_d2_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3218(.data_in(wire_d2_17),.data_out(wire_d2_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3219(.data_in(wire_d2_18),.data_out(wire_d2_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3220(.data_in(wire_d2_19),.data_out(wire_d2_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3221(.data_in(wire_d2_20),.data_out(wire_d2_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3222(.data_in(wire_d2_21),.data_out(wire_d2_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3223(.data_in(wire_d2_22),.data_out(wire_d2_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3224(.data_in(wire_d2_23),.data_out(wire_d2_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3225(.data_in(wire_d2_24),.data_out(wire_d2_25),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3226(.data_in(wire_d2_25),.data_out(wire_d2_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3227(.data_in(wire_d2_26),.data_out(wire_d2_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3228(.data_in(wire_d2_27),.data_out(wire_d2_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3229(.data_in(wire_d2_28),.data_out(wire_d2_29),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3230(.data_in(wire_d2_29),.data_out(wire_d2_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3231(.data_in(wire_d2_30),.data_out(wire_d2_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3232(.data_in(wire_d2_31),.data_out(wire_d2_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3233(.data_in(wire_d2_32),.data_out(wire_d2_33),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3234(.data_in(wire_d2_33),.data_out(wire_d2_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3235(.data_in(wire_d2_34),.data_out(wire_d2_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3236(.data_in(wire_d2_35),.data_out(wire_d2_36),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3237(.data_in(wire_d2_36),.data_out(wire_d2_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3238(.data_in(wire_d2_37),.data_out(wire_d2_38),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3239(.data_in(wire_d2_38),.data_out(wire_d2_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3240(.data_in(wire_d2_39),.data_out(wire_d2_40),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3241(.data_in(wire_d2_40),.data_out(wire_d2_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3242(.data_in(wire_d2_41),.data_out(wire_d2_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3243(.data_in(wire_d2_42),.data_out(wire_d2_43),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3244(.data_in(wire_d2_43),.data_out(wire_d2_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3245(.data_in(wire_d2_44),.data_out(wire_d2_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3246(.data_in(wire_d2_45),.data_out(wire_d2_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3247(.data_in(wire_d2_46),.data_out(wire_d2_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3248(.data_in(wire_d2_47),.data_out(wire_d2_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3249(.data_in(wire_d2_48),.data_out(wire_d2_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3250(.data_in(wire_d2_49),.data_out(wire_d2_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3251(.data_in(wire_d2_50),.data_out(wire_d2_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3252(.data_in(wire_d2_51),.data_out(wire_d2_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3253(.data_in(wire_d2_52),.data_out(wire_d2_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3254(.data_in(wire_d2_53),.data_out(wire_d2_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3255(.data_in(wire_d2_54),.data_out(wire_d2_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3256(.data_in(wire_d2_55),.data_out(wire_d2_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3257(.data_in(wire_d2_56),.data_out(wire_d2_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3258(.data_in(wire_d2_57),.data_out(wire_d2_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3259(.data_in(wire_d2_58),.data_out(wire_d2_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3260(.data_in(wire_d2_59),.data_out(wire_d2_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3261(.data_in(wire_d2_60),.data_out(wire_d2_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3262(.data_in(wire_d2_61),.data_out(wire_d2_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3263(.data_in(wire_d2_62),.data_out(wire_d2_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3264(.data_in(wire_d2_63),.data_out(wire_d2_64),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3265(.data_in(wire_d2_64),.data_out(wire_d2_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3266(.data_in(wire_d2_65),.data_out(wire_d2_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3267(.data_in(wire_d2_66),.data_out(wire_d2_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3268(.data_in(wire_d2_67),.data_out(wire_d2_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3269(.data_in(wire_d2_68),.data_out(wire_d2_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3270(.data_in(wire_d2_69),.data_out(wire_d2_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3271(.data_in(wire_d2_70),.data_out(wire_d2_71),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3272(.data_in(wire_d2_71),.data_out(wire_d2_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3273(.data_in(wire_d2_72),.data_out(wire_d2_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3274(.data_in(wire_d2_73),.data_out(wire_d2_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3275(.data_in(wire_d2_74),.data_out(wire_d2_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3276(.data_in(wire_d2_75),.data_out(wire_d2_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3277(.data_in(wire_d2_76),.data_out(wire_d2_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3278(.data_in(wire_d2_77),.data_out(wire_d2_78),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3279(.data_in(wire_d2_78),.data_out(wire_d2_79),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3280(.data_in(wire_d2_79),.data_out(wire_d2_80),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3281(.data_in(wire_d2_80),.data_out(wire_d2_81),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3282(.data_in(wire_d2_81),.data_out(wire_d2_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3283(.data_in(wire_d2_82),.data_out(wire_d2_83),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3284(.data_in(wire_d2_83),.data_out(wire_d2_84),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3285(.data_in(wire_d2_84),.data_out(wire_d2_85),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3286(.data_in(wire_d2_85),.data_out(wire_d2_86),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3287(.data_in(wire_d2_86),.data_out(wire_d2_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3288(.data_in(wire_d2_87),.data_out(wire_d2_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3289(.data_in(wire_d2_88),.data_out(wire_d2_89),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3290(.data_in(wire_d2_89),.data_out(wire_d2_90),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3291(.data_in(wire_d2_90),.data_out(wire_d2_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3292(.data_in(wire_d2_91),.data_out(wire_d2_92),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3293(.data_in(wire_d2_92),.data_out(wire_d2_93),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3294(.data_in(wire_d2_93),.data_out(wire_d2_94),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3295(.data_in(wire_d2_94),.data_out(wire_d2_95),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3296(.data_in(wire_d2_95),.data_out(wire_d2_96),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3297(.data_in(wire_d2_96),.data_out(wire_d2_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3298(.data_in(wire_d2_97),.data_out(wire_d2_98),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3299(.data_in(wire_d2_98),.data_out(wire_d2_99),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance32100(.data_in(wire_d2_99),.data_out(wire_d2_100),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance32101(.data_in(wire_d2_100),.data_out(wire_d2_101),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance32102(.data_in(wire_d2_101),.data_out(wire_d2_102),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance32103(.data_in(wire_d2_102),.data_out(wire_d2_103),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance32104(.data_in(wire_d2_103),.data_out(wire_d2_104),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance32105(.data_in(wire_d2_104),.data_out(wire_d2_105),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance32106(.data_in(wire_d2_105),.data_out(wire_d2_106),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance32107(.data_in(wire_d2_106),.data_out(wire_d2_107),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance32108(.data_in(wire_d2_107),.data_out(wire_d2_108),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance32109(.data_in(wire_d2_108),.data_out(wire_d2_109),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance32110(.data_in(wire_d2_109),.data_out(wire_d2_110),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance32111(.data_in(wire_d2_110),.data_out(wire_d2_111),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance32112(.data_in(wire_d2_111),.data_out(wire_d2_112),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance32113(.data_in(wire_d2_112),.data_out(wire_d2_113),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance32114(.data_in(wire_d2_113),.data_out(wire_d2_114),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance32115(.data_in(wire_d2_114),.data_out(wire_d2_115),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance32116(.data_in(wire_d2_115),.data_out(wire_d2_116),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance32117(.data_in(wire_d2_116),.data_out(wire_d2_117),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance32118(.data_in(wire_d2_117),.data_out(wire_d2_118),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance32119(.data_in(wire_d2_118),.data_out(d_out2),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance430(.data_in(d_in3),.data_out(wire_d3_0),.clk(clk),.rst(rst));            //channel 4
	encoder #(.WIDTH(WIDTH)) encoder_instance431(.data_in(wire_d3_0),.data_out(wire_d3_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance432(.data_in(wire_d3_1),.data_out(wire_d3_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance433(.data_in(wire_d3_2),.data_out(wire_d3_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance434(.data_in(wire_d3_3),.data_out(wire_d3_4),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance435(.data_in(wire_d3_4),.data_out(wire_d3_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance436(.data_in(wire_d3_5),.data_out(wire_d3_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance437(.data_in(wire_d3_6),.data_out(wire_d3_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance438(.data_in(wire_d3_7),.data_out(wire_d3_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance439(.data_in(wire_d3_8),.data_out(wire_d3_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4310(.data_in(wire_d3_9),.data_out(wire_d3_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4311(.data_in(wire_d3_10),.data_out(wire_d3_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4312(.data_in(wire_d3_11),.data_out(wire_d3_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4313(.data_in(wire_d3_12),.data_out(wire_d3_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4314(.data_in(wire_d3_13),.data_out(wire_d3_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4315(.data_in(wire_d3_14),.data_out(wire_d3_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4316(.data_in(wire_d3_15),.data_out(wire_d3_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4317(.data_in(wire_d3_16),.data_out(wire_d3_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4318(.data_in(wire_d3_17),.data_out(wire_d3_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4319(.data_in(wire_d3_18),.data_out(wire_d3_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4320(.data_in(wire_d3_19),.data_out(wire_d3_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4321(.data_in(wire_d3_20),.data_out(wire_d3_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4322(.data_in(wire_d3_21),.data_out(wire_d3_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4323(.data_in(wire_d3_22),.data_out(wire_d3_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4324(.data_in(wire_d3_23),.data_out(wire_d3_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4325(.data_in(wire_d3_24),.data_out(wire_d3_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4326(.data_in(wire_d3_25),.data_out(wire_d3_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4327(.data_in(wire_d3_26),.data_out(wire_d3_27),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4328(.data_in(wire_d3_27),.data_out(wire_d3_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4329(.data_in(wire_d3_28),.data_out(wire_d3_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4330(.data_in(wire_d3_29),.data_out(wire_d3_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4331(.data_in(wire_d3_30),.data_out(wire_d3_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4332(.data_in(wire_d3_31),.data_out(wire_d3_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4333(.data_in(wire_d3_32),.data_out(wire_d3_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4334(.data_in(wire_d3_33),.data_out(wire_d3_34),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4335(.data_in(wire_d3_34),.data_out(wire_d3_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4336(.data_in(wire_d3_35),.data_out(wire_d3_36),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4337(.data_in(wire_d3_36),.data_out(wire_d3_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4338(.data_in(wire_d3_37),.data_out(wire_d3_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4339(.data_in(wire_d3_38),.data_out(wire_d3_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4340(.data_in(wire_d3_39),.data_out(wire_d3_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4341(.data_in(wire_d3_40),.data_out(wire_d3_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4342(.data_in(wire_d3_41),.data_out(wire_d3_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4343(.data_in(wire_d3_42),.data_out(wire_d3_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4344(.data_in(wire_d3_43),.data_out(wire_d3_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4345(.data_in(wire_d3_44),.data_out(wire_d3_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4346(.data_in(wire_d3_45),.data_out(wire_d3_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4347(.data_in(wire_d3_46),.data_out(wire_d3_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4348(.data_in(wire_d3_47),.data_out(wire_d3_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4349(.data_in(wire_d3_48),.data_out(wire_d3_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4350(.data_in(wire_d3_49),.data_out(wire_d3_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4351(.data_in(wire_d3_50),.data_out(wire_d3_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4352(.data_in(wire_d3_51),.data_out(wire_d3_52),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4353(.data_in(wire_d3_52),.data_out(wire_d3_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4354(.data_in(wire_d3_53),.data_out(wire_d3_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4355(.data_in(wire_d3_54),.data_out(wire_d3_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4356(.data_in(wire_d3_55),.data_out(wire_d3_56),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4357(.data_in(wire_d3_56),.data_out(wire_d3_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4358(.data_in(wire_d3_57),.data_out(wire_d3_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4359(.data_in(wire_d3_58),.data_out(wire_d3_59),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4360(.data_in(wire_d3_59),.data_out(wire_d3_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4361(.data_in(wire_d3_60),.data_out(wire_d3_61),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4362(.data_in(wire_d3_61),.data_out(wire_d3_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4363(.data_in(wire_d3_62),.data_out(wire_d3_63),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4364(.data_in(wire_d3_63),.data_out(wire_d3_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4365(.data_in(wire_d3_64),.data_out(wire_d3_65),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4366(.data_in(wire_d3_65),.data_out(wire_d3_66),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4367(.data_in(wire_d3_66),.data_out(wire_d3_67),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4368(.data_in(wire_d3_67),.data_out(wire_d3_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4369(.data_in(wire_d3_68),.data_out(wire_d3_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4370(.data_in(wire_d3_69),.data_out(wire_d3_70),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4371(.data_in(wire_d3_70),.data_out(wire_d3_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4372(.data_in(wire_d3_71),.data_out(wire_d3_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4373(.data_in(wire_d3_72),.data_out(wire_d3_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4374(.data_in(wire_d3_73),.data_out(wire_d3_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4375(.data_in(wire_d3_74),.data_out(wire_d3_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4376(.data_in(wire_d3_75),.data_out(wire_d3_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4377(.data_in(wire_d3_76),.data_out(wire_d3_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4378(.data_in(wire_d3_77),.data_out(wire_d3_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4379(.data_in(wire_d3_78),.data_out(wire_d3_79),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4380(.data_in(wire_d3_79),.data_out(wire_d3_80),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4381(.data_in(wire_d3_80),.data_out(wire_d3_81),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4382(.data_in(wire_d3_81),.data_out(wire_d3_82),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4383(.data_in(wire_d3_82),.data_out(wire_d3_83),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4384(.data_in(wire_d3_83),.data_out(wire_d3_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4385(.data_in(wire_d3_84),.data_out(wire_d3_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4386(.data_in(wire_d3_85),.data_out(wire_d3_86),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4387(.data_in(wire_d3_86),.data_out(wire_d3_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4388(.data_in(wire_d3_87),.data_out(wire_d3_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4389(.data_in(wire_d3_88),.data_out(wire_d3_89),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4390(.data_in(wire_d3_89),.data_out(wire_d3_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4391(.data_in(wire_d3_90),.data_out(wire_d3_91),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4392(.data_in(wire_d3_91),.data_out(wire_d3_92),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4393(.data_in(wire_d3_92),.data_out(wire_d3_93),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4394(.data_in(wire_d3_93),.data_out(wire_d3_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4395(.data_in(wire_d3_94),.data_out(wire_d3_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4396(.data_in(wire_d3_95),.data_out(wire_d3_96),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4397(.data_in(wire_d3_96),.data_out(wire_d3_97),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4398(.data_in(wire_d3_97),.data_out(wire_d3_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4399(.data_in(wire_d3_98),.data_out(wire_d3_99),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance43100(.data_in(wire_d3_99),.data_out(wire_d3_100),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance43101(.data_in(wire_d3_100),.data_out(wire_d3_101),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance43102(.data_in(wire_d3_101),.data_out(wire_d3_102),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance43103(.data_in(wire_d3_102),.data_out(wire_d3_103),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance43104(.data_in(wire_d3_103),.data_out(wire_d3_104),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance43105(.data_in(wire_d3_104),.data_out(wire_d3_105),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance43106(.data_in(wire_d3_105),.data_out(wire_d3_106),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance43107(.data_in(wire_d3_106),.data_out(wire_d3_107),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance43108(.data_in(wire_d3_107),.data_out(wire_d3_108),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance43109(.data_in(wire_d3_108),.data_out(wire_d3_109),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance43110(.data_in(wire_d3_109),.data_out(wire_d3_110),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance43111(.data_in(wire_d3_110),.data_out(wire_d3_111),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance43112(.data_in(wire_d3_111),.data_out(wire_d3_112),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance43113(.data_in(wire_d3_112),.data_out(wire_d3_113),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance43114(.data_in(wire_d3_113),.data_out(wire_d3_114),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance43115(.data_in(wire_d3_114),.data_out(wire_d3_115),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance43116(.data_in(wire_d3_115),.data_out(wire_d3_116),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance43117(.data_in(wire_d3_116),.data_out(wire_d3_117),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance43118(.data_in(wire_d3_117),.data_out(wire_d3_118),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance43119(.data_in(wire_d3_118),.data_out(d_out3),.clk(clk),.rst(rst));

	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance540(.data_in(d_in4),.data_out(wire_d4_0),.clk(clk),.rst(rst));            //channel 5
	decoder_top #(.WIDTH(WIDTH)) decoder_instance541(.data_in(wire_d4_0),.data_out(wire_d4_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance542(.data_in(wire_d4_1),.data_out(wire_d4_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance543(.data_in(wire_d4_2),.data_out(wire_d4_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance544(.data_in(wire_d4_3),.data_out(wire_d4_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance545(.data_in(wire_d4_4),.data_out(wire_d4_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance546(.data_in(wire_d4_5),.data_out(wire_d4_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance547(.data_in(wire_d4_6),.data_out(wire_d4_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance548(.data_in(wire_d4_7),.data_out(wire_d4_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance549(.data_in(wire_d4_8),.data_out(wire_d4_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5410(.data_in(wire_d4_9),.data_out(wire_d4_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5411(.data_in(wire_d4_10),.data_out(wire_d4_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5412(.data_in(wire_d4_11),.data_out(wire_d4_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5413(.data_in(wire_d4_12),.data_out(wire_d4_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5414(.data_in(wire_d4_13),.data_out(wire_d4_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5415(.data_in(wire_d4_14),.data_out(wire_d4_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5416(.data_in(wire_d4_15),.data_out(wire_d4_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5417(.data_in(wire_d4_16),.data_out(wire_d4_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5418(.data_in(wire_d4_17),.data_out(wire_d4_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5419(.data_in(wire_d4_18),.data_out(wire_d4_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5420(.data_in(wire_d4_19),.data_out(wire_d4_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5421(.data_in(wire_d4_20),.data_out(wire_d4_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5422(.data_in(wire_d4_21),.data_out(wire_d4_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5423(.data_in(wire_d4_22),.data_out(wire_d4_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5424(.data_in(wire_d4_23),.data_out(wire_d4_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5425(.data_in(wire_d4_24),.data_out(wire_d4_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5426(.data_in(wire_d4_25),.data_out(wire_d4_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5427(.data_in(wire_d4_26),.data_out(wire_d4_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5428(.data_in(wire_d4_27),.data_out(wire_d4_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5429(.data_in(wire_d4_28),.data_out(wire_d4_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5430(.data_in(wire_d4_29),.data_out(wire_d4_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5431(.data_in(wire_d4_30),.data_out(wire_d4_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5432(.data_in(wire_d4_31),.data_out(wire_d4_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5433(.data_in(wire_d4_32),.data_out(wire_d4_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5434(.data_in(wire_d4_33),.data_out(wire_d4_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5435(.data_in(wire_d4_34),.data_out(wire_d4_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5436(.data_in(wire_d4_35),.data_out(wire_d4_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5437(.data_in(wire_d4_36),.data_out(wire_d4_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5438(.data_in(wire_d4_37),.data_out(wire_d4_38),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5439(.data_in(wire_d4_38),.data_out(wire_d4_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5440(.data_in(wire_d4_39),.data_out(wire_d4_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5441(.data_in(wire_d4_40),.data_out(wire_d4_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5442(.data_in(wire_d4_41),.data_out(wire_d4_42),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5443(.data_in(wire_d4_42),.data_out(wire_d4_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5444(.data_in(wire_d4_43),.data_out(wire_d4_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5445(.data_in(wire_d4_44),.data_out(wire_d4_45),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5446(.data_in(wire_d4_45),.data_out(wire_d4_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5447(.data_in(wire_d4_46),.data_out(wire_d4_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5448(.data_in(wire_d4_47),.data_out(wire_d4_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5449(.data_in(wire_d4_48),.data_out(wire_d4_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5450(.data_in(wire_d4_49),.data_out(wire_d4_50),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5451(.data_in(wire_d4_50),.data_out(wire_d4_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5452(.data_in(wire_d4_51),.data_out(wire_d4_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5453(.data_in(wire_d4_52),.data_out(wire_d4_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5454(.data_in(wire_d4_53),.data_out(wire_d4_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5455(.data_in(wire_d4_54),.data_out(wire_d4_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5456(.data_in(wire_d4_55),.data_out(wire_d4_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5457(.data_in(wire_d4_56),.data_out(wire_d4_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5458(.data_in(wire_d4_57),.data_out(wire_d4_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5459(.data_in(wire_d4_58),.data_out(wire_d4_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5460(.data_in(wire_d4_59),.data_out(wire_d4_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5461(.data_in(wire_d4_60),.data_out(wire_d4_61),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5462(.data_in(wire_d4_61),.data_out(wire_d4_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5463(.data_in(wire_d4_62),.data_out(wire_d4_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5464(.data_in(wire_d4_63),.data_out(wire_d4_64),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5465(.data_in(wire_d4_64),.data_out(wire_d4_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5466(.data_in(wire_d4_65),.data_out(wire_d4_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5467(.data_in(wire_d4_66),.data_out(wire_d4_67),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5468(.data_in(wire_d4_67),.data_out(wire_d4_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5469(.data_in(wire_d4_68),.data_out(wire_d4_69),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5470(.data_in(wire_d4_69),.data_out(wire_d4_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5471(.data_in(wire_d4_70),.data_out(wire_d4_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5472(.data_in(wire_d4_71),.data_out(wire_d4_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5473(.data_in(wire_d4_72),.data_out(wire_d4_73),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5474(.data_in(wire_d4_73),.data_out(wire_d4_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5475(.data_in(wire_d4_74),.data_out(wire_d4_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5476(.data_in(wire_d4_75),.data_out(wire_d4_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5477(.data_in(wire_d4_76),.data_out(wire_d4_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5478(.data_in(wire_d4_77),.data_out(wire_d4_78),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5479(.data_in(wire_d4_78),.data_out(wire_d4_79),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5480(.data_in(wire_d4_79),.data_out(wire_d4_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5481(.data_in(wire_d4_80),.data_out(wire_d4_81),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5482(.data_in(wire_d4_81),.data_out(wire_d4_82),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5483(.data_in(wire_d4_82),.data_out(wire_d4_83),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5484(.data_in(wire_d4_83),.data_out(wire_d4_84),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5485(.data_in(wire_d4_84),.data_out(wire_d4_85),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5486(.data_in(wire_d4_85),.data_out(wire_d4_86),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5487(.data_in(wire_d4_86),.data_out(wire_d4_87),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5488(.data_in(wire_d4_87),.data_out(wire_d4_88),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5489(.data_in(wire_d4_88),.data_out(wire_d4_89),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5490(.data_in(wire_d4_89),.data_out(wire_d4_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5491(.data_in(wire_d4_90),.data_out(wire_d4_91),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5492(.data_in(wire_d4_91),.data_out(wire_d4_92),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5493(.data_in(wire_d4_92),.data_out(wire_d4_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5494(.data_in(wire_d4_93),.data_out(wire_d4_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5495(.data_in(wire_d4_94),.data_out(wire_d4_95),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5496(.data_in(wire_d4_95),.data_out(wire_d4_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5497(.data_in(wire_d4_96),.data_out(wire_d4_97),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5498(.data_in(wire_d4_97),.data_out(wire_d4_98),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5499(.data_in(wire_d4_98),.data_out(wire_d4_99),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance54100(.data_in(wire_d4_99),.data_out(wire_d4_100),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance54101(.data_in(wire_d4_100),.data_out(wire_d4_101),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance54102(.data_in(wire_d4_101),.data_out(wire_d4_102),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance54103(.data_in(wire_d4_102),.data_out(wire_d4_103),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance54104(.data_in(wire_d4_103),.data_out(wire_d4_104),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance54105(.data_in(wire_d4_104),.data_out(wire_d4_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54106(.data_in(wire_d4_105),.data_out(wire_d4_106),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance54107(.data_in(wire_d4_106),.data_out(wire_d4_107),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance54108(.data_in(wire_d4_107),.data_out(wire_d4_108),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance54109(.data_in(wire_d4_108),.data_out(wire_d4_109),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance54110(.data_in(wire_d4_109),.data_out(wire_d4_110),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance54111(.data_in(wire_d4_110),.data_out(wire_d4_111),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance54112(.data_in(wire_d4_111),.data_out(wire_d4_112),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance54113(.data_in(wire_d4_112),.data_out(wire_d4_113),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance54114(.data_in(wire_d4_113),.data_out(wire_d4_114),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance54115(.data_in(wire_d4_114),.data_out(wire_d4_115),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance54116(.data_in(wire_d4_115),.data_out(wire_d4_116),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance54117(.data_in(wire_d4_116),.data_out(wire_d4_117),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance54118(.data_in(wire_d4_117),.data_out(wire_d4_118),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance54119(.data_in(wire_d4_118),.data_out(d_out4),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance650(.data_in(d_in5),.data_out(wire_d5_0),.clk(clk),.rst(rst));            //channel 6
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance651(.data_in(wire_d5_0),.data_out(wire_d5_1),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance652(.data_in(wire_d5_1),.data_out(wire_d5_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance653(.data_in(wire_d5_2),.data_out(wire_d5_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance654(.data_in(wire_d5_3),.data_out(wire_d5_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance655(.data_in(wire_d5_4),.data_out(wire_d5_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance656(.data_in(wire_d5_5),.data_out(wire_d5_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance657(.data_in(wire_d5_6),.data_out(wire_d5_7),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance658(.data_in(wire_d5_7),.data_out(wire_d5_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance659(.data_in(wire_d5_8),.data_out(wire_d5_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6510(.data_in(wire_d5_9),.data_out(wire_d5_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6511(.data_in(wire_d5_10),.data_out(wire_d5_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6512(.data_in(wire_d5_11),.data_out(wire_d5_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6513(.data_in(wire_d5_12),.data_out(wire_d5_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6514(.data_in(wire_d5_13),.data_out(wire_d5_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6515(.data_in(wire_d5_14),.data_out(wire_d5_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6516(.data_in(wire_d5_15),.data_out(wire_d5_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6517(.data_in(wire_d5_16),.data_out(wire_d5_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6518(.data_in(wire_d5_17),.data_out(wire_d5_18),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6519(.data_in(wire_d5_18),.data_out(wire_d5_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6520(.data_in(wire_d5_19),.data_out(wire_d5_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6521(.data_in(wire_d5_20),.data_out(wire_d5_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6522(.data_in(wire_d5_21),.data_out(wire_d5_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6523(.data_in(wire_d5_22),.data_out(wire_d5_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6524(.data_in(wire_d5_23),.data_out(wire_d5_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6525(.data_in(wire_d5_24),.data_out(wire_d5_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6526(.data_in(wire_d5_25),.data_out(wire_d5_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6527(.data_in(wire_d5_26),.data_out(wire_d5_27),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6528(.data_in(wire_d5_27),.data_out(wire_d5_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6529(.data_in(wire_d5_28),.data_out(wire_d5_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6530(.data_in(wire_d5_29),.data_out(wire_d5_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6531(.data_in(wire_d5_30),.data_out(wire_d5_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6532(.data_in(wire_d5_31),.data_out(wire_d5_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6533(.data_in(wire_d5_32),.data_out(wire_d5_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6534(.data_in(wire_d5_33),.data_out(wire_d5_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6535(.data_in(wire_d5_34),.data_out(wire_d5_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6536(.data_in(wire_d5_35),.data_out(wire_d5_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6537(.data_in(wire_d5_36),.data_out(wire_d5_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6538(.data_in(wire_d5_37),.data_out(wire_d5_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6539(.data_in(wire_d5_38),.data_out(wire_d5_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6540(.data_in(wire_d5_39),.data_out(wire_d5_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6541(.data_in(wire_d5_40),.data_out(wire_d5_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6542(.data_in(wire_d5_41),.data_out(wire_d5_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6543(.data_in(wire_d5_42),.data_out(wire_d5_43),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6544(.data_in(wire_d5_43),.data_out(wire_d5_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6545(.data_in(wire_d5_44),.data_out(wire_d5_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6546(.data_in(wire_d5_45),.data_out(wire_d5_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6547(.data_in(wire_d5_46),.data_out(wire_d5_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6548(.data_in(wire_d5_47),.data_out(wire_d5_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6549(.data_in(wire_d5_48),.data_out(wire_d5_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6550(.data_in(wire_d5_49),.data_out(wire_d5_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6551(.data_in(wire_d5_50),.data_out(wire_d5_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6552(.data_in(wire_d5_51),.data_out(wire_d5_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6553(.data_in(wire_d5_52),.data_out(wire_d5_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6554(.data_in(wire_d5_53),.data_out(wire_d5_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6555(.data_in(wire_d5_54),.data_out(wire_d5_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6556(.data_in(wire_d5_55),.data_out(wire_d5_56),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6557(.data_in(wire_d5_56),.data_out(wire_d5_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6558(.data_in(wire_d5_57),.data_out(wire_d5_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6559(.data_in(wire_d5_58),.data_out(wire_d5_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6560(.data_in(wire_d5_59),.data_out(wire_d5_60),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6561(.data_in(wire_d5_60),.data_out(wire_d5_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6562(.data_in(wire_d5_61),.data_out(wire_d5_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6563(.data_in(wire_d5_62),.data_out(wire_d5_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6564(.data_in(wire_d5_63),.data_out(wire_d5_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6565(.data_in(wire_d5_64),.data_out(wire_d5_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6566(.data_in(wire_d5_65),.data_out(wire_d5_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6567(.data_in(wire_d5_66),.data_out(wire_d5_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6568(.data_in(wire_d5_67),.data_out(wire_d5_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6569(.data_in(wire_d5_68),.data_out(wire_d5_69),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6570(.data_in(wire_d5_69),.data_out(wire_d5_70),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6571(.data_in(wire_d5_70),.data_out(wire_d5_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6572(.data_in(wire_d5_71),.data_out(wire_d5_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6573(.data_in(wire_d5_72),.data_out(wire_d5_73),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6574(.data_in(wire_d5_73),.data_out(wire_d5_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6575(.data_in(wire_d5_74),.data_out(wire_d5_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6576(.data_in(wire_d5_75),.data_out(wire_d5_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6577(.data_in(wire_d5_76),.data_out(wire_d5_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6578(.data_in(wire_d5_77),.data_out(wire_d5_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6579(.data_in(wire_d5_78),.data_out(wire_d5_79),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6580(.data_in(wire_d5_79),.data_out(wire_d5_80),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6581(.data_in(wire_d5_80),.data_out(wire_d5_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6582(.data_in(wire_d5_81),.data_out(wire_d5_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6583(.data_in(wire_d5_82),.data_out(wire_d5_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6584(.data_in(wire_d5_83),.data_out(wire_d5_84),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6585(.data_in(wire_d5_84),.data_out(wire_d5_85),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6586(.data_in(wire_d5_85),.data_out(wire_d5_86),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6587(.data_in(wire_d5_86),.data_out(wire_d5_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6588(.data_in(wire_d5_87),.data_out(wire_d5_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6589(.data_in(wire_d5_88),.data_out(wire_d5_89),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6590(.data_in(wire_d5_89),.data_out(wire_d5_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6591(.data_in(wire_d5_90),.data_out(wire_d5_91),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6592(.data_in(wire_d5_91),.data_out(wire_d5_92),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6593(.data_in(wire_d5_92),.data_out(wire_d5_93),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6594(.data_in(wire_d5_93),.data_out(wire_d5_94),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6595(.data_in(wire_d5_94),.data_out(wire_d5_95),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6596(.data_in(wire_d5_95),.data_out(wire_d5_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6597(.data_in(wire_d5_96),.data_out(wire_d5_97),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6598(.data_in(wire_d5_97),.data_out(wire_d5_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6599(.data_in(wire_d5_98),.data_out(wire_d5_99),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance65100(.data_in(wire_d5_99),.data_out(wire_d5_100),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance65101(.data_in(wire_d5_100),.data_out(wire_d5_101),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance65102(.data_in(wire_d5_101),.data_out(wire_d5_102),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65103(.data_in(wire_d5_102),.data_out(wire_d5_103),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance65104(.data_in(wire_d5_103),.data_out(wire_d5_104),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance65105(.data_in(wire_d5_104),.data_out(wire_d5_105),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance65106(.data_in(wire_d5_105),.data_out(wire_d5_106),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance65107(.data_in(wire_d5_106),.data_out(wire_d5_107),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance65108(.data_in(wire_d5_107),.data_out(wire_d5_108),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance65109(.data_in(wire_d5_108),.data_out(wire_d5_109),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance65110(.data_in(wire_d5_109),.data_out(wire_d5_110),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance65111(.data_in(wire_d5_110),.data_out(wire_d5_111),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance65112(.data_in(wire_d5_111),.data_out(wire_d5_112),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance65113(.data_in(wire_d5_112),.data_out(wire_d5_113),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance65114(.data_in(wire_d5_113),.data_out(wire_d5_114),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance65115(.data_in(wire_d5_114),.data_out(wire_d5_115),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance65116(.data_in(wire_d5_115),.data_out(wire_d5_116),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance65117(.data_in(wire_d5_116),.data_out(wire_d5_117),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance65118(.data_in(wire_d5_117),.data_out(wire_d5_118),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance65119(.data_in(wire_d5_118),.data_out(d_out5),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance760(.data_in(d_in6),.data_out(wire_d6_0),.clk(clk),.rst(rst));            //channel 7
	large_mux #(.WIDTH(WIDTH)) large_mux_instance761(.data_in(wire_d6_0),.data_out(wire_d6_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance762(.data_in(wire_d6_1),.data_out(wire_d6_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance763(.data_in(wire_d6_2),.data_out(wire_d6_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance764(.data_in(wire_d6_3),.data_out(wire_d6_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance765(.data_in(wire_d6_4),.data_out(wire_d6_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance766(.data_in(wire_d6_5),.data_out(wire_d6_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767(.data_in(wire_d6_6),.data_out(wire_d6_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance768(.data_in(wire_d6_7),.data_out(wire_d6_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance769(.data_in(wire_d6_8),.data_out(wire_d6_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7610(.data_in(wire_d6_9),.data_out(wire_d6_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7611(.data_in(wire_d6_10),.data_out(wire_d6_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7612(.data_in(wire_d6_11),.data_out(wire_d6_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7613(.data_in(wire_d6_12),.data_out(wire_d6_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7614(.data_in(wire_d6_13),.data_out(wire_d6_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7615(.data_in(wire_d6_14),.data_out(wire_d6_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7616(.data_in(wire_d6_15),.data_out(wire_d6_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7617(.data_in(wire_d6_16),.data_out(wire_d6_17),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7618(.data_in(wire_d6_17),.data_out(wire_d6_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7619(.data_in(wire_d6_18),.data_out(wire_d6_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7620(.data_in(wire_d6_19),.data_out(wire_d6_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7621(.data_in(wire_d6_20),.data_out(wire_d6_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7622(.data_in(wire_d6_21),.data_out(wire_d6_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7623(.data_in(wire_d6_22),.data_out(wire_d6_23),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7624(.data_in(wire_d6_23),.data_out(wire_d6_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7625(.data_in(wire_d6_24),.data_out(wire_d6_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7626(.data_in(wire_d6_25),.data_out(wire_d6_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7627(.data_in(wire_d6_26),.data_out(wire_d6_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7628(.data_in(wire_d6_27),.data_out(wire_d6_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7629(.data_in(wire_d6_28),.data_out(wire_d6_29),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7630(.data_in(wire_d6_29),.data_out(wire_d6_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7631(.data_in(wire_d6_30),.data_out(wire_d6_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7632(.data_in(wire_d6_31),.data_out(wire_d6_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7633(.data_in(wire_d6_32),.data_out(wire_d6_33),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7634(.data_in(wire_d6_33),.data_out(wire_d6_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7635(.data_in(wire_d6_34),.data_out(wire_d6_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7636(.data_in(wire_d6_35),.data_out(wire_d6_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7637(.data_in(wire_d6_36),.data_out(wire_d6_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7638(.data_in(wire_d6_37),.data_out(wire_d6_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7639(.data_in(wire_d6_38),.data_out(wire_d6_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7640(.data_in(wire_d6_39),.data_out(wire_d6_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7641(.data_in(wire_d6_40),.data_out(wire_d6_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7642(.data_in(wire_d6_41),.data_out(wire_d6_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7643(.data_in(wire_d6_42),.data_out(wire_d6_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7644(.data_in(wire_d6_43),.data_out(wire_d6_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7645(.data_in(wire_d6_44),.data_out(wire_d6_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7646(.data_in(wire_d6_45),.data_out(wire_d6_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7647(.data_in(wire_d6_46),.data_out(wire_d6_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7648(.data_in(wire_d6_47),.data_out(wire_d6_48),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7649(.data_in(wire_d6_48),.data_out(wire_d6_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7650(.data_in(wire_d6_49),.data_out(wire_d6_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7651(.data_in(wire_d6_50),.data_out(wire_d6_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7652(.data_in(wire_d6_51),.data_out(wire_d6_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7653(.data_in(wire_d6_52),.data_out(wire_d6_53),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7654(.data_in(wire_d6_53),.data_out(wire_d6_54),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7655(.data_in(wire_d6_54),.data_out(wire_d6_55),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7656(.data_in(wire_d6_55),.data_out(wire_d6_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7657(.data_in(wire_d6_56),.data_out(wire_d6_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7658(.data_in(wire_d6_57),.data_out(wire_d6_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7659(.data_in(wire_d6_58),.data_out(wire_d6_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7660(.data_in(wire_d6_59),.data_out(wire_d6_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7661(.data_in(wire_d6_60),.data_out(wire_d6_61),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7662(.data_in(wire_d6_61),.data_out(wire_d6_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7663(.data_in(wire_d6_62),.data_out(wire_d6_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7664(.data_in(wire_d6_63),.data_out(wire_d6_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7665(.data_in(wire_d6_64),.data_out(wire_d6_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7666(.data_in(wire_d6_65),.data_out(wire_d6_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7667(.data_in(wire_d6_66),.data_out(wire_d6_67),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7668(.data_in(wire_d6_67),.data_out(wire_d6_68),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7669(.data_in(wire_d6_68),.data_out(wire_d6_69),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7670(.data_in(wire_d6_69),.data_out(wire_d6_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7671(.data_in(wire_d6_70),.data_out(wire_d6_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7672(.data_in(wire_d6_71),.data_out(wire_d6_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7673(.data_in(wire_d6_72),.data_out(wire_d6_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7674(.data_in(wire_d6_73),.data_out(wire_d6_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7675(.data_in(wire_d6_74),.data_out(wire_d6_75),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7676(.data_in(wire_d6_75),.data_out(wire_d6_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7677(.data_in(wire_d6_76),.data_out(wire_d6_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7678(.data_in(wire_d6_77),.data_out(wire_d6_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7679(.data_in(wire_d6_78),.data_out(wire_d6_79),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7680(.data_in(wire_d6_79),.data_out(wire_d6_80),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7681(.data_in(wire_d6_80),.data_out(wire_d6_81),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7682(.data_in(wire_d6_81),.data_out(wire_d6_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7683(.data_in(wire_d6_82),.data_out(wire_d6_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7684(.data_in(wire_d6_83),.data_out(wire_d6_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7685(.data_in(wire_d6_84),.data_out(wire_d6_85),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7686(.data_in(wire_d6_85),.data_out(wire_d6_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7687(.data_in(wire_d6_86),.data_out(wire_d6_87),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7688(.data_in(wire_d6_87),.data_out(wire_d6_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7689(.data_in(wire_d6_88),.data_out(wire_d6_89),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7690(.data_in(wire_d6_89),.data_out(wire_d6_90),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7691(.data_in(wire_d6_90),.data_out(wire_d6_91),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7692(.data_in(wire_d6_91),.data_out(wire_d6_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7693(.data_in(wire_d6_92),.data_out(wire_d6_93),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7694(.data_in(wire_d6_93),.data_out(wire_d6_94),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7695(.data_in(wire_d6_94),.data_out(wire_d6_95),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7696(.data_in(wire_d6_95),.data_out(wire_d6_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7697(.data_in(wire_d6_96),.data_out(wire_d6_97),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7698(.data_in(wire_d6_97),.data_out(wire_d6_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7699(.data_in(wire_d6_98),.data_out(wire_d6_99),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance76100(.data_in(wire_d6_99),.data_out(wire_d6_100),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance76101(.data_in(wire_d6_100),.data_out(wire_d6_101),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance76102(.data_in(wire_d6_101),.data_out(wire_d6_102),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance76103(.data_in(wire_d6_102),.data_out(wire_d6_103),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance76104(.data_in(wire_d6_103),.data_out(wire_d6_104),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance76105(.data_in(wire_d6_104),.data_out(wire_d6_105),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance76106(.data_in(wire_d6_105),.data_out(wire_d6_106),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76107(.data_in(wire_d6_106),.data_out(wire_d6_107),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance76108(.data_in(wire_d6_107),.data_out(wire_d6_108),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance76109(.data_in(wire_d6_108),.data_out(wire_d6_109),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance76110(.data_in(wire_d6_109),.data_out(wire_d6_110),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance76111(.data_in(wire_d6_110),.data_out(wire_d6_111),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance76112(.data_in(wire_d6_111),.data_out(wire_d6_112),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance76113(.data_in(wire_d6_112),.data_out(wire_d6_113),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance76114(.data_in(wire_d6_113),.data_out(wire_d6_114),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance76115(.data_in(wire_d6_114),.data_out(wire_d6_115),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance76116(.data_in(wire_d6_115),.data_out(wire_d6_116),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance76117(.data_in(wire_d6_116),.data_out(wire_d6_117),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance76118(.data_in(wire_d6_117),.data_out(wire_d6_118),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance76119(.data_in(wire_d6_118),.data_out(d_out6),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance870(.data_in(d_in7),.data_out(wire_d7_0),.clk(clk),.rst(rst));            //channel 8
	decoder_top #(.WIDTH(WIDTH)) decoder_instance871(.data_in(wire_d7_0),.data_out(wire_d7_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance872(.data_in(wire_d7_1),.data_out(wire_d7_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance873(.data_in(wire_d7_2),.data_out(wire_d7_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance874(.data_in(wire_d7_3),.data_out(wire_d7_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance875(.data_in(wire_d7_4),.data_out(wire_d7_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance876(.data_in(wire_d7_5),.data_out(wire_d7_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance877(.data_in(wire_d7_6),.data_out(wire_d7_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance878(.data_in(wire_d7_7),.data_out(wire_d7_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance879(.data_in(wire_d7_8),.data_out(wire_d7_9),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8710(.data_in(wire_d7_9),.data_out(wire_d7_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8711(.data_in(wire_d7_10),.data_out(wire_d7_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8712(.data_in(wire_d7_11),.data_out(wire_d7_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8713(.data_in(wire_d7_12),.data_out(wire_d7_13),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8714(.data_in(wire_d7_13),.data_out(wire_d7_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8715(.data_in(wire_d7_14),.data_out(wire_d7_15),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8716(.data_in(wire_d7_15),.data_out(wire_d7_16),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8717(.data_in(wire_d7_16),.data_out(wire_d7_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8718(.data_in(wire_d7_17),.data_out(wire_d7_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8719(.data_in(wire_d7_18),.data_out(wire_d7_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8720(.data_in(wire_d7_19),.data_out(wire_d7_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8721(.data_in(wire_d7_20),.data_out(wire_d7_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8722(.data_in(wire_d7_21),.data_out(wire_d7_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8723(.data_in(wire_d7_22),.data_out(wire_d7_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8724(.data_in(wire_d7_23),.data_out(wire_d7_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8725(.data_in(wire_d7_24),.data_out(wire_d7_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8726(.data_in(wire_d7_25),.data_out(wire_d7_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8727(.data_in(wire_d7_26),.data_out(wire_d7_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8728(.data_in(wire_d7_27),.data_out(wire_d7_28),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8729(.data_in(wire_d7_28),.data_out(wire_d7_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8730(.data_in(wire_d7_29),.data_out(wire_d7_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8731(.data_in(wire_d7_30),.data_out(wire_d7_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8732(.data_in(wire_d7_31),.data_out(wire_d7_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8733(.data_in(wire_d7_32),.data_out(wire_d7_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8734(.data_in(wire_d7_33),.data_out(wire_d7_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8735(.data_in(wire_d7_34),.data_out(wire_d7_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8736(.data_in(wire_d7_35),.data_out(wire_d7_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8737(.data_in(wire_d7_36),.data_out(wire_d7_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8738(.data_in(wire_d7_37),.data_out(wire_d7_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8739(.data_in(wire_d7_38),.data_out(wire_d7_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8740(.data_in(wire_d7_39),.data_out(wire_d7_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8741(.data_in(wire_d7_40),.data_out(wire_d7_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8742(.data_in(wire_d7_41),.data_out(wire_d7_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8743(.data_in(wire_d7_42),.data_out(wire_d7_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8744(.data_in(wire_d7_43),.data_out(wire_d7_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8745(.data_in(wire_d7_44),.data_out(wire_d7_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8746(.data_in(wire_d7_45),.data_out(wire_d7_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8747(.data_in(wire_d7_46),.data_out(wire_d7_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8748(.data_in(wire_d7_47),.data_out(wire_d7_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8749(.data_in(wire_d7_48),.data_out(wire_d7_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8750(.data_in(wire_d7_49),.data_out(wire_d7_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8751(.data_in(wire_d7_50),.data_out(wire_d7_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8752(.data_in(wire_d7_51),.data_out(wire_d7_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8753(.data_in(wire_d7_52),.data_out(wire_d7_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8754(.data_in(wire_d7_53),.data_out(wire_d7_54),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8755(.data_in(wire_d7_54),.data_out(wire_d7_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8756(.data_in(wire_d7_55),.data_out(wire_d7_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8757(.data_in(wire_d7_56),.data_out(wire_d7_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8758(.data_in(wire_d7_57),.data_out(wire_d7_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8759(.data_in(wire_d7_58),.data_out(wire_d7_59),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8760(.data_in(wire_d7_59),.data_out(wire_d7_60),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8761(.data_in(wire_d7_60),.data_out(wire_d7_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8762(.data_in(wire_d7_61),.data_out(wire_d7_62),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8763(.data_in(wire_d7_62),.data_out(wire_d7_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8764(.data_in(wire_d7_63),.data_out(wire_d7_64),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8765(.data_in(wire_d7_64),.data_out(wire_d7_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8766(.data_in(wire_d7_65),.data_out(wire_d7_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8767(.data_in(wire_d7_66),.data_out(wire_d7_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8768(.data_in(wire_d7_67),.data_out(wire_d7_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8769(.data_in(wire_d7_68),.data_out(wire_d7_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8770(.data_in(wire_d7_69),.data_out(wire_d7_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8771(.data_in(wire_d7_70),.data_out(wire_d7_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8772(.data_in(wire_d7_71),.data_out(wire_d7_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8773(.data_in(wire_d7_72),.data_out(wire_d7_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8774(.data_in(wire_d7_73),.data_out(wire_d7_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8775(.data_in(wire_d7_74),.data_out(wire_d7_75),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8776(.data_in(wire_d7_75),.data_out(wire_d7_76),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8777(.data_in(wire_d7_76),.data_out(wire_d7_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8778(.data_in(wire_d7_77),.data_out(wire_d7_78),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8779(.data_in(wire_d7_78),.data_out(wire_d7_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8780(.data_in(wire_d7_79),.data_out(wire_d7_80),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8781(.data_in(wire_d7_80),.data_out(wire_d7_81),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8782(.data_in(wire_d7_81),.data_out(wire_d7_82),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8783(.data_in(wire_d7_82),.data_out(wire_d7_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8784(.data_in(wire_d7_83),.data_out(wire_d7_84),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8785(.data_in(wire_d7_84),.data_out(wire_d7_85),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8786(.data_in(wire_d7_85),.data_out(wire_d7_86),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8787(.data_in(wire_d7_86),.data_out(wire_d7_87),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8788(.data_in(wire_d7_87),.data_out(wire_d7_88),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8789(.data_in(wire_d7_88),.data_out(wire_d7_89),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8790(.data_in(wire_d7_89),.data_out(wire_d7_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8791(.data_in(wire_d7_90),.data_out(wire_d7_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8792(.data_in(wire_d7_91),.data_out(wire_d7_92),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8793(.data_in(wire_d7_92),.data_out(wire_d7_93),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8794(.data_in(wire_d7_93),.data_out(wire_d7_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8795(.data_in(wire_d7_94),.data_out(wire_d7_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8796(.data_in(wire_d7_95),.data_out(wire_d7_96),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8797(.data_in(wire_d7_96),.data_out(wire_d7_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8798(.data_in(wire_d7_97),.data_out(wire_d7_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8799(.data_in(wire_d7_98),.data_out(wire_d7_99),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance87100(.data_in(wire_d7_99),.data_out(wire_d7_100),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance87101(.data_in(wire_d7_100),.data_out(wire_d7_101),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance87102(.data_in(wire_d7_101),.data_out(wire_d7_102),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance87103(.data_in(wire_d7_102),.data_out(wire_d7_103),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance87104(.data_in(wire_d7_103),.data_out(wire_d7_104),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87105(.data_in(wire_d7_104),.data_out(wire_d7_105),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance87106(.data_in(wire_d7_105),.data_out(wire_d7_106),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance87107(.data_in(wire_d7_106),.data_out(wire_d7_107),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance87108(.data_in(wire_d7_107),.data_out(wire_d7_108),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance87109(.data_in(wire_d7_108),.data_out(wire_d7_109),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance87110(.data_in(wire_d7_109),.data_out(wire_d7_110),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance87111(.data_in(wire_d7_110),.data_out(wire_d7_111),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance87112(.data_in(wire_d7_111),.data_out(wire_d7_112),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance87113(.data_in(wire_d7_112),.data_out(wire_d7_113),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance87114(.data_in(wire_d7_113),.data_out(wire_d7_114),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance87115(.data_in(wire_d7_114),.data_out(wire_d7_115),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance87116(.data_in(wire_d7_115),.data_out(wire_d7_116),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance87117(.data_in(wire_d7_116),.data_out(wire_d7_117),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance87118(.data_in(wire_d7_117),.data_out(wire_d7_118),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance87119(.data_in(wire_d7_118),.data_out(d_out7),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance980(.data_in(d_in8),.data_out(wire_d8_0),.clk(clk),.rst(rst));            //channel 9
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance981(.data_in(wire_d8_0),.data_out(wire_d8_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance982(.data_in(wire_d8_1),.data_out(wire_d8_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance983(.data_in(wire_d8_2),.data_out(wire_d8_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance984(.data_in(wire_d8_3),.data_out(wire_d8_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance985(.data_in(wire_d8_4),.data_out(wire_d8_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance986(.data_in(wire_d8_5),.data_out(wire_d8_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance987(.data_in(wire_d8_6),.data_out(wire_d8_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance988(.data_in(wire_d8_7),.data_out(wire_d8_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance989(.data_in(wire_d8_8),.data_out(wire_d8_9),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9810(.data_in(wire_d8_9),.data_out(wire_d8_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9811(.data_in(wire_d8_10),.data_out(wire_d8_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9812(.data_in(wire_d8_11),.data_out(wire_d8_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9813(.data_in(wire_d8_12),.data_out(wire_d8_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9814(.data_in(wire_d8_13),.data_out(wire_d8_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9815(.data_in(wire_d8_14),.data_out(wire_d8_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9816(.data_in(wire_d8_15),.data_out(wire_d8_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9817(.data_in(wire_d8_16),.data_out(wire_d8_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9818(.data_in(wire_d8_17),.data_out(wire_d8_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9819(.data_in(wire_d8_18),.data_out(wire_d8_19),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9820(.data_in(wire_d8_19),.data_out(wire_d8_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9821(.data_in(wire_d8_20),.data_out(wire_d8_21),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9822(.data_in(wire_d8_21),.data_out(wire_d8_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9823(.data_in(wire_d8_22),.data_out(wire_d8_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9824(.data_in(wire_d8_23),.data_out(wire_d8_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9825(.data_in(wire_d8_24),.data_out(wire_d8_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9826(.data_in(wire_d8_25),.data_out(wire_d8_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9827(.data_in(wire_d8_26),.data_out(wire_d8_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9828(.data_in(wire_d8_27),.data_out(wire_d8_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9829(.data_in(wire_d8_28),.data_out(wire_d8_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9830(.data_in(wire_d8_29),.data_out(wire_d8_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9831(.data_in(wire_d8_30),.data_out(wire_d8_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9832(.data_in(wire_d8_31),.data_out(wire_d8_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9833(.data_in(wire_d8_32),.data_out(wire_d8_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9834(.data_in(wire_d8_33),.data_out(wire_d8_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9835(.data_in(wire_d8_34),.data_out(wire_d8_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9836(.data_in(wire_d8_35),.data_out(wire_d8_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9837(.data_in(wire_d8_36),.data_out(wire_d8_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9838(.data_in(wire_d8_37),.data_out(wire_d8_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9839(.data_in(wire_d8_38),.data_out(wire_d8_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9840(.data_in(wire_d8_39),.data_out(wire_d8_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9841(.data_in(wire_d8_40),.data_out(wire_d8_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9842(.data_in(wire_d8_41),.data_out(wire_d8_42),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9843(.data_in(wire_d8_42),.data_out(wire_d8_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9844(.data_in(wire_d8_43),.data_out(wire_d8_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9845(.data_in(wire_d8_44),.data_out(wire_d8_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9846(.data_in(wire_d8_45),.data_out(wire_d8_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9847(.data_in(wire_d8_46),.data_out(wire_d8_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9848(.data_in(wire_d8_47),.data_out(wire_d8_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9849(.data_in(wire_d8_48),.data_out(wire_d8_49),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9850(.data_in(wire_d8_49),.data_out(wire_d8_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9851(.data_in(wire_d8_50),.data_out(wire_d8_51),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9852(.data_in(wire_d8_51),.data_out(wire_d8_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9853(.data_in(wire_d8_52),.data_out(wire_d8_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9854(.data_in(wire_d8_53),.data_out(wire_d8_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9855(.data_in(wire_d8_54),.data_out(wire_d8_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9856(.data_in(wire_d8_55),.data_out(wire_d8_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9857(.data_in(wire_d8_56),.data_out(wire_d8_57),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9858(.data_in(wire_d8_57),.data_out(wire_d8_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9859(.data_in(wire_d8_58),.data_out(wire_d8_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9860(.data_in(wire_d8_59),.data_out(wire_d8_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9861(.data_in(wire_d8_60),.data_out(wire_d8_61),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9862(.data_in(wire_d8_61),.data_out(wire_d8_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9863(.data_in(wire_d8_62),.data_out(wire_d8_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9864(.data_in(wire_d8_63),.data_out(wire_d8_64),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9865(.data_in(wire_d8_64),.data_out(wire_d8_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9866(.data_in(wire_d8_65),.data_out(wire_d8_66),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9867(.data_in(wire_d8_66),.data_out(wire_d8_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9868(.data_in(wire_d8_67),.data_out(wire_d8_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9869(.data_in(wire_d8_68),.data_out(wire_d8_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9870(.data_in(wire_d8_69),.data_out(wire_d8_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9871(.data_in(wire_d8_70),.data_out(wire_d8_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9872(.data_in(wire_d8_71),.data_out(wire_d8_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9873(.data_in(wire_d8_72),.data_out(wire_d8_73),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9874(.data_in(wire_d8_73),.data_out(wire_d8_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9875(.data_in(wire_d8_74),.data_out(wire_d8_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9876(.data_in(wire_d8_75),.data_out(wire_d8_76),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9877(.data_in(wire_d8_76),.data_out(wire_d8_77),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9878(.data_in(wire_d8_77),.data_out(wire_d8_78),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9879(.data_in(wire_d8_78),.data_out(wire_d8_79),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9880(.data_in(wire_d8_79),.data_out(wire_d8_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9881(.data_in(wire_d8_80),.data_out(wire_d8_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9882(.data_in(wire_d8_81),.data_out(wire_d8_82),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9883(.data_in(wire_d8_82),.data_out(wire_d8_83),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9884(.data_in(wire_d8_83),.data_out(wire_d8_84),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9885(.data_in(wire_d8_84),.data_out(wire_d8_85),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9886(.data_in(wire_d8_85),.data_out(wire_d8_86),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9887(.data_in(wire_d8_86),.data_out(wire_d8_87),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9888(.data_in(wire_d8_87),.data_out(wire_d8_88),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9889(.data_in(wire_d8_88),.data_out(wire_d8_89),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9890(.data_in(wire_d8_89),.data_out(wire_d8_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9891(.data_in(wire_d8_90),.data_out(wire_d8_91),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9892(.data_in(wire_d8_91),.data_out(wire_d8_92),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9893(.data_in(wire_d8_92),.data_out(wire_d8_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9894(.data_in(wire_d8_93),.data_out(wire_d8_94),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9895(.data_in(wire_d8_94),.data_out(wire_d8_95),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9896(.data_in(wire_d8_95),.data_out(wire_d8_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9897(.data_in(wire_d8_96),.data_out(wire_d8_97),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9898(.data_in(wire_d8_97),.data_out(wire_d8_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9899(.data_in(wire_d8_98),.data_out(wire_d8_99),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance98100(.data_in(wire_d8_99),.data_out(wire_d8_100),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance98101(.data_in(wire_d8_100),.data_out(wire_d8_101),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance98102(.data_in(wire_d8_101),.data_out(wire_d8_102),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance98103(.data_in(wire_d8_102),.data_out(wire_d8_103),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance98104(.data_in(wire_d8_103),.data_out(wire_d8_104),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance98105(.data_in(wire_d8_104),.data_out(wire_d8_105),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance98106(.data_in(wire_d8_105),.data_out(wire_d8_106),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance98107(.data_in(wire_d8_106),.data_out(wire_d8_107),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance98108(.data_in(wire_d8_107),.data_out(wire_d8_108),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance98109(.data_in(wire_d8_108),.data_out(wire_d8_109),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance98110(.data_in(wire_d8_109),.data_out(wire_d8_110),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance98111(.data_in(wire_d8_110),.data_out(wire_d8_111),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance98112(.data_in(wire_d8_111),.data_out(wire_d8_112),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance98113(.data_in(wire_d8_112),.data_out(wire_d8_113),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance98114(.data_in(wire_d8_113),.data_out(wire_d8_114),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance98115(.data_in(wire_d8_114),.data_out(wire_d8_115),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance98116(.data_in(wire_d8_115),.data_out(wire_d8_116),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance98117(.data_in(wire_d8_116),.data_out(wire_d8_117),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance98118(.data_in(wire_d8_117),.data_out(wire_d8_118),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance98119(.data_in(wire_d8_118),.data_out(d_out8),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance10090(.data_in(d_in9),.data_out(wire_d9_0),.clk(clk),.rst(rst));            //channel 10
	decoder_top #(.WIDTH(WIDTH)) decoder_instance10091(.data_in(wire_d9_0),.data_out(wire_d9_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10092(.data_in(wire_d9_1),.data_out(wire_d9_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10093(.data_in(wire_d9_2),.data_out(wire_d9_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance10094(.data_in(wire_d9_3),.data_out(wire_d9_4),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance10095(.data_in(wire_d9_4),.data_out(wire_d9_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance10096(.data_in(wire_d9_5),.data_out(wire_d9_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance10097(.data_in(wire_d9_6),.data_out(wire_d9_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance10098(.data_in(wire_d9_7),.data_out(wire_d9_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10099(.data_in(wire_d9_8),.data_out(wire_d9_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100910(.data_in(wire_d9_9),.data_out(wire_d9_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance100911(.data_in(wire_d9_10),.data_out(wire_d9_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100912(.data_in(wire_d9_11),.data_out(wire_d9_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100913(.data_in(wire_d9_12),.data_out(wire_d9_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100914(.data_in(wire_d9_13),.data_out(wire_d9_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance100915(.data_in(wire_d9_14),.data_out(wire_d9_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100916(.data_in(wire_d9_15),.data_out(wire_d9_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance100917(.data_in(wire_d9_16),.data_out(wire_d9_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance100918(.data_in(wire_d9_17),.data_out(wire_d9_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100919(.data_in(wire_d9_18),.data_out(wire_d9_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100920(.data_in(wire_d9_19),.data_out(wire_d9_20),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100921(.data_in(wire_d9_20),.data_out(wire_d9_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100922(.data_in(wire_d9_21),.data_out(wire_d9_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100923(.data_in(wire_d9_22),.data_out(wire_d9_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100924(.data_in(wire_d9_23),.data_out(wire_d9_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100925(.data_in(wire_d9_24),.data_out(wire_d9_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100926(.data_in(wire_d9_25),.data_out(wire_d9_26),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance100927(.data_in(wire_d9_26),.data_out(wire_d9_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance100928(.data_in(wire_d9_27),.data_out(wire_d9_28),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100929(.data_in(wire_d9_28),.data_out(wire_d9_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance100930(.data_in(wire_d9_29),.data_out(wire_d9_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance100931(.data_in(wire_d9_30),.data_out(wire_d9_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100932(.data_in(wire_d9_31),.data_out(wire_d9_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100933(.data_in(wire_d9_32),.data_out(wire_d9_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100934(.data_in(wire_d9_33),.data_out(wire_d9_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100935(.data_in(wire_d9_34),.data_out(wire_d9_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100936(.data_in(wire_d9_35),.data_out(wire_d9_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100937(.data_in(wire_d9_36),.data_out(wire_d9_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100938(.data_in(wire_d9_37),.data_out(wire_d9_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100939(.data_in(wire_d9_38),.data_out(wire_d9_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100940(.data_in(wire_d9_39),.data_out(wire_d9_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100941(.data_in(wire_d9_40),.data_out(wire_d9_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100942(.data_in(wire_d9_41),.data_out(wire_d9_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100943(.data_in(wire_d9_42),.data_out(wire_d9_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance100944(.data_in(wire_d9_43),.data_out(wire_d9_44),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100945(.data_in(wire_d9_44),.data_out(wire_d9_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance100946(.data_in(wire_d9_45),.data_out(wire_d9_46),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance100947(.data_in(wire_d9_46),.data_out(wire_d9_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance100948(.data_in(wire_d9_47),.data_out(wire_d9_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100949(.data_in(wire_d9_48),.data_out(wire_d9_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100950(.data_in(wire_d9_49),.data_out(wire_d9_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100951(.data_in(wire_d9_50),.data_out(wire_d9_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100952(.data_in(wire_d9_51),.data_out(wire_d9_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100953(.data_in(wire_d9_52),.data_out(wire_d9_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100954(.data_in(wire_d9_53),.data_out(wire_d9_54),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100955(.data_in(wire_d9_54),.data_out(wire_d9_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100956(.data_in(wire_d9_55),.data_out(wire_d9_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100957(.data_in(wire_d9_56),.data_out(wire_d9_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance100958(.data_in(wire_d9_57),.data_out(wire_d9_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100959(.data_in(wire_d9_58),.data_out(wire_d9_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100960(.data_in(wire_d9_59),.data_out(wire_d9_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100961(.data_in(wire_d9_60),.data_out(wire_d9_61),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance100962(.data_in(wire_d9_61),.data_out(wire_d9_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100963(.data_in(wire_d9_62),.data_out(wire_d9_63),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance100964(.data_in(wire_d9_63),.data_out(wire_d9_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100965(.data_in(wire_d9_64),.data_out(wire_d9_65),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100966(.data_in(wire_d9_65),.data_out(wire_d9_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100967(.data_in(wire_d9_66),.data_out(wire_d9_67),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100968(.data_in(wire_d9_67),.data_out(wire_d9_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100969(.data_in(wire_d9_68),.data_out(wire_d9_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100970(.data_in(wire_d9_69),.data_out(wire_d9_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100971(.data_in(wire_d9_70),.data_out(wire_d9_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100972(.data_in(wire_d9_71),.data_out(wire_d9_72),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance100973(.data_in(wire_d9_72),.data_out(wire_d9_73),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance100974(.data_in(wire_d9_73),.data_out(wire_d9_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100975(.data_in(wire_d9_74),.data_out(wire_d9_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100976(.data_in(wire_d9_75),.data_out(wire_d9_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100977(.data_in(wire_d9_76),.data_out(wire_d9_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100978(.data_in(wire_d9_77),.data_out(wire_d9_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100979(.data_in(wire_d9_78),.data_out(wire_d9_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100980(.data_in(wire_d9_79),.data_out(wire_d9_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100981(.data_in(wire_d9_80),.data_out(wire_d9_81),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance100982(.data_in(wire_d9_81),.data_out(wire_d9_82),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100983(.data_in(wire_d9_82),.data_out(wire_d9_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance100984(.data_in(wire_d9_83),.data_out(wire_d9_84),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100985(.data_in(wire_d9_84),.data_out(wire_d9_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100986(.data_in(wire_d9_85),.data_out(wire_d9_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance100987(.data_in(wire_d9_86),.data_out(wire_d9_87),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100988(.data_in(wire_d9_87),.data_out(wire_d9_88),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100989(.data_in(wire_d9_88),.data_out(wire_d9_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100990(.data_in(wire_d9_89),.data_out(wire_d9_90),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100991(.data_in(wire_d9_90),.data_out(wire_d9_91),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance100992(.data_in(wire_d9_91),.data_out(wire_d9_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100993(.data_in(wire_d9_92),.data_out(wire_d9_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100994(.data_in(wire_d9_93),.data_out(wire_d9_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100995(.data_in(wire_d9_94),.data_out(wire_d9_95),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100996(.data_in(wire_d9_95),.data_out(wire_d9_96),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100997(.data_in(wire_d9_96),.data_out(wire_d9_97),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100998(.data_in(wire_d9_97),.data_out(wire_d9_98),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100999(.data_in(wire_d9_98),.data_out(wire_d9_99),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1009100(.data_in(wire_d9_99),.data_out(wire_d9_100),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1009101(.data_in(wire_d9_100),.data_out(wire_d9_101),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009102(.data_in(wire_d9_101),.data_out(wire_d9_102),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1009103(.data_in(wire_d9_102),.data_out(wire_d9_103),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1009104(.data_in(wire_d9_103),.data_out(wire_d9_104),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1009105(.data_in(wire_d9_104),.data_out(wire_d9_105),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1009106(.data_in(wire_d9_105),.data_out(wire_d9_106),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1009107(.data_in(wire_d9_106),.data_out(wire_d9_107),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1009108(.data_in(wire_d9_107),.data_out(wire_d9_108),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1009109(.data_in(wire_d9_108),.data_out(wire_d9_109),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1009110(.data_in(wire_d9_109),.data_out(wire_d9_110),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1009111(.data_in(wire_d9_110),.data_out(wire_d9_111),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1009112(.data_in(wire_d9_111),.data_out(wire_d9_112),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1009113(.data_in(wire_d9_112),.data_out(wire_d9_113),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1009114(.data_in(wire_d9_113),.data_out(wire_d9_114),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1009115(.data_in(wire_d9_114),.data_out(wire_d9_115),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1009116(.data_in(wire_d9_115),.data_out(wire_d9_116),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1009117(.data_in(wire_d9_116),.data_out(wire_d9_117),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1009118(.data_in(wire_d9_117),.data_out(wire_d9_118),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1009119(.data_in(wire_d9_118),.data_out(d_out9),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance110100(.data_in(d_in10),.data_out(wire_d10_0),.clk(clk),.rst(rst));            //channel 11
	large_adder #(.WIDTH(WIDTH)) large_adder_instance110101(.data_in(wire_d10_0),.data_out(wire_d10_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance110102(.data_in(wire_d10_1),.data_out(wire_d10_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance110103(.data_in(wire_d10_2),.data_out(wire_d10_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance110104(.data_in(wire_d10_3),.data_out(wire_d10_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance110105(.data_in(wire_d10_4),.data_out(wire_d10_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance110106(.data_in(wire_d10_5),.data_out(wire_d10_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance110107(.data_in(wire_d10_6),.data_out(wire_d10_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance110108(.data_in(wire_d10_7),.data_out(wire_d10_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance110109(.data_in(wire_d10_8),.data_out(wire_d10_9),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101010(.data_in(wire_d10_9),.data_out(wire_d10_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1101011(.data_in(wire_d10_10),.data_out(wire_d10_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101012(.data_in(wire_d10_11),.data_out(wire_d10_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101013(.data_in(wire_d10_12),.data_out(wire_d10_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1101014(.data_in(wire_d10_13),.data_out(wire_d10_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101015(.data_in(wire_d10_14),.data_out(wire_d10_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101016(.data_in(wire_d10_15),.data_out(wire_d10_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101017(.data_in(wire_d10_16),.data_out(wire_d10_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101018(.data_in(wire_d10_17),.data_out(wire_d10_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1101019(.data_in(wire_d10_18),.data_out(wire_d10_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101020(.data_in(wire_d10_19),.data_out(wire_d10_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1101021(.data_in(wire_d10_20),.data_out(wire_d10_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101022(.data_in(wire_d10_21),.data_out(wire_d10_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1101023(.data_in(wire_d10_22),.data_out(wire_d10_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101024(.data_in(wire_d10_23),.data_out(wire_d10_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1101025(.data_in(wire_d10_24),.data_out(wire_d10_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1101026(.data_in(wire_d10_25),.data_out(wire_d10_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101027(.data_in(wire_d10_26),.data_out(wire_d10_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1101028(.data_in(wire_d10_27),.data_out(wire_d10_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1101029(.data_in(wire_d10_28),.data_out(wire_d10_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101030(.data_in(wire_d10_29),.data_out(wire_d10_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101031(.data_in(wire_d10_30),.data_out(wire_d10_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101032(.data_in(wire_d10_31),.data_out(wire_d10_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101033(.data_in(wire_d10_32),.data_out(wire_d10_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1101034(.data_in(wire_d10_33),.data_out(wire_d10_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101035(.data_in(wire_d10_34),.data_out(wire_d10_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101036(.data_in(wire_d10_35),.data_out(wire_d10_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1101037(.data_in(wire_d10_36),.data_out(wire_d10_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101038(.data_in(wire_d10_37),.data_out(wire_d10_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101039(.data_in(wire_d10_38),.data_out(wire_d10_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101040(.data_in(wire_d10_39),.data_out(wire_d10_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101041(.data_in(wire_d10_40),.data_out(wire_d10_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101042(.data_in(wire_d10_41),.data_out(wire_d10_42),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1101043(.data_in(wire_d10_42),.data_out(wire_d10_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1101044(.data_in(wire_d10_43),.data_out(wire_d10_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1101045(.data_in(wire_d10_44),.data_out(wire_d10_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101046(.data_in(wire_d10_45),.data_out(wire_d10_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101047(.data_in(wire_d10_46),.data_out(wire_d10_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1101048(.data_in(wire_d10_47),.data_out(wire_d10_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101049(.data_in(wire_d10_48),.data_out(wire_d10_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101050(.data_in(wire_d10_49),.data_out(wire_d10_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101051(.data_in(wire_d10_50),.data_out(wire_d10_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101052(.data_in(wire_d10_51),.data_out(wire_d10_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101053(.data_in(wire_d10_52),.data_out(wire_d10_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101054(.data_in(wire_d10_53),.data_out(wire_d10_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101055(.data_in(wire_d10_54),.data_out(wire_d10_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101056(.data_in(wire_d10_55),.data_out(wire_d10_56),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1101057(.data_in(wire_d10_56),.data_out(wire_d10_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101058(.data_in(wire_d10_57),.data_out(wire_d10_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101059(.data_in(wire_d10_58),.data_out(wire_d10_59),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101060(.data_in(wire_d10_59),.data_out(wire_d10_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1101061(.data_in(wire_d10_60),.data_out(wire_d10_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1101062(.data_in(wire_d10_61),.data_out(wire_d10_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101063(.data_in(wire_d10_62),.data_out(wire_d10_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1101064(.data_in(wire_d10_63),.data_out(wire_d10_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1101065(.data_in(wire_d10_64),.data_out(wire_d10_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101066(.data_in(wire_d10_65),.data_out(wire_d10_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101067(.data_in(wire_d10_66),.data_out(wire_d10_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101068(.data_in(wire_d10_67),.data_out(wire_d10_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1101069(.data_in(wire_d10_68),.data_out(wire_d10_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101070(.data_in(wire_d10_69),.data_out(wire_d10_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1101071(.data_in(wire_d10_70),.data_out(wire_d10_71),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101072(.data_in(wire_d10_71),.data_out(wire_d10_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101073(.data_in(wire_d10_72),.data_out(wire_d10_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101074(.data_in(wire_d10_73),.data_out(wire_d10_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1101075(.data_in(wire_d10_74),.data_out(wire_d10_75),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1101076(.data_in(wire_d10_75),.data_out(wire_d10_76),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1101077(.data_in(wire_d10_76),.data_out(wire_d10_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1101078(.data_in(wire_d10_77),.data_out(wire_d10_78),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1101079(.data_in(wire_d10_78),.data_out(wire_d10_79),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101080(.data_in(wire_d10_79),.data_out(wire_d10_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1101081(.data_in(wire_d10_80),.data_out(wire_d10_81),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101082(.data_in(wire_d10_81),.data_out(wire_d10_82),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101083(.data_in(wire_d10_82),.data_out(wire_d10_83),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101084(.data_in(wire_d10_83),.data_out(wire_d10_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1101085(.data_in(wire_d10_84),.data_out(wire_d10_85),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101086(.data_in(wire_d10_85),.data_out(wire_d10_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1101087(.data_in(wire_d10_86),.data_out(wire_d10_87),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101088(.data_in(wire_d10_87),.data_out(wire_d10_88),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101089(.data_in(wire_d10_88),.data_out(wire_d10_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1101090(.data_in(wire_d10_89),.data_out(wire_d10_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1101091(.data_in(wire_d10_90),.data_out(wire_d10_91),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1101092(.data_in(wire_d10_91),.data_out(wire_d10_92),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101093(.data_in(wire_d10_92),.data_out(wire_d10_93),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101094(.data_in(wire_d10_93),.data_out(wire_d10_94),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101095(.data_in(wire_d10_94),.data_out(wire_d10_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1101096(.data_in(wire_d10_95),.data_out(wire_d10_96),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101097(.data_in(wire_d10_96),.data_out(wire_d10_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1101098(.data_in(wire_d10_97),.data_out(wire_d10_98),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101099(.data_in(wire_d10_98),.data_out(wire_d10_99),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance11010100(.data_in(wire_d10_99),.data_out(wire_d10_100),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance11010101(.data_in(wire_d10_100),.data_out(wire_d10_101),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance11010102(.data_in(wire_d10_101),.data_out(wire_d10_102),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance11010103(.data_in(wire_d10_102),.data_out(wire_d10_103),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance11010104(.data_in(wire_d10_103),.data_out(wire_d10_104),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance11010105(.data_in(wire_d10_104),.data_out(wire_d10_105),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance11010106(.data_in(wire_d10_105),.data_out(wire_d10_106),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance11010107(.data_in(wire_d10_106),.data_out(wire_d10_107),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance11010108(.data_in(wire_d10_107),.data_out(wire_d10_108),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance11010109(.data_in(wire_d10_108),.data_out(wire_d10_109),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance11010110(.data_in(wire_d10_109),.data_out(wire_d10_110),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance11010111(.data_in(wire_d10_110),.data_out(wire_d10_111),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance11010112(.data_in(wire_d10_111),.data_out(wire_d10_112),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance11010113(.data_in(wire_d10_112),.data_out(wire_d10_113),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance11010114(.data_in(wire_d10_113),.data_out(wire_d10_114),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance11010115(.data_in(wire_d10_114),.data_out(wire_d10_115),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance11010116(.data_in(wire_d10_115),.data_out(wire_d10_116),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance11010117(.data_in(wire_d10_116),.data_out(wire_d10_117),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance11010118(.data_in(wire_d10_117),.data_out(wire_d10_118),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance11010119(.data_in(wire_d10_118),.data_out(d_out10),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance120110(.data_in(d_in11),.data_out(wire_d11_0),.clk(clk),.rst(rst));            //channel 12
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance120111(.data_in(wire_d11_0),.data_out(wire_d11_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance120112(.data_in(wire_d11_1),.data_out(wire_d11_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance120113(.data_in(wire_d11_2),.data_out(wire_d11_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance120114(.data_in(wire_d11_3),.data_out(wire_d11_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance120115(.data_in(wire_d11_4),.data_out(wire_d11_5),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance120116(.data_in(wire_d11_5),.data_out(wire_d11_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance120117(.data_in(wire_d11_6),.data_out(wire_d11_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance120118(.data_in(wire_d11_7),.data_out(wire_d11_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance120119(.data_in(wire_d11_8),.data_out(wire_d11_9),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201110(.data_in(wire_d11_9),.data_out(wire_d11_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1201111(.data_in(wire_d11_10),.data_out(wire_d11_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1201112(.data_in(wire_d11_11),.data_out(wire_d11_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201113(.data_in(wire_d11_12),.data_out(wire_d11_13),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201114(.data_in(wire_d11_13),.data_out(wire_d11_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201115(.data_in(wire_d11_14),.data_out(wire_d11_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1201116(.data_in(wire_d11_15),.data_out(wire_d11_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1201117(.data_in(wire_d11_16),.data_out(wire_d11_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1201118(.data_in(wire_d11_17),.data_out(wire_d11_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201119(.data_in(wire_d11_18),.data_out(wire_d11_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201120(.data_in(wire_d11_19),.data_out(wire_d11_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201121(.data_in(wire_d11_20),.data_out(wire_d11_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201122(.data_in(wire_d11_21),.data_out(wire_d11_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201123(.data_in(wire_d11_22),.data_out(wire_d11_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201124(.data_in(wire_d11_23),.data_out(wire_d11_24),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1201125(.data_in(wire_d11_24),.data_out(wire_d11_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201126(.data_in(wire_d11_25),.data_out(wire_d11_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201127(.data_in(wire_d11_26),.data_out(wire_d11_27),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1201128(.data_in(wire_d11_27),.data_out(wire_d11_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1201129(.data_in(wire_d11_28),.data_out(wire_d11_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201130(.data_in(wire_d11_29),.data_out(wire_d11_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1201131(.data_in(wire_d11_30),.data_out(wire_d11_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201132(.data_in(wire_d11_31),.data_out(wire_d11_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201133(.data_in(wire_d11_32),.data_out(wire_d11_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1201134(.data_in(wire_d11_33),.data_out(wire_d11_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201135(.data_in(wire_d11_34),.data_out(wire_d11_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201136(.data_in(wire_d11_35),.data_out(wire_d11_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201137(.data_in(wire_d11_36),.data_out(wire_d11_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1201138(.data_in(wire_d11_37),.data_out(wire_d11_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201139(.data_in(wire_d11_38),.data_out(wire_d11_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201140(.data_in(wire_d11_39),.data_out(wire_d11_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201141(.data_in(wire_d11_40),.data_out(wire_d11_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201142(.data_in(wire_d11_41),.data_out(wire_d11_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201143(.data_in(wire_d11_42),.data_out(wire_d11_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201144(.data_in(wire_d11_43),.data_out(wire_d11_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201145(.data_in(wire_d11_44),.data_out(wire_d11_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201146(.data_in(wire_d11_45),.data_out(wire_d11_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201147(.data_in(wire_d11_46),.data_out(wire_d11_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1201148(.data_in(wire_d11_47),.data_out(wire_d11_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201149(.data_in(wire_d11_48),.data_out(wire_d11_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201150(.data_in(wire_d11_49),.data_out(wire_d11_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201151(.data_in(wire_d11_50),.data_out(wire_d11_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201152(.data_in(wire_d11_51),.data_out(wire_d11_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1201153(.data_in(wire_d11_52),.data_out(wire_d11_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201154(.data_in(wire_d11_53),.data_out(wire_d11_54),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1201155(.data_in(wire_d11_54),.data_out(wire_d11_55),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1201156(.data_in(wire_d11_55),.data_out(wire_d11_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201157(.data_in(wire_d11_56),.data_out(wire_d11_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201158(.data_in(wire_d11_57),.data_out(wire_d11_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1201159(.data_in(wire_d11_58),.data_out(wire_d11_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201160(.data_in(wire_d11_59),.data_out(wire_d11_60),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201161(.data_in(wire_d11_60),.data_out(wire_d11_61),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201162(.data_in(wire_d11_61),.data_out(wire_d11_62),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201163(.data_in(wire_d11_62),.data_out(wire_d11_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1201164(.data_in(wire_d11_63),.data_out(wire_d11_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1201165(.data_in(wire_d11_64),.data_out(wire_d11_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201166(.data_in(wire_d11_65),.data_out(wire_d11_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201167(.data_in(wire_d11_66),.data_out(wire_d11_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201168(.data_in(wire_d11_67),.data_out(wire_d11_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201169(.data_in(wire_d11_68),.data_out(wire_d11_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1201170(.data_in(wire_d11_69),.data_out(wire_d11_70),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201171(.data_in(wire_d11_70),.data_out(wire_d11_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1201172(.data_in(wire_d11_71),.data_out(wire_d11_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201173(.data_in(wire_d11_72),.data_out(wire_d11_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201174(.data_in(wire_d11_73),.data_out(wire_d11_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201175(.data_in(wire_d11_74),.data_out(wire_d11_75),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1201176(.data_in(wire_d11_75),.data_out(wire_d11_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201177(.data_in(wire_d11_76),.data_out(wire_d11_77),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201178(.data_in(wire_d11_77),.data_out(wire_d11_78),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201179(.data_in(wire_d11_78),.data_out(wire_d11_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1201180(.data_in(wire_d11_79),.data_out(wire_d11_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201181(.data_in(wire_d11_80),.data_out(wire_d11_81),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1201182(.data_in(wire_d11_81),.data_out(wire_d11_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1201183(.data_in(wire_d11_82),.data_out(wire_d11_83),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201184(.data_in(wire_d11_83),.data_out(wire_d11_84),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201185(.data_in(wire_d11_84),.data_out(wire_d11_85),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201186(.data_in(wire_d11_85),.data_out(wire_d11_86),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201187(.data_in(wire_d11_86),.data_out(wire_d11_87),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1201188(.data_in(wire_d11_87),.data_out(wire_d11_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201189(.data_in(wire_d11_88),.data_out(wire_d11_89),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1201190(.data_in(wire_d11_89),.data_out(wire_d11_90),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201191(.data_in(wire_d11_90),.data_out(wire_d11_91),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1201192(.data_in(wire_d11_91),.data_out(wire_d11_92),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201193(.data_in(wire_d11_92),.data_out(wire_d11_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201194(.data_in(wire_d11_93),.data_out(wire_d11_94),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1201195(.data_in(wire_d11_94),.data_out(wire_d11_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1201196(.data_in(wire_d11_95),.data_out(wire_d11_96),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1201197(.data_in(wire_d11_96),.data_out(wire_d11_97),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201198(.data_in(wire_d11_97),.data_out(wire_d11_98),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201199(.data_in(wire_d11_98),.data_out(wire_d11_99),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance12011100(.data_in(wire_d11_99),.data_out(wire_d11_100),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance12011101(.data_in(wire_d11_100),.data_out(wire_d11_101),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance12011102(.data_in(wire_d11_101),.data_out(wire_d11_102),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance12011103(.data_in(wire_d11_102),.data_out(wire_d11_103),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance12011104(.data_in(wire_d11_103),.data_out(wire_d11_104),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance12011105(.data_in(wire_d11_104),.data_out(wire_d11_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance12011106(.data_in(wire_d11_105),.data_out(wire_d11_106),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance12011107(.data_in(wire_d11_106),.data_out(wire_d11_107),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance12011108(.data_in(wire_d11_107),.data_out(wire_d11_108),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance12011109(.data_in(wire_d11_108),.data_out(wire_d11_109),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance12011110(.data_in(wire_d11_109),.data_out(wire_d11_110),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance12011111(.data_in(wire_d11_110),.data_out(wire_d11_111),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance12011112(.data_in(wire_d11_111),.data_out(wire_d11_112),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance12011113(.data_in(wire_d11_112),.data_out(wire_d11_113),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance12011114(.data_in(wire_d11_113),.data_out(wire_d11_114),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance12011115(.data_in(wire_d11_114),.data_out(wire_d11_115),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance12011116(.data_in(wire_d11_115),.data_out(wire_d11_116),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance12011117(.data_in(wire_d11_116),.data_out(wire_d11_117),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance12011118(.data_in(wire_d11_117),.data_out(wire_d11_118),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance12011119(.data_in(wire_d11_118),.data_out(d_out11),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance130120(.data_in(d_in12),.data_out(wire_d12_0),.clk(clk),.rst(rst));            //channel 13
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance130121(.data_in(wire_d12_0),.data_out(wire_d12_1),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance130122(.data_in(wire_d12_1),.data_out(wire_d12_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance130123(.data_in(wire_d12_2),.data_out(wire_d12_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance130124(.data_in(wire_d12_3),.data_out(wire_d12_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance130125(.data_in(wire_d12_4),.data_out(wire_d12_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance130126(.data_in(wire_d12_5),.data_out(wire_d12_6),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance130127(.data_in(wire_d12_6),.data_out(wire_d12_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance130128(.data_in(wire_d12_7),.data_out(wire_d12_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance130129(.data_in(wire_d12_8),.data_out(wire_d12_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301210(.data_in(wire_d12_9),.data_out(wire_d12_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301211(.data_in(wire_d12_10),.data_out(wire_d12_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301212(.data_in(wire_d12_11),.data_out(wire_d12_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1301213(.data_in(wire_d12_12),.data_out(wire_d12_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301214(.data_in(wire_d12_13),.data_out(wire_d12_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301215(.data_in(wire_d12_14),.data_out(wire_d12_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301216(.data_in(wire_d12_15),.data_out(wire_d12_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301217(.data_in(wire_d12_16),.data_out(wire_d12_17),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1301218(.data_in(wire_d12_17),.data_out(wire_d12_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301219(.data_in(wire_d12_18),.data_out(wire_d12_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301220(.data_in(wire_d12_19),.data_out(wire_d12_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301221(.data_in(wire_d12_20),.data_out(wire_d12_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1301222(.data_in(wire_d12_21),.data_out(wire_d12_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301223(.data_in(wire_d12_22),.data_out(wire_d12_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1301224(.data_in(wire_d12_23),.data_out(wire_d12_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1301225(.data_in(wire_d12_24),.data_out(wire_d12_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301226(.data_in(wire_d12_25),.data_out(wire_d12_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301227(.data_in(wire_d12_26),.data_out(wire_d12_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301228(.data_in(wire_d12_27),.data_out(wire_d12_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301229(.data_in(wire_d12_28),.data_out(wire_d12_29),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301230(.data_in(wire_d12_29),.data_out(wire_d12_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1301231(.data_in(wire_d12_30),.data_out(wire_d12_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301232(.data_in(wire_d12_31),.data_out(wire_d12_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1301233(.data_in(wire_d12_32),.data_out(wire_d12_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301234(.data_in(wire_d12_33),.data_out(wire_d12_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1301235(.data_in(wire_d12_34),.data_out(wire_d12_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301236(.data_in(wire_d12_35),.data_out(wire_d12_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1301237(.data_in(wire_d12_36),.data_out(wire_d12_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1301238(.data_in(wire_d12_37),.data_out(wire_d12_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301239(.data_in(wire_d12_38),.data_out(wire_d12_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301240(.data_in(wire_d12_39),.data_out(wire_d12_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301241(.data_in(wire_d12_40),.data_out(wire_d12_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1301242(.data_in(wire_d12_41),.data_out(wire_d12_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301243(.data_in(wire_d12_42),.data_out(wire_d12_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301244(.data_in(wire_d12_43),.data_out(wire_d12_44),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301245(.data_in(wire_d12_44),.data_out(wire_d12_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301246(.data_in(wire_d12_45),.data_out(wire_d12_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301247(.data_in(wire_d12_46),.data_out(wire_d12_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301248(.data_in(wire_d12_47),.data_out(wire_d12_48),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1301249(.data_in(wire_d12_48),.data_out(wire_d12_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301250(.data_in(wire_d12_49),.data_out(wire_d12_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301251(.data_in(wire_d12_50),.data_out(wire_d12_51),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1301252(.data_in(wire_d12_51),.data_out(wire_d12_52),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1301253(.data_in(wire_d12_52),.data_out(wire_d12_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301254(.data_in(wire_d12_53),.data_out(wire_d12_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1301255(.data_in(wire_d12_54),.data_out(wire_d12_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1301256(.data_in(wire_d12_55),.data_out(wire_d12_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301257(.data_in(wire_d12_56),.data_out(wire_d12_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301258(.data_in(wire_d12_57),.data_out(wire_d12_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1301259(.data_in(wire_d12_58),.data_out(wire_d12_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1301260(.data_in(wire_d12_59),.data_out(wire_d12_60),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301261(.data_in(wire_d12_60),.data_out(wire_d12_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301262(.data_in(wire_d12_61),.data_out(wire_d12_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1301263(.data_in(wire_d12_62),.data_out(wire_d12_63),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301264(.data_in(wire_d12_63),.data_out(wire_d12_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1301265(.data_in(wire_d12_64),.data_out(wire_d12_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1301266(.data_in(wire_d12_65),.data_out(wire_d12_66),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301267(.data_in(wire_d12_66),.data_out(wire_d12_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301268(.data_in(wire_d12_67),.data_out(wire_d12_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301269(.data_in(wire_d12_68),.data_out(wire_d12_69),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1301270(.data_in(wire_d12_69),.data_out(wire_d12_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301271(.data_in(wire_d12_70),.data_out(wire_d12_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301272(.data_in(wire_d12_71),.data_out(wire_d12_72),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1301273(.data_in(wire_d12_72),.data_out(wire_d12_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301274(.data_in(wire_d12_73),.data_out(wire_d12_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1301275(.data_in(wire_d12_74),.data_out(wire_d12_75),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301276(.data_in(wire_d12_75),.data_out(wire_d12_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301277(.data_in(wire_d12_76),.data_out(wire_d12_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301278(.data_in(wire_d12_77),.data_out(wire_d12_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1301279(.data_in(wire_d12_78),.data_out(wire_d12_79),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301280(.data_in(wire_d12_79),.data_out(wire_d12_80),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301281(.data_in(wire_d12_80),.data_out(wire_d12_81),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301282(.data_in(wire_d12_81),.data_out(wire_d12_82),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301283(.data_in(wire_d12_82),.data_out(wire_d12_83),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301284(.data_in(wire_d12_83),.data_out(wire_d12_84),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1301285(.data_in(wire_d12_84),.data_out(wire_d12_85),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1301286(.data_in(wire_d12_85),.data_out(wire_d12_86),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301287(.data_in(wire_d12_86),.data_out(wire_d12_87),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1301288(.data_in(wire_d12_87),.data_out(wire_d12_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1301289(.data_in(wire_d12_88),.data_out(wire_d12_89),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301290(.data_in(wire_d12_89),.data_out(wire_d12_90),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301291(.data_in(wire_d12_90),.data_out(wire_d12_91),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301292(.data_in(wire_d12_91),.data_out(wire_d12_92),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301293(.data_in(wire_d12_92),.data_out(wire_d12_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1301294(.data_in(wire_d12_93),.data_out(wire_d12_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301295(.data_in(wire_d12_94),.data_out(wire_d12_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1301296(.data_in(wire_d12_95),.data_out(wire_d12_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1301297(.data_in(wire_d12_96),.data_out(wire_d12_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1301298(.data_in(wire_d12_97),.data_out(wire_d12_98),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1301299(.data_in(wire_d12_98),.data_out(wire_d12_99),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance13012100(.data_in(wire_d12_99),.data_out(wire_d12_100),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance13012101(.data_in(wire_d12_100),.data_out(wire_d12_101),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance13012102(.data_in(wire_d12_101),.data_out(wire_d12_102),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance13012103(.data_in(wire_d12_102),.data_out(wire_d12_103),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance13012104(.data_in(wire_d12_103),.data_out(wire_d12_104),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance13012105(.data_in(wire_d12_104),.data_out(wire_d12_105),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance13012106(.data_in(wire_d12_105),.data_out(wire_d12_106),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance13012107(.data_in(wire_d12_106),.data_out(wire_d12_107),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance13012108(.data_in(wire_d12_107),.data_out(wire_d12_108),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance13012109(.data_in(wire_d12_108),.data_out(wire_d12_109),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance13012110(.data_in(wire_d12_109),.data_out(wire_d12_110),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance13012111(.data_in(wire_d12_110),.data_out(wire_d12_111),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance13012112(.data_in(wire_d12_111),.data_out(wire_d12_112),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance13012113(.data_in(wire_d12_112),.data_out(wire_d12_113),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance13012114(.data_in(wire_d12_113),.data_out(wire_d12_114),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance13012115(.data_in(wire_d12_114),.data_out(wire_d12_115),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance13012116(.data_in(wire_d12_115),.data_out(wire_d12_116),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance13012117(.data_in(wire_d12_116),.data_out(wire_d12_117),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance13012118(.data_in(wire_d12_117),.data_out(wire_d12_118),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance13012119(.data_in(wire_d12_118),.data_out(d_out12),.clk(clk),.rst(rst));

	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance140130(.data_in(d_in13),.data_out(wire_d13_0),.clk(clk),.rst(rst));            //channel 14
	decoder_top #(.WIDTH(WIDTH)) decoder_instance140131(.data_in(wire_d13_0),.data_out(wire_d13_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance140132(.data_in(wire_d13_1),.data_out(wire_d13_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance140133(.data_in(wire_d13_2),.data_out(wire_d13_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance140134(.data_in(wire_d13_3),.data_out(wire_d13_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance140135(.data_in(wire_d13_4),.data_out(wire_d13_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance140136(.data_in(wire_d13_5),.data_out(wire_d13_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance140137(.data_in(wire_d13_6),.data_out(wire_d13_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance140138(.data_in(wire_d13_7),.data_out(wire_d13_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance140139(.data_in(wire_d13_8),.data_out(wire_d13_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401310(.data_in(wire_d13_9),.data_out(wire_d13_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401311(.data_in(wire_d13_10),.data_out(wire_d13_11),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1401312(.data_in(wire_d13_11),.data_out(wire_d13_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1401313(.data_in(wire_d13_12),.data_out(wire_d13_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401314(.data_in(wire_d13_13),.data_out(wire_d13_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401315(.data_in(wire_d13_14),.data_out(wire_d13_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401316(.data_in(wire_d13_15),.data_out(wire_d13_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401317(.data_in(wire_d13_16),.data_out(wire_d13_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1401318(.data_in(wire_d13_17),.data_out(wire_d13_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401319(.data_in(wire_d13_18),.data_out(wire_d13_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401320(.data_in(wire_d13_19),.data_out(wire_d13_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401321(.data_in(wire_d13_20),.data_out(wire_d13_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1401322(.data_in(wire_d13_21),.data_out(wire_d13_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401323(.data_in(wire_d13_22),.data_out(wire_d13_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401324(.data_in(wire_d13_23),.data_out(wire_d13_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401325(.data_in(wire_d13_24),.data_out(wire_d13_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401326(.data_in(wire_d13_25),.data_out(wire_d13_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401327(.data_in(wire_d13_26),.data_out(wire_d13_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401328(.data_in(wire_d13_27),.data_out(wire_d13_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401329(.data_in(wire_d13_28),.data_out(wire_d13_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401330(.data_in(wire_d13_29),.data_out(wire_d13_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401331(.data_in(wire_d13_30),.data_out(wire_d13_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401332(.data_in(wire_d13_31),.data_out(wire_d13_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401333(.data_in(wire_d13_32),.data_out(wire_d13_33),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1401334(.data_in(wire_d13_33),.data_out(wire_d13_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401335(.data_in(wire_d13_34),.data_out(wire_d13_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401336(.data_in(wire_d13_35),.data_out(wire_d13_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1401337(.data_in(wire_d13_36),.data_out(wire_d13_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401338(.data_in(wire_d13_37),.data_out(wire_d13_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1401339(.data_in(wire_d13_38),.data_out(wire_d13_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1401340(.data_in(wire_d13_39),.data_out(wire_d13_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1401341(.data_in(wire_d13_40),.data_out(wire_d13_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1401342(.data_in(wire_d13_41),.data_out(wire_d13_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1401343(.data_in(wire_d13_42),.data_out(wire_d13_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401344(.data_in(wire_d13_43),.data_out(wire_d13_44),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1401345(.data_in(wire_d13_44),.data_out(wire_d13_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401346(.data_in(wire_d13_45),.data_out(wire_d13_46),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401347(.data_in(wire_d13_46),.data_out(wire_d13_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401348(.data_in(wire_d13_47),.data_out(wire_d13_48),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1401349(.data_in(wire_d13_48),.data_out(wire_d13_49),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1401350(.data_in(wire_d13_49),.data_out(wire_d13_50),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1401351(.data_in(wire_d13_50),.data_out(wire_d13_51),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1401352(.data_in(wire_d13_51),.data_out(wire_d13_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401353(.data_in(wire_d13_52),.data_out(wire_d13_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401354(.data_in(wire_d13_53),.data_out(wire_d13_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401355(.data_in(wire_d13_54),.data_out(wire_d13_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401356(.data_in(wire_d13_55),.data_out(wire_d13_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1401357(.data_in(wire_d13_56),.data_out(wire_d13_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401358(.data_in(wire_d13_57),.data_out(wire_d13_58),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1401359(.data_in(wire_d13_58),.data_out(wire_d13_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401360(.data_in(wire_d13_59),.data_out(wire_d13_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1401361(.data_in(wire_d13_60),.data_out(wire_d13_61),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1401362(.data_in(wire_d13_61),.data_out(wire_d13_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401363(.data_in(wire_d13_62),.data_out(wire_d13_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401364(.data_in(wire_d13_63),.data_out(wire_d13_64),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1401365(.data_in(wire_d13_64),.data_out(wire_d13_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401366(.data_in(wire_d13_65),.data_out(wire_d13_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401367(.data_in(wire_d13_66),.data_out(wire_d13_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401368(.data_in(wire_d13_67),.data_out(wire_d13_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401369(.data_in(wire_d13_68),.data_out(wire_d13_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401370(.data_in(wire_d13_69),.data_out(wire_d13_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401371(.data_in(wire_d13_70),.data_out(wire_d13_71),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1401372(.data_in(wire_d13_71),.data_out(wire_d13_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401373(.data_in(wire_d13_72),.data_out(wire_d13_73),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401374(.data_in(wire_d13_73),.data_out(wire_d13_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401375(.data_in(wire_d13_74),.data_out(wire_d13_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401376(.data_in(wire_d13_75),.data_out(wire_d13_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1401377(.data_in(wire_d13_76),.data_out(wire_d13_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1401378(.data_in(wire_d13_77),.data_out(wire_d13_78),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401379(.data_in(wire_d13_78),.data_out(wire_d13_79),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1401380(.data_in(wire_d13_79),.data_out(wire_d13_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401381(.data_in(wire_d13_80),.data_out(wire_d13_81),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401382(.data_in(wire_d13_81),.data_out(wire_d13_82),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1401383(.data_in(wire_d13_82),.data_out(wire_d13_83),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401384(.data_in(wire_d13_83),.data_out(wire_d13_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1401385(.data_in(wire_d13_84),.data_out(wire_d13_85),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401386(.data_in(wire_d13_85),.data_out(wire_d13_86),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401387(.data_in(wire_d13_86),.data_out(wire_d13_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401388(.data_in(wire_d13_87),.data_out(wire_d13_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1401389(.data_in(wire_d13_88),.data_out(wire_d13_89),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1401390(.data_in(wire_d13_89),.data_out(wire_d13_90),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401391(.data_in(wire_d13_90),.data_out(wire_d13_91),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401392(.data_in(wire_d13_91),.data_out(wire_d13_92),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401393(.data_in(wire_d13_92),.data_out(wire_d13_93),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401394(.data_in(wire_d13_93),.data_out(wire_d13_94),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401395(.data_in(wire_d13_94),.data_out(wire_d13_95),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1401396(.data_in(wire_d13_95),.data_out(wire_d13_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401397(.data_in(wire_d13_96),.data_out(wire_d13_97),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1401398(.data_in(wire_d13_97),.data_out(wire_d13_98),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401399(.data_in(wire_d13_98),.data_out(wire_d13_99),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance14013100(.data_in(wire_d13_99),.data_out(wire_d13_100),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance14013101(.data_in(wire_d13_100),.data_out(wire_d13_101),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance14013102(.data_in(wire_d13_101),.data_out(wire_d13_102),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance14013103(.data_in(wire_d13_102),.data_out(wire_d13_103),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance14013104(.data_in(wire_d13_103),.data_out(wire_d13_104),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance14013105(.data_in(wire_d13_104),.data_out(wire_d13_105),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance14013106(.data_in(wire_d13_105),.data_out(wire_d13_106),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance14013107(.data_in(wire_d13_106),.data_out(wire_d13_107),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance14013108(.data_in(wire_d13_107),.data_out(wire_d13_108),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance14013109(.data_in(wire_d13_108),.data_out(wire_d13_109),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance14013110(.data_in(wire_d13_109),.data_out(wire_d13_110),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance14013111(.data_in(wire_d13_110),.data_out(wire_d13_111),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance14013112(.data_in(wire_d13_111),.data_out(wire_d13_112),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance14013113(.data_in(wire_d13_112),.data_out(wire_d13_113),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance14013114(.data_in(wire_d13_113),.data_out(wire_d13_114),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance14013115(.data_in(wire_d13_114),.data_out(wire_d13_115),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance14013116(.data_in(wire_d13_115),.data_out(wire_d13_116),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance14013117(.data_in(wire_d13_116),.data_out(wire_d13_117),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance14013118(.data_in(wire_d13_117),.data_out(wire_d13_118),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance14013119(.data_in(wire_d13_118),.data_out(d_out13),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance150140(.data_in(d_in14),.data_out(wire_d14_0),.clk(clk),.rst(rst));            //channel 15
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance150141(.data_in(wire_d14_0),.data_out(wire_d14_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance150142(.data_in(wire_d14_1),.data_out(wire_d14_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance150143(.data_in(wire_d14_2),.data_out(wire_d14_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance150144(.data_in(wire_d14_3),.data_out(wire_d14_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance150145(.data_in(wire_d14_4),.data_out(wire_d14_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance150146(.data_in(wire_d14_5),.data_out(wire_d14_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance150147(.data_in(wire_d14_6),.data_out(wire_d14_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance150148(.data_in(wire_d14_7),.data_out(wire_d14_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance150149(.data_in(wire_d14_8),.data_out(wire_d14_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501410(.data_in(wire_d14_9),.data_out(wire_d14_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1501411(.data_in(wire_d14_10),.data_out(wire_d14_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501412(.data_in(wire_d14_11),.data_out(wire_d14_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501413(.data_in(wire_d14_12),.data_out(wire_d14_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501414(.data_in(wire_d14_13),.data_out(wire_d14_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1501415(.data_in(wire_d14_14),.data_out(wire_d14_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1501416(.data_in(wire_d14_15),.data_out(wire_d14_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1501417(.data_in(wire_d14_16),.data_out(wire_d14_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501418(.data_in(wire_d14_17),.data_out(wire_d14_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1501419(.data_in(wire_d14_18),.data_out(wire_d14_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501420(.data_in(wire_d14_19),.data_out(wire_d14_20),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1501421(.data_in(wire_d14_20),.data_out(wire_d14_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501422(.data_in(wire_d14_21),.data_out(wire_d14_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501423(.data_in(wire_d14_22),.data_out(wire_d14_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1501424(.data_in(wire_d14_23),.data_out(wire_d14_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1501425(.data_in(wire_d14_24),.data_out(wire_d14_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501426(.data_in(wire_d14_25),.data_out(wire_d14_26),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1501427(.data_in(wire_d14_26),.data_out(wire_d14_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501428(.data_in(wire_d14_27),.data_out(wire_d14_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501429(.data_in(wire_d14_28),.data_out(wire_d14_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1501430(.data_in(wire_d14_29),.data_out(wire_d14_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1501431(.data_in(wire_d14_30),.data_out(wire_d14_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501432(.data_in(wire_d14_31),.data_out(wire_d14_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501433(.data_in(wire_d14_32),.data_out(wire_d14_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1501434(.data_in(wire_d14_33),.data_out(wire_d14_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1501435(.data_in(wire_d14_34),.data_out(wire_d14_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501436(.data_in(wire_d14_35),.data_out(wire_d14_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501437(.data_in(wire_d14_36),.data_out(wire_d14_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501438(.data_in(wire_d14_37),.data_out(wire_d14_38),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1501439(.data_in(wire_d14_38),.data_out(wire_d14_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1501440(.data_in(wire_d14_39),.data_out(wire_d14_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501441(.data_in(wire_d14_40),.data_out(wire_d14_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1501442(.data_in(wire_d14_41),.data_out(wire_d14_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501443(.data_in(wire_d14_42),.data_out(wire_d14_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1501444(.data_in(wire_d14_43),.data_out(wire_d14_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1501445(.data_in(wire_d14_44),.data_out(wire_d14_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501446(.data_in(wire_d14_45),.data_out(wire_d14_46),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1501447(.data_in(wire_d14_46),.data_out(wire_d14_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501448(.data_in(wire_d14_47),.data_out(wire_d14_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501449(.data_in(wire_d14_48),.data_out(wire_d14_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1501450(.data_in(wire_d14_49),.data_out(wire_d14_50),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501451(.data_in(wire_d14_50),.data_out(wire_d14_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501452(.data_in(wire_d14_51),.data_out(wire_d14_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1501453(.data_in(wire_d14_52),.data_out(wire_d14_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1501454(.data_in(wire_d14_53),.data_out(wire_d14_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1501455(.data_in(wire_d14_54),.data_out(wire_d14_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1501456(.data_in(wire_d14_55),.data_out(wire_d14_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1501457(.data_in(wire_d14_56),.data_out(wire_d14_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501458(.data_in(wire_d14_57),.data_out(wire_d14_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1501459(.data_in(wire_d14_58),.data_out(wire_d14_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501460(.data_in(wire_d14_59),.data_out(wire_d14_60),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501461(.data_in(wire_d14_60),.data_out(wire_d14_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501462(.data_in(wire_d14_61),.data_out(wire_d14_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1501463(.data_in(wire_d14_62),.data_out(wire_d14_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501464(.data_in(wire_d14_63),.data_out(wire_d14_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501465(.data_in(wire_d14_64),.data_out(wire_d14_65),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1501466(.data_in(wire_d14_65),.data_out(wire_d14_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1501467(.data_in(wire_d14_66),.data_out(wire_d14_67),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1501468(.data_in(wire_d14_67),.data_out(wire_d14_68),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1501469(.data_in(wire_d14_68),.data_out(wire_d14_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501470(.data_in(wire_d14_69),.data_out(wire_d14_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501471(.data_in(wire_d14_70),.data_out(wire_d14_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1501472(.data_in(wire_d14_71),.data_out(wire_d14_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501473(.data_in(wire_d14_72),.data_out(wire_d14_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501474(.data_in(wire_d14_73),.data_out(wire_d14_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1501475(.data_in(wire_d14_74),.data_out(wire_d14_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501476(.data_in(wire_d14_75),.data_out(wire_d14_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1501477(.data_in(wire_d14_76),.data_out(wire_d14_77),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501478(.data_in(wire_d14_77),.data_out(wire_d14_78),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501479(.data_in(wire_d14_78),.data_out(wire_d14_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1501480(.data_in(wire_d14_79),.data_out(wire_d14_80),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1501481(.data_in(wire_d14_80),.data_out(wire_d14_81),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501482(.data_in(wire_d14_81),.data_out(wire_d14_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501483(.data_in(wire_d14_82),.data_out(wire_d14_83),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1501484(.data_in(wire_d14_83),.data_out(wire_d14_84),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1501485(.data_in(wire_d14_84),.data_out(wire_d14_85),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501486(.data_in(wire_d14_85),.data_out(wire_d14_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1501487(.data_in(wire_d14_86),.data_out(wire_d14_87),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501488(.data_in(wire_d14_87),.data_out(wire_d14_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501489(.data_in(wire_d14_88),.data_out(wire_d14_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501490(.data_in(wire_d14_89),.data_out(wire_d14_90),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1501491(.data_in(wire_d14_90),.data_out(wire_d14_91),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1501492(.data_in(wire_d14_91),.data_out(wire_d14_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501493(.data_in(wire_d14_92),.data_out(wire_d14_93),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1501494(.data_in(wire_d14_93),.data_out(wire_d14_94),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1501495(.data_in(wire_d14_94),.data_out(wire_d14_95),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501496(.data_in(wire_d14_95),.data_out(wire_d14_96),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1501497(.data_in(wire_d14_96),.data_out(wire_d14_97),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501498(.data_in(wire_d14_97),.data_out(wire_d14_98),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1501499(.data_in(wire_d14_98),.data_out(wire_d14_99),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance15014100(.data_in(wire_d14_99),.data_out(wire_d14_100),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance15014101(.data_in(wire_d14_100),.data_out(wire_d14_101),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance15014102(.data_in(wire_d14_101),.data_out(wire_d14_102),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance15014103(.data_in(wire_d14_102),.data_out(wire_d14_103),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance15014104(.data_in(wire_d14_103),.data_out(wire_d14_104),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance15014105(.data_in(wire_d14_104),.data_out(wire_d14_105),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance15014106(.data_in(wire_d14_105),.data_out(wire_d14_106),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance15014107(.data_in(wire_d14_106),.data_out(wire_d14_107),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance15014108(.data_in(wire_d14_107),.data_out(wire_d14_108),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance15014109(.data_in(wire_d14_108),.data_out(wire_d14_109),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance15014110(.data_in(wire_d14_109),.data_out(wire_d14_110),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance15014111(.data_in(wire_d14_110),.data_out(wire_d14_111),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance15014112(.data_in(wire_d14_111),.data_out(wire_d14_112),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance15014113(.data_in(wire_d14_112),.data_out(wire_d14_113),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance15014114(.data_in(wire_d14_113),.data_out(wire_d14_114),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance15014115(.data_in(wire_d14_114),.data_out(wire_d14_115),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance15014116(.data_in(wire_d14_115),.data_out(wire_d14_116),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance15014117(.data_in(wire_d14_116),.data_out(wire_d14_117),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance15014118(.data_in(wire_d14_117),.data_out(wire_d14_118),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance15014119(.data_in(wire_d14_118),.data_out(d_out14),.clk(clk),.rst(rst));

	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance160150(.data_in(d_in15),.data_out(wire_d15_0),.clk(clk),.rst(rst));            //channel 16
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance160151(.data_in(wire_d15_0),.data_out(wire_d15_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance160152(.data_in(wire_d15_1),.data_out(wire_d15_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance160153(.data_in(wire_d15_2),.data_out(wire_d15_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance160154(.data_in(wire_d15_3),.data_out(wire_d15_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance160155(.data_in(wire_d15_4),.data_out(wire_d15_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance160156(.data_in(wire_d15_5),.data_out(wire_d15_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance160157(.data_in(wire_d15_6),.data_out(wire_d15_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance160158(.data_in(wire_d15_7),.data_out(wire_d15_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance160159(.data_in(wire_d15_8),.data_out(wire_d15_9),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1601510(.data_in(wire_d15_9),.data_out(wire_d15_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601511(.data_in(wire_d15_10),.data_out(wire_d15_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1601512(.data_in(wire_d15_11),.data_out(wire_d15_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1601513(.data_in(wire_d15_12),.data_out(wire_d15_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601514(.data_in(wire_d15_13),.data_out(wire_d15_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601515(.data_in(wire_d15_14),.data_out(wire_d15_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1601516(.data_in(wire_d15_15),.data_out(wire_d15_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601517(.data_in(wire_d15_16),.data_out(wire_d15_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1601518(.data_in(wire_d15_17),.data_out(wire_d15_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1601519(.data_in(wire_d15_18),.data_out(wire_d15_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601520(.data_in(wire_d15_19),.data_out(wire_d15_20),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601521(.data_in(wire_d15_20),.data_out(wire_d15_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1601522(.data_in(wire_d15_21),.data_out(wire_d15_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1601523(.data_in(wire_d15_22),.data_out(wire_d15_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1601524(.data_in(wire_d15_23),.data_out(wire_d15_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601525(.data_in(wire_d15_24),.data_out(wire_d15_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601526(.data_in(wire_d15_25),.data_out(wire_d15_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601527(.data_in(wire_d15_26),.data_out(wire_d15_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601528(.data_in(wire_d15_27),.data_out(wire_d15_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1601529(.data_in(wire_d15_28),.data_out(wire_d15_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1601530(.data_in(wire_d15_29),.data_out(wire_d15_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1601531(.data_in(wire_d15_30),.data_out(wire_d15_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1601532(.data_in(wire_d15_31),.data_out(wire_d15_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601533(.data_in(wire_d15_32),.data_out(wire_d15_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601534(.data_in(wire_d15_33),.data_out(wire_d15_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601535(.data_in(wire_d15_34),.data_out(wire_d15_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601536(.data_in(wire_d15_35),.data_out(wire_d15_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1601537(.data_in(wire_d15_36),.data_out(wire_d15_37),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1601538(.data_in(wire_d15_37),.data_out(wire_d15_38),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601539(.data_in(wire_d15_38),.data_out(wire_d15_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1601540(.data_in(wire_d15_39),.data_out(wire_d15_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601541(.data_in(wire_d15_40),.data_out(wire_d15_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601542(.data_in(wire_d15_41),.data_out(wire_d15_42),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601543(.data_in(wire_d15_42),.data_out(wire_d15_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601544(.data_in(wire_d15_43),.data_out(wire_d15_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601545(.data_in(wire_d15_44),.data_out(wire_d15_45),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601546(.data_in(wire_d15_45),.data_out(wire_d15_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601547(.data_in(wire_d15_46),.data_out(wire_d15_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601548(.data_in(wire_d15_47),.data_out(wire_d15_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601549(.data_in(wire_d15_48),.data_out(wire_d15_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1601550(.data_in(wire_d15_49),.data_out(wire_d15_50),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1601551(.data_in(wire_d15_50),.data_out(wire_d15_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601552(.data_in(wire_d15_51),.data_out(wire_d15_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1601553(.data_in(wire_d15_52),.data_out(wire_d15_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1601554(.data_in(wire_d15_53),.data_out(wire_d15_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601555(.data_in(wire_d15_54),.data_out(wire_d15_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1601556(.data_in(wire_d15_55),.data_out(wire_d15_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601557(.data_in(wire_d15_56),.data_out(wire_d15_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601558(.data_in(wire_d15_57),.data_out(wire_d15_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1601559(.data_in(wire_d15_58),.data_out(wire_d15_59),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1601560(.data_in(wire_d15_59),.data_out(wire_d15_60),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601561(.data_in(wire_d15_60),.data_out(wire_d15_61),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601562(.data_in(wire_d15_61),.data_out(wire_d15_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601563(.data_in(wire_d15_62),.data_out(wire_d15_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1601564(.data_in(wire_d15_63),.data_out(wire_d15_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601565(.data_in(wire_d15_64),.data_out(wire_d15_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601566(.data_in(wire_d15_65),.data_out(wire_d15_66),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1601567(.data_in(wire_d15_66),.data_out(wire_d15_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601568(.data_in(wire_d15_67),.data_out(wire_d15_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601569(.data_in(wire_d15_68),.data_out(wire_d15_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601570(.data_in(wire_d15_69),.data_out(wire_d15_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1601571(.data_in(wire_d15_70),.data_out(wire_d15_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601572(.data_in(wire_d15_71),.data_out(wire_d15_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601573(.data_in(wire_d15_72),.data_out(wire_d15_73),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601574(.data_in(wire_d15_73),.data_out(wire_d15_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601575(.data_in(wire_d15_74),.data_out(wire_d15_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601576(.data_in(wire_d15_75),.data_out(wire_d15_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1601577(.data_in(wire_d15_76),.data_out(wire_d15_77),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601578(.data_in(wire_d15_77),.data_out(wire_d15_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601579(.data_in(wire_d15_78),.data_out(wire_d15_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601580(.data_in(wire_d15_79),.data_out(wire_d15_80),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601581(.data_in(wire_d15_80),.data_out(wire_d15_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601582(.data_in(wire_d15_81),.data_out(wire_d15_82),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601583(.data_in(wire_d15_82),.data_out(wire_d15_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1601584(.data_in(wire_d15_83),.data_out(wire_d15_84),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1601585(.data_in(wire_d15_84),.data_out(wire_d15_85),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601586(.data_in(wire_d15_85),.data_out(wire_d15_86),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1601587(.data_in(wire_d15_86),.data_out(wire_d15_87),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601588(.data_in(wire_d15_87),.data_out(wire_d15_88),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601589(.data_in(wire_d15_88),.data_out(wire_d15_89),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1601590(.data_in(wire_d15_89),.data_out(wire_d15_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1601591(.data_in(wire_d15_90),.data_out(wire_d15_91),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601592(.data_in(wire_d15_91),.data_out(wire_d15_92),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1601593(.data_in(wire_d15_92),.data_out(wire_d15_93),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1601594(.data_in(wire_d15_93),.data_out(wire_d15_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1601595(.data_in(wire_d15_94),.data_out(wire_d15_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601596(.data_in(wire_d15_95),.data_out(wire_d15_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601597(.data_in(wire_d15_96),.data_out(wire_d15_97),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1601598(.data_in(wire_d15_97),.data_out(wire_d15_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601599(.data_in(wire_d15_98),.data_out(wire_d15_99),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance16015100(.data_in(wire_d15_99),.data_out(wire_d15_100),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance16015101(.data_in(wire_d15_100),.data_out(wire_d15_101),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance16015102(.data_in(wire_d15_101),.data_out(wire_d15_102),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance16015103(.data_in(wire_d15_102),.data_out(wire_d15_103),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance16015104(.data_in(wire_d15_103),.data_out(wire_d15_104),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance16015105(.data_in(wire_d15_104),.data_out(wire_d15_105),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance16015106(.data_in(wire_d15_105),.data_out(wire_d15_106),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance16015107(.data_in(wire_d15_106),.data_out(wire_d15_107),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance16015108(.data_in(wire_d15_107),.data_out(wire_d15_108),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance16015109(.data_in(wire_d15_108),.data_out(wire_d15_109),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance16015110(.data_in(wire_d15_109),.data_out(wire_d15_110),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance16015111(.data_in(wire_d15_110),.data_out(wire_d15_111),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance16015112(.data_in(wire_d15_111),.data_out(wire_d15_112),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance16015113(.data_in(wire_d15_112),.data_out(wire_d15_113),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance16015114(.data_in(wire_d15_113),.data_out(wire_d15_114),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance16015115(.data_in(wire_d15_114),.data_out(wire_d15_115),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance16015116(.data_in(wire_d15_115),.data_out(wire_d15_116),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance16015117(.data_in(wire_d15_116),.data_out(wire_d15_117),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance16015118(.data_in(wire_d15_117),.data_out(wire_d15_118),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance16015119(.data_in(wire_d15_118),.data_out(d_out15),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance170160(.data_in(d_in16),.data_out(wire_d16_0),.clk(clk),.rst(rst));            //channel 17
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance170161(.data_in(wire_d16_0),.data_out(wire_d16_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance170162(.data_in(wire_d16_1),.data_out(wire_d16_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance170163(.data_in(wire_d16_2),.data_out(wire_d16_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance170164(.data_in(wire_d16_3),.data_out(wire_d16_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance170165(.data_in(wire_d16_4),.data_out(wire_d16_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance170166(.data_in(wire_d16_5),.data_out(wire_d16_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance170167(.data_in(wire_d16_6),.data_out(wire_d16_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance170168(.data_in(wire_d16_7),.data_out(wire_d16_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance170169(.data_in(wire_d16_8),.data_out(wire_d16_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701610(.data_in(wire_d16_9),.data_out(wire_d16_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701611(.data_in(wire_d16_10),.data_out(wire_d16_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701612(.data_in(wire_d16_11),.data_out(wire_d16_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701613(.data_in(wire_d16_12),.data_out(wire_d16_13),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1701614(.data_in(wire_d16_13),.data_out(wire_d16_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701615(.data_in(wire_d16_14),.data_out(wire_d16_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1701616(.data_in(wire_d16_15),.data_out(wire_d16_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701617(.data_in(wire_d16_16),.data_out(wire_d16_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701618(.data_in(wire_d16_17),.data_out(wire_d16_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1701619(.data_in(wire_d16_18),.data_out(wire_d16_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701620(.data_in(wire_d16_19),.data_out(wire_d16_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701621(.data_in(wire_d16_20),.data_out(wire_d16_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1701622(.data_in(wire_d16_21),.data_out(wire_d16_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1701623(.data_in(wire_d16_22),.data_out(wire_d16_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1701624(.data_in(wire_d16_23),.data_out(wire_d16_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701625(.data_in(wire_d16_24),.data_out(wire_d16_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1701626(.data_in(wire_d16_25),.data_out(wire_d16_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701627(.data_in(wire_d16_26),.data_out(wire_d16_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701628(.data_in(wire_d16_27),.data_out(wire_d16_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701629(.data_in(wire_d16_28),.data_out(wire_d16_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1701630(.data_in(wire_d16_29),.data_out(wire_d16_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1701631(.data_in(wire_d16_30),.data_out(wire_d16_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1701632(.data_in(wire_d16_31),.data_out(wire_d16_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701633(.data_in(wire_d16_32),.data_out(wire_d16_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701634(.data_in(wire_d16_33),.data_out(wire_d16_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1701635(.data_in(wire_d16_34),.data_out(wire_d16_35),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1701636(.data_in(wire_d16_35),.data_out(wire_d16_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701637(.data_in(wire_d16_36),.data_out(wire_d16_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701638(.data_in(wire_d16_37),.data_out(wire_d16_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701639(.data_in(wire_d16_38),.data_out(wire_d16_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701640(.data_in(wire_d16_39),.data_out(wire_d16_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701641(.data_in(wire_d16_40),.data_out(wire_d16_41),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1701642(.data_in(wire_d16_41),.data_out(wire_d16_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1701643(.data_in(wire_d16_42),.data_out(wire_d16_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1701644(.data_in(wire_d16_43),.data_out(wire_d16_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701645(.data_in(wire_d16_44),.data_out(wire_d16_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701646(.data_in(wire_d16_45),.data_out(wire_d16_46),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1701647(.data_in(wire_d16_46),.data_out(wire_d16_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701648(.data_in(wire_d16_47),.data_out(wire_d16_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701649(.data_in(wire_d16_48),.data_out(wire_d16_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1701650(.data_in(wire_d16_49),.data_out(wire_d16_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701651(.data_in(wire_d16_50),.data_out(wire_d16_51),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1701652(.data_in(wire_d16_51),.data_out(wire_d16_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701653(.data_in(wire_d16_52),.data_out(wire_d16_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1701654(.data_in(wire_d16_53),.data_out(wire_d16_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701655(.data_in(wire_d16_54),.data_out(wire_d16_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1701656(.data_in(wire_d16_55),.data_out(wire_d16_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1701657(.data_in(wire_d16_56),.data_out(wire_d16_57),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1701658(.data_in(wire_d16_57),.data_out(wire_d16_58),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1701659(.data_in(wire_d16_58),.data_out(wire_d16_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701660(.data_in(wire_d16_59),.data_out(wire_d16_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1701661(.data_in(wire_d16_60),.data_out(wire_d16_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701662(.data_in(wire_d16_61),.data_out(wire_d16_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1701663(.data_in(wire_d16_62),.data_out(wire_d16_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701664(.data_in(wire_d16_63),.data_out(wire_d16_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701665(.data_in(wire_d16_64),.data_out(wire_d16_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701666(.data_in(wire_d16_65),.data_out(wire_d16_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701667(.data_in(wire_d16_66),.data_out(wire_d16_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701668(.data_in(wire_d16_67),.data_out(wire_d16_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1701669(.data_in(wire_d16_68),.data_out(wire_d16_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701670(.data_in(wire_d16_69),.data_out(wire_d16_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1701671(.data_in(wire_d16_70),.data_out(wire_d16_71),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701672(.data_in(wire_d16_71),.data_out(wire_d16_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701673(.data_in(wire_d16_72),.data_out(wire_d16_73),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1701674(.data_in(wire_d16_73),.data_out(wire_d16_74),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701675(.data_in(wire_d16_74),.data_out(wire_d16_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701676(.data_in(wire_d16_75),.data_out(wire_d16_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701677(.data_in(wire_d16_76),.data_out(wire_d16_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701678(.data_in(wire_d16_77),.data_out(wire_d16_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701679(.data_in(wire_d16_78),.data_out(wire_d16_79),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1701680(.data_in(wire_d16_79),.data_out(wire_d16_80),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1701681(.data_in(wire_d16_80),.data_out(wire_d16_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1701682(.data_in(wire_d16_81),.data_out(wire_d16_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1701683(.data_in(wire_d16_82),.data_out(wire_d16_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701684(.data_in(wire_d16_83),.data_out(wire_d16_84),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701685(.data_in(wire_d16_84),.data_out(wire_d16_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1701686(.data_in(wire_d16_85),.data_out(wire_d16_86),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1701687(.data_in(wire_d16_86),.data_out(wire_d16_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1701688(.data_in(wire_d16_87),.data_out(wire_d16_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701689(.data_in(wire_d16_88),.data_out(wire_d16_89),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701690(.data_in(wire_d16_89),.data_out(wire_d16_90),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701691(.data_in(wire_d16_90),.data_out(wire_d16_91),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701692(.data_in(wire_d16_91),.data_out(wire_d16_92),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701693(.data_in(wire_d16_92),.data_out(wire_d16_93),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1701694(.data_in(wire_d16_93),.data_out(wire_d16_94),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1701695(.data_in(wire_d16_94),.data_out(wire_d16_95),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701696(.data_in(wire_d16_95),.data_out(wire_d16_96),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701697(.data_in(wire_d16_96),.data_out(wire_d16_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701698(.data_in(wire_d16_97),.data_out(wire_d16_98),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1701699(.data_in(wire_d16_98),.data_out(wire_d16_99),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance17016100(.data_in(wire_d16_99),.data_out(wire_d16_100),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance17016101(.data_in(wire_d16_100),.data_out(wire_d16_101),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance17016102(.data_in(wire_d16_101),.data_out(wire_d16_102),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance17016103(.data_in(wire_d16_102),.data_out(wire_d16_103),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance17016104(.data_in(wire_d16_103),.data_out(wire_d16_104),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance17016105(.data_in(wire_d16_104),.data_out(wire_d16_105),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance17016106(.data_in(wire_d16_105),.data_out(wire_d16_106),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance17016107(.data_in(wire_d16_106),.data_out(wire_d16_107),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance17016108(.data_in(wire_d16_107),.data_out(wire_d16_108),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance17016109(.data_in(wire_d16_108),.data_out(wire_d16_109),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance17016110(.data_in(wire_d16_109),.data_out(wire_d16_110),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance17016111(.data_in(wire_d16_110),.data_out(wire_d16_111),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance17016112(.data_in(wire_d16_111),.data_out(wire_d16_112),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance17016113(.data_in(wire_d16_112),.data_out(wire_d16_113),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance17016114(.data_in(wire_d16_113),.data_out(wire_d16_114),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance17016115(.data_in(wire_d16_114),.data_out(wire_d16_115),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance17016116(.data_in(wire_d16_115),.data_out(wire_d16_116),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance17016117(.data_in(wire_d16_116),.data_out(wire_d16_117),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance17016118(.data_in(wire_d16_117),.data_out(wire_d16_118),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance17016119(.data_in(wire_d16_118),.data_out(d_out16),.clk(clk),.rst(rst));

	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance180170(.data_in(d_in17),.data_out(wire_d17_0),.clk(clk),.rst(rst));            //channel 18
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance180171(.data_in(wire_d17_0),.data_out(wire_d17_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance180172(.data_in(wire_d17_1),.data_out(wire_d17_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance180173(.data_in(wire_d17_2),.data_out(wire_d17_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance180174(.data_in(wire_d17_3),.data_out(wire_d17_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance180175(.data_in(wire_d17_4),.data_out(wire_d17_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance180176(.data_in(wire_d17_5),.data_out(wire_d17_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance180177(.data_in(wire_d17_6),.data_out(wire_d17_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance180178(.data_in(wire_d17_7),.data_out(wire_d17_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance180179(.data_in(wire_d17_8),.data_out(wire_d17_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801710(.data_in(wire_d17_9),.data_out(wire_d17_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801711(.data_in(wire_d17_10),.data_out(wire_d17_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801712(.data_in(wire_d17_11),.data_out(wire_d17_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801713(.data_in(wire_d17_12),.data_out(wire_d17_13),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801714(.data_in(wire_d17_13),.data_out(wire_d17_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801715(.data_in(wire_d17_14),.data_out(wire_d17_15),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1801716(.data_in(wire_d17_15),.data_out(wire_d17_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801717(.data_in(wire_d17_16),.data_out(wire_d17_17),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801718(.data_in(wire_d17_17),.data_out(wire_d17_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801719(.data_in(wire_d17_18),.data_out(wire_d17_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1801720(.data_in(wire_d17_19),.data_out(wire_d17_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801721(.data_in(wire_d17_20),.data_out(wire_d17_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1801722(.data_in(wire_d17_21),.data_out(wire_d17_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801723(.data_in(wire_d17_22),.data_out(wire_d17_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1801724(.data_in(wire_d17_23),.data_out(wire_d17_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801725(.data_in(wire_d17_24),.data_out(wire_d17_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801726(.data_in(wire_d17_25),.data_out(wire_d17_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801727(.data_in(wire_d17_26),.data_out(wire_d17_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1801728(.data_in(wire_d17_27),.data_out(wire_d17_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801729(.data_in(wire_d17_28),.data_out(wire_d17_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801730(.data_in(wire_d17_29),.data_out(wire_d17_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801731(.data_in(wire_d17_30),.data_out(wire_d17_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801732(.data_in(wire_d17_31),.data_out(wire_d17_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801733(.data_in(wire_d17_32),.data_out(wire_d17_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801734(.data_in(wire_d17_33),.data_out(wire_d17_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1801735(.data_in(wire_d17_34),.data_out(wire_d17_35),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1801736(.data_in(wire_d17_35),.data_out(wire_d17_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801737(.data_in(wire_d17_36),.data_out(wire_d17_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801738(.data_in(wire_d17_37),.data_out(wire_d17_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801739(.data_in(wire_d17_38),.data_out(wire_d17_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801740(.data_in(wire_d17_39),.data_out(wire_d17_40),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801741(.data_in(wire_d17_40),.data_out(wire_d17_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801742(.data_in(wire_d17_41),.data_out(wire_d17_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1801743(.data_in(wire_d17_42),.data_out(wire_d17_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801744(.data_in(wire_d17_43),.data_out(wire_d17_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801745(.data_in(wire_d17_44),.data_out(wire_d17_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801746(.data_in(wire_d17_45),.data_out(wire_d17_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801747(.data_in(wire_d17_46),.data_out(wire_d17_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801748(.data_in(wire_d17_47),.data_out(wire_d17_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801749(.data_in(wire_d17_48),.data_out(wire_d17_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801750(.data_in(wire_d17_49),.data_out(wire_d17_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801751(.data_in(wire_d17_50),.data_out(wire_d17_51),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801752(.data_in(wire_d17_51),.data_out(wire_d17_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1801753(.data_in(wire_d17_52),.data_out(wire_d17_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1801754(.data_in(wire_d17_53),.data_out(wire_d17_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1801755(.data_in(wire_d17_54),.data_out(wire_d17_55),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801756(.data_in(wire_d17_55),.data_out(wire_d17_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801757(.data_in(wire_d17_56),.data_out(wire_d17_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801758(.data_in(wire_d17_57),.data_out(wire_d17_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801759(.data_in(wire_d17_58),.data_out(wire_d17_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801760(.data_in(wire_d17_59),.data_out(wire_d17_60),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801761(.data_in(wire_d17_60),.data_out(wire_d17_61),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1801762(.data_in(wire_d17_61),.data_out(wire_d17_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801763(.data_in(wire_d17_62),.data_out(wire_d17_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1801764(.data_in(wire_d17_63),.data_out(wire_d17_64),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801765(.data_in(wire_d17_64),.data_out(wire_d17_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801766(.data_in(wire_d17_65),.data_out(wire_d17_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1801767(.data_in(wire_d17_66),.data_out(wire_d17_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801768(.data_in(wire_d17_67),.data_out(wire_d17_68),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801769(.data_in(wire_d17_68),.data_out(wire_d17_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1801770(.data_in(wire_d17_69),.data_out(wire_d17_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801771(.data_in(wire_d17_70),.data_out(wire_d17_71),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801772(.data_in(wire_d17_71),.data_out(wire_d17_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801773(.data_in(wire_d17_72),.data_out(wire_d17_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1801774(.data_in(wire_d17_73),.data_out(wire_d17_74),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801775(.data_in(wire_d17_74),.data_out(wire_d17_75),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1801776(.data_in(wire_d17_75),.data_out(wire_d17_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801777(.data_in(wire_d17_76),.data_out(wire_d17_77),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1801778(.data_in(wire_d17_77),.data_out(wire_d17_78),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1801779(.data_in(wire_d17_78),.data_out(wire_d17_79),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801780(.data_in(wire_d17_79),.data_out(wire_d17_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1801781(.data_in(wire_d17_80),.data_out(wire_d17_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1801782(.data_in(wire_d17_81),.data_out(wire_d17_82),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801783(.data_in(wire_d17_82),.data_out(wire_d17_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1801784(.data_in(wire_d17_83),.data_out(wire_d17_84),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801785(.data_in(wire_d17_84),.data_out(wire_d17_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1801786(.data_in(wire_d17_85),.data_out(wire_d17_86),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801787(.data_in(wire_d17_86),.data_out(wire_d17_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801788(.data_in(wire_d17_87),.data_out(wire_d17_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1801789(.data_in(wire_d17_88),.data_out(wire_d17_89),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801790(.data_in(wire_d17_89),.data_out(wire_d17_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1801791(.data_in(wire_d17_90),.data_out(wire_d17_91),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801792(.data_in(wire_d17_91),.data_out(wire_d17_92),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801793(.data_in(wire_d17_92),.data_out(wire_d17_93),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801794(.data_in(wire_d17_93),.data_out(wire_d17_94),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1801795(.data_in(wire_d17_94),.data_out(wire_d17_95),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801796(.data_in(wire_d17_95),.data_out(wire_d17_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1801797(.data_in(wire_d17_96),.data_out(wire_d17_97),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801798(.data_in(wire_d17_97),.data_out(wire_d17_98),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801799(.data_in(wire_d17_98),.data_out(wire_d17_99),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance18017100(.data_in(wire_d17_99),.data_out(wire_d17_100),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance18017101(.data_in(wire_d17_100),.data_out(wire_d17_101),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance18017102(.data_in(wire_d17_101),.data_out(wire_d17_102),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance18017103(.data_in(wire_d17_102),.data_out(wire_d17_103),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance18017104(.data_in(wire_d17_103),.data_out(wire_d17_104),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance18017105(.data_in(wire_d17_104),.data_out(wire_d17_105),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance18017106(.data_in(wire_d17_105),.data_out(wire_d17_106),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance18017107(.data_in(wire_d17_106),.data_out(wire_d17_107),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance18017108(.data_in(wire_d17_107),.data_out(wire_d17_108),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance18017109(.data_in(wire_d17_108),.data_out(wire_d17_109),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance18017110(.data_in(wire_d17_109),.data_out(wire_d17_110),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance18017111(.data_in(wire_d17_110),.data_out(wire_d17_111),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance18017112(.data_in(wire_d17_111),.data_out(wire_d17_112),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance18017113(.data_in(wire_d17_112),.data_out(wire_d17_113),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance18017114(.data_in(wire_d17_113),.data_out(wire_d17_114),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance18017115(.data_in(wire_d17_114),.data_out(wire_d17_115),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance18017116(.data_in(wire_d17_115),.data_out(wire_d17_116),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance18017117(.data_in(wire_d17_116),.data_out(wire_d17_117),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance18017118(.data_in(wire_d17_117),.data_out(wire_d17_118),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance18017119(.data_in(wire_d17_118),.data_out(d_out17),.clk(clk),.rst(rst));

	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance190180(.data_in(d_in18),.data_out(wire_d18_0),.clk(clk),.rst(rst));            //channel 19
	decoder_top #(.WIDTH(WIDTH)) decoder_instance190181(.data_in(wire_d18_0),.data_out(wire_d18_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance190182(.data_in(wire_d18_1),.data_out(wire_d18_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance190183(.data_in(wire_d18_2),.data_out(wire_d18_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance190184(.data_in(wire_d18_3),.data_out(wire_d18_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance190185(.data_in(wire_d18_4),.data_out(wire_d18_5),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance190186(.data_in(wire_d18_5),.data_out(wire_d18_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance190187(.data_in(wire_d18_6),.data_out(wire_d18_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance190188(.data_in(wire_d18_7),.data_out(wire_d18_8),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance190189(.data_in(wire_d18_8),.data_out(wire_d18_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901810(.data_in(wire_d18_9),.data_out(wire_d18_10),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1901811(.data_in(wire_d18_10),.data_out(wire_d18_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1901812(.data_in(wire_d18_11),.data_out(wire_d18_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901813(.data_in(wire_d18_12),.data_out(wire_d18_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901814(.data_in(wire_d18_13),.data_out(wire_d18_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901815(.data_in(wire_d18_14),.data_out(wire_d18_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901816(.data_in(wire_d18_15),.data_out(wire_d18_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901817(.data_in(wire_d18_16),.data_out(wire_d18_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1901818(.data_in(wire_d18_17),.data_out(wire_d18_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901819(.data_in(wire_d18_18),.data_out(wire_d18_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901820(.data_in(wire_d18_19),.data_out(wire_d18_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1901821(.data_in(wire_d18_20),.data_out(wire_d18_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901822(.data_in(wire_d18_21),.data_out(wire_d18_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1901823(.data_in(wire_d18_22),.data_out(wire_d18_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1901824(.data_in(wire_d18_23),.data_out(wire_d18_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1901825(.data_in(wire_d18_24),.data_out(wire_d18_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901826(.data_in(wire_d18_25),.data_out(wire_d18_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901827(.data_in(wire_d18_26),.data_out(wire_d18_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901828(.data_in(wire_d18_27),.data_out(wire_d18_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901829(.data_in(wire_d18_28),.data_out(wire_d18_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901830(.data_in(wire_d18_29),.data_out(wire_d18_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1901831(.data_in(wire_d18_30),.data_out(wire_d18_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1901832(.data_in(wire_d18_31),.data_out(wire_d18_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901833(.data_in(wire_d18_32),.data_out(wire_d18_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901834(.data_in(wire_d18_33),.data_out(wire_d18_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901835(.data_in(wire_d18_34),.data_out(wire_d18_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1901836(.data_in(wire_d18_35),.data_out(wire_d18_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901837(.data_in(wire_d18_36),.data_out(wire_d18_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901838(.data_in(wire_d18_37),.data_out(wire_d18_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901839(.data_in(wire_d18_38),.data_out(wire_d18_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901840(.data_in(wire_d18_39),.data_out(wire_d18_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901841(.data_in(wire_d18_40),.data_out(wire_d18_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901842(.data_in(wire_d18_41),.data_out(wire_d18_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901843(.data_in(wire_d18_42),.data_out(wire_d18_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901844(.data_in(wire_d18_43),.data_out(wire_d18_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1901845(.data_in(wire_d18_44),.data_out(wire_d18_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901846(.data_in(wire_d18_45),.data_out(wire_d18_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901847(.data_in(wire_d18_46),.data_out(wire_d18_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1901848(.data_in(wire_d18_47),.data_out(wire_d18_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901849(.data_in(wire_d18_48),.data_out(wire_d18_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901850(.data_in(wire_d18_49),.data_out(wire_d18_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901851(.data_in(wire_d18_50),.data_out(wire_d18_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1901852(.data_in(wire_d18_51),.data_out(wire_d18_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1901853(.data_in(wire_d18_52),.data_out(wire_d18_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901854(.data_in(wire_d18_53),.data_out(wire_d18_54),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1901855(.data_in(wire_d18_54),.data_out(wire_d18_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901856(.data_in(wire_d18_55),.data_out(wire_d18_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901857(.data_in(wire_d18_56),.data_out(wire_d18_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901858(.data_in(wire_d18_57),.data_out(wire_d18_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901859(.data_in(wire_d18_58),.data_out(wire_d18_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901860(.data_in(wire_d18_59),.data_out(wire_d18_60),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1901861(.data_in(wire_d18_60),.data_out(wire_d18_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901862(.data_in(wire_d18_61),.data_out(wire_d18_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901863(.data_in(wire_d18_62),.data_out(wire_d18_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901864(.data_in(wire_d18_63),.data_out(wire_d18_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901865(.data_in(wire_d18_64),.data_out(wire_d18_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901866(.data_in(wire_d18_65),.data_out(wire_d18_66),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1901867(.data_in(wire_d18_66),.data_out(wire_d18_67),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1901868(.data_in(wire_d18_67),.data_out(wire_d18_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1901869(.data_in(wire_d18_68),.data_out(wire_d18_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901870(.data_in(wire_d18_69),.data_out(wire_d18_70),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901871(.data_in(wire_d18_70),.data_out(wire_d18_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901872(.data_in(wire_d18_71),.data_out(wire_d18_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901873(.data_in(wire_d18_72),.data_out(wire_d18_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901874(.data_in(wire_d18_73),.data_out(wire_d18_74),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901875(.data_in(wire_d18_74),.data_out(wire_d18_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1901876(.data_in(wire_d18_75),.data_out(wire_d18_76),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1901877(.data_in(wire_d18_76),.data_out(wire_d18_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901878(.data_in(wire_d18_77),.data_out(wire_d18_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1901879(.data_in(wire_d18_78),.data_out(wire_d18_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1901880(.data_in(wire_d18_79),.data_out(wire_d18_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901881(.data_in(wire_d18_80),.data_out(wire_d18_81),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901882(.data_in(wire_d18_81),.data_out(wire_d18_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1901883(.data_in(wire_d18_82),.data_out(wire_d18_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901884(.data_in(wire_d18_83),.data_out(wire_d18_84),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901885(.data_in(wire_d18_84),.data_out(wire_d18_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901886(.data_in(wire_d18_85),.data_out(wire_d18_86),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901887(.data_in(wire_d18_86),.data_out(wire_d18_87),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901888(.data_in(wire_d18_87),.data_out(wire_d18_88),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901889(.data_in(wire_d18_88),.data_out(wire_d18_89),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1901890(.data_in(wire_d18_89),.data_out(wire_d18_90),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901891(.data_in(wire_d18_90),.data_out(wire_d18_91),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901892(.data_in(wire_d18_91),.data_out(wire_d18_92),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901893(.data_in(wire_d18_92),.data_out(wire_d18_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1901894(.data_in(wire_d18_93),.data_out(wire_d18_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1901895(.data_in(wire_d18_94),.data_out(wire_d18_95),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901896(.data_in(wire_d18_95),.data_out(wire_d18_96),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901897(.data_in(wire_d18_96),.data_out(wire_d18_97),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1901898(.data_in(wire_d18_97),.data_out(wire_d18_98),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901899(.data_in(wire_d18_98),.data_out(wire_d18_99),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance19018100(.data_in(wire_d18_99),.data_out(wire_d18_100),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance19018101(.data_in(wire_d18_100),.data_out(wire_d18_101),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance19018102(.data_in(wire_d18_101),.data_out(wire_d18_102),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance19018103(.data_in(wire_d18_102),.data_out(wire_d18_103),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance19018104(.data_in(wire_d18_103),.data_out(wire_d18_104),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance19018105(.data_in(wire_d18_104),.data_out(wire_d18_105),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance19018106(.data_in(wire_d18_105),.data_out(wire_d18_106),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance19018107(.data_in(wire_d18_106),.data_out(wire_d18_107),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance19018108(.data_in(wire_d18_107),.data_out(wire_d18_108),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance19018109(.data_in(wire_d18_108),.data_out(wire_d18_109),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance19018110(.data_in(wire_d18_109),.data_out(wire_d18_110),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance19018111(.data_in(wire_d18_110),.data_out(wire_d18_111),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance19018112(.data_in(wire_d18_111),.data_out(wire_d18_112),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance19018113(.data_in(wire_d18_112),.data_out(wire_d18_113),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance19018114(.data_in(wire_d18_113),.data_out(wire_d18_114),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance19018115(.data_in(wire_d18_114),.data_out(wire_d18_115),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance19018116(.data_in(wire_d18_115),.data_out(wire_d18_116),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance19018117(.data_in(wire_d18_116),.data_out(wire_d18_117),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance19018118(.data_in(wire_d18_117),.data_out(wire_d18_118),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance19018119(.data_in(wire_d18_118),.data_out(d_out18),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance200190(.data_in(d_in19),.data_out(wire_d19_0),.clk(clk),.rst(rst));            //channel 20
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance200191(.data_in(wire_d19_0),.data_out(wire_d19_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance200192(.data_in(wire_d19_1),.data_out(wire_d19_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance200193(.data_in(wire_d19_2),.data_out(wire_d19_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance200194(.data_in(wire_d19_3),.data_out(wire_d19_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance200195(.data_in(wire_d19_4),.data_out(wire_d19_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance200196(.data_in(wire_d19_5),.data_out(wire_d19_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance200197(.data_in(wire_d19_6),.data_out(wire_d19_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance200198(.data_in(wire_d19_7),.data_out(wire_d19_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance200199(.data_in(wire_d19_8),.data_out(wire_d19_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2001910(.data_in(wire_d19_9),.data_out(wire_d19_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001911(.data_in(wire_d19_10),.data_out(wire_d19_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001912(.data_in(wire_d19_11),.data_out(wire_d19_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001913(.data_in(wire_d19_12),.data_out(wire_d19_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2001914(.data_in(wire_d19_13),.data_out(wire_d19_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001915(.data_in(wire_d19_14),.data_out(wire_d19_15),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2001916(.data_in(wire_d19_15),.data_out(wire_d19_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001917(.data_in(wire_d19_16),.data_out(wire_d19_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2001918(.data_in(wire_d19_17),.data_out(wire_d19_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001919(.data_in(wire_d19_18),.data_out(wire_d19_19),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2001920(.data_in(wire_d19_19),.data_out(wire_d19_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001921(.data_in(wire_d19_20),.data_out(wire_d19_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2001922(.data_in(wire_d19_21),.data_out(wire_d19_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2001923(.data_in(wire_d19_22),.data_out(wire_d19_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001924(.data_in(wire_d19_23),.data_out(wire_d19_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001925(.data_in(wire_d19_24),.data_out(wire_d19_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2001926(.data_in(wire_d19_25),.data_out(wire_d19_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2001927(.data_in(wire_d19_26),.data_out(wire_d19_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001928(.data_in(wire_d19_27),.data_out(wire_d19_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001929(.data_in(wire_d19_28),.data_out(wire_d19_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001930(.data_in(wire_d19_29),.data_out(wire_d19_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001931(.data_in(wire_d19_30),.data_out(wire_d19_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001932(.data_in(wire_d19_31),.data_out(wire_d19_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001933(.data_in(wire_d19_32),.data_out(wire_d19_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2001934(.data_in(wire_d19_33),.data_out(wire_d19_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001935(.data_in(wire_d19_34),.data_out(wire_d19_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2001936(.data_in(wire_d19_35),.data_out(wire_d19_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001937(.data_in(wire_d19_36),.data_out(wire_d19_37),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001938(.data_in(wire_d19_37),.data_out(wire_d19_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2001939(.data_in(wire_d19_38),.data_out(wire_d19_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001940(.data_in(wire_d19_39),.data_out(wire_d19_40),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2001941(.data_in(wire_d19_40),.data_out(wire_d19_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001942(.data_in(wire_d19_41),.data_out(wire_d19_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001943(.data_in(wire_d19_42),.data_out(wire_d19_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2001944(.data_in(wire_d19_43),.data_out(wire_d19_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001945(.data_in(wire_d19_44),.data_out(wire_d19_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2001946(.data_in(wire_d19_45),.data_out(wire_d19_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2001947(.data_in(wire_d19_46),.data_out(wire_d19_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001948(.data_in(wire_d19_47),.data_out(wire_d19_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001949(.data_in(wire_d19_48),.data_out(wire_d19_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001950(.data_in(wire_d19_49),.data_out(wire_d19_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001951(.data_in(wire_d19_50),.data_out(wire_d19_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001952(.data_in(wire_d19_51),.data_out(wire_d19_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001953(.data_in(wire_d19_52),.data_out(wire_d19_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001954(.data_in(wire_d19_53),.data_out(wire_d19_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2001955(.data_in(wire_d19_54),.data_out(wire_d19_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2001956(.data_in(wire_d19_55),.data_out(wire_d19_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001957(.data_in(wire_d19_56),.data_out(wire_d19_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2001958(.data_in(wire_d19_57),.data_out(wire_d19_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001959(.data_in(wire_d19_58),.data_out(wire_d19_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001960(.data_in(wire_d19_59),.data_out(wire_d19_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001961(.data_in(wire_d19_60),.data_out(wire_d19_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001962(.data_in(wire_d19_61),.data_out(wire_d19_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2001963(.data_in(wire_d19_62),.data_out(wire_d19_63),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2001964(.data_in(wire_d19_63),.data_out(wire_d19_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001965(.data_in(wire_d19_64),.data_out(wire_d19_65),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2001966(.data_in(wire_d19_65),.data_out(wire_d19_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2001967(.data_in(wire_d19_66),.data_out(wire_d19_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001968(.data_in(wire_d19_67),.data_out(wire_d19_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2001969(.data_in(wire_d19_68),.data_out(wire_d19_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2001970(.data_in(wire_d19_69),.data_out(wire_d19_70),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001971(.data_in(wire_d19_70),.data_out(wire_d19_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2001972(.data_in(wire_d19_71),.data_out(wire_d19_72),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2001973(.data_in(wire_d19_72),.data_out(wire_d19_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2001974(.data_in(wire_d19_73),.data_out(wire_d19_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2001975(.data_in(wire_d19_74),.data_out(wire_d19_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001976(.data_in(wire_d19_75),.data_out(wire_d19_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2001977(.data_in(wire_d19_76),.data_out(wire_d19_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001978(.data_in(wire_d19_77),.data_out(wire_d19_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2001979(.data_in(wire_d19_78),.data_out(wire_d19_79),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2001980(.data_in(wire_d19_79),.data_out(wire_d19_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001981(.data_in(wire_d19_80),.data_out(wire_d19_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001982(.data_in(wire_d19_81),.data_out(wire_d19_82),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2001983(.data_in(wire_d19_82),.data_out(wire_d19_83),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001984(.data_in(wire_d19_83),.data_out(wire_d19_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2001985(.data_in(wire_d19_84),.data_out(wire_d19_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2001986(.data_in(wire_d19_85),.data_out(wire_d19_86),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001987(.data_in(wire_d19_86),.data_out(wire_d19_87),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001988(.data_in(wire_d19_87),.data_out(wire_d19_88),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001989(.data_in(wire_d19_88),.data_out(wire_d19_89),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2001990(.data_in(wire_d19_89),.data_out(wire_d19_90),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001991(.data_in(wire_d19_90),.data_out(wire_d19_91),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001992(.data_in(wire_d19_91),.data_out(wire_d19_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2001993(.data_in(wire_d19_92),.data_out(wire_d19_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2001994(.data_in(wire_d19_93),.data_out(wire_d19_94),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2001995(.data_in(wire_d19_94),.data_out(wire_d19_95),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001996(.data_in(wire_d19_95),.data_out(wire_d19_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001997(.data_in(wire_d19_96),.data_out(wire_d19_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2001998(.data_in(wire_d19_97),.data_out(wire_d19_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001999(.data_in(wire_d19_98),.data_out(wire_d19_99),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance20019100(.data_in(wire_d19_99),.data_out(wire_d19_100),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance20019101(.data_in(wire_d19_100),.data_out(wire_d19_101),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance20019102(.data_in(wire_d19_101),.data_out(wire_d19_102),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance20019103(.data_in(wire_d19_102),.data_out(wire_d19_103),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance20019104(.data_in(wire_d19_103),.data_out(wire_d19_104),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance20019105(.data_in(wire_d19_104),.data_out(wire_d19_105),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance20019106(.data_in(wire_d19_105),.data_out(wire_d19_106),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance20019107(.data_in(wire_d19_106),.data_out(wire_d19_107),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance20019108(.data_in(wire_d19_107),.data_out(wire_d19_108),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance20019109(.data_in(wire_d19_108),.data_out(wire_d19_109),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance20019110(.data_in(wire_d19_109),.data_out(wire_d19_110),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance20019111(.data_in(wire_d19_110),.data_out(wire_d19_111),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance20019112(.data_in(wire_d19_111),.data_out(wire_d19_112),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance20019113(.data_in(wire_d19_112),.data_out(wire_d19_113),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance20019114(.data_in(wire_d19_113),.data_out(wire_d19_114),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance20019115(.data_in(wire_d19_114),.data_out(wire_d19_115),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance20019116(.data_in(wire_d19_115),.data_out(wire_d19_116),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance20019117(.data_in(wire_d19_116),.data_out(wire_d19_117),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance20019118(.data_in(wire_d19_117),.data_out(wire_d19_118),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance20019119(.data_in(wire_d19_118),.data_out(d_out19),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance210200(.data_in(d_in20),.data_out(wire_d20_0),.clk(clk),.rst(rst));            //channel 21
	large_adder #(.WIDTH(WIDTH)) large_adder_instance210201(.data_in(wire_d20_0),.data_out(wire_d20_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance210202(.data_in(wire_d20_1),.data_out(wire_d20_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance210203(.data_in(wire_d20_2),.data_out(wire_d20_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance210204(.data_in(wire_d20_3),.data_out(wire_d20_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance210205(.data_in(wire_d20_4),.data_out(wire_d20_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance210206(.data_in(wire_d20_5),.data_out(wire_d20_6),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance210207(.data_in(wire_d20_6),.data_out(wire_d20_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance210208(.data_in(wire_d20_7),.data_out(wire_d20_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance210209(.data_in(wire_d20_8),.data_out(wire_d20_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102010(.data_in(wire_d20_9),.data_out(wire_d20_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102011(.data_in(wire_d20_10),.data_out(wire_d20_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102012(.data_in(wire_d20_11),.data_out(wire_d20_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2102013(.data_in(wire_d20_12),.data_out(wire_d20_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2102014(.data_in(wire_d20_13),.data_out(wire_d20_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2102015(.data_in(wire_d20_14),.data_out(wire_d20_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102016(.data_in(wire_d20_15),.data_out(wire_d20_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102017(.data_in(wire_d20_16),.data_out(wire_d20_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102018(.data_in(wire_d20_17),.data_out(wire_d20_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2102019(.data_in(wire_d20_18),.data_out(wire_d20_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102020(.data_in(wire_d20_19),.data_out(wire_d20_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102021(.data_in(wire_d20_20),.data_out(wire_d20_21),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102022(.data_in(wire_d20_21),.data_out(wire_d20_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2102023(.data_in(wire_d20_22),.data_out(wire_d20_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2102024(.data_in(wire_d20_23),.data_out(wire_d20_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2102025(.data_in(wire_d20_24),.data_out(wire_d20_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102026(.data_in(wire_d20_25),.data_out(wire_d20_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102027(.data_in(wire_d20_26),.data_out(wire_d20_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102028(.data_in(wire_d20_27),.data_out(wire_d20_28),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102029(.data_in(wire_d20_28),.data_out(wire_d20_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102030(.data_in(wire_d20_29),.data_out(wire_d20_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102031(.data_in(wire_d20_30),.data_out(wire_d20_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102032(.data_in(wire_d20_31),.data_out(wire_d20_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102033(.data_in(wire_d20_32),.data_out(wire_d20_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102034(.data_in(wire_d20_33),.data_out(wire_d20_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102035(.data_in(wire_d20_34),.data_out(wire_d20_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2102036(.data_in(wire_d20_35),.data_out(wire_d20_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102037(.data_in(wire_d20_36),.data_out(wire_d20_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102038(.data_in(wire_d20_37),.data_out(wire_d20_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102039(.data_in(wire_d20_38),.data_out(wire_d20_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102040(.data_in(wire_d20_39),.data_out(wire_d20_40),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102041(.data_in(wire_d20_40),.data_out(wire_d20_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102042(.data_in(wire_d20_41),.data_out(wire_d20_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2102043(.data_in(wire_d20_42),.data_out(wire_d20_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2102044(.data_in(wire_d20_43),.data_out(wire_d20_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2102045(.data_in(wire_d20_44),.data_out(wire_d20_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2102046(.data_in(wire_d20_45),.data_out(wire_d20_46),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2102047(.data_in(wire_d20_46),.data_out(wire_d20_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102048(.data_in(wire_d20_47),.data_out(wire_d20_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102049(.data_in(wire_d20_48),.data_out(wire_d20_49),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2102050(.data_in(wire_d20_49),.data_out(wire_d20_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102051(.data_in(wire_d20_50),.data_out(wire_d20_51),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2102052(.data_in(wire_d20_51),.data_out(wire_d20_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2102053(.data_in(wire_d20_52),.data_out(wire_d20_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102054(.data_in(wire_d20_53),.data_out(wire_d20_54),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2102055(.data_in(wire_d20_54),.data_out(wire_d20_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2102056(.data_in(wire_d20_55),.data_out(wire_d20_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102057(.data_in(wire_d20_56),.data_out(wire_d20_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102058(.data_in(wire_d20_57),.data_out(wire_d20_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2102059(.data_in(wire_d20_58),.data_out(wire_d20_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2102060(.data_in(wire_d20_59),.data_out(wire_d20_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2102061(.data_in(wire_d20_60),.data_out(wire_d20_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102062(.data_in(wire_d20_61),.data_out(wire_d20_62),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102063(.data_in(wire_d20_62),.data_out(wire_d20_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2102064(.data_in(wire_d20_63),.data_out(wire_d20_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102065(.data_in(wire_d20_64),.data_out(wire_d20_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102066(.data_in(wire_d20_65),.data_out(wire_d20_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102067(.data_in(wire_d20_66),.data_out(wire_d20_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102068(.data_in(wire_d20_67),.data_out(wire_d20_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2102069(.data_in(wire_d20_68),.data_out(wire_d20_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102070(.data_in(wire_d20_69),.data_out(wire_d20_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102071(.data_in(wire_d20_70),.data_out(wire_d20_71),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2102072(.data_in(wire_d20_71),.data_out(wire_d20_72),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102073(.data_in(wire_d20_72),.data_out(wire_d20_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2102074(.data_in(wire_d20_73),.data_out(wire_d20_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2102075(.data_in(wire_d20_74),.data_out(wire_d20_75),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102076(.data_in(wire_d20_75),.data_out(wire_d20_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102077(.data_in(wire_d20_76),.data_out(wire_d20_77),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102078(.data_in(wire_d20_77),.data_out(wire_d20_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102079(.data_in(wire_d20_78),.data_out(wire_d20_79),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2102080(.data_in(wire_d20_79),.data_out(wire_d20_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102081(.data_in(wire_d20_80),.data_out(wire_d20_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2102082(.data_in(wire_d20_81),.data_out(wire_d20_82),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102083(.data_in(wire_d20_82),.data_out(wire_d20_83),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102084(.data_in(wire_d20_83),.data_out(wire_d20_84),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102085(.data_in(wire_d20_84),.data_out(wire_d20_85),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2102086(.data_in(wire_d20_85),.data_out(wire_d20_86),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2102087(.data_in(wire_d20_86),.data_out(wire_d20_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102088(.data_in(wire_d20_87),.data_out(wire_d20_88),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2102089(.data_in(wire_d20_88),.data_out(wire_d20_89),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102090(.data_in(wire_d20_89),.data_out(wire_d20_90),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2102091(.data_in(wire_d20_90),.data_out(wire_d20_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2102092(.data_in(wire_d20_91),.data_out(wire_d20_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102093(.data_in(wire_d20_92),.data_out(wire_d20_93),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2102094(.data_in(wire_d20_93),.data_out(wire_d20_94),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102095(.data_in(wire_d20_94),.data_out(wire_d20_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2102096(.data_in(wire_d20_95),.data_out(wire_d20_96),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2102097(.data_in(wire_d20_96),.data_out(wire_d20_97),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102098(.data_in(wire_d20_97),.data_out(wire_d20_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2102099(.data_in(wire_d20_98),.data_out(wire_d20_99),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance21020100(.data_in(wire_d20_99),.data_out(wire_d20_100),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21020101(.data_in(wire_d20_100),.data_out(wire_d20_101),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance21020102(.data_in(wire_d20_101),.data_out(wire_d20_102),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance21020103(.data_in(wire_d20_102),.data_out(wire_d20_103),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance21020104(.data_in(wire_d20_103),.data_out(wire_d20_104),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance21020105(.data_in(wire_d20_104),.data_out(wire_d20_105),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance21020106(.data_in(wire_d20_105),.data_out(wire_d20_106),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance21020107(.data_in(wire_d20_106),.data_out(wire_d20_107),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance21020108(.data_in(wire_d20_107),.data_out(wire_d20_108),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance21020109(.data_in(wire_d20_108),.data_out(wire_d20_109),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance21020110(.data_in(wire_d20_109),.data_out(wire_d20_110),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance21020111(.data_in(wire_d20_110),.data_out(wire_d20_111),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance21020112(.data_in(wire_d20_111),.data_out(wire_d20_112),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance21020113(.data_in(wire_d20_112),.data_out(wire_d20_113),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance21020114(.data_in(wire_d20_113),.data_out(wire_d20_114),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance21020115(.data_in(wire_d20_114),.data_out(wire_d20_115),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance21020116(.data_in(wire_d20_115),.data_out(wire_d20_116),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance21020117(.data_in(wire_d20_116),.data_out(wire_d20_117),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance21020118(.data_in(wire_d20_117),.data_out(wire_d20_118),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance21020119(.data_in(wire_d20_118),.data_out(d_out20),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance220210(.data_in(d_in21),.data_out(wire_d21_0),.clk(clk),.rst(rst));            //channel 22
	large_mux #(.WIDTH(WIDTH)) large_mux_instance220211(.data_in(wire_d21_0),.data_out(wire_d21_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance220212(.data_in(wire_d21_1),.data_out(wire_d21_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance220213(.data_in(wire_d21_2),.data_out(wire_d21_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance220214(.data_in(wire_d21_3),.data_out(wire_d21_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance220215(.data_in(wire_d21_4),.data_out(wire_d21_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance220216(.data_in(wire_d21_5),.data_out(wire_d21_6),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance220217(.data_in(wire_d21_6),.data_out(wire_d21_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance220218(.data_in(wire_d21_7),.data_out(wire_d21_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance220219(.data_in(wire_d21_8),.data_out(wire_d21_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2202110(.data_in(wire_d21_9),.data_out(wire_d21_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202111(.data_in(wire_d21_10),.data_out(wire_d21_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2202112(.data_in(wire_d21_11),.data_out(wire_d21_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2202113(.data_in(wire_d21_12),.data_out(wire_d21_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2202114(.data_in(wire_d21_13),.data_out(wire_d21_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2202115(.data_in(wire_d21_14),.data_out(wire_d21_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202116(.data_in(wire_d21_15),.data_out(wire_d21_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2202117(.data_in(wire_d21_16),.data_out(wire_d21_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2202118(.data_in(wire_d21_17),.data_out(wire_d21_18),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202119(.data_in(wire_d21_18),.data_out(wire_d21_19),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2202120(.data_in(wire_d21_19),.data_out(wire_d21_20),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2202121(.data_in(wire_d21_20),.data_out(wire_d21_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2202122(.data_in(wire_d21_21),.data_out(wire_d21_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202123(.data_in(wire_d21_22),.data_out(wire_d21_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202124(.data_in(wire_d21_23),.data_out(wire_d21_24),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2202125(.data_in(wire_d21_24),.data_out(wire_d21_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2202126(.data_in(wire_d21_25),.data_out(wire_d21_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2202127(.data_in(wire_d21_26),.data_out(wire_d21_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2202128(.data_in(wire_d21_27),.data_out(wire_d21_28),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202129(.data_in(wire_d21_28),.data_out(wire_d21_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2202130(.data_in(wire_d21_29),.data_out(wire_d21_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2202131(.data_in(wire_d21_30),.data_out(wire_d21_31),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2202132(.data_in(wire_d21_31),.data_out(wire_d21_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2202133(.data_in(wire_d21_32),.data_out(wire_d21_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202134(.data_in(wire_d21_33),.data_out(wire_d21_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202135(.data_in(wire_d21_34),.data_out(wire_d21_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202136(.data_in(wire_d21_35),.data_out(wire_d21_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2202137(.data_in(wire_d21_36),.data_out(wire_d21_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202138(.data_in(wire_d21_37),.data_out(wire_d21_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202139(.data_in(wire_d21_38),.data_out(wire_d21_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202140(.data_in(wire_d21_39),.data_out(wire_d21_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202141(.data_in(wire_d21_40),.data_out(wire_d21_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202142(.data_in(wire_d21_41),.data_out(wire_d21_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202143(.data_in(wire_d21_42),.data_out(wire_d21_43),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202144(.data_in(wire_d21_43),.data_out(wire_d21_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202145(.data_in(wire_d21_44),.data_out(wire_d21_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202146(.data_in(wire_d21_45),.data_out(wire_d21_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2202147(.data_in(wire_d21_46),.data_out(wire_d21_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202148(.data_in(wire_d21_47),.data_out(wire_d21_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2202149(.data_in(wire_d21_48),.data_out(wire_d21_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2202150(.data_in(wire_d21_49),.data_out(wire_d21_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2202151(.data_in(wire_d21_50),.data_out(wire_d21_51),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202152(.data_in(wire_d21_51),.data_out(wire_d21_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202153(.data_in(wire_d21_52),.data_out(wire_d21_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202154(.data_in(wire_d21_53),.data_out(wire_d21_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2202155(.data_in(wire_d21_54),.data_out(wire_d21_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202156(.data_in(wire_d21_55),.data_out(wire_d21_56),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2202157(.data_in(wire_d21_56),.data_out(wire_d21_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2202158(.data_in(wire_d21_57),.data_out(wire_d21_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2202159(.data_in(wire_d21_58),.data_out(wire_d21_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202160(.data_in(wire_d21_59),.data_out(wire_d21_60),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202161(.data_in(wire_d21_60),.data_out(wire_d21_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2202162(.data_in(wire_d21_61),.data_out(wire_d21_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2202163(.data_in(wire_d21_62),.data_out(wire_d21_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2202164(.data_in(wire_d21_63),.data_out(wire_d21_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202165(.data_in(wire_d21_64),.data_out(wire_d21_65),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202166(.data_in(wire_d21_65),.data_out(wire_d21_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2202167(.data_in(wire_d21_66),.data_out(wire_d21_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202168(.data_in(wire_d21_67),.data_out(wire_d21_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202169(.data_in(wire_d21_68),.data_out(wire_d21_69),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202170(.data_in(wire_d21_69),.data_out(wire_d21_70),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202171(.data_in(wire_d21_70),.data_out(wire_d21_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202172(.data_in(wire_d21_71),.data_out(wire_d21_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2202173(.data_in(wire_d21_72),.data_out(wire_d21_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2202174(.data_in(wire_d21_73),.data_out(wire_d21_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2202175(.data_in(wire_d21_74),.data_out(wire_d21_75),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2202176(.data_in(wire_d21_75),.data_out(wire_d21_76),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2202177(.data_in(wire_d21_76),.data_out(wire_d21_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2202178(.data_in(wire_d21_77),.data_out(wire_d21_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202179(.data_in(wire_d21_78),.data_out(wire_d21_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202180(.data_in(wire_d21_79),.data_out(wire_d21_80),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202181(.data_in(wire_d21_80),.data_out(wire_d21_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2202182(.data_in(wire_d21_81),.data_out(wire_d21_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202183(.data_in(wire_d21_82),.data_out(wire_d21_83),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202184(.data_in(wire_d21_83),.data_out(wire_d21_84),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2202185(.data_in(wire_d21_84),.data_out(wire_d21_85),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202186(.data_in(wire_d21_85),.data_out(wire_d21_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2202187(.data_in(wire_d21_86),.data_out(wire_d21_87),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202188(.data_in(wire_d21_87),.data_out(wire_d21_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202189(.data_in(wire_d21_88),.data_out(wire_d21_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2202190(.data_in(wire_d21_89),.data_out(wire_d21_90),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202191(.data_in(wire_d21_90),.data_out(wire_d21_91),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202192(.data_in(wire_d21_91),.data_out(wire_d21_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2202193(.data_in(wire_d21_92),.data_out(wire_d21_93),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202194(.data_in(wire_d21_93),.data_out(wire_d21_94),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202195(.data_in(wire_d21_94),.data_out(wire_d21_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2202196(.data_in(wire_d21_95),.data_out(wire_d21_96),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202197(.data_in(wire_d21_96),.data_out(wire_d21_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2202198(.data_in(wire_d21_97),.data_out(wire_d21_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202199(.data_in(wire_d21_98),.data_out(wire_d21_99),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance22021100(.data_in(wire_d21_99),.data_out(wire_d21_100),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance22021101(.data_in(wire_d21_100),.data_out(wire_d21_101),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance22021102(.data_in(wire_d21_101),.data_out(wire_d21_102),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance22021103(.data_in(wire_d21_102),.data_out(wire_d21_103),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance22021104(.data_in(wire_d21_103),.data_out(wire_d21_104),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance22021105(.data_in(wire_d21_104),.data_out(wire_d21_105),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance22021106(.data_in(wire_d21_105),.data_out(wire_d21_106),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance22021107(.data_in(wire_d21_106),.data_out(wire_d21_107),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance22021108(.data_in(wire_d21_107),.data_out(wire_d21_108),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance22021109(.data_in(wire_d21_108),.data_out(wire_d21_109),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance22021110(.data_in(wire_d21_109),.data_out(wire_d21_110),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance22021111(.data_in(wire_d21_110),.data_out(wire_d21_111),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance22021112(.data_in(wire_d21_111),.data_out(wire_d21_112),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance22021113(.data_in(wire_d21_112),.data_out(wire_d21_113),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance22021114(.data_in(wire_d21_113),.data_out(wire_d21_114),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance22021115(.data_in(wire_d21_114),.data_out(wire_d21_115),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance22021116(.data_in(wire_d21_115),.data_out(wire_d21_116),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance22021117(.data_in(wire_d21_116),.data_out(wire_d21_117),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance22021118(.data_in(wire_d21_117),.data_out(wire_d21_118),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance22021119(.data_in(wire_d21_118),.data_out(d_out21),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance230220(.data_in(d_in22),.data_out(wire_d22_0),.clk(clk),.rst(rst));            //channel 23
	register #(.WIDTH(WIDTH)) register_instance230221(.data_in(wire_d22_0),.data_out(wire_d22_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance230222(.data_in(wire_d22_1),.data_out(wire_d22_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance230223(.data_in(wire_d22_2),.data_out(wire_d22_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance230224(.data_in(wire_d22_3),.data_out(wire_d22_4),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance230225(.data_in(wire_d22_4),.data_out(wire_d22_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance230226(.data_in(wire_d22_5),.data_out(wire_d22_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance230227(.data_in(wire_d22_6),.data_out(wire_d22_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance230228(.data_in(wire_d22_7),.data_out(wire_d22_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance230229(.data_in(wire_d22_8),.data_out(wire_d22_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302210(.data_in(wire_d22_9),.data_out(wire_d22_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302211(.data_in(wire_d22_10),.data_out(wire_d22_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302212(.data_in(wire_d22_11),.data_out(wire_d22_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302213(.data_in(wire_d22_12),.data_out(wire_d22_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302214(.data_in(wire_d22_13),.data_out(wire_d22_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2302215(.data_in(wire_d22_14),.data_out(wire_d22_15),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2302216(.data_in(wire_d22_15),.data_out(wire_d22_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302217(.data_in(wire_d22_16),.data_out(wire_d22_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302218(.data_in(wire_d22_17),.data_out(wire_d22_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2302219(.data_in(wire_d22_18),.data_out(wire_d22_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302220(.data_in(wire_d22_19),.data_out(wire_d22_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302221(.data_in(wire_d22_20),.data_out(wire_d22_21),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2302222(.data_in(wire_d22_21),.data_out(wire_d22_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2302223(.data_in(wire_d22_22),.data_out(wire_d22_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302224(.data_in(wire_d22_23),.data_out(wire_d22_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2302225(.data_in(wire_d22_24),.data_out(wire_d22_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302226(.data_in(wire_d22_25),.data_out(wire_d22_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302227(.data_in(wire_d22_26),.data_out(wire_d22_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302228(.data_in(wire_d22_27),.data_out(wire_d22_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2302229(.data_in(wire_d22_28),.data_out(wire_d22_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302230(.data_in(wire_d22_29),.data_out(wire_d22_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302231(.data_in(wire_d22_30),.data_out(wire_d22_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302232(.data_in(wire_d22_31),.data_out(wire_d22_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302233(.data_in(wire_d22_32),.data_out(wire_d22_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302234(.data_in(wire_d22_33),.data_out(wire_d22_34),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2302235(.data_in(wire_d22_34),.data_out(wire_d22_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302236(.data_in(wire_d22_35),.data_out(wire_d22_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302237(.data_in(wire_d22_36),.data_out(wire_d22_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302238(.data_in(wire_d22_37),.data_out(wire_d22_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2302239(.data_in(wire_d22_38),.data_out(wire_d22_39),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2302240(.data_in(wire_d22_39),.data_out(wire_d22_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2302241(.data_in(wire_d22_40),.data_out(wire_d22_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302242(.data_in(wire_d22_41),.data_out(wire_d22_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302243(.data_in(wire_d22_42),.data_out(wire_d22_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302244(.data_in(wire_d22_43),.data_out(wire_d22_44),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302245(.data_in(wire_d22_44),.data_out(wire_d22_45),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2302246(.data_in(wire_d22_45),.data_out(wire_d22_46),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2302247(.data_in(wire_d22_46),.data_out(wire_d22_47),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302248(.data_in(wire_d22_47),.data_out(wire_d22_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2302249(.data_in(wire_d22_48),.data_out(wire_d22_49),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302250(.data_in(wire_d22_49),.data_out(wire_d22_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2302251(.data_in(wire_d22_50),.data_out(wire_d22_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302252(.data_in(wire_d22_51),.data_out(wire_d22_52),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2302253(.data_in(wire_d22_52),.data_out(wire_d22_53),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2302254(.data_in(wire_d22_53),.data_out(wire_d22_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2302255(.data_in(wire_d22_54),.data_out(wire_d22_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302256(.data_in(wire_d22_55),.data_out(wire_d22_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302257(.data_in(wire_d22_56),.data_out(wire_d22_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302258(.data_in(wire_d22_57),.data_out(wire_d22_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302259(.data_in(wire_d22_58),.data_out(wire_d22_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2302260(.data_in(wire_d22_59),.data_out(wire_d22_60),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302261(.data_in(wire_d22_60),.data_out(wire_d22_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302262(.data_in(wire_d22_61),.data_out(wire_d22_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302263(.data_in(wire_d22_62),.data_out(wire_d22_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302264(.data_in(wire_d22_63),.data_out(wire_d22_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302265(.data_in(wire_d22_64),.data_out(wire_d22_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302266(.data_in(wire_d22_65),.data_out(wire_d22_66),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302267(.data_in(wire_d22_66),.data_out(wire_d22_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302268(.data_in(wire_d22_67),.data_out(wire_d22_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302269(.data_in(wire_d22_68),.data_out(wire_d22_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2302270(.data_in(wire_d22_69),.data_out(wire_d22_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2302271(.data_in(wire_d22_70),.data_out(wire_d22_71),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302272(.data_in(wire_d22_71),.data_out(wire_d22_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2302273(.data_in(wire_d22_72),.data_out(wire_d22_73),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302274(.data_in(wire_d22_73),.data_out(wire_d22_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302275(.data_in(wire_d22_74),.data_out(wire_d22_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2302276(.data_in(wire_d22_75),.data_out(wire_d22_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302277(.data_in(wire_d22_76),.data_out(wire_d22_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302278(.data_in(wire_d22_77),.data_out(wire_d22_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2302279(.data_in(wire_d22_78),.data_out(wire_d22_79),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302280(.data_in(wire_d22_79),.data_out(wire_d22_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302281(.data_in(wire_d22_80),.data_out(wire_d22_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2302282(.data_in(wire_d22_81),.data_out(wire_d22_82),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302283(.data_in(wire_d22_82),.data_out(wire_d22_83),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302284(.data_in(wire_d22_83),.data_out(wire_d22_84),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302285(.data_in(wire_d22_84),.data_out(wire_d22_85),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302286(.data_in(wire_d22_85),.data_out(wire_d22_86),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302287(.data_in(wire_d22_86),.data_out(wire_d22_87),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2302288(.data_in(wire_d22_87),.data_out(wire_d22_88),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302289(.data_in(wire_d22_88),.data_out(wire_d22_89),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302290(.data_in(wire_d22_89),.data_out(wire_d22_90),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302291(.data_in(wire_d22_90),.data_out(wire_d22_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302292(.data_in(wire_d22_91),.data_out(wire_d22_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2302293(.data_in(wire_d22_92),.data_out(wire_d22_93),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302294(.data_in(wire_d22_93),.data_out(wire_d22_94),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2302295(.data_in(wire_d22_94),.data_out(wire_d22_95),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2302296(.data_in(wire_d22_95),.data_out(wire_d22_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2302297(.data_in(wire_d22_96),.data_out(wire_d22_97),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302298(.data_in(wire_d22_97),.data_out(wire_d22_98),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302299(.data_in(wire_d22_98),.data_out(wire_d22_99),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance23022100(.data_in(wire_d22_99),.data_out(wire_d22_100),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance23022101(.data_in(wire_d22_100),.data_out(wire_d22_101),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance23022102(.data_in(wire_d22_101),.data_out(wire_d22_102),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance23022103(.data_in(wire_d22_102),.data_out(wire_d22_103),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance23022104(.data_in(wire_d22_103),.data_out(wire_d22_104),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance23022105(.data_in(wire_d22_104),.data_out(wire_d22_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance23022106(.data_in(wire_d22_105),.data_out(wire_d22_106),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance23022107(.data_in(wire_d22_106),.data_out(wire_d22_107),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance23022108(.data_in(wire_d22_107),.data_out(wire_d22_108),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance23022109(.data_in(wire_d22_108),.data_out(wire_d22_109),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance23022110(.data_in(wire_d22_109),.data_out(wire_d22_110),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance23022111(.data_in(wire_d22_110),.data_out(wire_d22_111),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance23022112(.data_in(wire_d22_111),.data_out(wire_d22_112),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance23022113(.data_in(wire_d22_112),.data_out(wire_d22_113),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance23022114(.data_in(wire_d22_113),.data_out(wire_d22_114),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance23022115(.data_in(wire_d22_114),.data_out(wire_d22_115),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance23022116(.data_in(wire_d22_115),.data_out(wire_d22_116),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance23022117(.data_in(wire_d22_116),.data_out(wire_d22_117),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance23022118(.data_in(wire_d22_117),.data_out(wire_d22_118),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance23022119(.data_in(wire_d22_118),.data_out(d_out22),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance240230(.data_in(d_in23),.data_out(wire_d23_0),.clk(clk),.rst(rst));            //channel 24
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance240231(.data_in(wire_d23_0),.data_out(wire_d23_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance240232(.data_in(wire_d23_1),.data_out(wire_d23_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance240233(.data_in(wire_d23_2),.data_out(wire_d23_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance240234(.data_in(wire_d23_3),.data_out(wire_d23_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance240235(.data_in(wire_d23_4),.data_out(wire_d23_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance240236(.data_in(wire_d23_5),.data_out(wire_d23_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance240237(.data_in(wire_d23_6),.data_out(wire_d23_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance240238(.data_in(wire_d23_7),.data_out(wire_d23_8),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance240239(.data_in(wire_d23_8),.data_out(wire_d23_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402310(.data_in(wire_d23_9),.data_out(wire_d23_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402311(.data_in(wire_d23_10),.data_out(wire_d23_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2402312(.data_in(wire_d23_11),.data_out(wire_d23_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402313(.data_in(wire_d23_12),.data_out(wire_d23_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402314(.data_in(wire_d23_13),.data_out(wire_d23_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402315(.data_in(wire_d23_14),.data_out(wire_d23_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402316(.data_in(wire_d23_15),.data_out(wire_d23_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402317(.data_in(wire_d23_16),.data_out(wire_d23_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2402318(.data_in(wire_d23_17),.data_out(wire_d23_18),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2402319(.data_in(wire_d23_18),.data_out(wire_d23_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402320(.data_in(wire_d23_19),.data_out(wire_d23_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2402321(.data_in(wire_d23_20),.data_out(wire_d23_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2402322(.data_in(wire_d23_21),.data_out(wire_d23_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402323(.data_in(wire_d23_22),.data_out(wire_d23_23),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2402324(.data_in(wire_d23_23),.data_out(wire_d23_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2402325(.data_in(wire_d23_24),.data_out(wire_d23_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2402326(.data_in(wire_d23_25),.data_out(wire_d23_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2402327(.data_in(wire_d23_26),.data_out(wire_d23_27),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2402328(.data_in(wire_d23_27),.data_out(wire_d23_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402329(.data_in(wire_d23_28),.data_out(wire_d23_29),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402330(.data_in(wire_d23_29),.data_out(wire_d23_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402331(.data_in(wire_d23_30),.data_out(wire_d23_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402332(.data_in(wire_d23_31),.data_out(wire_d23_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402333(.data_in(wire_d23_32),.data_out(wire_d23_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402334(.data_in(wire_d23_33),.data_out(wire_d23_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402335(.data_in(wire_d23_34),.data_out(wire_d23_35),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2402336(.data_in(wire_d23_35),.data_out(wire_d23_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402337(.data_in(wire_d23_36),.data_out(wire_d23_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402338(.data_in(wire_d23_37),.data_out(wire_d23_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402339(.data_in(wire_d23_38),.data_out(wire_d23_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402340(.data_in(wire_d23_39),.data_out(wire_d23_40),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2402341(.data_in(wire_d23_40),.data_out(wire_d23_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402342(.data_in(wire_d23_41),.data_out(wire_d23_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2402343(.data_in(wire_d23_42),.data_out(wire_d23_43),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402344(.data_in(wire_d23_43),.data_out(wire_d23_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402345(.data_in(wire_d23_44),.data_out(wire_d23_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402346(.data_in(wire_d23_45),.data_out(wire_d23_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2402347(.data_in(wire_d23_46),.data_out(wire_d23_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2402348(.data_in(wire_d23_47),.data_out(wire_d23_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402349(.data_in(wire_d23_48),.data_out(wire_d23_49),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402350(.data_in(wire_d23_49),.data_out(wire_d23_50),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402351(.data_in(wire_d23_50),.data_out(wire_d23_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2402352(.data_in(wire_d23_51),.data_out(wire_d23_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2402353(.data_in(wire_d23_52),.data_out(wire_d23_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402354(.data_in(wire_d23_53),.data_out(wire_d23_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402355(.data_in(wire_d23_54),.data_out(wire_d23_55),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2402356(.data_in(wire_d23_55),.data_out(wire_d23_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402357(.data_in(wire_d23_56),.data_out(wire_d23_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402358(.data_in(wire_d23_57),.data_out(wire_d23_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402359(.data_in(wire_d23_58),.data_out(wire_d23_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402360(.data_in(wire_d23_59),.data_out(wire_d23_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2402361(.data_in(wire_d23_60),.data_out(wire_d23_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2402362(.data_in(wire_d23_61),.data_out(wire_d23_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402363(.data_in(wire_d23_62),.data_out(wire_d23_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402364(.data_in(wire_d23_63),.data_out(wire_d23_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402365(.data_in(wire_d23_64),.data_out(wire_d23_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2402366(.data_in(wire_d23_65),.data_out(wire_d23_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402367(.data_in(wire_d23_66),.data_out(wire_d23_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402368(.data_in(wire_d23_67),.data_out(wire_d23_68),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402369(.data_in(wire_d23_68),.data_out(wire_d23_69),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402370(.data_in(wire_d23_69),.data_out(wire_d23_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402371(.data_in(wire_d23_70),.data_out(wire_d23_71),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402372(.data_in(wire_d23_71),.data_out(wire_d23_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2402373(.data_in(wire_d23_72),.data_out(wire_d23_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2402374(.data_in(wire_d23_73),.data_out(wire_d23_74),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2402375(.data_in(wire_d23_74),.data_out(wire_d23_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402376(.data_in(wire_d23_75),.data_out(wire_d23_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2402377(.data_in(wire_d23_76),.data_out(wire_d23_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2402378(.data_in(wire_d23_77),.data_out(wire_d23_78),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402379(.data_in(wire_d23_78),.data_out(wire_d23_79),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402380(.data_in(wire_d23_79),.data_out(wire_d23_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402381(.data_in(wire_d23_80),.data_out(wire_d23_81),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2402382(.data_in(wire_d23_81),.data_out(wire_d23_82),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402383(.data_in(wire_d23_82),.data_out(wire_d23_83),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402384(.data_in(wire_d23_83),.data_out(wire_d23_84),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402385(.data_in(wire_d23_84),.data_out(wire_d23_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2402386(.data_in(wire_d23_85),.data_out(wire_d23_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402387(.data_in(wire_d23_86),.data_out(wire_d23_87),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402388(.data_in(wire_d23_87),.data_out(wire_d23_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2402389(.data_in(wire_d23_88),.data_out(wire_d23_89),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402390(.data_in(wire_d23_89),.data_out(wire_d23_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402391(.data_in(wire_d23_90),.data_out(wire_d23_91),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402392(.data_in(wire_d23_91),.data_out(wire_d23_92),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2402393(.data_in(wire_d23_92),.data_out(wire_d23_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2402394(.data_in(wire_d23_93),.data_out(wire_d23_94),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402395(.data_in(wire_d23_94),.data_out(wire_d23_95),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402396(.data_in(wire_d23_95),.data_out(wire_d23_96),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402397(.data_in(wire_d23_96),.data_out(wire_d23_97),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402398(.data_in(wire_d23_97),.data_out(wire_d23_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2402399(.data_in(wire_d23_98),.data_out(wire_d23_99),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance24023100(.data_in(wire_d23_99),.data_out(wire_d23_100),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance24023101(.data_in(wire_d23_100),.data_out(wire_d23_101),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance24023102(.data_in(wire_d23_101),.data_out(wire_d23_102),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance24023103(.data_in(wire_d23_102),.data_out(wire_d23_103),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance24023104(.data_in(wire_d23_103),.data_out(wire_d23_104),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance24023105(.data_in(wire_d23_104),.data_out(wire_d23_105),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance24023106(.data_in(wire_d23_105),.data_out(wire_d23_106),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance24023107(.data_in(wire_d23_106),.data_out(wire_d23_107),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance24023108(.data_in(wire_d23_107),.data_out(wire_d23_108),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance24023109(.data_in(wire_d23_108),.data_out(wire_d23_109),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance24023110(.data_in(wire_d23_109),.data_out(wire_d23_110),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance24023111(.data_in(wire_d23_110),.data_out(wire_d23_111),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance24023112(.data_in(wire_d23_111),.data_out(wire_d23_112),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance24023113(.data_in(wire_d23_112),.data_out(wire_d23_113),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance24023114(.data_in(wire_d23_113),.data_out(wire_d23_114),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance24023115(.data_in(wire_d23_114),.data_out(wire_d23_115),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance24023116(.data_in(wire_d23_115),.data_out(wire_d23_116),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance24023117(.data_in(wire_d23_116),.data_out(wire_d23_117),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance24023118(.data_in(wire_d23_117),.data_out(wire_d23_118),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance24023119(.data_in(wire_d23_118),.data_out(d_out23),.clk(clk),.rst(rst));

	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance250240(.data_in(d_in24),.data_out(wire_d24_0),.clk(clk),.rst(rst));            //channel 25
	decoder_top #(.WIDTH(WIDTH)) decoder_instance250241(.data_in(wire_d24_0),.data_out(wire_d24_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance250242(.data_in(wire_d24_1),.data_out(wire_d24_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance250243(.data_in(wire_d24_2),.data_out(wire_d24_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance250244(.data_in(wire_d24_3),.data_out(wire_d24_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance250245(.data_in(wire_d24_4),.data_out(wire_d24_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance250246(.data_in(wire_d24_5),.data_out(wire_d24_6),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance250247(.data_in(wire_d24_6),.data_out(wire_d24_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance250248(.data_in(wire_d24_7),.data_out(wire_d24_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance250249(.data_in(wire_d24_8),.data_out(wire_d24_9),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502410(.data_in(wire_d24_9),.data_out(wire_d24_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502411(.data_in(wire_d24_10),.data_out(wire_d24_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502412(.data_in(wire_d24_11),.data_out(wire_d24_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2502413(.data_in(wire_d24_12),.data_out(wire_d24_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502414(.data_in(wire_d24_13),.data_out(wire_d24_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502415(.data_in(wire_d24_14),.data_out(wire_d24_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502416(.data_in(wire_d24_15),.data_out(wire_d24_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502417(.data_in(wire_d24_16),.data_out(wire_d24_17),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2502418(.data_in(wire_d24_17),.data_out(wire_d24_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502419(.data_in(wire_d24_18),.data_out(wire_d24_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2502420(.data_in(wire_d24_19),.data_out(wire_d24_20),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502421(.data_in(wire_d24_20),.data_out(wire_d24_21),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502422(.data_in(wire_d24_21),.data_out(wire_d24_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502423(.data_in(wire_d24_22),.data_out(wire_d24_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502424(.data_in(wire_d24_23),.data_out(wire_d24_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2502425(.data_in(wire_d24_24),.data_out(wire_d24_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2502426(.data_in(wire_d24_25),.data_out(wire_d24_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502427(.data_in(wire_d24_26),.data_out(wire_d24_27),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2502428(.data_in(wire_d24_27),.data_out(wire_d24_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2502429(.data_in(wire_d24_28),.data_out(wire_d24_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502430(.data_in(wire_d24_29),.data_out(wire_d24_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2502431(.data_in(wire_d24_30),.data_out(wire_d24_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2502432(.data_in(wire_d24_31),.data_out(wire_d24_32),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502433(.data_in(wire_d24_32),.data_out(wire_d24_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502434(.data_in(wire_d24_33),.data_out(wire_d24_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502435(.data_in(wire_d24_34),.data_out(wire_d24_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2502436(.data_in(wire_d24_35),.data_out(wire_d24_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2502437(.data_in(wire_d24_36),.data_out(wire_d24_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502438(.data_in(wire_d24_37),.data_out(wire_d24_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2502439(.data_in(wire_d24_38),.data_out(wire_d24_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2502440(.data_in(wire_d24_39),.data_out(wire_d24_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2502441(.data_in(wire_d24_40),.data_out(wire_d24_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502442(.data_in(wire_d24_41),.data_out(wire_d24_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502443(.data_in(wire_d24_42),.data_out(wire_d24_43),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2502444(.data_in(wire_d24_43),.data_out(wire_d24_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502445(.data_in(wire_d24_44),.data_out(wire_d24_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502446(.data_in(wire_d24_45),.data_out(wire_d24_46),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2502447(.data_in(wire_d24_46),.data_out(wire_d24_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2502448(.data_in(wire_d24_47),.data_out(wire_d24_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2502449(.data_in(wire_d24_48),.data_out(wire_d24_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2502450(.data_in(wire_d24_49),.data_out(wire_d24_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502451(.data_in(wire_d24_50),.data_out(wire_d24_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502452(.data_in(wire_d24_51),.data_out(wire_d24_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2502453(.data_in(wire_d24_52),.data_out(wire_d24_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502454(.data_in(wire_d24_53),.data_out(wire_d24_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2502455(.data_in(wire_d24_54),.data_out(wire_d24_55),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2502456(.data_in(wire_d24_55),.data_out(wire_d24_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502457(.data_in(wire_d24_56),.data_out(wire_d24_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2502458(.data_in(wire_d24_57),.data_out(wire_d24_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502459(.data_in(wire_d24_58),.data_out(wire_d24_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2502460(.data_in(wire_d24_59),.data_out(wire_d24_60),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502461(.data_in(wire_d24_60),.data_out(wire_d24_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502462(.data_in(wire_d24_61),.data_out(wire_d24_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2502463(.data_in(wire_d24_62),.data_out(wire_d24_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502464(.data_in(wire_d24_63),.data_out(wire_d24_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502465(.data_in(wire_d24_64),.data_out(wire_d24_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2502466(.data_in(wire_d24_65),.data_out(wire_d24_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502467(.data_in(wire_d24_66),.data_out(wire_d24_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2502468(.data_in(wire_d24_67),.data_out(wire_d24_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502469(.data_in(wire_d24_68),.data_out(wire_d24_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2502470(.data_in(wire_d24_69),.data_out(wire_d24_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502471(.data_in(wire_d24_70),.data_out(wire_d24_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2502472(.data_in(wire_d24_71),.data_out(wire_d24_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502473(.data_in(wire_d24_72),.data_out(wire_d24_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2502474(.data_in(wire_d24_73),.data_out(wire_d24_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2502475(.data_in(wire_d24_74),.data_out(wire_d24_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2502476(.data_in(wire_d24_75),.data_out(wire_d24_76),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502477(.data_in(wire_d24_76),.data_out(wire_d24_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2502478(.data_in(wire_d24_77),.data_out(wire_d24_78),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502479(.data_in(wire_d24_78),.data_out(wire_d24_79),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502480(.data_in(wire_d24_79),.data_out(wire_d24_80),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502481(.data_in(wire_d24_80),.data_out(wire_d24_81),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502482(.data_in(wire_d24_81),.data_out(wire_d24_82),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502483(.data_in(wire_d24_82),.data_out(wire_d24_83),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2502484(.data_in(wire_d24_83),.data_out(wire_d24_84),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502485(.data_in(wire_d24_84),.data_out(wire_d24_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2502486(.data_in(wire_d24_85),.data_out(wire_d24_86),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502487(.data_in(wire_d24_86),.data_out(wire_d24_87),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2502488(.data_in(wire_d24_87),.data_out(wire_d24_88),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502489(.data_in(wire_d24_88),.data_out(wire_d24_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2502490(.data_in(wire_d24_89),.data_out(wire_d24_90),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502491(.data_in(wire_d24_90),.data_out(wire_d24_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2502492(.data_in(wire_d24_91),.data_out(wire_d24_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2502493(.data_in(wire_d24_92),.data_out(wire_d24_93),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2502494(.data_in(wire_d24_93),.data_out(wire_d24_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2502495(.data_in(wire_d24_94),.data_out(wire_d24_95),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502496(.data_in(wire_d24_95),.data_out(wire_d24_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502497(.data_in(wire_d24_96),.data_out(wire_d24_97),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502498(.data_in(wire_d24_97),.data_out(wire_d24_98),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502499(.data_in(wire_d24_98),.data_out(wire_d24_99),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance25024100(.data_in(wire_d24_99),.data_out(wire_d24_100),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance25024101(.data_in(wire_d24_100),.data_out(wire_d24_101),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance25024102(.data_in(wire_d24_101),.data_out(wire_d24_102),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance25024103(.data_in(wire_d24_102),.data_out(wire_d24_103),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance25024104(.data_in(wire_d24_103),.data_out(wire_d24_104),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance25024105(.data_in(wire_d24_104),.data_out(wire_d24_105),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance25024106(.data_in(wire_d24_105),.data_out(wire_d24_106),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance25024107(.data_in(wire_d24_106),.data_out(wire_d24_107),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance25024108(.data_in(wire_d24_107),.data_out(wire_d24_108),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance25024109(.data_in(wire_d24_108),.data_out(wire_d24_109),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance25024110(.data_in(wire_d24_109),.data_out(wire_d24_110),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance25024111(.data_in(wire_d24_110),.data_out(wire_d24_111),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance25024112(.data_in(wire_d24_111),.data_out(wire_d24_112),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance25024113(.data_in(wire_d24_112),.data_out(wire_d24_113),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance25024114(.data_in(wire_d24_113),.data_out(wire_d24_114),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance25024115(.data_in(wire_d24_114),.data_out(wire_d24_115),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance25024116(.data_in(wire_d24_115),.data_out(wire_d24_116),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance25024117(.data_in(wire_d24_116),.data_out(wire_d24_117),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance25024118(.data_in(wire_d24_117),.data_out(wire_d24_118),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance25024119(.data_in(wire_d24_118),.data_out(d_out24),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance260250(.data_in(d_in25),.data_out(wire_d25_0),.clk(clk),.rst(rst));            //channel 26
	encoder #(.WIDTH(WIDTH)) encoder_instance260251(.data_in(wire_d25_0),.data_out(wire_d25_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance260252(.data_in(wire_d25_1),.data_out(wire_d25_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance260253(.data_in(wire_d25_2),.data_out(wire_d25_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance260254(.data_in(wire_d25_3),.data_out(wire_d25_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance260255(.data_in(wire_d25_4),.data_out(wire_d25_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance260256(.data_in(wire_d25_5),.data_out(wire_d25_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance260257(.data_in(wire_d25_6),.data_out(wire_d25_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance260258(.data_in(wire_d25_7),.data_out(wire_d25_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance260259(.data_in(wire_d25_8),.data_out(wire_d25_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602510(.data_in(wire_d25_9),.data_out(wire_d25_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602511(.data_in(wire_d25_10),.data_out(wire_d25_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602512(.data_in(wire_d25_11),.data_out(wire_d25_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602513(.data_in(wire_d25_12),.data_out(wire_d25_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2602514(.data_in(wire_d25_13),.data_out(wire_d25_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602515(.data_in(wire_d25_14),.data_out(wire_d25_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602516(.data_in(wire_d25_15),.data_out(wire_d25_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602517(.data_in(wire_d25_16),.data_out(wire_d25_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602518(.data_in(wire_d25_17),.data_out(wire_d25_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602519(.data_in(wire_d25_18),.data_out(wire_d25_19),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2602520(.data_in(wire_d25_19),.data_out(wire_d25_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602521(.data_in(wire_d25_20),.data_out(wire_d25_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2602522(.data_in(wire_d25_21),.data_out(wire_d25_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602523(.data_in(wire_d25_22),.data_out(wire_d25_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602524(.data_in(wire_d25_23),.data_out(wire_d25_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602525(.data_in(wire_d25_24),.data_out(wire_d25_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2602526(.data_in(wire_d25_25),.data_out(wire_d25_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2602527(.data_in(wire_d25_26),.data_out(wire_d25_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2602528(.data_in(wire_d25_27),.data_out(wire_d25_28),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602529(.data_in(wire_d25_28),.data_out(wire_d25_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602530(.data_in(wire_d25_29),.data_out(wire_d25_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2602531(.data_in(wire_d25_30),.data_out(wire_d25_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2602532(.data_in(wire_d25_31),.data_out(wire_d25_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602533(.data_in(wire_d25_32),.data_out(wire_d25_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602534(.data_in(wire_d25_33),.data_out(wire_d25_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2602535(.data_in(wire_d25_34),.data_out(wire_d25_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602536(.data_in(wire_d25_35),.data_out(wire_d25_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2602537(.data_in(wire_d25_36),.data_out(wire_d25_37),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2602538(.data_in(wire_d25_37),.data_out(wire_d25_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602539(.data_in(wire_d25_38),.data_out(wire_d25_39),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2602540(.data_in(wire_d25_39),.data_out(wire_d25_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602541(.data_in(wire_d25_40),.data_out(wire_d25_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602542(.data_in(wire_d25_41),.data_out(wire_d25_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2602543(.data_in(wire_d25_42),.data_out(wire_d25_43),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602544(.data_in(wire_d25_43),.data_out(wire_d25_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2602545(.data_in(wire_d25_44),.data_out(wire_d25_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602546(.data_in(wire_d25_45),.data_out(wire_d25_46),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602547(.data_in(wire_d25_46),.data_out(wire_d25_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602548(.data_in(wire_d25_47),.data_out(wire_d25_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602549(.data_in(wire_d25_48),.data_out(wire_d25_49),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602550(.data_in(wire_d25_49),.data_out(wire_d25_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602551(.data_in(wire_d25_50),.data_out(wire_d25_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2602552(.data_in(wire_d25_51),.data_out(wire_d25_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602553(.data_in(wire_d25_52),.data_out(wire_d25_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2602554(.data_in(wire_d25_53),.data_out(wire_d25_54),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602555(.data_in(wire_d25_54),.data_out(wire_d25_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602556(.data_in(wire_d25_55),.data_out(wire_d25_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602557(.data_in(wire_d25_56),.data_out(wire_d25_57),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2602558(.data_in(wire_d25_57),.data_out(wire_d25_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602559(.data_in(wire_d25_58),.data_out(wire_d25_59),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2602560(.data_in(wire_d25_59),.data_out(wire_d25_60),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2602561(.data_in(wire_d25_60),.data_out(wire_d25_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602562(.data_in(wire_d25_61),.data_out(wire_d25_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602563(.data_in(wire_d25_62),.data_out(wire_d25_63),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602564(.data_in(wire_d25_63),.data_out(wire_d25_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2602565(.data_in(wire_d25_64),.data_out(wire_d25_65),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602566(.data_in(wire_d25_65),.data_out(wire_d25_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2602567(.data_in(wire_d25_66),.data_out(wire_d25_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602568(.data_in(wire_d25_67),.data_out(wire_d25_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602569(.data_in(wire_d25_68),.data_out(wire_d25_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2602570(.data_in(wire_d25_69),.data_out(wire_d25_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2602571(.data_in(wire_d25_70),.data_out(wire_d25_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2602572(.data_in(wire_d25_71),.data_out(wire_d25_72),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2602573(.data_in(wire_d25_72),.data_out(wire_d25_73),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2602574(.data_in(wire_d25_73),.data_out(wire_d25_74),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2602575(.data_in(wire_d25_74),.data_out(wire_d25_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602576(.data_in(wire_d25_75),.data_out(wire_d25_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602577(.data_in(wire_d25_76),.data_out(wire_d25_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602578(.data_in(wire_d25_77),.data_out(wire_d25_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2602579(.data_in(wire_d25_78),.data_out(wire_d25_79),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2602580(.data_in(wire_d25_79),.data_out(wire_d25_80),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602581(.data_in(wire_d25_80),.data_out(wire_d25_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2602582(.data_in(wire_d25_81),.data_out(wire_d25_82),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602583(.data_in(wire_d25_82),.data_out(wire_d25_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2602584(.data_in(wire_d25_83),.data_out(wire_d25_84),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602585(.data_in(wire_d25_84),.data_out(wire_d25_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2602586(.data_in(wire_d25_85),.data_out(wire_d25_86),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2602587(.data_in(wire_d25_86),.data_out(wire_d25_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2602588(.data_in(wire_d25_87),.data_out(wire_d25_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2602589(.data_in(wire_d25_88),.data_out(wire_d25_89),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602590(.data_in(wire_d25_89),.data_out(wire_d25_90),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602591(.data_in(wire_d25_90),.data_out(wire_d25_91),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602592(.data_in(wire_d25_91),.data_out(wire_d25_92),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602593(.data_in(wire_d25_92),.data_out(wire_d25_93),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602594(.data_in(wire_d25_93),.data_out(wire_d25_94),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602595(.data_in(wire_d25_94),.data_out(wire_d25_95),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2602596(.data_in(wire_d25_95),.data_out(wire_d25_96),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602597(.data_in(wire_d25_96),.data_out(wire_d25_97),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602598(.data_in(wire_d25_97),.data_out(wire_d25_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2602599(.data_in(wire_d25_98),.data_out(wire_d25_99),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance26025100(.data_in(wire_d25_99),.data_out(wire_d25_100),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance26025101(.data_in(wire_d25_100),.data_out(wire_d25_101),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance26025102(.data_in(wire_d25_101),.data_out(wire_d25_102),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance26025103(.data_in(wire_d25_102),.data_out(wire_d25_103),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance26025104(.data_in(wire_d25_103),.data_out(wire_d25_104),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance26025105(.data_in(wire_d25_104),.data_out(wire_d25_105),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance26025106(.data_in(wire_d25_105),.data_out(wire_d25_106),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance26025107(.data_in(wire_d25_106),.data_out(wire_d25_107),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance26025108(.data_in(wire_d25_107),.data_out(wire_d25_108),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance26025109(.data_in(wire_d25_108),.data_out(wire_d25_109),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance26025110(.data_in(wire_d25_109),.data_out(wire_d25_110),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance26025111(.data_in(wire_d25_110),.data_out(wire_d25_111),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance26025112(.data_in(wire_d25_111),.data_out(wire_d25_112),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance26025113(.data_in(wire_d25_112),.data_out(wire_d25_113),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance26025114(.data_in(wire_d25_113),.data_out(wire_d25_114),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance26025115(.data_in(wire_d25_114),.data_out(wire_d25_115),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance26025116(.data_in(wire_d25_115),.data_out(wire_d25_116),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance26025117(.data_in(wire_d25_116),.data_out(wire_d25_117),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance26025118(.data_in(wire_d25_117),.data_out(wire_d25_118),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance26025119(.data_in(wire_d25_118),.data_out(d_out25),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance270260(.data_in(d_in26),.data_out(wire_d26_0),.clk(clk),.rst(rst));            //channel 27
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance270261(.data_in(wire_d26_0),.data_out(wire_d26_1),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance270262(.data_in(wire_d26_1),.data_out(wire_d26_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance270263(.data_in(wire_d26_2),.data_out(wire_d26_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance270264(.data_in(wire_d26_3),.data_out(wire_d26_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance270265(.data_in(wire_d26_4),.data_out(wire_d26_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance270266(.data_in(wire_d26_5),.data_out(wire_d26_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance270267(.data_in(wire_d26_6),.data_out(wire_d26_7),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance270268(.data_in(wire_d26_7),.data_out(wire_d26_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance270269(.data_in(wire_d26_8),.data_out(wire_d26_9),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2702610(.data_in(wire_d26_9),.data_out(wire_d26_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2702611(.data_in(wire_d26_10),.data_out(wire_d26_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702612(.data_in(wire_d26_11),.data_out(wire_d26_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702613(.data_in(wire_d26_12),.data_out(wire_d26_13),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702614(.data_in(wire_d26_13),.data_out(wire_d26_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2702615(.data_in(wire_d26_14),.data_out(wire_d26_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2702616(.data_in(wire_d26_15),.data_out(wire_d26_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702617(.data_in(wire_d26_16),.data_out(wire_d26_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702618(.data_in(wire_d26_17),.data_out(wire_d26_18),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702619(.data_in(wire_d26_18),.data_out(wire_d26_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2702620(.data_in(wire_d26_19),.data_out(wire_d26_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702621(.data_in(wire_d26_20),.data_out(wire_d26_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2702622(.data_in(wire_d26_21),.data_out(wire_d26_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702623(.data_in(wire_d26_22),.data_out(wire_d26_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2702624(.data_in(wire_d26_23),.data_out(wire_d26_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702625(.data_in(wire_d26_24),.data_out(wire_d26_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2702626(.data_in(wire_d26_25),.data_out(wire_d26_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702627(.data_in(wire_d26_26),.data_out(wire_d26_27),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2702628(.data_in(wire_d26_27),.data_out(wire_d26_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702629(.data_in(wire_d26_28),.data_out(wire_d26_29),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2702630(.data_in(wire_d26_29),.data_out(wire_d26_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2702631(.data_in(wire_d26_30),.data_out(wire_d26_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702632(.data_in(wire_d26_31),.data_out(wire_d26_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702633(.data_in(wire_d26_32),.data_out(wire_d26_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702634(.data_in(wire_d26_33),.data_out(wire_d26_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702635(.data_in(wire_d26_34),.data_out(wire_d26_35),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2702636(.data_in(wire_d26_35),.data_out(wire_d26_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2702637(.data_in(wire_d26_36),.data_out(wire_d26_37),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2702638(.data_in(wire_d26_37),.data_out(wire_d26_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702639(.data_in(wire_d26_38),.data_out(wire_d26_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702640(.data_in(wire_d26_39),.data_out(wire_d26_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2702641(.data_in(wire_d26_40),.data_out(wire_d26_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702642(.data_in(wire_d26_41),.data_out(wire_d26_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702643(.data_in(wire_d26_42),.data_out(wire_d26_43),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2702644(.data_in(wire_d26_43),.data_out(wire_d26_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702645(.data_in(wire_d26_44),.data_out(wire_d26_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2702646(.data_in(wire_d26_45),.data_out(wire_d26_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702647(.data_in(wire_d26_46),.data_out(wire_d26_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2702648(.data_in(wire_d26_47),.data_out(wire_d26_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702649(.data_in(wire_d26_48),.data_out(wire_d26_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2702650(.data_in(wire_d26_49),.data_out(wire_d26_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702651(.data_in(wire_d26_50),.data_out(wire_d26_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2702652(.data_in(wire_d26_51),.data_out(wire_d26_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2702653(.data_in(wire_d26_52),.data_out(wire_d26_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2702654(.data_in(wire_d26_53),.data_out(wire_d26_54),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2702655(.data_in(wire_d26_54),.data_out(wire_d26_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702656(.data_in(wire_d26_55),.data_out(wire_d26_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2702657(.data_in(wire_d26_56),.data_out(wire_d26_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702658(.data_in(wire_d26_57),.data_out(wire_d26_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2702659(.data_in(wire_d26_58),.data_out(wire_d26_59),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702660(.data_in(wire_d26_59),.data_out(wire_d26_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702661(.data_in(wire_d26_60),.data_out(wire_d26_61),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702662(.data_in(wire_d26_61),.data_out(wire_d26_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702663(.data_in(wire_d26_62),.data_out(wire_d26_63),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2702664(.data_in(wire_d26_63),.data_out(wire_d26_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702665(.data_in(wire_d26_64),.data_out(wire_d26_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2702666(.data_in(wire_d26_65),.data_out(wire_d26_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2702667(.data_in(wire_d26_66),.data_out(wire_d26_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702668(.data_in(wire_d26_67),.data_out(wire_d26_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2702669(.data_in(wire_d26_68),.data_out(wire_d26_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702670(.data_in(wire_d26_69),.data_out(wire_d26_70),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2702671(.data_in(wire_d26_70),.data_out(wire_d26_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2702672(.data_in(wire_d26_71),.data_out(wire_d26_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702673(.data_in(wire_d26_72),.data_out(wire_d26_73),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2702674(.data_in(wire_d26_73),.data_out(wire_d26_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702675(.data_in(wire_d26_74),.data_out(wire_d26_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702676(.data_in(wire_d26_75),.data_out(wire_d26_76),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2702677(.data_in(wire_d26_76),.data_out(wire_d26_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702678(.data_in(wire_d26_77),.data_out(wire_d26_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702679(.data_in(wire_d26_78),.data_out(wire_d26_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702680(.data_in(wire_d26_79),.data_out(wire_d26_80),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702681(.data_in(wire_d26_80),.data_out(wire_d26_81),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702682(.data_in(wire_d26_81),.data_out(wire_d26_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702683(.data_in(wire_d26_82),.data_out(wire_d26_83),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2702684(.data_in(wire_d26_83),.data_out(wire_d26_84),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702685(.data_in(wire_d26_84),.data_out(wire_d26_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2702686(.data_in(wire_d26_85),.data_out(wire_d26_86),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702687(.data_in(wire_d26_86),.data_out(wire_d26_87),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2702688(.data_in(wire_d26_87),.data_out(wire_d26_88),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702689(.data_in(wire_d26_88),.data_out(wire_d26_89),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2702690(.data_in(wire_d26_89),.data_out(wire_d26_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702691(.data_in(wire_d26_90),.data_out(wire_d26_91),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2702692(.data_in(wire_d26_91),.data_out(wire_d26_92),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702693(.data_in(wire_d26_92),.data_out(wire_d26_93),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702694(.data_in(wire_d26_93),.data_out(wire_d26_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702695(.data_in(wire_d26_94),.data_out(wire_d26_95),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702696(.data_in(wire_d26_95),.data_out(wire_d26_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702697(.data_in(wire_d26_96),.data_out(wire_d26_97),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702698(.data_in(wire_d26_97),.data_out(wire_d26_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2702699(.data_in(wire_d26_98),.data_out(wire_d26_99),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance27026100(.data_in(wire_d26_99),.data_out(wire_d26_100),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance27026101(.data_in(wire_d26_100),.data_out(wire_d26_101),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance27026102(.data_in(wire_d26_101),.data_out(wire_d26_102),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance27026103(.data_in(wire_d26_102),.data_out(wire_d26_103),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance27026104(.data_in(wire_d26_103),.data_out(wire_d26_104),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance27026105(.data_in(wire_d26_104),.data_out(wire_d26_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance27026106(.data_in(wire_d26_105),.data_out(wire_d26_106),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance27026107(.data_in(wire_d26_106),.data_out(wire_d26_107),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance27026108(.data_in(wire_d26_107),.data_out(wire_d26_108),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance27026109(.data_in(wire_d26_108),.data_out(wire_d26_109),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance27026110(.data_in(wire_d26_109),.data_out(wire_d26_110),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance27026111(.data_in(wire_d26_110),.data_out(wire_d26_111),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance27026112(.data_in(wire_d26_111),.data_out(wire_d26_112),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance27026113(.data_in(wire_d26_112),.data_out(wire_d26_113),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance27026114(.data_in(wire_d26_113),.data_out(wire_d26_114),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance27026115(.data_in(wire_d26_114),.data_out(wire_d26_115),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance27026116(.data_in(wire_d26_115),.data_out(wire_d26_116),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance27026117(.data_in(wire_d26_116),.data_out(wire_d26_117),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance27026118(.data_in(wire_d26_117),.data_out(wire_d26_118),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance27026119(.data_in(wire_d26_118),.data_out(d_out26),.clk(clk),.rst(rst));

	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance280270(.data_in(d_in27),.data_out(wire_d27_0),.clk(clk),.rst(rst));            //channel 28
	encoder #(.WIDTH(WIDTH)) encoder_instance280271(.data_in(wire_d27_0),.data_out(wire_d27_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance280272(.data_in(wire_d27_1),.data_out(wire_d27_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance280273(.data_in(wire_d27_2),.data_out(wire_d27_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance280274(.data_in(wire_d27_3),.data_out(wire_d27_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance280275(.data_in(wire_d27_4),.data_out(wire_d27_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance280276(.data_in(wire_d27_5),.data_out(wire_d27_6),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance280277(.data_in(wire_d27_6),.data_out(wire_d27_7),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance280278(.data_in(wire_d27_7),.data_out(wire_d27_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance280279(.data_in(wire_d27_8),.data_out(wire_d27_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802710(.data_in(wire_d27_9),.data_out(wire_d27_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802711(.data_in(wire_d27_10),.data_out(wire_d27_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802712(.data_in(wire_d27_11),.data_out(wire_d27_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802713(.data_in(wire_d27_12),.data_out(wire_d27_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802714(.data_in(wire_d27_13),.data_out(wire_d27_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802715(.data_in(wire_d27_14),.data_out(wire_d27_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2802716(.data_in(wire_d27_15),.data_out(wire_d27_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802717(.data_in(wire_d27_16),.data_out(wire_d27_17),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2802718(.data_in(wire_d27_17),.data_out(wire_d27_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802719(.data_in(wire_d27_18),.data_out(wire_d27_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802720(.data_in(wire_d27_19),.data_out(wire_d27_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2802721(.data_in(wire_d27_20),.data_out(wire_d27_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802722(.data_in(wire_d27_21),.data_out(wire_d27_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2802723(.data_in(wire_d27_22),.data_out(wire_d27_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802724(.data_in(wire_d27_23),.data_out(wire_d27_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802725(.data_in(wire_d27_24),.data_out(wire_d27_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802726(.data_in(wire_d27_25),.data_out(wire_d27_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802727(.data_in(wire_d27_26),.data_out(wire_d27_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802728(.data_in(wire_d27_27),.data_out(wire_d27_28),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802729(.data_in(wire_d27_28),.data_out(wire_d27_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802730(.data_in(wire_d27_29),.data_out(wire_d27_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802731(.data_in(wire_d27_30),.data_out(wire_d27_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802732(.data_in(wire_d27_31),.data_out(wire_d27_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802733(.data_in(wire_d27_32),.data_out(wire_d27_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802734(.data_in(wire_d27_33),.data_out(wire_d27_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802735(.data_in(wire_d27_34),.data_out(wire_d27_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802736(.data_in(wire_d27_35),.data_out(wire_d27_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802737(.data_in(wire_d27_36),.data_out(wire_d27_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802738(.data_in(wire_d27_37),.data_out(wire_d27_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802739(.data_in(wire_d27_38),.data_out(wire_d27_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802740(.data_in(wire_d27_39),.data_out(wire_d27_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2802741(.data_in(wire_d27_40),.data_out(wire_d27_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802742(.data_in(wire_d27_41),.data_out(wire_d27_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2802743(.data_in(wire_d27_42),.data_out(wire_d27_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802744(.data_in(wire_d27_43),.data_out(wire_d27_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802745(.data_in(wire_d27_44),.data_out(wire_d27_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802746(.data_in(wire_d27_45),.data_out(wire_d27_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802747(.data_in(wire_d27_46),.data_out(wire_d27_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802748(.data_in(wire_d27_47),.data_out(wire_d27_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2802749(.data_in(wire_d27_48),.data_out(wire_d27_49),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802750(.data_in(wire_d27_49),.data_out(wire_d27_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802751(.data_in(wire_d27_50),.data_out(wire_d27_51),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802752(.data_in(wire_d27_51),.data_out(wire_d27_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802753(.data_in(wire_d27_52),.data_out(wire_d27_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2802754(.data_in(wire_d27_53),.data_out(wire_d27_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802755(.data_in(wire_d27_54),.data_out(wire_d27_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802756(.data_in(wire_d27_55),.data_out(wire_d27_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802757(.data_in(wire_d27_56),.data_out(wire_d27_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802758(.data_in(wire_d27_57),.data_out(wire_d27_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802759(.data_in(wire_d27_58),.data_out(wire_d27_59),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2802760(.data_in(wire_d27_59),.data_out(wire_d27_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802761(.data_in(wire_d27_60),.data_out(wire_d27_61),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2802762(.data_in(wire_d27_61),.data_out(wire_d27_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802763(.data_in(wire_d27_62),.data_out(wire_d27_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802764(.data_in(wire_d27_63),.data_out(wire_d27_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802765(.data_in(wire_d27_64),.data_out(wire_d27_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802766(.data_in(wire_d27_65),.data_out(wire_d27_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802767(.data_in(wire_d27_66),.data_out(wire_d27_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802768(.data_in(wire_d27_67),.data_out(wire_d27_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2802769(.data_in(wire_d27_68),.data_out(wire_d27_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802770(.data_in(wire_d27_69),.data_out(wire_d27_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802771(.data_in(wire_d27_70),.data_out(wire_d27_71),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802772(.data_in(wire_d27_71),.data_out(wire_d27_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802773(.data_in(wire_d27_72),.data_out(wire_d27_73),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802774(.data_in(wire_d27_73),.data_out(wire_d27_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802775(.data_in(wire_d27_74),.data_out(wire_d27_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2802776(.data_in(wire_d27_75),.data_out(wire_d27_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802777(.data_in(wire_d27_76),.data_out(wire_d27_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802778(.data_in(wire_d27_77),.data_out(wire_d27_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802779(.data_in(wire_d27_78),.data_out(wire_d27_79),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802780(.data_in(wire_d27_79),.data_out(wire_d27_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2802781(.data_in(wire_d27_80),.data_out(wire_d27_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2802782(.data_in(wire_d27_81),.data_out(wire_d27_82),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802783(.data_in(wire_d27_82),.data_out(wire_d27_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802784(.data_in(wire_d27_83),.data_out(wire_d27_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2802785(.data_in(wire_d27_84),.data_out(wire_d27_85),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2802786(.data_in(wire_d27_85),.data_out(wire_d27_86),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802787(.data_in(wire_d27_86),.data_out(wire_d27_87),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802788(.data_in(wire_d27_87),.data_out(wire_d27_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2802789(.data_in(wire_d27_88),.data_out(wire_d27_89),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802790(.data_in(wire_d27_89),.data_out(wire_d27_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2802791(.data_in(wire_d27_90),.data_out(wire_d27_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802792(.data_in(wire_d27_91),.data_out(wire_d27_92),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802793(.data_in(wire_d27_92),.data_out(wire_d27_93),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802794(.data_in(wire_d27_93),.data_out(wire_d27_94),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802795(.data_in(wire_d27_94),.data_out(wire_d27_95),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2802796(.data_in(wire_d27_95),.data_out(wire_d27_96),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802797(.data_in(wire_d27_96),.data_out(wire_d27_97),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802798(.data_in(wire_d27_97),.data_out(wire_d27_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802799(.data_in(wire_d27_98),.data_out(wire_d27_99),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance28027100(.data_in(wire_d27_99),.data_out(wire_d27_100),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance28027101(.data_in(wire_d27_100),.data_out(wire_d27_101),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance28027102(.data_in(wire_d27_101),.data_out(wire_d27_102),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance28027103(.data_in(wire_d27_102),.data_out(wire_d27_103),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance28027104(.data_in(wire_d27_103),.data_out(wire_d27_104),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance28027105(.data_in(wire_d27_104),.data_out(wire_d27_105),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance28027106(.data_in(wire_d27_105),.data_out(wire_d27_106),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance28027107(.data_in(wire_d27_106),.data_out(wire_d27_107),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance28027108(.data_in(wire_d27_107),.data_out(wire_d27_108),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance28027109(.data_in(wire_d27_108),.data_out(wire_d27_109),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance28027110(.data_in(wire_d27_109),.data_out(wire_d27_110),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance28027111(.data_in(wire_d27_110),.data_out(wire_d27_111),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance28027112(.data_in(wire_d27_111),.data_out(wire_d27_112),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance28027113(.data_in(wire_d27_112),.data_out(wire_d27_113),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance28027114(.data_in(wire_d27_113),.data_out(wire_d27_114),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance28027115(.data_in(wire_d27_114),.data_out(wire_d27_115),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance28027116(.data_in(wire_d27_115),.data_out(wire_d27_116),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance28027117(.data_in(wire_d27_116),.data_out(wire_d27_117),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance28027118(.data_in(wire_d27_117),.data_out(wire_d27_118),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance28027119(.data_in(wire_d27_118),.data_out(d_out27),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance290280(.data_in(d_in28),.data_out(wire_d28_0),.clk(clk),.rst(rst));            //channel 29
	encoder #(.WIDTH(WIDTH)) encoder_instance290281(.data_in(wire_d28_0),.data_out(wire_d28_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance290282(.data_in(wire_d28_1),.data_out(wire_d28_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance290283(.data_in(wire_d28_2),.data_out(wire_d28_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance290284(.data_in(wire_d28_3),.data_out(wire_d28_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance290285(.data_in(wire_d28_4),.data_out(wire_d28_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance290286(.data_in(wire_d28_5),.data_out(wire_d28_6),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance290287(.data_in(wire_d28_6),.data_out(wire_d28_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance290288(.data_in(wire_d28_7),.data_out(wire_d28_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance290289(.data_in(wire_d28_8),.data_out(wire_d28_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2902810(.data_in(wire_d28_9),.data_out(wire_d28_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902811(.data_in(wire_d28_10),.data_out(wire_d28_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2902812(.data_in(wire_d28_11),.data_out(wire_d28_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902813(.data_in(wire_d28_12),.data_out(wire_d28_13),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2902814(.data_in(wire_d28_13),.data_out(wire_d28_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902815(.data_in(wire_d28_14),.data_out(wire_d28_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902816(.data_in(wire_d28_15),.data_out(wire_d28_16),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902817(.data_in(wire_d28_16),.data_out(wire_d28_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902818(.data_in(wire_d28_17),.data_out(wire_d28_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902819(.data_in(wire_d28_18),.data_out(wire_d28_19),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2902820(.data_in(wire_d28_19),.data_out(wire_d28_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902821(.data_in(wire_d28_20),.data_out(wire_d28_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2902822(.data_in(wire_d28_21),.data_out(wire_d28_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902823(.data_in(wire_d28_22),.data_out(wire_d28_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902824(.data_in(wire_d28_23),.data_out(wire_d28_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902825(.data_in(wire_d28_24),.data_out(wire_d28_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902826(.data_in(wire_d28_25),.data_out(wire_d28_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902827(.data_in(wire_d28_26),.data_out(wire_d28_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902828(.data_in(wire_d28_27),.data_out(wire_d28_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902829(.data_in(wire_d28_28),.data_out(wire_d28_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902830(.data_in(wire_d28_29),.data_out(wire_d28_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902831(.data_in(wire_d28_30),.data_out(wire_d28_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902832(.data_in(wire_d28_31),.data_out(wire_d28_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2902833(.data_in(wire_d28_32),.data_out(wire_d28_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902834(.data_in(wire_d28_33),.data_out(wire_d28_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902835(.data_in(wire_d28_34),.data_out(wire_d28_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902836(.data_in(wire_d28_35),.data_out(wire_d28_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902837(.data_in(wire_d28_36),.data_out(wire_d28_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2902838(.data_in(wire_d28_37),.data_out(wire_d28_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902839(.data_in(wire_d28_38),.data_out(wire_d28_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2902840(.data_in(wire_d28_39),.data_out(wire_d28_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2902841(.data_in(wire_d28_40),.data_out(wire_d28_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902842(.data_in(wire_d28_41),.data_out(wire_d28_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902843(.data_in(wire_d28_42),.data_out(wire_d28_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902844(.data_in(wire_d28_43),.data_out(wire_d28_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902845(.data_in(wire_d28_44),.data_out(wire_d28_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902846(.data_in(wire_d28_45),.data_out(wire_d28_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902847(.data_in(wire_d28_46),.data_out(wire_d28_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902848(.data_in(wire_d28_47),.data_out(wire_d28_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902849(.data_in(wire_d28_48),.data_out(wire_d28_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902850(.data_in(wire_d28_49),.data_out(wire_d28_50),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902851(.data_in(wire_d28_50),.data_out(wire_d28_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902852(.data_in(wire_d28_51),.data_out(wire_d28_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2902853(.data_in(wire_d28_52),.data_out(wire_d28_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902854(.data_in(wire_d28_53),.data_out(wire_d28_54),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2902855(.data_in(wire_d28_54),.data_out(wire_d28_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2902856(.data_in(wire_d28_55),.data_out(wire_d28_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902857(.data_in(wire_d28_56),.data_out(wire_d28_57),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902858(.data_in(wire_d28_57),.data_out(wire_d28_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2902859(.data_in(wire_d28_58),.data_out(wire_d28_59),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2902860(.data_in(wire_d28_59),.data_out(wire_d28_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902861(.data_in(wire_d28_60),.data_out(wire_d28_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2902862(.data_in(wire_d28_61),.data_out(wire_d28_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2902863(.data_in(wire_d28_62),.data_out(wire_d28_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902864(.data_in(wire_d28_63),.data_out(wire_d28_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902865(.data_in(wire_d28_64),.data_out(wire_d28_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2902866(.data_in(wire_d28_65),.data_out(wire_d28_66),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902867(.data_in(wire_d28_66),.data_out(wire_d28_67),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2902868(.data_in(wire_d28_67),.data_out(wire_d28_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902869(.data_in(wire_d28_68),.data_out(wire_d28_69),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902870(.data_in(wire_d28_69),.data_out(wire_d28_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902871(.data_in(wire_d28_70),.data_out(wire_d28_71),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902872(.data_in(wire_d28_71),.data_out(wire_d28_72),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2902873(.data_in(wire_d28_72),.data_out(wire_d28_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902874(.data_in(wire_d28_73),.data_out(wire_d28_74),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2902875(.data_in(wire_d28_74),.data_out(wire_d28_75),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2902876(.data_in(wire_d28_75),.data_out(wire_d28_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902877(.data_in(wire_d28_76),.data_out(wire_d28_77),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902878(.data_in(wire_d28_77),.data_out(wire_d28_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902879(.data_in(wire_d28_78),.data_out(wire_d28_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2902880(.data_in(wire_d28_79),.data_out(wire_d28_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902881(.data_in(wire_d28_80),.data_out(wire_d28_81),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902882(.data_in(wire_d28_81),.data_out(wire_d28_82),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902883(.data_in(wire_d28_82),.data_out(wire_d28_83),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2902884(.data_in(wire_d28_83),.data_out(wire_d28_84),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902885(.data_in(wire_d28_84),.data_out(wire_d28_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2902886(.data_in(wire_d28_85),.data_out(wire_d28_86),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902887(.data_in(wire_d28_86),.data_out(wire_d28_87),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902888(.data_in(wire_d28_87),.data_out(wire_d28_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2902889(.data_in(wire_d28_88),.data_out(wire_d28_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2902890(.data_in(wire_d28_89),.data_out(wire_d28_90),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902891(.data_in(wire_d28_90),.data_out(wire_d28_91),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2902892(.data_in(wire_d28_91),.data_out(wire_d28_92),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902893(.data_in(wire_d28_92),.data_out(wire_d28_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2902894(.data_in(wire_d28_93),.data_out(wire_d28_94),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902895(.data_in(wire_d28_94),.data_out(wire_d28_95),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902896(.data_in(wire_d28_95),.data_out(wire_d28_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902897(.data_in(wire_d28_96),.data_out(wire_d28_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2902898(.data_in(wire_d28_97),.data_out(wire_d28_98),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902899(.data_in(wire_d28_98),.data_out(wire_d28_99),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance29028100(.data_in(wire_d28_99),.data_out(wire_d28_100),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance29028101(.data_in(wire_d28_100),.data_out(wire_d28_101),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance29028102(.data_in(wire_d28_101),.data_out(wire_d28_102),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance29028103(.data_in(wire_d28_102),.data_out(wire_d28_103),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance29028104(.data_in(wire_d28_103),.data_out(wire_d28_104),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance29028105(.data_in(wire_d28_104),.data_out(wire_d28_105),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance29028106(.data_in(wire_d28_105),.data_out(wire_d28_106),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance29028107(.data_in(wire_d28_106),.data_out(wire_d28_107),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance29028108(.data_in(wire_d28_107),.data_out(wire_d28_108),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance29028109(.data_in(wire_d28_108),.data_out(wire_d28_109),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance29028110(.data_in(wire_d28_109),.data_out(wire_d28_110),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance29028111(.data_in(wire_d28_110),.data_out(wire_d28_111),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance29028112(.data_in(wire_d28_111),.data_out(wire_d28_112),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance29028113(.data_in(wire_d28_112),.data_out(wire_d28_113),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance29028114(.data_in(wire_d28_113),.data_out(wire_d28_114),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance29028115(.data_in(wire_d28_114),.data_out(wire_d28_115),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance29028116(.data_in(wire_d28_115),.data_out(wire_d28_116),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance29028117(.data_in(wire_d28_116),.data_out(wire_d28_117),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance29028118(.data_in(wire_d28_117),.data_out(wire_d28_118),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance29028119(.data_in(wire_d28_118),.data_out(d_out28),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance300290(.data_in(d_in29),.data_out(wire_d29_0),.clk(clk),.rst(rst));            //channel 30
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance300291(.data_in(wire_d29_0),.data_out(wire_d29_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance300292(.data_in(wire_d29_1),.data_out(wire_d29_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance300293(.data_in(wire_d29_2),.data_out(wire_d29_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance300294(.data_in(wire_d29_3),.data_out(wire_d29_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance300295(.data_in(wire_d29_4),.data_out(wire_d29_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance300296(.data_in(wire_d29_5),.data_out(wire_d29_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance300297(.data_in(wire_d29_6),.data_out(wire_d29_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance300298(.data_in(wire_d29_7),.data_out(wire_d29_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance300299(.data_in(wire_d29_8),.data_out(wire_d29_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002910(.data_in(wire_d29_9),.data_out(wire_d29_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002911(.data_in(wire_d29_10),.data_out(wire_d29_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002912(.data_in(wire_d29_11),.data_out(wire_d29_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002913(.data_in(wire_d29_12),.data_out(wire_d29_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002914(.data_in(wire_d29_13),.data_out(wire_d29_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002915(.data_in(wire_d29_14),.data_out(wire_d29_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002916(.data_in(wire_d29_15),.data_out(wire_d29_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002917(.data_in(wire_d29_16),.data_out(wire_d29_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3002918(.data_in(wire_d29_17),.data_out(wire_d29_18),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002919(.data_in(wire_d29_18),.data_out(wire_d29_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002920(.data_in(wire_d29_19),.data_out(wire_d29_20),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002921(.data_in(wire_d29_20),.data_out(wire_d29_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002922(.data_in(wire_d29_21),.data_out(wire_d29_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002923(.data_in(wire_d29_22),.data_out(wire_d29_23),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3002924(.data_in(wire_d29_23),.data_out(wire_d29_24),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3002925(.data_in(wire_d29_24),.data_out(wire_d29_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002926(.data_in(wire_d29_25),.data_out(wire_d29_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002927(.data_in(wire_d29_26),.data_out(wire_d29_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3002928(.data_in(wire_d29_27),.data_out(wire_d29_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3002929(.data_in(wire_d29_28),.data_out(wire_d29_29),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3002930(.data_in(wire_d29_29),.data_out(wire_d29_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002931(.data_in(wire_d29_30),.data_out(wire_d29_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002932(.data_in(wire_d29_31),.data_out(wire_d29_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3002933(.data_in(wire_d29_32),.data_out(wire_d29_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002934(.data_in(wire_d29_33),.data_out(wire_d29_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3002935(.data_in(wire_d29_34),.data_out(wire_d29_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002936(.data_in(wire_d29_35),.data_out(wire_d29_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002937(.data_in(wire_d29_36),.data_out(wire_d29_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002938(.data_in(wire_d29_37),.data_out(wire_d29_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002939(.data_in(wire_d29_38),.data_out(wire_d29_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002940(.data_in(wire_d29_39),.data_out(wire_d29_40),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3002941(.data_in(wire_d29_40),.data_out(wire_d29_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002942(.data_in(wire_d29_41),.data_out(wire_d29_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3002943(.data_in(wire_d29_42),.data_out(wire_d29_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002944(.data_in(wire_d29_43),.data_out(wire_d29_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002945(.data_in(wire_d29_44),.data_out(wire_d29_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002946(.data_in(wire_d29_45),.data_out(wire_d29_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002947(.data_in(wire_d29_46),.data_out(wire_d29_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002948(.data_in(wire_d29_47),.data_out(wire_d29_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002949(.data_in(wire_d29_48),.data_out(wire_d29_49),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002950(.data_in(wire_d29_49),.data_out(wire_d29_50),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3002951(.data_in(wire_d29_50),.data_out(wire_d29_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002952(.data_in(wire_d29_51),.data_out(wire_d29_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002953(.data_in(wire_d29_52),.data_out(wire_d29_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002954(.data_in(wire_d29_53),.data_out(wire_d29_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3002955(.data_in(wire_d29_54),.data_out(wire_d29_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3002956(.data_in(wire_d29_55),.data_out(wire_d29_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002957(.data_in(wire_d29_56),.data_out(wire_d29_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002958(.data_in(wire_d29_57),.data_out(wire_d29_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002959(.data_in(wire_d29_58),.data_out(wire_d29_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3002960(.data_in(wire_d29_59),.data_out(wire_d29_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002961(.data_in(wire_d29_60),.data_out(wire_d29_61),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002962(.data_in(wire_d29_61),.data_out(wire_d29_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002963(.data_in(wire_d29_62),.data_out(wire_d29_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3002964(.data_in(wire_d29_63),.data_out(wire_d29_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002965(.data_in(wire_d29_64),.data_out(wire_d29_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002966(.data_in(wire_d29_65),.data_out(wire_d29_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002967(.data_in(wire_d29_66),.data_out(wire_d29_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3002968(.data_in(wire_d29_67),.data_out(wire_d29_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3002969(.data_in(wire_d29_68),.data_out(wire_d29_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002970(.data_in(wire_d29_69),.data_out(wire_d29_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002971(.data_in(wire_d29_70),.data_out(wire_d29_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002972(.data_in(wire_d29_71),.data_out(wire_d29_72),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3002973(.data_in(wire_d29_72),.data_out(wire_d29_73),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3002974(.data_in(wire_d29_73),.data_out(wire_d29_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002975(.data_in(wire_d29_74),.data_out(wire_d29_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002976(.data_in(wire_d29_75),.data_out(wire_d29_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3002977(.data_in(wire_d29_76),.data_out(wire_d29_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3002978(.data_in(wire_d29_77),.data_out(wire_d29_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002979(.data_in(wire_d29_78),.data_out(wire_d29_79),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002980(.data_in(wire_d29_79),.data_out(wire_d29_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3002981(.data_in(wire_d29_80),.data_out(wire_d29_81),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3002982(.data_in(wire_d29_81),.data_out(wire_d29_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002983(.data_in(wire_d29_82),.data_out(wire_d29_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3002984(.data_in(wire_d29_83),.data_out(wire_d29_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002985(.data_in(wire_d29_84),.data_out(wire_d29_85),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002986(.data_in(wire_d29_85),.data_out(wire_d29_86),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002987(.data_in(wire_d29_86),.data_out(wire_d29_87),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002988(.data_in(wire_d29_87),.data_out(wire_d29_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3002989(.data_in(wire_d29_88),.data_out(wire_d29_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3002990(.data_in(wire_d29_89),.data_out(wire_d29_90),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002991(.data_in(wire_d29_90),.data_out(wire_d29_91),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002992(.data_in(wire_d29_91),.data_out(wire_d29_92),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002993(.data_in(wire_d29_92),.data_out(wire_d29_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3002994(.data_in(wire_d29_93),.data_out(wire_d29_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002995(.data_in(wire_d29_94),.data_out(wire_d29_95),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002996(.data_in(wire_d29_95),.data_out(wire_d29_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002997(.data_in(wire_d29_96),.data_out(wire_d29_97),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002998(.data_in(wire_d29_97),.data_out(wire_d29_98),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002999(.data_in(wire_d29_98),.data_out(wire_d29_99),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance30029100(.data_in(wire_d29_99),.data_out(wire_d29_100),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance30029101(.data_in(wire_d29_100),.data_out(wire_d29_101),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance30029102(.data_in(wire_d29_101),.data_out(wire_d29_102),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance30029103(.data_in(wire_d29_102),.data_out(wire_d29_103),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance30029104(.data_in(wire_d29_103),.data_out(wire_d29_104),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance30029105(.data_in(wire_d29_104),.data_out(wire_d29_105),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance30029106(.data_in(wire_d29_105),.data_out(wire_d29_106),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance30029107(.data_in(wire_d29_106),.data_out(wire_d29_107),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance30029108(.data_in(wire_d29_107),.data_out(wire_d29_108),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance30029109(.data_in(wire_d29_108),.data_out(wire_d29_109),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance30029110(.data_in(wire_d29_109),.data_out(wire_d29_110),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance30029111(.data_in(wire_d29_110),.data_out(wire_d29_111),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance30029112(.data_in(wire_d29_111),.data_out(wire_d29_112),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance30029113(.data_in(wire_d29_112),.data_out(wire_d29_113),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance30029114(.data_in(wire_d29_113),.data_out(wire_d29_114),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance30029115(.data_in(wire_d29_114),.data_out(wire_d29_115),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance30029116(.data_in(wire_d29_115),.data_out(wire_d29_116),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance30029117(.data_in(wire_d29_116),.data_out(wire_d29_117),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance30029118(.data_in(wire_d29_117),.data_out(wire_d29_118),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance30029119(.data_in(wire_d29_118),.data_out(d_out29),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance310300(.data_in(d_in30),.data_out(wire_d30_0),.clk(clk),.rst(rst));            //channel 31
	decoder_top #(.WIDTH(WIDTH)) decoder_instance310301(.data_in(wire_d30_0),.data_out(wire_d30_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance310302(.data_in(wire_d30_1),.data_out(wire_d30_2),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance310303(.data_in(wire_d30_2),.data_out(wire_d30_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance310304(.data_in(wire_d30_3),.data_out(wire_d30_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance310305(.data_in(wire_d30_4),.data_out(wire_d30_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance310306(.data_in(wire_d30_5),.data_out(wire_d30_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance310307(.data_in(wire_d30_6),.data_out(wire_d30_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance310308(.data_in(wire_d30_7),.data_out(wire_d30_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance310309(.data_in(wire_d30_8),.data_out(wire_d30_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3103010(.data_in(wire_d30_9),.data_out(wire_d30_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3103011(.data_in(wire_d30_10),.data_out(wire_d30_11),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3103012(.data_in(wire_d30_11),.data_out(wire_d30_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103013(.data_in(wire_d30_12),.data_out(wire_d30_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103014(.data_in(wire_d30_13),.data_out(wire_d30_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103015(.data_in(wire_d30_14),.data_out(wire_d30_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103016(.data_in(wire_d30_15),.data_out(wire_d30_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103017(.data_in(wire_d30_16),.data_out(wire_d30_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103018(.data_in(wire_d30_17),.data_out(wire_d30_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103019(.data_in(wire_d30_18),.data_out(wire_d30_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103020(.data_in(wire_d30_19),.data_out(wire_d30_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103021(.data_in(wire_d30_20),.data_out(wire_d30_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103022(.data_in(wire_d30_21),.data_out(wire_d30_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103023(.data_in(wire_d30_22),.data_out(wire_d30_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3103024(.data_in(wire_d30_23),.data_out(wire_d30_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3103025(.data_in(wire_d30_24),.data_out(wire_d30_25),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3103026(.data_in(wire_d30_25),.data_out(wire_d30_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3103027(.data_in(wire_d30_26),.data_out(wire_d30_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3103028(.data_in(wire_d30_27),.data_out(wire_d30_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103029(.data_in(wire_d30_28),.data_out(wire_d30_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103030(.data_in(wire_d30_29),.data_out(wire_d30_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3103031(.data_in(wire_d30_30),.data_out(wire_d30_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103032(.data_in(wire_d30_31),.data_out(wire_d30_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3103033(.data_in(wire_d30_32),.data_out(wire_d30_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103034(.data_in(wire_d30_33),.data_out(wire_d30_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103035(.data_in(wire_d30_34),.data_out(wire_d30_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103036(.data_in(wire_d30_35),.data_out(wire_d30_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3103037(.data_in(wire_d30_36),.data_out(wire_d30_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103038(.data_in(wire_d30_37),.data_out(wire_d30_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103039(.data_in(wire_d30_38),.data_out(wire_d30_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103040(.data_in(wire_d30_39),.data_out(wire_d30_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3103041(.data_in(wire_d30_40),.data_out(wire_d30_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103042(.data_in(wire_d30_41),.data_out(wire_d30_42),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3103043(.data_in(wire_d30_42),.data_out(wire_d30_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103044(.data_in(wire_d30_43),.data_out(wire_d30_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3103045(.data_in(wire_d30_44),.data_out(wire_d30_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103046(.data_in(wire_d30_45),.data_out(wire_d30_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103047(.data_in(wire_d30_46),.data_out(wire_d30_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103048(.data_in(wire_d30_47),.data_out(wire_d30_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3103049(.data_in(wire_d30_48),.data_out(wire_d30_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103050(.data_in(wire_d30_49),.data_out(wire_d30_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103051(.data_in(wire_d30_50),.data_out(wire_d30_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3103052(.data_in(wire_d30_51),.data_out(wire_d30_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103053(.data_in(wire_d30_52),.data_out(wire_d30_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3103054(.data_in(wire_d30_53),.data_out(wire_d30_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3103055(.data_in(wire_d30_54),.data_out(wire_d30_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3103056(.data_in(wire_d30_55),.data_out(wire_d30_56),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103057(.data_in(wire_d30_56),.data_out(wire_d30_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3103058(.data_in(wire_d30_57),.data_out(wire_d30_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103059(.data_in(wire_d30_58),.data_out(wire_d30_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103060(.data_in(wire_d30_59),.data_out(wire_d30_60),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103061(.data_in(wire_d30_60),.data_out(wire_d30_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103062(.data_in(wire_d30_61),.data_out(wire_d30_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103063(.data_in(wire_d30_62),.data_out(wire_d30_63),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103064(.data_in(wire_d30_63),.data_out(wire_d30_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103065(.data_in(wire_d30_64),.data_out(wire_d30_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3103066(.data_in(wire_d30_65),.data_out(wire_d30_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103067(.data_in(wire_d30_66),.data_out(wire_d30_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3103068(.data_in(wire_d30_67),.data_out(wire_d30_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3103069(.data_in(wire_d30_68),.data_out(wire_d30_69),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3103070(.data_in(wire_d30_69),.data_out(wire_d30_70),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103071(.data_in(wire_d30_70),.data_out(wire_d30_71),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103072(.data_in(wire_d30_71),.data_out(wire_d30_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103073(.data_in(wire_d30_72),.data_out(wire_d30_73),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3103074(.data_in(wire_d30_73),.data_out(wire_d30_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3103075(.data_in(wire_d30_74),.data_out(wire_d30_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3103076(.data_in(wire_d30_75),.data_out(wire_d30_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103077(.data_in(wire_d30_76),.data_out(wire_d30_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103078(.data_in(wire_d30_77),.data_out(wire_d30_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3103079(.data_in(wire_d30_78),.data_out(wire_d30_79),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103080(.data_in(wire_d30_79),.data_out(wire_d30_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103081(.data_in(wire_d30_80),.data_out(wire_d30_81),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3103082(.data_in(wire_d30_81),.data_out(wire_d30_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3103083(.data_in(wire_d30_82),.data_out(wire_d30_83),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103084(.data_in(wire_d30_83),.data_out(wire_d30_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103085(.data_in(wire_d30_84),.data_out(wire_d30_85),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103086(.data_in(wire_d30_85),.data_out(wire_d30_86),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103087(.data_in(wire_d30_86),.data_out(wire_d30_87),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103088(.data_in(wire_d30_87),.data_out(wire_d30_88),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103089(.data_in(wire_d30_88),.data_out(wire_d30_89),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103090(.data_in(wire_d30_89),.data_out(wire_d30_90),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103091(.data_in(wire_d30_90),.data_out(wire_d30_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3103092(.data_in(wire_d30_91),.data_out(wire_d30_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103093(.data_in(wire_d30_92),.data_out(wire_d30_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3103094(.data_in(wire_d30_93),.data_out(wire_d30_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3103095(.data_in(wire_d30_94),.data_out(wire_d30_95),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103096(.data_in(wire_d30_95),.data_out(wire_d30_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3103097(.data_in(wire_d30_96),.data_out(wire_d30_97),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103098(.data_in(wire_d30_97),.data_out(wire_d30_98),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103099(.data_in(wire_d30_98),.data_out(wire_d30_99),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance31030100(.data_in(wire_d30_99),.data_out(wire_d30_100),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance31030101(.data_in(wire_d30_100),.data_out(wire_d30_101),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance31030102(.data_in(wire_d30_101),.data_out(wire_d30_102),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance31030103(.data_in(wire_d30_102),.data_out(wire_d30_103),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance31030104(.data_in(wire_d30_103),.data_out(wire_d30_104),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance31030105(.data_in(wire_d30_104),.data_out(wire_d30_105),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance31030106(.data_in(wire_d30_105),.data_out(wire_d30_106),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance31030107(.data_in(wire_d30_106),.data_out(wire_d30_107),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance31030108(.data_in(wire_d30_107),.data_out(wire_d30_108),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance31030109(.data_in(wire_d30_108),.data_out(wire_d30_109),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance31030110(.data_in(wire_d30_109),.data_out(wire_d30_110),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance31030111(.data_in(wire_d30_110),.data_out(wire_d30_111),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance31030112(.data_in(wire_d30_111),.data_out(wire_d30_112),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance31030113(.data_in(wire_d30_112),.data_out(wire_d30_113),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance31030114(.data_in(wire_d30_113),.data_out(wire_d30_114),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance31030115(.data_in(wire_d30_114),.data_out(wire_d30_115),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance31030116(.data_in(wire_d30_115),.data_out(wire_d30_116),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance31030117(.data_in(wire_d30_116),.data_out(wire_d30_117),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance31030118(.data_in(wire_d30_117),.data_out(wire_d30_118),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance31030119(.data_in(wire_d30_118),.data_out(d_out30),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance320310(.data_in(d_in31),.data_out(wire_d31_0),.clk(clk),.rst(rst));            //channel 32
	large_mux #(.WIDTH(WIDTH)) large_mux_instance320311(.data_in(wire_d31_0),.data_out(wire_d31_1),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance320312(.data_in(wire_d31_1),.data_out(wire_d31_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance320313(.data_in(wire_d31_2),.data_out(wire_d31_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance320314(.data_in(wire_d31_3),.data_out(wire_d31_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance320315(.data_in(wire_d31_4),.data_out(wire_d31_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance320316(.data_in(wire_d31_5),.data_out(wire_d31_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance320317(.data_in(wire_d31_6),.data_out(wire_d31_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance320318(.data_in(wire_d31_7),.data_out(wire_d31_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance320319(.data_in(wire_d31_8),.data_out(wire_d31_9),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3203110(.data_in(wire_d31_9),.data_out(wire_d31_10),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3203111(.data_in(wire_d31_10),.data_out(wire_d31_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203112(.data_in(wire_d31_11),.data_out(wire_d31_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203113(.data_in(wire_d31_12),.data_out(wire_d31_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203114(.data_in(wire_d31_13),.data_out(wire_d31_14),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203115(.data_in(wire_d31_14),.data_out(wire_d31_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203116(.data_in(wire_d31_15),.data_out(wire_d31_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203117(.data_in(wire_d31_16),.data_out(wire_d31_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203118(.data_in(wire_d31_17),.data_out(wire_d31_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203119(.data_in(wire_d31_18),.data_out(wire_d31_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203120(.data_in(wire_d31_19),.data_out(wire_d31_20),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203121(.data_in(wire_d31_20),.data_out(wire_d31_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203122(.data_in(wire_d31_21),.data_out(wire_d31_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203123(.data_in(wire_d31_22),.data_out(wire_d31_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203124(.data_in(wire_d31_23),.data_out(wire_d31_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203125(.data_in(wire_d31_24),.data_out(wire_d31_25),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3203126(.data_in(wire_d31_25),.data_out(wire_d31_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203127(.data_in(wire_d31_26),.data_out(wire_d31_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203128(.data_in(wire_d31_27),.data_out(wire_d31_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3203129(.data_in(wire_d31_28),.data_out(wire_d31_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203130(.data_in(wire_d31_29),.data_out(wire_d31_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3203131(.data_in(wire_d31_30),.data_out(wire_d31_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203132(.data_in(wire_d31_31),.data_out(wire_d31_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203133(.data_in(wire_d31_32),.data_out(wire_d31_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203134(.data_in(wire_d31_33),.data_out(wire_d31_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203135(.data_in(wire_d31_34),.data_out(wire_d31_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203136(.data_in(wire_d31_35),.data_out(wire_d31_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203137(.data_in(wire_d31_36),.data_out(wire_d31_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203138(.data_in(wire_d31_37),.data_out(wire_d31_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203139(.data_in(wire_d31_38),.data_out(wire_d31_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203140(.data_in(wire_d31_39),.data_out(wire_d31_40),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203141(.data_in(wire_d31_40),.data_out(wire_d31_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203142(.data_in(wire_d31_41),.data_out(wire_d31_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203143(.data_in(wire_d31_42),.data_out(wire_d31_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203144(.data_in(wire_d31_43),.data_out(wire_d31_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203145(.data_in(wire_d31_44),.data_out(wire_d31_45),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3203146(.data_in(wire_d31_45),.data_out(wire_d31_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3203147(.data_in(wire_d31_46),.data_out(wire_d31_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203148(.data_in(wire_d31_47),.data_out(wire_d31_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3203149(.data_in(wire_d31_48),.data_out(wire_d31_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203150(.data_in(wire_d31_49),.data_out(wire_d31_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203151(.data_in(wire_d31_50),.data_out(wire_d31_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203152(.data_in(wire_d31_51),.data_out(wire_d31_52),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3203153(.data_in(wire_d31_52),.data_out(wire_d31_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203154(.data_in(wire_d31_53),.data_out(wire_d31_54),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203155(.data_in(wire_d31_54),.data_out(wire_d31_55),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3203156(.data_in(wire_d31_55),.data_out(wire_d31_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203157(.data_in(wire_d31_56),.data_out(wire_d31_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203158(.data_in(wire_d31_57),.data_out(wire_d31_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203159(.data_in(wire_d31_58),.data_out(wire_d31_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203160(.data_in(wire_d31_59),.data_out(wire_d31_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3203161(.data_in(wire_d31_60),.data_out(wire_d31_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3203162(.data_in(wire_d31_61),.data_out(wire_d31_62),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203163(.data_in(wire_d31_62),.data_out(wire_d31_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203164(.data_in(wire_d31_63),.data_out(wire_d31_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203165(.data_in(wire_d31_64),.data_out(wire_d31_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203166(.data_in(wire_d31_65),.data_out(wire_d31_66),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3203167(.data_in(wire_d31_66),.data_out(wire_d31_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203168(.data_in(wire_d31_67),.data_out(wire_d31_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3203169(.data_in(wire_d31_68),.data_out(wire_d31_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203170(.data_in(wire_d31_69),.data_out(wire_d31_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203171(.data_in(wire_d31_70),.data_out(wire_d31_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203172(.data_in(wire_d31_71),.data_out(wire_d31_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3203173(.data_in(wire_d31_72),.data_out(wire_d31_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203174(.data_in(wire_d31_73),.data_out(wire_d31_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203175(.data_in(wire_d31_74),.data_out(wire_d31_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203176(.data_in(wire_d31_75),.data_out(wire_d31_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203177(.data_in(wire_d31_76),.data_out(wire_d31_77),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203178(.data_in(wire_d31_77),.data_out(wire_d31_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3203179(.data_in(wire_d31_78),.data_out(wire_d31_79),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203180(.data_in(wire_d31_79),.data_out(wire_d31_80),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203181(.data_in(wire_d31_80),.data_out(wire_d31_81),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203182(.data_in(wire_d31_81),.data_out(wire_d31_82),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203183(.data_in(wire_d31_82),.data_out(wire_d31_83),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3203184(.data_in(wire_d31_83),.data_out(wire_d31_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3203185(.data_in(wire_d31_84),.data_out(wire_d31_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3203186(.data_in(wire_d31_85),.data_out(wire_d31_86),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203187(.data_in(wire_d31_86),.data_out(wire_d31_87),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203188(.data_in(wire_d31_87),.data_out(wire_d31_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203189(.data_in(wire_d31_88),.data_out(wire_d31_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3203190(.data_in(wire_d31_89),.data_out(wire_d31_90),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203191(.data_in(wire_d31_90),.data_out(wire_d31_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203192(.data_in(wire_d31_91),.data_out(wire_d31_92),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203193(.data_in(wire_d31_92),.data_out(wire_d31_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203194(.data_in(wire_d31_93),.data_out(wire_d31_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3203195(.data_in(wire_d31_94),.data_out(wire_d31_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3203196(.data_in(wire_d31_95),.data_out(wire_d31_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203197(.data_in(wire_d31_96),.data_out(wire_d31_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3203198(.data_in(wire_d31_97),.data_out(wire_d31_98),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203199(.data_in(wire_d31_98),.data_out(wire_d31_99),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance32031100(.data_in(wire_d31_99),.data_out(wire_d31_100),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance32031101(.data_in(wire_d31_100),.data_out(wire_d31_101),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance32031102(.data_in(wire_d31_101),.data_out(wire_d31_102),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance32031103(.data_in(wire_d31_102),.data_out(wire_d31_103),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance32031104(.data_in(wire_d31_103),.data_out(wire_d31_104),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance32031105(.data_in(wire_d31_104),.data_out(wire_d31_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32031106(.data_in(wire_d31_105),.data_out(wire_d31_106),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance32031107(.data_in(wire_d31_106),.data_out(wire_d31_107),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance32031108(.data_in(wire_d31_107),.data_out(wire_d31_108),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance32031109(.data_in(wire_d31_108),.data_out(wire_d31_109),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance32031110(.data_in(wire_d31_109),.data_out(wire_d31_110),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance32031111(.data_in(wire_d31_110),.data_out(wire_d31_111),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32031112(.data_in(wire_d31_111),.data_out(wire_d31_112),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance32031113(.data_in(wire_d31_112),.data_out(wire_d31_113),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance32031114(.data_in(wire_d31_113),.data_out(wire_d31_114),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance32031115(.data_in(wire_d31_114),.data_out(wire_d31_115),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance32031116(.data_in(wire_d31_115),.data_out(wire_d31_116),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance32031117(.data_in(wire_d31_116),.data_out(wire_d31_117),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance32031118(.data_in(wire_d31_117),.data_out(wire_d31_118),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance32031119(.data_in(wire_d31_118),.data_out(d_out31),.clk(clk),.rst(rst));

	large_adder #(.WIDTH(WIDTH)) large_adder_instance330320(.data_in(d_in32),.data_out(wire_d32_0),.clk(clk),.rst(rst));            //channel 33
	large_adder #(.WIDTH(WIDTH)) large_adder_instance330321(.data_in(wire_d32_0),.data_out(wire_d32_1),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance330322(.data_in(wire_d32_1),.data_out(wire_d32_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance330323(.data_in(wire_d32_2),.data_out(wire_d32_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance330324(.data_in(wire_d32_3),.data_out(wire_d32_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance330325(.data_in(wire_d32_4),.data_out(wire_d32_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance330326(.data_in(wire_d32_5),.data_out(wire_d32_6),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance330327(.data_in(wire_d32_6),.data_out(wire_d32_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance330328(.data_in(wire_d32_7),.data_out(wire_d32_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance330329(.data_in(wire_d32_8),.data_out(wire_d32_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303210(.data_in(wire_d32_9),.data_out(wire_d32_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3303211(.data_in(wire_d32_10),.data_out(wire_d32_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303212(.data_in(wire_d32_11),.data_out(wire_d32_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303213(.data_in(wire_d32_12),.data_out(wire_d32_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3303214(.data_in(wire_d32_13),.data_out(wire_d32_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3303215(.data_in(wire_d32_14),.data_out(wire_d32_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3303216(.data_in(wire_d32_15),.data_out(wire_d32_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303217(.data_in(wire_d32_16),.data_out(wire_d32_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303218(.data_in(wire_d32_17),.data_out(wire_d32_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303219(.data_in(wire_d32_18),.data_out(wire_d32_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303220(.data_in(wire_d32_19),.data_out(wire_d32_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303221(.data_in(wire_d32_20),.data_out(wire_d32_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303222(.data_in(wire_d32_21),.data_out(wire_d32_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303223(.data_in(wire_d32_22),.data_out(wire_d32_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303224(.data_in(wire_d32_23),.data_out(wire_d32_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303225(.data_in(wire_d32_24),.data_out(wire_d32_25),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3303226(.data_in(wire_d32_25),.data_out(wire_d32_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303227(.data_in(wire_d32_26),.data_out(wire_d32_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303228(.data_in(wire_d32_27),.data_out(wire_d32_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303229(.data_in(wire_d32_28),.data_out(wire_d32_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303230(.data_in(wire_d32_29),.data_out(wire_d32_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303231(.data_in(wire_d32_30),.data_out(wire_d32_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3303232(.data_in(wire_d32_31),.data_out(wire_d32_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3303233(.data_in(wire_d32_32),.data_out(wire_d32_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303234(.data_in(wire_d32_33),.data_out(wire_d32_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303235(.data_in(wire_d32_34),.data_out(wire_d32_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303236(.data_in(wire_d32_35),.data_out(wire_d32_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303237(.data_in(wire_d32_36),.data_out(wire_d32_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3303238(.data_in(wire_d32_37),.data_out(wire_d32_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303239(.data_in(wire_d32_38),.data_out(wire_d32_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303240(.data_in(wire_d32_39),.data_out(wire_d32_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303241(.data_in(wire_d32_40),.data_out(wire_d32_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303242(.data_in(wire_d32_41),.data_out(wire_d32_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3303243(.data_in(wire_d32_42),.data_out(wire_d32_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303244(.data_in(wire_d32_43),.data_out(wire_d32_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3303245(.data_in(wire_d32_44),.data_out(wire_d32_45),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303246(.data_in(wire_d32_45),.data_out(wire_d32_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3303247(.data_in(wire_d32_46),.data_out(wire_d32_47),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303248(.data_in(wire_d32_47),.data_out(wire_d32_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303249(.data_in(wire_d32_48),.data_out(wire_d32_49),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3303250(.data_in(wire_d32_49),.data_out(wire_d32_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303251(.data_in(wire_d32_50),.data_out(wire_d32_51),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303252(.data_in(wire_d32_51),.data_out(wire_d32_52),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3303253(.data_in(wire_d32_52),.data_out(wire_d32_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303254(.data_in(wire_d32_53),.data_out(wire_d32_54),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3303255(.data_in(wire_d32_54),.data_out(wire_d32_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303256(.data_in(wire_d32_55),.data_out(wire_d32_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303257(.data_in(wire_d32_56),.data_out(wire_d32_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303258(.data_in(wire_d32_57),.data_out(wire_d32_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303259(.data_in(wire_d32_58),.data_out(wire_d32_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303260(.data_in(wire_d32_59),.data_out(wire_d32_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303261(.data_in(wire_d32_60),.data_out(wire_d32_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303262(.data_in(wire_d32_61),.data_out(wire_d32_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303263(.data_in(wire_d32_62),.data_out(wire_d32_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3303264(.data_in(wire_d32_63),.data_out(wire_d32_64),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303265(.data_in(wire_d32_64),.data_out(wire_d32_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3303266(.data_in(wire_d32_65),.data_out(wire_d32_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303267(.data_in(wire_d32_66),.data_out(wire_d32_67),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3303268(.data_in(wire_d32_67),.data_out(wire_d32_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3303269(.data_in(wire_d32_68),.data_out(wire_d32_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3303270(.data_in(wire_d32_69),.data_out(wire_d32_70),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303271(.data_in(wire_d32_70),.data_out(wire_d32_71),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303272(.data_in(wire_d32_71),.data_out(wire_d32_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303273(.data_in(wire_d32_72),.data_out(wire_d32_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303274(.data_in(wire_d32_73),.data_out(wire_d32_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303275(.data_in(wire_d32_74),.data_out(wire_d32_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3303276(.data_in(wire_d32_75),.data_out(wire_d32_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3303277(.data_in(wire_d32_76),.data_out(wire_d32_77),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3303278(.data_in(wire_d32_77),.data_out(wire_d32_78),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303279(.data_in(wire_d32_78),.data_out(wire_d32_79),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303280(.data_in(wire_d32_79),.data_out(wire_d32_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3303281(.data_in(wire_d32_80),.data_out(wire_d32_81),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303282(.data_in(wire_d32_81),.data_out(wire_d32_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303283(.data_in(wire_d32_82),.data_out(wire_d32_83),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303284(.data_in(wire_d32_83),.data_out(wire_d32_84),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303285(.data_in(wire_d32_84),.data_out(wire_d32_85),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303286(.data_in(wire_d32_85),.data_out(wire_d32_86),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303287(.data_in(wire_d32_86),.data_out(wire_d32_87),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303288(.data_in(wire_d32_87),.data_out(wire_d32_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3303289(.data_in(wire_d32_88),.data_out(wire_d32_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3303290(.data_in(wire_d32_89),.data_out(wire_d32_90),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303291(.data_in(wire_d32_90),.data_out(wire_d32_91),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303292(.data_in(wire_d32_91),.data_out(wire_d32_92),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303293(.data_in(wire_d32_92),.data_out(wire_d32_93),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303294(.data_in(wire_d32_93),.data_out(wire_d32_94),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303295(.data_in(wire_d32_94),.data_out(wire_d32_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3303296(.data_in(wire_d32_95),.data_out(wire_d32_96),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3303297(.data_in(wire_d32_96),.data_out(wire_d32_97),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303298(.data_in(wire_d32_97),.data_out(wire_d32_98),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3303299(.data_in(wire_d32_98),.data_out(wire_d32_99),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance33032100(.data_in(wire_d32_99),.data_out(wire_d32_100),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance33032101(.data_in(wire_d32_100),.data_out(wire_d32_101),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance33032102(.data_in(wire_d32_101),.data_out(wire_d32_102),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance33032103(.data_in(wire_d32_102),.data_out(wire_d32_103),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance33032104(.data_in(wire_d32_103),.data_out(wire_d32_104),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance33032105(.data_in(wire_d32_104),.data_out(wire_d32_105),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance33032106(.data_in(wire_d32_105),.data_out(wire_d32_106),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance33032107(.data_in(wire_d32_106),.data_out(wire_d32_107),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance33032108(.data_in(wire_d32_107),.data_out(wire_d32_108),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance33032109(.data_in(wire_d32_108),.data_out(wire_d32_109),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance33032110(.data_in(wire_d32_109),.data_out(wire_d32_110),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance33032111(.data_in(wire_d32_110),.data_out(wire_d32_111),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance33032112(.data_in(wire_d32_111),.data_out(wire_d32_112),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance33032113(.data_in(wire_d32_112),.data_out(wire_d32_113),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance33032114(.data_in(wire_d32_113),.data_out(wire_d32_114),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance33032115(.data_in(wire_d32_114),.data_out(wire_d32_115),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance33032116(.data_in(wire_d32_115),.data_out(wire_d32_116),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance33032117(.data_in(wire_d32_116),.data_out(wire_d32_117),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance33032118(.data_in(wire_d32_117),.data_out(wire_d32_118),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance33032119(.data_in(wire_d32_118),.data_out(d_out32),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance340330(.data_in(d_in33),.data_out(wire_d33_0),.clk(clk),.rst(rst));            //channel 34
	large_adder #(.WIDTH(WIDTH)) large_adder_instance340331(.data_in(wire_d33_0),.data_out(wire_d33_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance340332(.data_in(wire_d33_1),.data_out(wire_d33_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance340333(.data_in(wire_d33_2),.data_out(wire_d33_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance340334(.data_in(wire_d33_3),.data_out(wire_d33_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance340335(.data_in(wire_d33_4),.data_out(wire_d33_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance340336(.data_in(wire_d33_5),.data_out(wire_d33_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance340337(.data_in(wire_d33_6),.data_out(wire_d33_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance340338(.data_in(wire_d33_7),.data_out(wire_d33_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance340339(.data_in(wire_d33_8),.data_out(wire_d33_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3403310(.data_in(wire_d33_9),.data_out(wire_d33_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403311(.data_in(wire_d33_10),.data_out(wire_d33_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3403312(.data_in(wire_d33_11),.data_out(wire_d33_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3403313(.data_in(wire_d33_12),.data_out(wire_d33_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403314(.data_in(wire_d33_13),.data_out(wire_d33_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403315(.data_in(wire_d33_14),.data_out(wire_d33_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403316(.data_in(wire_d33_15),.data_out(wire_d33_16),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3403317(.data_in(wire_d33_16),.data_out(wire_d33_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403318(.data_in(wire_d33_17),.data_out(wire_d33_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403319(.data_in(wire_d33_18),.data_out(wire_d33_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3403320(.data_in(wire_d33_19),.data_out(wire_d33_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3403321(.data_in(wire_d33_20),.data_out(wire_d33_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3403322(.data_in(wire_d33_21),.data_out(wire_d33_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403323(.data_in(wire_d33_22),.data_out(wire_d33_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403324(.data_in(wire_d33_23),.data_out(wire_d33_24),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3403325(.data_in(wire_d33_24),.data_out(wire_d33_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3403326(.data_in(wire_d33_25),.data_out(wire_d33_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3403327(.data_in(wire_d33_26),.data_out(wire_d33_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3403328(.data_in(wire_d33_27),.data_out(wire_d33_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3403329(.data_in(wire_d33_28),.data_out(wire_d33_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403330(.data_in(wire_d33_29),.data_out(wire_d33_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403331(.data_in(wire_d33_30),.data_out(wire_d33_31),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3403332(.data_in(wire_d33_31),.data_out(wire_d33_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403333(.data_in(wire_d33_32),.data_out(wire_d33_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403334(.data_in(wire_d33_33),.data_out(wire_d33_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3403335(.data_in(wire_d33_34),.data_out(wire_d33_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3403336(.data_in(wire_d33_35),.data_out(wire_d33_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403337(.data_in(wire_d33_36),.data_out(wire_d33_37),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3403338(.data_in(wire_d33_37),.data_out(wire_d33_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3403339(.data_in(wire_d33_38),.data_out(wire_d33_39),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3403340(.data_in(wire_d33_39),.data_out(wire_d33_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403341(.data_in(wire_d33_40),.data_out(wire_d33_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403342(.data_in(wire_d33_41),.data_out(wire_d33_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403343(.data_in(wire_d33_42),.data_out(wire_d33_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403344(.data_in(wire_d33_43),.data_out(wire_d33_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403345(.data_in(wire_d33_44),.data_out(wire_d33_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403346(.data_in(wire_d33_45),.data_out(wire_d33_46),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3403347(.data_in(wire_d33_46),.data_out(wire_d33_47),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3403348(.data_in(wire_d33_47),.data_out(wire_d33_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403349(.data_in(wire_d33_48),.data_out(wire_d33_49),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3403350(.data_in(wire_d33_49),.data_out(wire_d33_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3403351(.data_in(wire_d33_50),.data_out(wire_d33_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3403352(.data_in(wire_d33_51),.data_out(wire_d33_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3403353(.data_in(wire_d33_52),.data_out(wire_d33_53),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3403354(.data_in(wire_d33_53),.data_out(wire_d33_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3403355(.data_in(wire_d33_54),.data_out(wire_d33_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403356(.data_in(wire_d33_55),.data_out(wire_d33_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403357(.data_in(wire_d33_56),.data_out(wire_d33_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403358(.data_in(wire_d33_57),.data_out(wire_d33_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3403359(.data_in(wire_d33_58),.data_out(wire_d33_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403360(.data_in(wire_d33_59),.data_out(wire_d33_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3403361(.data_in(wire_d33_60),.data_out(wire_d33_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3403362(.data_in(wire_d33_61),.data_out(wire_d33_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403363(.data_in(wire_d33_62),.data_out(wire_d33_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3403364(.data_in(wire_d33_63),.data_out(wire_d33_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403365(.data_in(wire_d33_64),.data_out(wire_d33_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3403366(.data_in(wire_d33_65),.data_out(wire_d33_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3403367(.data_in(wire_d33_66),.data_out(wire_d33_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3403368(.data_in(wire_d33_67),.data_out(wire_d33_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403369(.data_in(wire_d33_68),.data_out(wire_d33_69),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3403370(.data_in(wire_d33_69),.data_out(wire_d33_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3403371(.data_in(wire_d33_70),.data_out(wire_d33_71),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403372(.data_in(wire_d33_71),.data_out(wire_d33_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3403373(.data_in(wire_d33_72),.data_out(wire_d33_73),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403374(.data_in(wire_d33_73),.data_out(wire_d33_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403375(.data_in(wire_d33_74),.data_out(wire_d33_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3403376(.data_in(wire_d33_75),.data_out(wire_d33_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3403377(.data_in(wire_d33_76),.data_out(wire_d33_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3403378(.data_in(wire_d33_77),.data_out(wire_d33_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3403379(.data_in(wire_d33_78),.data_out(wire_d33_79),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403380(.data_in(wire_d33_79),.data_out(wire_d33_80),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403381(.data_in(wire_d33_80),.data_out(wire_d33_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3403382(.data_in(wire_d33_81),.data_out(wire_d33_82),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403383(.data_in(wire_d33_82),.data_out(wire_d33_83),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403384(.data_in(wire_d33_83),.data_out(wire_d33_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3403385(.data_in(wire_d33_84),.data_out(wire_d33_85),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403386(.data_in(wire_d33_85),.data_out(wire_d33_86),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3403387(.data_in(wire_d33_86),.data_out(wire_d33_87),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3403388(.data_in(wire_d33_87),.data_out(wire_d33_88),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403389(.data_in(wire_d33_88),.data_out(wire_d33_89),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403390(.data_in(wire_d33_89),.data_out(wire_d33_90),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3403391(.data_in(wire_d33_90),.data_out(wire_d33_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3403392(.data_in(wire_d33_91),.data_out(wire_d33_92),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3403393(.data_in(wire_d33_92),.data_out(wire_d33_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3403394(.data_in(wire_d33_93),.data_out(wire_d33_94),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3403395(.data_in(wire_d33_94),.data_out(wire_d33_95),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3403396(.data_in(wire_d33_95),.data_out(wire_d33_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3403397(.data_in(wire_d33_96),.data_out(wire_d33_97),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3403398(.data_in(wire_d33_97),.data_out(wire_d33_98),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3403399(.data_in(wire_d33_98),.data_out(wire_d33_99),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance34033100(.data_in(wire_d33_99),.data_out(wire_d33_100),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance34033101(.data_in(wire_d33_100),.data_out(wire_d33_101),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance34033102(.data_in(wire_d33_101),.data_out(wire_d33_102),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance34033103(.data_in(wire_d33_102),.data_out(wire_d33_103),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance34033104(.data_in(wire_d33_103),.data_out(wire_d33_104),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance34033105(.data_in(wire_d33_104),.data_out(wire_d33_105),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance34033106(.data_in(wire_d33_105),.data_out(wire_d33_106),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance34033107(.data_in(wire_d33_106),.data_out(wire_d33_107),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance34033108(.data_in(wire_d33_107),.data_out(wire_d33_108),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance34033109(.data_in(wire_d33_108),.data_out(wire_d33_109),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance34033110(.data_in(wire_d33_109),.data_out(wire_d33_110),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance34033111(.data_in(wire_d33_110),.data_out(wire_d33_111),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance34033112(.data_in(wire_d33_111),.data_out(wire_d33_112),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance34033113(.data_in(wire_d33_112),.data_out(wire_d33_113),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance34033114(.data_in(wire_d33_113),.data_out(wire_d33_114),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance34033115(.data_in(wire_d33_114),.data_out(wire_d33_115),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance34033116(.data_in(wire_d33_115),.data_out(wire_d33_116),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance34033117(.data_in(wire_d33_116),.data_out(wire_d33_117),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance34033118(.data_in(wire_d33_117),.data_out(wire_d33_118),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance34033119(.data_in(wire_d33_118),.data_out(d_out33),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance350340(.data_in(d_in34),.data_out(wire_d34_0),.clk(clk),.rst(rst));            //channel 35
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance350341(.data_in(wire_d34_0),.data_out(wire_d34_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance350342(.data_in(wire_d34_1),.data_out(wire_d34_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance350343(.data_in(wire_d34_2),.data_out(wire_d34_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance350344(.data_in(wire_d34_3),.data_out(wire_d34_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance350345(.data_in(wire_d34_4),.data_out(wire_d34_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance350346(.data_in(wire_d34_5),.data_out(wire_d34_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance350347(.data_in(wire_d34_6),.data_out(wire_d34_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance350348(.data_in(wire_d34_7),.data_out(wire_d34_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance350349(.data_in(wire_d34_8),.data_out(wire_d34_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503410(.data_in(wire_d34_9),.data_out(wire_d34_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503411(.data_in(wire_d34_10),.data_out(wire_d34_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503412(.data_in(wire_d34_11),.data_out(wire_d34_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503413(.data_in(wire_d34_12),.data_out(wire_d34_13),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3503414(.data_in(wire_d34_13),.data_out(wire_d34_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503415(.data_in(wire_d34_14),.data_out(wire_d34_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503416(.data_in(wire_d34_15),.data_out(wire_d34_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503417(.data_in(wire_d34_16),.data_out(wire_d34_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503418(.data_in(wire_d34_17),.data_out(wire_d34_18),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503419(.data_in(wire_d34_18),.data_out(wire_d34_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503420(.data_in(wire_d34_19),.data_out(wire_d34_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3503421(.data_in(wire_d34_20),.data_out(wire_d34_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3503422(.data_in(wire_d34_21),.data_out(wire_d34_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3503423(.data_in(wire_d34_22),.data_out(wire_d34_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3503424(.data_in(wire_d34_23),.data_out(wire_d34_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503425(.data_in(wire_d34_24),.data_out(wire_d34_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503426(.data_in(wire_d34_25),.data_out(wire_d34_26),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3503427(.data_in(wire_d34_26),.data_out(wire_d34_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503428(.data_in(wire_d34_27),.data_out(wire_d34_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503429(.data_in(wire_d34_28),.data_out(wire_d34_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3503430(.data_in(wire_d34_29),.data_out(wire_d34_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503431(.data_in(wire_d34_30),.data_out(wire_d34_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503432(.data_in(wire_d34_31),.data_out(wire_d34_32),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3503433(.data_in(wire_d34_32),.data_out(wire_d34_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503434(.data_in(wire_d34_33),.data_out(wire_d34_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3503435(.data_in(wire_d34_34),.data_out(wire_d34_35),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3503436(.data_in(wire_d34_35),.data_out(wire_d34_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3503437(.data_in(wire_d34_36),.data_out(wire_d34_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503438(.data_in(wire_d34_37),.data_out(wire_d34_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503439(.data_in(wire_d34_38),.data_out(wire_d34_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503440(.data_in(wire_d34_39),.data_out(wire_d34_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503441(.data_in(wire_d34_40),.data_out(wire_d34_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503442(.data_in(wire_d34_41),.data_out(wire_d34_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503443(.data_in(wire_d34_42),.data_out(wire_d34_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503444(.data_in(wire_d34_43),.data_out(wire_d34_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503445(.data_in(wire_d34_44),.data_out(wire_d34_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503446(.data_in(wire_d34_45),.data_out(wire_d34_46),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3503447(.data_in(wire_d34_46),.data_out(wire_d34_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503448(.data_in(wire_d34_47),.data_out(wire_d34_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503449(.data_in(wire_d34_48),.data_out(wire_d34_49),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503450(.data_in(wire_d34_49),.data_out(wire_d34_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503451(.data_in(wire_d34_50),.data_out(wire_d34_51),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503452(.data_in(wire_d34_51),.data_out(wire_d34_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3503453(.data_in(wire_d34_52),.data_out(wire_d34_53),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503454(.data_in(wire_d34_53),.data_out(wire_d34_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503455(.data_in(wire_d34_54),.data_out(wire_d34_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503456(.data_in(wire_d34_55),.data_out(wire_d34_56),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503457(.data_in(wire_d34_56),.data_out(wire_d34_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503458(.data_in(wire_d34_57),.data_out(wire_d34_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503459(.data_in(wire_d34_58),.data_out(wire_d34_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3503460(.data_in(wire_d34_59),.data_out(wire_d34_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503461(.data_in(wire_d34_60),.data_out(wire_d34_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503462(.data_in(wire_d34_61),.data_out(wire_d34_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3503463(.data_in(wire_d34_62),.data_out(wire_d34_63),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3503464(.data_in(wire_d34_63),.data_out(wire_d34_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503465(.data_in(wire_d34_64),.data_out(wire_d34_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503466(.data_in(wire_d34_65),.data_out(wire_d34_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503467(.data_in(wire_d34_66),.data_out(wire_d34_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3503468(.data_in(wire_d34_67),.data_out(wire_d34_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503469(.data_in(wire_d34_68),.data_out(wire_d34_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503470(.data_in(wire_d34_69),.data_out(wire_d34_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503471(.data_in(wire_d34_70),.data_out(wire_d34_71),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3503472(.data_in(wire_d34_71),.data_out(wire_d34_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3503473(.data_in(wire_d34_72),.data_out(wire_d34_73),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503474(.data_in(wire_d34_73),.data_out(wire_d34_74),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503475(.data_in(wire_d34_74),.data_out(wire_d34_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503476(.data_in(wire_d34_75),.data_out(wire_d34_76),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503477(.data_in(wire_d34_76),.data_out(wire_d34_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503478(.data_in(wire_d34_77),.data_out(wire_d34_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503479(.data_in(wire_d34_78),.data_out(wire_d34_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3503480(.data_in(wire_d34_79),.data_out(wire_d34_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3503481(.data_in(wire_d34_80),.data_out(wire_d34_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3503482(.data_in(wire_d34_81),.data_out(wire_d34_82),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3503483(.data_in(wire_d34_82),.data_out(wire_d34_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503484(.data_in(wire_d34_83),.data_out(wire_d34_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3503485(.data_in(wire_d34_84),.data_out(wire_d34_85),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503486(.data_in(wire_d34_85),.data_out(wire_d34_86),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503487(.data_in(wire_d34_86),.data_out(wire_d34_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3503488(.data_in(wire_d34_87),.data_out(wire_d34_88),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503489(.data_in(wire_d34_88),.data_out(wire_d34_89),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503490(.data_in(wire_d34_89),.data_out(wire_d34_90),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503491(.data_in(wire_d34_90),.data_out(wire_d34_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3503492(.data_in(wire_d34_91),.data_out(wire_d34_92),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3503493(.data_in(wire_d34_92),.data_out(wire_d34_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3503494(.data_in(wire_d34_93),.data_out(wire_d34_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3503495(.data_in(wire_d34_94),.data_out(wire_d34_95),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503496(.data_in(wire_d34_95),.data_out(wire_d34_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3503497(.data_in(wire_d34_96),.data_out(wire_d34_97),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503498(.data_in(wire_d34_97),.data_out(wire_d34_98),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503499(.data_in(wire_d34_98),.data_out(wire_d34_99),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance35034100(.data_in(wire_d34_99),.data_out(wire_d34_100),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance35034101(.data_in(wire_d34_100),.data_out(wire_d34_101),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance35034102(.data_in(wire_d34_101),.data_out(wire_d34_102),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance35034103(.data_in(wire_d34_102),.data_out(wire_d34_103),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance35034104(.data_in(wire_d34_103),.data_out(wire_d34_104),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance35034105(.data_in(wire_d34_104),.data_out(wire_d34_105),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance35034106(.data_in(wire_d34_105),.data_out(wire_d34_106),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance35034107(.data_in(wire_d34_106),.data_out(wire_d34_107),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance35034108(.data_in(wire_d34_107),.data_out(wire_d34_108),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance35034109(.data_in(wire_d34_108),.data_out(wire_d34_109),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance35034110(.data_in(wire_d34_109),.data_out(wire_d34_110),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance35034111(.data_in(wire_d34_110),.data_out(wire_d34_111),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance35034112(.data_in(wire_d34_111),.data_out(wire_d34_112),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance35034113(.data_in(wire_d34_112),.data_out(wire_d34_113),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance35034114(.data_in(wire_d34_113),.data_out(wire_d34_114),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance35034115(.data_in(wire_d34_114),.data_out(wire_d34_115),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance35034116(.data_in(wire_d34_115),.data_out(wire_d34_116),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance35034117(.data_in(wire_d34_116),.data_out(wire_d34_117),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance35034118(.data_in(wire_d34_117),.data_out(wire_d34_118),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance35034119(.data_in(wire_d34_118),.data_out(d_out34),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance360350(.data_in(d_in35),.data_out(wire_d35_0),.clk(clk),.rst(rst));            //channel 36
	invertion #(.WIDTH(WIDTH)) invertion_instance360351(.data_in(wire_d35_0),.data_out(wire_d35_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance360352(.data_in(wire_d35_1),.data_out(wire_d35_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance360353(.data_in(wire_d35_2),.data_out(wire_d35_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance360354(.data_in(wire_d35_3),.data_out(wire_d35_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance360355(.data_in(wire_d35_4),.data_out(wire_d35_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance360356(.data_in(wire_d35_5),.data_out(wire_d35_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance360357(.data_in(wire_d35_6),.data_out(wire_d35_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance360358(.data_in(wire_d35_7),.data_out(wire_d35_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance360359(.data_in(wire_d35_8),.data_out(wire_d35_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603510(.data_in(wire_d35_9),.data_out(wire_d35_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603511(.data_in(wire_d35_10),.data_out(wire_d35_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3603512(.data_in(wire_d35_11),.data_out(wire_d35_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603513(.data_in(wire_d35_12),.data_out(wire_d35_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603514(.data_in(wire_d35_13),.data_out(wire_d35_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603515(.data_in(wire_d35_14),.data_out(wire_d35_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603516(.data_in(wire_d35_15),.data_out(wire_d35_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3603517(.data_in(wire_d35_16),.data_out(wire_d35_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603518(.data_in(wire_d35_17),.data_out(wire_d35_18),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603519(.data_in(wire_d35_18),.data_out(wire_d35_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603520(.data_in(wire_d35_19),.data_out(wire_d35_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603521(.data_in(wire_d35_20),.data_out(wire_d35_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603522(.data_in(wire_d35_21),.data_out(wire_d35_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603523(.data_in(wire_d35_22),.data_out(wire_d35_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603524(.data_in(wire_d35_23),.data_out(wire_d35_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603525(.data_in(wire_d35_24),.data_out(wire_d35_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603526(.data_in(wire_d35_25),.data_out(wire_d35_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603527(.data_in(wire_d35_26),.data_out(wire_d35_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603528(.data_in(wire_d35_27),.data_out(wire_d35_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603529(.data_in(wire_d35_28),.data_out(wire_d35_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603530(.data_in(wire_d35_29),.data_out(wire_d35_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603531(.data_in(wire_d35_30),.data_out(wire_d35_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603532(.data_in(wire_d35_31),.data_out(wire_d35_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3603533(.data_in(wire_d35_32),.data_out(wire_d35_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3603534(.data_in(wire_d35_33),.data_out(wire_d35_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603535(.data_in(wire_d35_34),.data_out(wire_d35_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603536(.data_in(wire_d35_35),.data_out(wire_d35_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603537(.data_in(wire_d35_36),.data_out(wire_d35_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603538(.data_in(wire_d35_37),.data_out(wire_d35_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603539(.data_in(wire_d35_38),.data_out(wire_d35_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3603540(.data_in(wire_d35_39),.data_out(wire_d35_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3603541(.data_in(wire_d35_40),.data_out(wire_d35_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603542(.data_in(wire_d35_41),.data_out(wire_d35_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603543(.data_in(wire_d35_42),.data_out(wire_d35_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3603544(.data_in(wire_d35_43),.data_out(wire_d35_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603545(.data_in(wire_d35_44),.data_out(wire_d35_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603546(.data_in(wire_d35_45),.data_out(wire_d35_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603547(.data_in(wire_d35_46),.data_out(wire_d35_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603548(.data_in(wire_d35_47),.data_out(wire_d35_48),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3603549(.data_in(wire_d35_48),.data_out(wire_d35_49),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3603550(.data_in(wire_d35_49),.data_out(wire_d35_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3603551(.data_in(wire_d35_50),.data_out(wire_d35_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603552(.data_in(wire_d35_51),.data_out(wire_d35_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603553(.data_in(wire_d35_52),.data_out(wire_d35_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603554(.data_in(wire_d35_53),.data_out(wire_d35_54),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3603555(.data_in(wire_d35_54),.data_out(wire_d35_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603556(.data_in(wire_d35_55),.data_out(wire_d35_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603557(.data_in(wire_d35_56),.data_out(wire_d35_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603558(.data_in(wire_d35_57),.data_out(wire_d35_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603559(.data_in(wire_d35_58),.data_out(wire_d35_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603560(.data_in(wire_d35_59),.data_out(wire_d35_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603561(.data_in(wire_d35_60),.data_out(wire_d35_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603562(.data_in(wire_d35_61),.data_out(wire_d35_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603563(.data_in(wire_d35_62),.data_out(wire_d35_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603564(.data_in(wire_d35_63),.data_out(wire_d35_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603565(.data_in(wire_d35_64),.data_out(wire_d35_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603566(.data_in(wire_d35_65),.data_out(wire_d35_66),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603567(.data_in(wire_d35_66),.data_out(wire_d35_67),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603568(.data_in(wire_d35_67),.data_out(wire_d35_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3603569(.data_in(wire_d35_68),.data_out(wire_d35_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3603570(.data_in(wire_d35_69),.data_out(wire_d35_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603571(.data_in(wire_d35_70),.data_out(wire_d35_71),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603572(.data_in(wire_d35_71),.data_out(wire_d35_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603573(.data_in(wire_d35_72),.data_out(wire_d35_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603574(.data_in(wire_d35_73),.data_out(wire_d35_74),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603575(.data_in(wire_d35_74),.data_out(wire_d35_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3603576(.data_in(wire_d35_75),.data_out(wire_d35_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603577(.data_in(wire_d35_76),.data_out(wire_d35_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603578(.data_in(wire_d35_77),.data_out(wire_d35_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603579(.data_in(wire_d35_78),.data_out(wire_d35_79),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603580(.data_in(wire_d35_79),.data_out(wire_d35_80),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3603581(.data_in(wire_d35_80),.data_out(wire_d35_81),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603582(.data_in(wire_d35_81),.data_out(wire_d35_82),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603583(.data_in(wire_d35_82),.data_out(wire_d35_83),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3603584(.data_in(wire_d35_83),.data_out(wire_d35_84),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603585(.data_in(wire_d35_84),.data_out(wire_d35_85),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603586(.data_in(wire_d35_85),.data_out(wire_d35_86),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3603587(.data_in(wire_d35_86),.data_out(wire_d35_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3603588(.data_in(wire_d35_87),.data_out(wire_d35_88),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603589(.data_in(wire_d35_88),.data_out(wire_d35_89),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603590(.data_in(wire_d35_89),.data_out(wire_d35_90),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603591(.data_in(wire_d35_90),.data_out(wire_d35_91),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603592(.data_in(wire_d35_91),.data_out(wire_d35_92),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603593(.data_in(wire_d35_92),.data_out(wire_d35_93),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3603594(.data_in(wire_d35_93),.data_out(wire_d35_94),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603595(.data_in(wire_d35_94),.data_out(wire_d35_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3603596(.data_in(wire_d35_95),.data_out(wire_d35_96),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603597(.data_in(wire_d35_96),.data_out(wire_d35_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603598(.data_in(wire_d35_97),.data_out(wire_d35_98),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603599(.data_in(wire_d35_98),.data_out(wire_d35_99),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance36035100(.data_in(wire_d35_99),.data_out(wire_d35_100),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance36035101(.data_in(wire_d35_100),.data_out(wire_d35_101),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance36035102(.data_in(wire_d35_101),.data_out(wire_d35_102),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance36035103(.data_in(wire_d35_102),.data_out(wire_d35_103),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance36035104(.data_in(wire_d35_103),.data_out(wire_d35_104),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance36035105(.data_in(wire_d35_104),.data_out(wire_d35_105),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance36035106(.data_in(wire_d35_105),.data_out(wire_d35_106),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance36035107(.data_in(wire_d35_106),.data_out(wire_d35_107),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance36035108(.data_in(wire_d35_107),.data_out(wire_d35_108),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance36035109(.data_in(wire_d35_108),.data_out(wire_d35_109),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance36035110(.data_in(wire_d35_109),.data_out(wire_d35_110),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance36035111(.data_in(wire_d35_110),.data_out(wire_d35_111),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance36035112(.data_in(wire_d35_111),.data_out(wire_d35_112),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance36035113(.data_in(wire_d35_112),.data_out(wire_d35_113),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance36035114(.data_in(wire_d35_113),.data_out(wire_d35_114),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance36035115(.data_in(wire_d35_114),.data_out(wire_d35_115),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance36035116(.data_in(wire_d35_115),.data_out(wire_d35_116),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance36035117(.data_in(wire_d35_116),.data_out(wire_d35_117),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance36035118(.data_in(wire_d35_117),.data_out(wire_d35_118),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance36035119(.data_in(wire_d35_118),.data_out(d_out35),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance370360(.data_in(d_in36),.data_out(wire_d36_0),.clk(clk),.rst(rst));            //channel 37
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance370361(.data_in(wire_d36_0),.data_out(wire_d36_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance370362(.data_in(wire_d36_1),.data_out(wire_d36_2),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance370363(.data_in(wire_d36_2),.data_out(wire_d36_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance370364(.data_in(wire_d36_3),.data_out(wire_d36_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance370365(.data_in(wire_d36_4),.data_out(wire_d36_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance370366(.data_in(wire_d36_5),.data_out(wire_d36_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance370367(.data_in(wire_d36_6),.data_out(wire_d36_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance370368(.data_in(wire_d36_7),.data_out(wire_d36_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance370369(.data_in(wire_d36_8),.data_out(wire_d36_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703610(.data_in(wire_d36_9),.data_out(wire_d36_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3703611(.data_in(wire_d36_10),.data_out(wire_d36_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3703612(.data_in(wire_d36_11),.data_out(wire_d36_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703613(.data_in(wire_d36_12),.data_out(wire_d36_13),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3703614(.data_in(wire_d36_13),.data_out(wire_d36_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703615(.data_in(wire_d36_14),.data_out(wire_d36_15),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3703616(.data_in(wire_d36_15),.data_out(wire_d36_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3703617(.data_in(wire_d36_16),.data_out(wire_d36_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703618(.data_in(wire_d36_17),.data_out(wire_d36_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3703619(.data_in(wire_d36_18),.data_out(wire_d36_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703620(.data_in(wire_d36_19),.data_out(wire_d36_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3703621(.data_in(wire_d36_20),.data_out(wire_d36_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703622(.data_in(wire_d36_21),.data_out(wire_d36_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3703623(.data_in(wire_d36_22),.data_out(wire_d36_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3703624(.data_in(wire_d36_23),.data_out(wire_d36_24),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3703625(.data_in(wire_d36_24),.data_out(wire_d36_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703626(.data_in(wire_d36_25),.data_out(wire_d36_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3703627(.data_in(wire_d36_26),.data_out(wire_d36_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703628(.data_in(wire_d36_27),.data_out(wire_d36_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3703629(.data_in(wire_d36_28),.data_out(wire_d36_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703630(.data_in(wire_d36_29),.data_out(wire_d36_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3703631(.data_in(wire_d36_30),.data_out(wire_d36_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703632(.data_in(wire_d36_31),.data_out(wire_d36_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703633(.data_in(wire_d36_32),.data_out(wire_d36_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703634(.data_in(wire_d36_33),.data_out(wire_d36_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703635(.data_in(wire_d36_34),.data_out(wire_d36_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703636(.data_in(wire_d36_35),.data_out(wire_d36_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703637(.data_in(wire_d36_36),.data_out(wire_d36_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703638(.data_in(wire_d36_37),.data_out(wire_d36_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703639(.data_in(wire_d36_38),.data_out(wire_d36_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703640(.data_in(wire_d36_39),.data_out(wire_d36_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3703641(.data_in(wire_d36_40),.data_out(wire_d36_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703642(.data_in(wire_d36_41),.data_out(wire_d36_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3703643(.data_in(wire_d36_42),.data_out(wire_d36_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703644(.data_in(wire_d36_43),.data_out(wire_d36_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3703645(.data_in(wire_d36_44),.data_out(wire_d36_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3703646(.data_in(wire_d36_45),.data_out(wire_d36_46),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703647(.data_in(wire_d36_46),.data_out(wire_d36_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3703648(.data_in(wire_d36_47),.data_out(wire_d36_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703649(.data_in(wire_d36_48),.data_out(wire_d36_49),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3703650(.data_in(wire_d36_49),.data_out(wire_d36_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703651(.data_in(wire_d36_50),.data_out(wire_d36_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3703652(.data_in(wire_d36_51),.data_out(wire_d36_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703653(.data_in(wire_d36_52),.data_out(wire_d36_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703654(.data_in(wire_d36_53),.data_out(wire_d36_54),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3703655(.data_in(wire_d36_54),.data_out(wire_d36_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3703656(.data_in(wire_d36_55),.data_out(wire_d36_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703657(.data_in(wire_d36_56),.data_out(wire_d36_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703658(.data_in(wire_d36_57),.data_out(wire_d36_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3703659(.data_in(wire_d36_58),.data_out(wire_d36_59),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703660(.data_in(wire_d36_59),.data_out(wire_d36_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703661(.data_in(wire_d36_60),.data_out(wire_d36_61),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703662(.data_in(wire_d36_61),.data_out(wire_d36_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703663(.data_in(wire_d36_62),.data_out(wire_d36_63),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3703664(.data_in(wire_d36_63),.data_out(wire_d36_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3703665(.data_in(wire_d36_64),.data_out(wire_d36_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3703666(.data_in(wire_d36_65),.data_out(wire_d36_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3703667(.data_in(wire_d36_66),.data_out(wire_d36_67),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3703668(.data_in(wire_d36_67),.data_out(wire_d36_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3703669(.data_in(wire_d36_68),.data_out(wire_d36_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703670(.data_in(wire_d36_69),.data_out(wire_d36_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3703671(.data_in(wire_d36_70),.data_out(wire_d36_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703672(.data_in(wire_d36_71),.data_out(wire_d36_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3703673(.data_in(wire_d36_72),.data_out(wire_d36_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703674(.data_in(wire_d36_73),.data_out(wire_d36_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3703675(.data_in(wire_d36_74),.data_out(wire_d36_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703676(.data_in(wire_d36_75),.data_out(wire_d36_76),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3703677(.data_in(wire_d36_76),.data_out(wire_d36_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703678(.data_in(wire_d36_77),.data_out(wire_d36_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703679(.data_in(wire_d36_78),.data_out(wire_d36_79),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703680(.data_in(wire_d36_79),.data_out(wire_d36_80),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703681(.data_in(wire_d36_80),.data_out(wire_d36_81),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3703682(.data_in(wire_d36_81),.data_out(wire_d36_82),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703683(.data_in(wire_d36_82),.data_out(wire_d36_83),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703684(.data_in(wire_d36_83),.data_out(wire_d36_84),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703685(.data_in(wire_d36_84),.data_out(wire_d36_85),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703686(.data_in(wire_d36_85),.data_out(wire_d36_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703687(.data_in(wire_d36_86),.data_out(wire_d36_87),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703688(.data_in(wire_d36_87),.data_out(wire_d36_88),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703689(.data_in(wire_d36_88),.data_out(wire_d36_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3703690(.data_in(wire_d36_89),.data_out(wire_d36_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3703691(.data_in(wire_d36_90),.data_out(wire_d36_91),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703692(.data_in(wire_d36_91),.data_out(wire_d36_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3703693(.data_in(wire_d36_92),.data_out(wire_d36_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3703694(.data_in(wire_d36_93),.data_out(wire_d36_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3703695(.data_in(wire_d36_94),.data_out(wire_d36_95),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3703696(.data_in(wire_d36_95),.data_out(wire_d36_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3703697(.data_in(wire_d36_96),.data_out(wire_d36_97),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3703698(.data_in(wire_d36_97),.data_out(wire_d36_98),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703699(.data_in(wire_d36_98),.data_out(wire_d36_99),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance37036100(.data_in(wire_d36_99),.data_out(wire_d36_100),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance37036101(.data_in(wire_d36_100),.data_out(wire_d36_101),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance37036102(.data_in(wire_d36_101),.data_out(wire_d36_102),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance37036103(.data_in(wire_d36_102),.data_out(wire_d36_103),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance37036104(.data_in(wire_d36_103),.data_out(wire_d36_104),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance37036105(.data_in(wire_d36_104),.data_out(wire_d36_105),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance37036106(.data_in(wire_d36_105),.data_out(wire_d36_106),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance37036107(.data_in(wire_d36_106),.data_out(wire_d36_107),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance37036108(.data_in(wire_d36_107),.data_out(wire_d36_108),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance37036109(.data_in(wire_d36_108),.data_out(wire_d36_109),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance37036110(.data_in(wire_d36_109),.data_out(wire_d36_110),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance37036111(.data_in(wire_d36_110),.data_out(wire_d36_111),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance37036112(.data_in(wire_d36_111),.data_out(wire_d36_112),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance37036113(.data_in(wire_d36_112),.data_out(wire_d36_113),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance37036114(.data_in(wire_d36_113),.data_out(wire_d36_114),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance37036115(.data_in(wire_d36_114),.data_out(wire_d36_115),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance37036116(.data_in(wire_d36_115),.data_out(wire_d36_116),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance37036117(.data_in(wire_d36_116),.data_out(wire_d36_117),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance37036118(.data_in(wire_d36_117),.data_out(wire_d36_118),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance37036119(.data_in(wire_d36_118),.data_out(d_out36),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance380370(.data_in(d_in37),.data_out(wire_d37_0),.clk(clk),.rst(rst));            //channel 38
	large_adder #(.WIDTH(WIDTH)) large_adder_instance380371(.data_in(wire_d37_0),.data_out(wire_d37_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance380372(.data_in(wire_d37_1),.data_out(wire_d37_2),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance380373(.data_in(wire_d37_2),.data_out(wire_d37_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance380374(.data_in(wire_d37_3),.data_out(wire_d37_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance380375(.data_in(wire_d37_4),.data_out(wire_d37_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance380376(.data_in(wire_d37_5),.data_out(wire_d37_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance380377(.data_in(wire_d37_6),.data_out(wire_d37_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance380378(.data_in(wire_d37_7),.data_out(wire_d37_8),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance380379(.data_in(wire_d37_8),.data_out(wire_d37_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803710(.data_in(wire_d37_9),.data_out(wire_d37_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803711(.data_in(wire_d37_10),.data_out(wire_d37_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3803712(.data_in(wire_d37_11),.data_out(wire_d37_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803713(.data_in(wire_d37_12),.data_out(wire_d37_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803714(.data_in(wire_d37_13),.data_out(wire_d37_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803715(.data_in(wire_d37_14),.data_out(wire_d37_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803716(.data_in(wire_d37_15),.data_out(wire_d37_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803717(.data_in(wire_d37_16),.data_out(wire_d37_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803718(.data_in(wire_d37_17),.data_out(wire_d37_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803719(.data_in(wire_d37_18),.data_out(wire_d37_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803720(.data_in(wire_d37_19),.data_out(wire_d37_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803721(.data_in(wire_d37_20),.data_out(wire_d37_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803722(.data_in(wire_d37_21),.data_out(wire_d37_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803723(.data_in(wire_d37_22),.data_out(wire_d37_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803724(.data_in(wire_d37_23),.data_out(wire_d37_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803725(.data_in(wire_d37_24),.data_out(wire_d37_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803726(.data_in(wire_d37_25),.data_out(wire_d37_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803727(.data_in(wire_d37_26),.data_out(wire_d37_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803728(.data_in(wire_d37_27),.data_out(wire_d37_28),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3803729(.data_in(wire_d37_28),.data_out(wire_d37_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3803730(.data_in(wire_d37_29),.data_out(wire_d37_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803731(.data_in(wire_d37_30),.data_out(wire_d37_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803732(.data_in(wire_d37_31),.data_out(wire_d37_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803733(.data_in(wire_d37_32),.data_out(wire_d37_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803734(.data_in(wire_d37_33),.data_out(wire_d37_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3803735(.data_in(wire_d37_34),.data_out(wire_d37_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3803736(.data_in(wire_d37_35),.data_out(wire_d37_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803737(.data_in(wire_d37_36),.data_out(wire_d37_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803738(.data_in(wire_d37_37),.data_out(wire_d37_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803739(.data_in(wire_d37_38),.data_out(wire_d37_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803740(.data_in(wire_d37_39),.data_out(wire_d37_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803741(.data_in(wire_d37_40),.data_out(wire_d37_41),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3803742(.data_in(wire_d37_41),.data_out(wire_d37_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3803743(.data_in(wire_d37_42),.data_out(wire_d37_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3803744(.data_in(wire_d37_43),.data_out(wire_d37_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803745(.data_in(wire_d37_44),.data_out(wire_d37_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803746(.data_in(wire_d37_45),.data_out(wire_d37_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3803747(.data_in(wire_d37_46),.data_out(wire_d37_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803748(.data_in(wire_d37_47),.data_out(wire_d37_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803749(.data_in(wire_d37_48),.data_out(wire_d37_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803750(.data_in(wire_d37_49),.data_out(wire_d37_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3803751(.data_in(wire_d37_50),.data_out(wire_d37_51),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3803752(.data_in(wire_d37_51),.data_out(wire_d37_52),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3803753(.data_in(wire_d37_52),.data_out(wire_d37_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803754(.data_in(wire_d37_53),.data_out(wire_d37_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3803755(.data_in(wire_d37_54),.data_out(wire_d37_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803756(.data_in(wire_d37_55),.data_out(wire_d37_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3803757(.data_in(wire_d37_56),.data_out(wire_d37_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803758(.data_in(wire_d37_57),.data_out(wire_d37_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3803759(.data_in(wire_d37_58),.data_out(wire_d37_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803760(.data_in(wire_d37_59),.data_out(wire_d37_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3803761(.data_in(wire_d37_60),.data_out(wire_d37_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803762(.data_in(wire_d37_61),.data_out(wire_d37_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803763(.data_in(wire_d37_62),.data_out(wire_d37_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803764(.data_in(wire_d37_63),.data_out(wire_d37_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803765(.data_in(wire_d37_64),.data_out(wire_d37_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803766(.data_in(wire_d37_65),.data_out(wire_d37_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803767(.data_in(wire_d37_66),.data_out(wire_d37_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803768(.data_in(wire_d37_67),.data_out(wire_d37_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803769(.data_in(wire_d37_68),.data_out(wire_d37_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803770(.data_in(wire_d37_69),.data_out(wire_d37_70),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803771(.data_in(wire_d37_70),.data_out(wire_d37_71),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3803772(.data_in(wire_d37_71),.data_out(wire_d37_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803773(.data_in(wire_d37_72),.data_out(wire_d37_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803774(.data_in(wire_d37_73),.data_out(wire_d37_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803775(.data_in(wire_d37_74),.data_out(wire_d37_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3803776(.data_in(wire_d37_75),.data_out(wire_d37_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3803777(.data_in(wire_d37_76),.data_out(wire_d37_77),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803778(.data_in(wire_d37_77),.data_out(wire_d37_78),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3803779(.data_in(wire_d37_78),.data_out(wire_d37_79),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803780(.data_in(wire_d37_79),.data_out(wire_d37_80),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803781(.data_in(wire_d37_80),.data_out(wire_d37_81),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803782(.data_in(wire_d37_81),.data_out(wire_d37_82),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803783(.data_in(wire_d37_82),.data_out(wire_d37_83),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3803784(.data_in(wire_d37_83),.data_out(wire_d37_84),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803785(.data_in(wire_d37_84),.data_out(wire_d37_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803786(.data_in(wire_d37_85),.data_out(wire_d37_86),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803787(.data_in(wire_d37_86),.data_out(wire_d37_87),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3803788(.data_in(wire_d37_87),.data_out(wire_d37_88),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803789(.data_in(wire_d37_88),.data_out(wire_d37_89),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803790(.data_in(wire_d37_89),.data_out(wire_d37_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803791(.data_in(wire_d37_90),.data_out(wire_d37_91),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803792(.data_in(wire_d37_91),.data_out(wire_d37_92),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3803793(.data_in(wire_d37_92),.data_out(wire_d37_93),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803794(.data_in(wire_d37_93),.data_out(wire_d37_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3803795(.data_in(wire_d37_94),.data_out(wire_d37_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803796(.data_in(wire_d37_95),.data_out(wire_d37_96),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803797(.data_in(wire_d37_96),.data_out(wire_d37_97),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803798(.data_in(wire_d37_97),.data_out(wire_d37_98),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803799(.data_in(wire_d37_98),.data_out(wire_d37_99),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance38037100(.data_in(wire_d37_99),.data_out(wire_d37_100),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance38037101(.data_in(wire_d37_100),.data_out(wire_d37_101),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance38037102(.data_in(wire_d37_101),.data_out(wire_d37_102),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance38037103(.data_in(wire_d37_102),.data_out(wire_d37_103),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance38037104(.data_in(wire_d37_103),.data_out(wire_d37_104),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance38037105(.data_in(wire_d37_104),.data_out(wire_d37_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance38037106(.data_in(wire_d37_105),.data_out(wire_d37_106),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance38037107(.data_in(wire_d37_106),.data_out(wire_d37_107),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance38037108(.data_in(wire_d37_107),.data_out(wire_d37_108),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance38037109(.data_in(wire_d37_108),.data_out(wire_d37_109),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance38037110(.data_in(wire_d37_109),.data_out(wire_d37_110),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance38037111(.data_in(wire_d37_110),.data_out(wire_d37_111),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance38037112(.data_in(wire_d37_111),.data_out(wire_d37_112),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance38037113(.data_in(wire_d37_112),.data_out(wire_d37_113),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance38037114(.data_in(wire_d37_113),.data_out(wire_d37_114),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance38037115(.data_in(wire_d37_114),.data_out(wire_d37_115),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance38037116(.data_in(wire_d37_115),.data_out(wire_d37_116),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance38037117(.data_in(wire_d37_116),.data_out(wire_d37_117),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance38037118(.data_in(wire_d37_117),.data_out(wire_d37_118),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance38037119(.data_in(wire_d37_118),.data_out(d_out37),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance390380(.data_in(d_in38),.data_out(wire_d38_0),.clk(clk),.rst(rst));            //channel 39
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance390381(.data_in(wire_d38_0),.data_out(wire_d38_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance390382(.data_in(wire_d38_1),.data_out(wire_d38_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance390383(.data_in(wire_d38_2),.data_out(wire_d38_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance390384(.data_in(wire_d38_3),.data_out(wire_d38_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance390385(.data_in(wire_d38_4),.data_out(wire_d38_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance390386(.data_in(wire_d38_5),.data_out(wire_d38_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance390387(.data_in(wire_d38_6),.data_out(wire_d38_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance390388(.data_in(wire_d38_7),.data_out(wire_d38_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance390389(.data_in(wire_d38_8),.data_out(wire_d38_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3903810(.data_in(wire_d38_9),.data_out(wire_d38_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3903811(.data_in(wire_d38_10),.data_out(wire_d38_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903812(.data_in(wire_d38_11),.data_out(wire_d38_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903813(.data_in(wire_d38_12),.data_out(wire_d38_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903814(.data_in(wire_d38_13),.data_out(wire_d38_14),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3903815(.data_in(wire_d38_14),.data_out(wire_d38_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3903816(.data_in(wire_d38_15),.data_out(wire_d38_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903817(.data_in(wire_d38_16),.data_out(wire_d38_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3903818(.data_in(wire_d38_17),.data_out(wire_d38_18),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3903819(.data_in(wire_d38_18),.data_out(wire_d38_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903820(.data_in(wire_d38_19),.data_out(wire_d38_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3903821(.data_in(wire_d38_20),.data_out(wire_d38_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903822(.data_in(wire_d38_21),.data_out(wire_d38_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903823(.data_in(wire_d38_22),.data_out(wire_d38_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903824(.data_in(wire_d38_23),.data_out(wire_d38_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3903825(.data_in(wire_d38_24),.data_out(wire_d38_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903826(.data_in(wire_d38_25),.data_out(wire_d38_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3903827(.data_in(wire_d38_26),.data_out(wire_d38_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903828(.data_in(wire_d38_27),.data_out(wire_d38_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3903829(.data_in(wire_d38_28),.data_out(wire_d38_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903830(.data_in(wire_d38_29),.data_out(wire_d38_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3903831(.data_in(wire_d38_30),.data_out(wire_d38_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3903832(.data_in(wire_d38_31),.data_out(wire_d38_32),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3903833(.data_in(wire_d38_32),.data_out(wire_d38_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903834(.data_in(wire_d38_33),.data_out(wire_d38_34),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3903835(.data_in(wire_d38_34),.data_out(wire_d38_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903836(.data_in(wire_d38_35),.data_out(wire_d38_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903837(.data_in(wire_d38_36),.data_out(wire_d38_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903838(.data_in(wire_d38_37),.data_out(wire_d38_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3903839(.data_in(wire_d38_38),.data_out(wire_d38_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903840(.data_in(wire_d38_39),.data_out(wire_d38_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3903841(.data_in(wire_d38_40),.data_out(wire_d38_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903842(.data_in(wire_d38_41),.data_out(wire_d38_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903843(.data_in(wire_d38_42),.data_out(wire_d38_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903844(.data_in(wire_d38_43),.data_out(wire_d38_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3903845(.data_in(wire_d38_44),.data_out(wire_d38_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903846(.data_in(wire_d38_45),.data_out(wire_d38_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3903847(.data_in(wire_d38_46),.data_out(wire_d38_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903848(.data_in(wire_d38_47),.data_out(wire_d38_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903849(.data_in(wire_d38_48),.data_out(wire_d38_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3903850(.data_in(wire_d38_49),.data_out(wire_d38_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903851(.data_in(wire_d38_50),.data_out(wire_d38_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3903852(.data_in(wire_d38_51),.data_out(wire_d38_52),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903853(.data_in(wire_d38_52),.data_out(wire_d38_53),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3903854(.data_in(wire_d38_53),.data_out(wire_d38_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3903855(.data_in(wire_d38_54),.data_out(wire_d38_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903856(.data_in(wire_d38_55),.data_out(wire_d38_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3903857(.data_in(wire_d38_56),.data_out(wire_d38_57),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903858(.data_in(wire_d38_57),.data_out(wire_d38_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903859(.data_in(wire_d38_58),.data_out(wire_d38_59),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3903860(.data_in(wire_d38_59),.data_out(wire_d38_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3903861(.data_in(wire_d38_60),.data_out(wire_d38_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3903862(.data_in(wire_d38_61),.data_out(wire_d38_62),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3903863(.data_in(wire_d38_62),.data_out(wire_d38_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3903864(.data_in(wire_d38_63),.data_out(wire_d38_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903865(.data_in(wire_d38_64),.data_out(wire_d38_65),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903866(.data_in(wire_d38_65),.data_out(wire_d38_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3903867(.data_in(wire_d38_66),.data_out(wire_d38_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903868(.data_in(wire_d38_67),.data_out(wire_d38_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3903869(.data_in(wire_d38_68),.data_out(wire_d38_69),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903870(.data_in(wire_d38_69),.data_out(wire_d38_70),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3903871(.data_in(wire_d38_70),.data_out(wire_d38_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3903872(.data_in(wire_d38_71),.data_out(wire_d38_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903873(.data_in(wire_d38_72),.data_out(wire_d38_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903874(.data_in(wire_d38_73),.data_out(wire_d38_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3903875(.data_in(wire_d38_74),.data_out(wire_d38_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3903876(.data_in(wire_d38_75),.data_out(wire_d38_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903877(.data_in(wire_d38_76),.data_out(wire_d38_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903878(.data_in(wire_d38_77),.data_out(wire_d38_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903879(.data_in(wire_d38_78),.data_out(wire_d38_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3903880(.data_in(wire_d38_79),.data_out(wire_d38_80),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3903881(.data_in(wire_d38_80),.data_out(wire_d38_81),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903882(.data_in(wire_d38_81),.data_out(wire_d38_82),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3903883(.data_in(wire_d38_82),.data_out(wire_d38_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3903884(.data_in(wire_d38_83),.data_out(wire_d38_84),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903885(.data_in(wire_d38_84),.data_out(wire_d38_85),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903886(.data_in(wire_d38_85),.data_out(wire_d38_86),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903887(.data_in(wire_d38_86),.data_out(wire_d38_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3903888(.data_in(wire_d38_87),.data_out(wire_d38_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3903889(.data_in(wire_d38_88),.data_out(wire_d38_89),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3903890(.data_in(wire_d38_89),.data_out(wire_d38_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903891(.data_in(wire_d38_90),.data_out(wire_d38_91),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903892(.data_in(wire_d38_91),.data_out(wire_d38_92),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903893(.data_in(wire_d38_92),.data_out(wire_d38_93),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3903894(.data_in(wire_d38_93),.data_out(wire_d38_94),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903895(.data_in(wire_d38_94),.data_out(wire_d38_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903896(.data_in(wire_d38_95),.data_out(wire_d38_96),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903897(.data_in(wire_d38_96),.data_out(wire_d38_97),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903898(.data_in(wire_d38_97),.data_out(wire_d38_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903899(.data_in(wire_d38_98),.data_out(wire_d38_99),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance39038100(.data_in(wire_d38_99),.data_out(wire_d38_100),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance39038101(.data_in(wire_d38_100),.data_out(wire_d38_101),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance39038102(.data_in(wire_d38_101),.data_out(wire_d38_102),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance39038103(.data_in(wire_d38_102),.data_out(wire_d38_103),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance39038104(.data_in(wire_d38_103),.data_out(wire_d38_104),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance39038105(.data_in(wire_d38_104),.data_out(wire_d38_105),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance39038106(.data_in(wire_d38_105),.data_out(wire_d38_106),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance39038107(.data_in(wire_d38_106),.data_out(wire_d38_107),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance39038108(.data_in(wire_d38_107),.data_out(wire_d38_108),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance39038109(.data_in(wire_d38_108),.data_out(wire_d38_109),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance39038110(.data_in(wire_d38_109),.data_out(wire_d38_110),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance39038111(.data_in(wire_d38_110),.data_out(wire_d38_111),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance39038112(.data_in(wire_d38_111),.data_out(wire_d38_112),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance39038113(.data_in(wire_d38_112),.data_out(wire_d38_113),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance39038114(.data_in(wire_d38_113),.data_out(wire_d38_114),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance39038115(.data_in(wire_d38_114),.data_out(wire_d38_115),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance39038116(.data_in(wire_d38_115),.data_out(wire_d38_116),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance39038117(.data_in(wire_d38_116),.data_out(wire_d38_117),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance39038118(.data_in(wire_d38_117),.data_out(wire_d38_118),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance39038119(.data_in(wire_d38_118),.data_out(d_out38),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance400390(.data_in(d_in39),.data_out(wire_d39_0),.clk(clk),.rst(rst));            //channel 40
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance400391(.data_in(wire_d39_0),.data_out(wire_d39_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance400392(.data_in(wire_d39_1),.data_out(wire_d39_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance400393(.data_in(wire_d39_2),.data_out(wire_d39_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance400394(.data_in(wire_d39_3),.data_out(wire_d39_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance400395(.data_in(wire_d39_4),.data_out(wire_d39_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance400396(.data_in(wire_d39_5),.data_out(wire_d39_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance400397(.data_in(wire_d39_6),.data_out(wire_d39_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance400398(.data_in(wire_d39_7),.data_out(wire_d39_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance400399(.data_in(wire_d39_8),.data_out(wire_d39_9),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003910(.data_in(wire_d39_9),.data_out(wire_d39_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4003911(.data_in(wire_d39_10),.data_out(wire_d39_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003912(.data_in(wire_d39_11),.data_out(wire_d39_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4003913(.data_in(wire_d39_12),.data_out(wire_d39_13),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4003914(.data_in(wire_d39_13),.data_out(wire_d39_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4003915(.data_in(wire_d39_14),.data_out(wire_d39_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003916(.data_in(wire_d39_15),.data_out(wire_d39_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4003917(.data_in(wire_d39_16),.data_out(wire_d39_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003918(.data_in(wire_d39_17),.data_out(wire_d39_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4003919(.data_in(wire_d39_18),.data_out(wire_d39_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003920(.data_in(wire_d39_19),.data_out(wire_d39_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003921(.data_in(wire_d39_20),.data_out(wire_d39_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003922(.data_in(wire_d39_21),.data_out(wire_d39_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003923(.data_in(wire_d39_22),.data_out(wire_d39_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003924(.data_in(wire_d39_23),.data_out(wire_d39_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4003925(.data_in(wire_d39_24),.data_out(wire_d39_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4003926(.data_in(wire_d39_25),.data_out(wire_d39_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003927(.data_in(wire_d39_26),.data_out(wire_d39_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4003928(.data_in(wire_d39_27),.data_out(wire_d39_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003929(.data_in(wire_d39_28),.data_out(wire_d39_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4003930(.data_in(wire_d39_29),.data_out(wire_d39_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003931(.data_in(wire_d39_30),.data_out(wire_d39_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003932(.data_in(wire_d39_31),.data_out(wire_d39_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003933(.data_in(wire_d39_32),.data_out(wire_d39_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4003934(.data_in(wire_d39_33),.data_out(wire_d39_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003935(.data_in(wire_d39_34),.data_out(wire_d39_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4003936(.data_in(wire_d39_35),.data_out(wire_d39_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4003937(.data_in(wire_d39_36),.data_out(wire_d39_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003938(.data_in(wire_d39_37),.data_out(wire_d39_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4003939(.data_in(wire_d39_38),.data_out(wire_d39_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003940(.data_in(wire_d39_39),.data_out(wire_d39_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4003941(.data_in(wire_d39_40),.data_out(wire_d39_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003942(.data_in(wire_d39_41),.data_out(wire_d39_42),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4003943(.data_in(wire_d39_42),.data_out(wire_d39_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003944(.data_in(wire_d39_43),.data_out(wire_d39_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4003945(.data_in(wire_d39_44),.data_out(wire_d39_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4003946(.data_in(wire_d39_45),.data_out(wire_d39_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003947(.data_in(wire_d39_46),.data_out(wire_d39_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003948(.data_in(wire_d39_47),.data_out(wire_d39_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4003949(.data_in(wire_d39_48),.data_out(wire_d39_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003950(.data_in(wire_d39_49),.data_out(wire_d39_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003951(.data_in(wire_d39_50),.data_out(wire_d39_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003952(.data_in(wire_d39_51),.data_out(wire_d39_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003953(.data_in(wire_d39_52),.data_out(wire_d39_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003954(.data_in(wire_d39_53),.data_out(wire_d39_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4003955(.data_in(wire_d39_54),.data_out(wire_d39_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003956(.data_in(wire_d39_55),.data_out(wire_d39_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003957(.data_in(wire_d39_56),.data_out(wire_d39_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4003958(.data_in(wire_d39_57),.data_out(wire_d39_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003959(.data_in(wire_d39_58),.data_out(wire_d39_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4003960(.data_in(wire_d39_59),.data_out(wire_d39_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003961(.data_in(wire_d39_60),.data_out(wire_d39_61),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003962(.data_in(wire_d39_61),.data_out(wire_d39_62),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4003963(.data_in(wire_d39_62),.data_out(wire_d39_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003964(.data_in(wire_d39_63),.data_out(wire_d39_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4003965(.data_in(wire_d39_64),.data_out(wire_d39_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003966(.data_in(wire_d39_65),.data_out(wire_d39_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003967(.data_in(wire_d39_66),.data_out(wire_d39_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4003968(.data_in(wire_d39_67),.data_out(wire_d39_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003969(.data_in(wire_d39_68),.data_out(wire_d39_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003970(.data_in(wire_d39_69),.data_out(wire_d39_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4003971(.data_in(wire_d39_70),.data_out(wire_d39_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003972(.data_in(wire_d39_71),.data_out(wire_d39_72),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4003973(.data_in(wire_d39_72),.data_out(wire_d39_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003974(.data_in(wire_d39_73),.data_out(wire_d39_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4003975(.data_in(wire_d39_74),.data_out(wire_d39_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4003976(.data_in(wire_d39_75),.data_out(wire_d39_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003977(.data_in(wire_d39_76),.data_out(wire_d39_77),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4003978(.data_in(wire_d39_77),.data_out(wire_d39_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4003979(.data_in(wire_d39_78),.data_out(wire_d39_79),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003980(.data_in(wire_d39_79),.data_out(wire_d39_80),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003981(.data_in(wire_d39_80),.data_out(wire_d39_81),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003982(.data_in(wire_d39_81),.data_out(wire_d39_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003983(.data_in(wire_d39_82),.data_out(wire_d39_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4003984(.data_in(wire_d39_83),.data_out(wire_d39_84),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4003985(.data_in(wire_d39_84),.data_out(wire_d39_85),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003986(.data_in(wire_d39_85),.data_out(wire_d39_86),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003987(.data_in(wire_d39_86),.data_out(wire_d39_87),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003988(.data_in(wire_d39_87),.data_out(wire_d39_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003989(.data_in(wire_d39_88),.data_out(wire_d39_89),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003990(.data_in(wire_d39_89),.data_out(wire_d39_90),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003991(.data_in(wire_d39_90),.data_out(wire_d39_91),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4003992(.data_in(wire_d39_91),.data_out(wire_d39_92),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003993(.data_in(wire_d39_92),.data_out(wire_d39_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003994(.data_in(wire_d39_93),.data_out(wire_d39_94),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003995(.data_in(wire_d39_94),.data_out(wire_d39_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003996(.data_in(wire_d39_95),.data_out(wire_d39_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4003997(.data_in(wire_d39_96),.data_out(wire_d39_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003998(.data_in(wire_d39_97),.data_out(wire_d39_98),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4003999(.data_in(wire_d39_98),.data_out(wire_d39_99),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance40039100(.data_in(wire_d39_99),.data_out(wire_d39_100),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance40039101(.data_in(wire_d39_100),.data_out(wire_d39_101),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance40039102(.data_in(wire_d39_101),.data_out(wire_d39_102),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance40039103(.data_in(wire_d39_102),.data_out(wire_d39_103),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance40039104(.data_in(wire_d39_103),.data_out(wire_d39_104),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance40039105(.data_in(wire_d39_104),.data_out(wire_d39_105),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance40039106(.data_in(wire_d39_105),.data_out(wire_d39_106),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance40039107(.data_in(wire_d39_106),.data_out(wire_d39_107),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance40039108(.data_in(wire_d39_107),.data_out(wire_d39_108),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance40039109(.data_in(wire_d39_108),.data_out(wire_d39_109),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance40039110(.data_in(wire_d39_109),.data_out(wire_d39_110),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance40039111(.data_in(wire_d39_110),.data_out(wire_d39_111),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance40039112(.data_in(wire_d39_111),.data_out(wire_d39_112),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance40039113(.data_in(wire_d39_112),.data_out(wire_d39_113),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance40039114(.data_in(wire_d39_113),.data_out(wire_d39_114),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance40039115(.data_in(wire_d39_114),.data_out(wire_d39_115),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance40039116(.data_in(wire_d39_115),.data_out(wire_d39_116),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance40039117(.data_in(wire_d39_116),.data_out(wire_d39_117),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance40039118(.data_in(wire_d39_117),.data_out(wire_d39_118),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance40039119(.data_in(wire_d39_118),.data_out(d_out39),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance410400(.data_in(d_in40),.data_out(wire_d40_0),.clk(clk),.rst(rst));            //channel 41
	large_adder #(.WIDTH(WIDTH)) large_adder_instance410401(.data_in(wire_d40_0),.data_out(wire_d40_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance410402(.data_in(wire_d40_1),.data_out(wire_d40_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance410403(.data_in(wire_d40_2),.data_out(wire_d40_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance410404(.data_in(wire_d40_3),.data_out(wire_d40_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance410405(.data_in(wire_d40_4),.data_out(wire_d40_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance410406(.data_in(wire_d40_5),.data_out(wire_d40_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance410407(.data_in(wire_d40_6),.data_out(wire_d40_7),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance410408(.data_in(wire_d40_7),.data_out(wire_d40_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance410409(.data_in(wire_d40_8),.data_out(wire_d40_9),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4104010(.data_in(wire_d40_9),.data_out(wire_d40_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104011(.data_in(wire_d40_10),.data_out(wire_d40_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4104012(.data_in(wire_d40_11),.data_out(wire_d40_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4104013(.data_in(wire_d40_12),.data_out(wire_d40_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4104014(.data_in(wire_d40_13),.data_out(wire_d40_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104015(.data_in(wire_d40_14),.data_out(wire_d40_15),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4104016(.data_in(wire_d40_15),.data_out(wire_d40_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104017(.data_in(wire_d40_16),.data_out(wire_d40_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104018(.data_in(wire_d40_17),.data_out(wire_d40_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4104019(.data_in(wire_d40_18),.data_out(wire_d40_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4104020(.data_in(wire_d40_19),.data_out(wire_d40_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104021(.data_in(wire_d40_20),.data_out(wire_d40_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104022(.data_in(wire_d40_21),.data_out(wire_d40_22),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4104023(.data_in(wire_d40_22),.data_out(wire_d40_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104024(.data_in(wire_d40_23),.data_out(wire_d40_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4104025(.data_in(wire_d40_24),.data_out(wire_d40_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4104026(.data_in(wire_d40_25),.data_out(wire_d40_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4104027(.data_in(wire_d40_26),.data_out(wire_d40_27),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4104028(.data_in(wire_d40_27),.data_out(wire_d40_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104029(.data_in(wire_d40_28),.data_out(wire_d40_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104030(.data_in(wire_d40_29),.data_out(wire_d40_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104031(.data_in(wire_d40_30),.data_out(wire_d40_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4104032(.data_in(wire_d40_31),.data_out(wire_d40_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104033(.data_in(wire_d40_32),.data_out(wire_d40_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104034(.data_in(wire_d40_33),.data_out(wire_d40_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104035(.data_in(wire_d40_34),.data_out(wire_d40_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104036(.data_in(wire_d40_35),.data_out(wire_d40_36),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104037(.data_in(wire_d40_36),.data_out(wire_d40_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4104038(.data_in(wire_d40_37),.data_out(wire_d40_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4104039(.data_in(wire_d40_38),.data_out(wire_d40_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104040(.data_in(wire_d40_39),.data_out(wire_d40_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4104041(.data_in(wire_d40_40),.data_out(wire_d40_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4104042(.data_in(wire_d40_41),.data_out(wire_d40_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104043(.data_in(wire_d40_42),.data_out(wire_d40_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104044(.data_in(wire_d40_43),.data_out(wire_d40_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104045(.data_in(wire_d40_44),.data_out(wire_d40_45),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104046(.data_in(wire_d40_45),.data_out(wire_d40_46),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104047(.data_in(wire_d40_46),.data_out(wire_d40_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104048(.data_in(wire_d40_47),.data_out(wire_d40_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4104049(.data_in(wire_d40_48),.data_out(wire_d40_49),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104050(.data_in(wire_d40_49),.data_out(wire_d40_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104051(.data_in(wire_d40_50),.data_out(wire_d40_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4104052(.data_in(wire_d40_51),.data_out(wire_d40_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104053(.data_in(wire_d40_52),.data_out(wire_d40_53),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4104054(.data_in(wire_d40_53),.data_out(wire_d40_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4104055(.data_in(wire_d40_54),.data_out(wire_d40_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104056(.data_in(wire_d40_55),.data_out(wire_d40_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104057(.data_in(wire_d40_56),.data_out(wire_d40_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104058(.data_in(wire_d40_57),.data_out(wire_d40_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4104059(.data_in(wire_d40_58),.data_out(wire_d40_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4104060(.data_in(wire_d40_59),.data_out(wire_d40_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104061(.data_in(wire_d40_60),.data_out(wire_d40_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104062(.data_in(wire_d40_61),.data_out(wire_d40_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4104063(.data_in(wire_d40_62),.data_out(wire_d40_63),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104064(.data_in(wire_d40_63),.data_out(wire_d40_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4104065(.data_in(wire_d40_64),.data_out(wire_d40_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4104066(.data_in(wire_d40_65),.data_out(wire_d40_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104067(.data_in(wire_d40_66),.data_out(wire_d40_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4104068(.data_in(wire_d40_67),.data_out(wire_d40_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4104069(.data_in(wire_d40_68),.data_out(wire_d40_69),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104070(.data_in(wire_d40_69),.data_out(wire_d40_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104071(.data_in(wire_d40_70),.data_out(wire_d40_71),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4104072(.data_in(wire_d40_71),.data_out(wire_d40_72),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104073(.data_in(wire_d40_72),.data_out(wire_d40_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104074(.data_in(wire_d40_73),.data_out(wire_d40_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104075(.data_in(wire_d40_74),.data_out(wire_d40_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4104076(.data_in(wire_d40_75),.data_out(wire_d40_76),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104077(.data_in(wire_d40_76),.data_out(wire_d40_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104078(.data_in(wire_d40_77),.data_out(wire_d40_78),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4104079(.data_in(wire_d40_78),.data_out(wire_d40_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104080(.data_in(wire_d40_79),.data_out(wire_d40_80),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4104081(.data_in(wire_d40_80),.data_out(wire_d40_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4104082(.data_in(wire_d40_81),.data_out(wire_d40_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4104083(.data_in(wire_d40_82),.data_out(wire_d40_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104084(.data_in(wire_d40_83),.data_out(wire_d40_84),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4104085(.data_in(wire_d40_84),.data_out(wire_d40_85),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104086(.data_in(wire_d40_85),.data_out(wire_d40_86),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4104087(.data_in(wire_d40_86),.data_out(wire_d40_87),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104088(.data_in(wire_d40_87),.data_out(wire_d40_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4104089(.data_in(wire_d40_88),.data_out(wire_d40_89),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104090(.data_in(wire_d40_89),.data_out(wire_d40_90),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104091(.data_in(wire_d40_90),.data_out(wire_d40_91),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104092(.data_in(wire_d40_91),.data_out(wire_d40_92),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4104093(.data_in(wire_d40_92),.data_out(wire_d40_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104094(.data_in(wire_d40_93),.data_out(wire_d40_94),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104095(.data_in(wire_d40_94),.data_out(wire_d40_95),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104096(.data_in(wire_d40_95),.data_out(wire_d40_96),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104097(.data_in(wire_d40_96),.data_out(wire_d40_97),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104098(.data_in(wire_d40_97),.data_out(wire_d40_98),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104099(.data_in(wire_d40_98),.data_out(wire_d40_99),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance41040100(.data_in(wire_d40_99),.data_out(wire_d40_100),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance41040101(.data_in(wire_d40_100),.data_out(wire_d40_101),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance41040102(.data_in(wire_d40_101),.data_out(wire_d40_102),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance41040103(.data_in(wire_d40_102),.data_out(wire_d40_103),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance41040104(.data_in(wire_d40_103),.data_out(wire_d40_104),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance41040105(.data_in(wire_d40_104),.data_out(wire_d40_105),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance41040106(.data_in(wire_d40_105),.data_out(wire_d40_106),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance41040107(.data_in(wire_d40_106),.data_out(wire_d40_107),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance41040108(.data_in(wire_d40_107),.data_out(wire_d40_108),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance41040109(.data_in(wire_d40_108),.data_out(wire_d40_109),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance41040110(.data_in(wire_d40_109),.data_out(wire_d40_110),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance41040111(.data_in(wire_d40_110),.data_out(wire_d40_111),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance41040112(.data_in(wire_d40_111),.data_out(wire_d40_112),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance41040113(.data_in(wire_d40_112),.data_out(wire_d40_113),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance41040114(.data_in(wire_d40_113),.data_out(wire_d40_114),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance41040115(.data_in(wire_d40_114),.data_out(wire_d40_115),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance41040116(.data_in(wire_d40_115),.data_out(wire_d40_116),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance41040117(.data_in(wire_d40_116),.data_out(wire_d40_117),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance41040118(.data_in(wire_d40_117),.data_out(wire_d40_118),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance41040119(.data_in(wire_d40_118),.data_out(d_out40),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance420410(.data_in(d_in41),.data_out(wire_d41_0),.clk(clk),.rst(rst));            //channel 42
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance420411(.data_in(wire_d41_0),.data_out(wire_d41_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance420412(.data_in(wire_d41_1),.data_out(wire_d41_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance420413(.data_in(wire_d41_2),.data_out(wire_d41_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance420414(.data_in(wire_d41_3),.data_out(wire_d41_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance420415(.data_in(wire_d41_4),.data_out(wire_d41_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance420416(.data_in(wire_d41_5),.data_out(wire_d41_6),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance420417(.data_in(wire_d41_6),.data_out(wire_d41_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance420418(.data_in(wire_d41_7),.data_out(wire_d41_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance420419(.data_in(wire_d41_8),.data_out(wire_d41_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204110(.data_in(wire_d41_9),.data_out(wire_d41_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4204111(.data_in(wire_d41_10),.data_out(wire_d41_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204112(.data_in(wire_d41_11),.data_out(wire_d41_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204113(.data_in(wire_d41_12),.data_out(wire_d41_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4204114(.data_in(wire_d41_13),.data_out(wire_d41_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204115(.data_in(wire_d41_14),.data_out(wire_d41_15),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4204116(.data_in(wire_d41_15),.data_out(wire_d41_16),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4204117(.data_in(wire_d41_16),.data_out(wire_d41_17),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4204118(.data_in(wire_d41_17),.data_out(wire_d41_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4204119(.data_in(wire_d41_18),.data_out(wire_d41_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204120(.data_in(wire_d41_19),.data_out(wire_d41_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4204121(.data_in(wire_d41_20),.data_out(wire_d41_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204122(.data_in(wire_d41_21),.data_out(wire_d41_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204123(.data_in(wire_d41_22),.data_out(wire_d41_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204124(.data_in(wire_d41_23),.data_out(wire_d41_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204125(.data_in(wire_d41_24),.data_out(wire_d41_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204126(.data_in(wire_d41_25),.data_out(wire_d41_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204127(.data_in(wire_d41_26),.data_out(wire_d41_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4204128(.data_in(wire_d41_27),.data_out(wire_d41_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204129(.data_in(wire_d41_28),.data_out(wire_d41_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4204130(.data_in(wire_d41_29),.data_out(wire_d41_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4204131(.data_in(wire_d41_30),.data_out(wire_d41_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204132(.data_in(wire_d41_31),.data_out(wire_d41_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4204133(.data_in(wire_d41_32),.data_out(wire_d41_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4204134(.data_in(wire_d41_33),.data_out(wire_d41_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204135(.data_in(wire_d41_34),.data_out(wire_d41_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4204136(.data_in(wire_d41_35),.data_out(wire_d41_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204137(.data_in(wire_d41_36),.data_out(wire_d41_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204138(.data_in(wire_d41_37),.data_out(wire_d41_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204139(.data_in(wire_d41_38),.data_out(wire_d41_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4204140(.data_in(wire_d41_39),.data_out(wire_d41_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204141(.data_in(wire_d41_40),.data_out(wire_d41_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4204142(.data_in(wire_d41_41),.data_out(wire_d41_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4204143(.data_in(wire_d41_42),.data_out(wire_d41_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204144(.data_in(wire_d41_43),.data_out(wire_d41_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204145(.data_in(wire_d41_44),.data_out(wire_d41_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4204146(.data_in(wire_d41_45),.data_out(wire_d41_46),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4204147(.data_in(wire_d41_46),.data_out(wire_d41_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204148(.data_in(wire_d41_47),.data_out(wire_d41_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204149(.data_in(wire_d41_48),.data_out(wire_d41_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204150(.data_in(wire_d41_49),.data_out(wire_d41_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204151(.data_in(wire_d41_50),.data_out(wire_d41_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204152(.data_in(wire_d41_51),.data_out(wire_d41_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204153(.data_in(wire_d41_52),.data_out(wire_d41_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4204154(.data_in(wire_d41_53),.data_out(wire_d41_54),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204155(.data_in(wire_d41_54),.data_out(wire_d41_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204156(.data_in(wire_d41_55),.data_out(wire_d41_56),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4204157(.data_in(wire_d41_56),.data_out(wire_d41_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204158(.data_in(wire_d41_57),.data_out(wire_d41_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4204159(.data_in(wire_d41_58),.data_out(wire_d41_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4204160(.data_in(wire_d41_59),.data_out(wire_d41_60),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204161(.data_in(wire_d41_60),.data_out(wire_d41_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4204162(.data_in(wire_d41_61),.data_out(wire_d41_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204163(.data_in(wire_d41_62),.data_out(wire_d41_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4204164(.data_in(wire_d41_63),.data_out(wire_d41_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204165(.data_in(wire_d41_64),.data_out(wire_d41_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204166(.data_in(wire_d41_65),.data_out(wire_d41_66),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204167(.data_in(wire_d41_66),.data_out(wire_d41_67),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4204168(.data_in(wire_d41_67),.data_out(wire_d41_68),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4204169(.data_in(wire_d41_68),.data_out(wire_d41_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204170(.data_in(wire_d41_69),.data_out(wire_d41_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4204171(.data_in(wire_d41_70),.data_out(wire_d41_71),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204172(.data_in(wire_d41_71),.data_out(wire_d41_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204173(.data_in(wire_d41_72),.data_out(wire_d41_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4204174(.data_in(wire_d41_73),.data_out(wire_d41_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4204175(.data_in(wire_d41_74),.data_out(wire_d41_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4204176(.data_in(wire_d41_75),.data_out(wire_d41_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204177(.data_in(wire_d41_76),.data_out(wire_d41_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204178(.data_in(wire_d41_77),.data_out(wire_d41_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4204179(.data_in(wire_d41_78),.data_out(wire_d41_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204180(.data_in(wire_d41_79),.data_out(wire_d41_80),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204181(.data_in(wire_d41_80),.data_out(wire_d41_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204182(.data_in(wire_d41_81),.data_out(wire_d41_82),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204183(.data_in(wire_d41_82),.data_out(wire_d41_83),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4204184(.data_in(wire_d41_83),.data_out(wire_d41_84),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204185(.data_in(wire_d41_84),.data_out(wire_d41_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4204186(.data_in(wire_d41_85),.data_out(wire_d41_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204187(.data_in(wire_d41_86),.data_out(wire_d41_87),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204188(.data_in(wire_d41_87),.data_out(wire_d41_88),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204189(.data_in(wire_d41_88),.data_out(wire_d41_89),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204190(.data_in(wire_d41_89),.data_out(wire_d41_90),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204191(.data_in(wire_d41_90),.data_out(wire_d41_91),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204192(.data_in(wire_d41_91),.data_out(wire_d41_92),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4204193(.data_in(wire_d41_92),.data_out(wire_d41_93),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204194(.data_in(wire_d41_93),.data_out(wire_d41_94),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204195(.data_in(wire_d41_94),.data_out(wire_d41_95),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204196(.data_in(wire_d41_95),.data_out(wire_d41_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4204197(.data_in(wire_d41_96),.data_out(wire_d41_97),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204198(.data_in(wire_d41_97),.data_out(wire_d41_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204199(.data_in(wire_d41_98),.data_out(wire_d41_99),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance42041100(.data_in(wire_d41_99),.data_out(wire_d41_100),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance42041101(.data_in(wire_d41_100),.data_out(wire_d41_101),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance42041102(.data_in(wire_d41_101),.data_out(wire_d41_102),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance42041103(.data_in(wire_d41_102),.data_out(wire_d41_103),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance42041104(.data_in(wire_d41_103),.data_out(wire_d41_104),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance42041105(.data_in(wire_d41_104),.data_out(wire_d41_105),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance42041106(.data_in(wire_d41_105),.data_out(wire_d41_106),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance42041107(.data_in(wire_d41_106),.data_out(wire_d41_107),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance42041108(.data_in(wire_d41_107),.data_out(wire_d41_108),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance42041109(.data_in(wire_d41_108),.data_out(wire_d41_109),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance42041110(.data_in(wire_d41_109),.data_out(wire_d41_110),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance42041111(.data_in(wire_d41_110),.data_out(wire_d41_111),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance42041112(.data_in(wire_d41_111),.data_out(wire_d41_112),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance42041113(.data_in(wire_d41_112),.data_out(wire_d41_113),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance42041114(.data_in(wire_d41_113),.data_out(wire_d41_114),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance42041115(.data_in(wire_d41_114),.data_out(wire_d41_115),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance42041116(.data_in(wire_d41_115),.data_out(wire_d41_116),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance42041117(.data_in(wire_d41_116),.data_out(wire_d41_117),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance42041118(.data_in(wire_d41_117),.data_out(wire_d41_118),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance42041119(.data_in(wire_d41_118),.data_out(d_out41),.clk(clk),.rst(rst));

	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance430420(.data_in(d_in42),.data_out(wire_d42_0),.clk(clk),.rst(rst));            //channel 43
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance430421(.data_in(wire_d42_0),.data_out(wire_d42_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance430422(.data_in(wire_d42_1),.data_out(wire_d42_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance430423(.data_in(wire_d42_2),.data_out(wire_d42_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance430424(.data_in(wire_d42_3),.data_out(wire_d42_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance430425(.data_in(wire_d42_4),.data_out(wire_d42_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance430426(.data_in(wire_d42_5),.data_out(wire_d42_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance430427(.data_in(wire_d42_6),.data_out(wire_d42_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance430428(.data_in(wire_d42_7),.data_out(wire_d42_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance430429(.data_in(wire_d42_8),.data_out(wire_d42_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304210(.data_in(wire_d42_9),.data_out(wire_d42_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304211(.data_in(wire_d42_10),.data_out(wire_d42_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304212(.data_in(wire_d42_11),.data_out(wire_d42_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304213(.data_in(wire_d42_12),.data_out(wire_d42_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304214(.data_in(wire_d42_13),.data_out(wire_d42_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4304215(.data_in(wire_d42_14),.data_out(wire_d42_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4304216(.data_in(wire_d42_15),.data_out(wire_d42_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304217(.data_in(wire_d42_16),.data_out(wire_d42_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304218(.data_in(wire_d42_17),.data_out(wire_d42_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304219(.data_in(wire_d42_18),.data_out(wire_d42_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4304220(.data_in(wire_d42_19),.data_out(wire_d42_20),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4304221(.data_in(wire_d42_20),.data_out(wire_d42_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304222(.data_in(wire_d42_21),.data_out(wire_d42_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4304223(.data_in(wire_d42_22),.data_out(wire_d42_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4304224(.data_in(wire_d42_23),.data_out(wire_d42_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4304225(.data_in(wire_d42_24),.data_out(wire_d42_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304226(.data_in(wire_d42_25),.data_out(wire_d42_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304227(.data_in(wire_d42_26),.data_out(wire_d42_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4304228(.data_in(wire_d42_27),.data_out(wire_d42_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304229(.data_in(wire_d42_28),.data_out(wire_d42_29),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304230(.data_in(wire_d42_29),.data_out(wire_d42_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304231(.data_in(wire_d42_30),.data_out(wire_d42_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304232(.data_in(wire_d42_31),.data_out(wire_d42_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304233(.data_in(wire_d42_32),.data_out(wire_d42_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4304234(.data_in(wire_d42_33),.data_out(wire_d42_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4304235(.data_in(wire_d42_34),.data_out(wire_d42_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304236(.data_in(wire_d42_35),.data_out(wire_d42_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304237(.data_in(wire_d42_36),.data_out(wire_d42_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304238(.data_in(wire_d42_37),.data_out(wire_d42_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304239(.data_in(wire_d42_38),.data_out(wire_d42_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304240(.data_in(wire_d42_39),.data_out(wire_d42_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304241(.data_in(wire_d42_40),.data_out(wire_d42_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304242(.data_in(wire_d42_41),.data_out(wire_d42_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304243(.data_in(wire_d42_42),.data_out(wire_d42_43),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4304244(.data_in(wire_d42_43),.data_out(wire_d42_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4304245(.data_in(wire_d42_44),.data_out(wire_d42_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304246(.data_in(wire_d42_45),.data_out(wire_d42_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304247(.data_in(wire_d42_46),.data_out(wire_d42_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304248(.data_in(wire_d42_47),.data_out(wire_d42_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304249(.data_in(wire_d42_48),.data_out(wire_d42_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304250(.data_in(wire_d42_49),.data_out(wire_d42_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304251(.data_in(wire_d42_50),.data_out(wire_d42_51),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4304252(.data_in(wire_d42_51),.data_out(wire_d42_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304253(.data_in(wire_d42_52),.data_out(wire_d42_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304254(.data_in(wire_d42_53),.data_out(wire_d42_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304255(.data_in(wire_d42_54),.data_out(wire_d42_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304256(.data_in(wire_d42_55),.data_out(wire_d42_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304257(.data_in(wire_d42_56),.data_out(wire_d42_57),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4304258(.data_in(wire_d42_57),.data_out(wire_d42_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304259(.data_in(wire_d42_58),.data_out(wire_d42_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304260(.data_in(wire_d42_59),.data_out(wire_d42_60),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304261(.data_in(wire_d42_60),.data_out(wire_d42_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4304262(.data_in(wire_d42_61),.data_out(wire_d42_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304263(.data_in(wire_d42_62),.data_out(wire_d42_63),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304264(.data_in(wire_d42_63),.data_out(wire_d42_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304265(.data_in(wire_d42_64),.data_out(wire_d42_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304266(.data_in(wire_d42_65),.data_out(wire_d42_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304267(.data_in(wire_d42_66),.data_out(wire_d42_67),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4304268(.data_in(wire_d42_67),.data_out(wire_d42_68),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4304269(.data_in(wire_d42_68),.data_out(wire_d42_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304270(.data_in(wire_d42_69),.data_out(wire_d42_70),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304271(.data_in(wire_d42_70),.data_out(wire_d42_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304272(.data_in(wire_d42_71),.data_out(wire_d42_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304273(.data_in(wire_d42_72),.data_out(wire_d42_73),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304274(.data_in(wire_d42_73),.data_out(wire_d42_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304275(.data_in(wire_d42_74),.data_out(wire_d42_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304276(.data_in(wire_d42_75),.data_out(wire_d42_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304277(.data_in(wire_d42_76),.data_out(wire_d42_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4304278(.data_in(wire_d42_77),.data_out(wire_d42_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4304279(.data_in(wire_d42_78),.data_out(wire_d42_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4304280(.data_in(wire_d42_79),.data_out(wire_d42_80),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304281(.data_in(wire_d42_80),.data_out(wire_d42_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4304282(.data_in(wire_d42_81),.data_out(wire_d42_82),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304283(.data_in(wire_d42_82),.data_out(wire_d42_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4304284(.data_in(wire_d42_83),.data_out(wire_d42_84),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304285(.data_in(wire_d42_84),.data_out(wire_d42_85),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304286(.data_in(wire_d42_85),.data_out(wire_d42_86),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304287(.data_in(wire_d42_86),.data_out(wire_d42_87),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304288(.data_in(wire_d42_87),.data_out(wire_d42_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4304289(.data_in(wire_d42_88),.data_out(wire_d42_89),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304290(.data_in(wire_d42_89),.data_out(wire_d42_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4304291(.data_in(wire_d42_90),.data_out(wire_d42_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4304292(.data_in(wire_d42_91),.data_out(wire_d42_92),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304293(.data_in(wire_d42_92),.data_out(wire_d42_93),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304294(.data_in(wire_d42_93),.data_out(wire_d42_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304295(.data_in(wire_d42_94),.data_out(wire_d42_95),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4304296(.data_in(wire_d42_95),.data_out(wire_d42_96),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304297(.data_in(wire_d42_96),.data_out(wire_d42_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304298(.data_in(wire_d42_97),.data_out(wire_d42_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4304299(.data_in(wire_d42_98),.data_out(wire_d42_99),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43042100(.data_in(wire_d42_99),.data_out(wire_d42_100),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance43042101(.data_in(wire_d42_100),.data_out(wire_d42_101),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance43042102(.data_in(wire_d42_101),.data_out(wire_d42_102),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance43042103(.data_in(wire_d42_102),.data_out(wire_d42_103),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance43042104(.data_in(wire_d42_103),.data_out(wire_d42_104),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance43042105(.data_in(wire_d42_104),.data_out(wire_d42_105),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance43042106(.data_in(wire_d42_105),.data_out(wire_d42_106),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance43042107(.data_in(wire_d42_106),.data_out(wire_d42_107),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance43042108(.data_in(wire_d42_107),.data_out(wire_d42_108),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance43042109(.data_in(wire_d42_108),.data_out(wire_d42_109),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance43042110(.data_in(wire_d42_109),.data_out(wire_d42_110),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43042111(.data_in(wire_d42_110),.data_out(wire_d42_111),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance43042112(.data_in(wire_d42_111),.data_out(wire_d42_112),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance43042113(.data_in(wire_d42_112),.data_out(wire_d42_113),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance43042114(.data_in(wire_d42_113),.data_out(wire_d42_114),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance43042115(.data_in(wire_d42_114),.data_out(wire_d42_115),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance43042116(.data_in(wire_d42_115),.data_out(wire_d42_116),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance43042117(.data_in(wire_d42_116),.data_out(wire_d42_117),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance43042118(.data_in(wire_d42_117),.data_out(wire_d42_118),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance43042119(.data_in(wire_d42_118),.data_out(d_out42),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance440430(.data_in(d_in43),.data_out(wire_d43_0),.clk(clk),.rst(rst));            //channel 44
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance440431(.data_in(wire_d43_0),.data_out(wire_d43_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance440432(.data_in(wire_d43_1),.data_out(wire_d43_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance440433(.data_in(wire_d43_2),.data_out(wire_d43_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance440434(.data_in(wire_d43_3),.data_out(wire_d43_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance440435(.data_in(wire_d43_4),.data_out(wire_d43_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance440436(.data_in(wire_d43_5),.data_out(wire_d43_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance440437(.data_in(wire_d43_6),.data_out(wire_d43_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance440438(.data_in(wire_d43_7),.data_out(wire_d43_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance440439(.data_in(wire_d43_8),.data_out(wire_d43_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404310(.data_in(wire_d43_9),.data_out(wire_d43_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404311(.data_in(wire_d43_10),.data_out(wire_d43_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404312(.data_in(wire_d43_11),.data_out(wire_d43_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404313(.data_in(wire_d43_12),.data_out(wire_d43_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404314(.data_in(wire_d43_13),.data_out(wire_d43_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404315(.data_in(wire_d43_14),.data_out(wire_d43_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404316(.data_in(wire_d43_15),.data_out(wire_d43_16),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4404317(.data_in(wire_d43_16),.data_out(wire_d43_17),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404318(.data_in(wire_d43_17),.data_out(wire_d43_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4404319(.data_in(wire_d43_18),.data_out(wire_d43_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404320(.data_in(wire_d43_19),.data_out(wire_d43_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4404321(.data_in(wire_d43_20),.data_out(wire_d43_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404322(.data_in(wire_d43_21),.data_out(wire_d43_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4404323(.data_in(wire_d43_22),.data_out(wire_d43_23),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4404324(.data_in(wire_d43_23),.data_out(wire_d43_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404325(.data_in(wire_d43_24),.data_out(wire_d43_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4404326(.data_in(wire_d43_25),.data_out(wire_d43_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4404327(.data_in(wire_d43_26),.data_out(wire_d43_27),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404328(.data_in(wire_d43_27),.data_out(wire_d43_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404329(.data_in(wire_d43_28),.data_out(wire_d43_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4404330(.data_in(wire_d43_29),.data_out(wire_d43_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404331(.data_in(wire_d43_30),.data_out(wire_d43_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404332(.data_in(wire_d43_31),.data_out(wire_d43_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4404333(.data_in(wire_d43_32),.data_out(wire_d43_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4404334(.data_in(wire_d43_33),.data_out(wire_d43_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404335(.data_in(wire_d43_34),.data_out(wire_d43_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404336(.data_in(wire_d43_35),.data_out(wire_d43_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4404337(.data_in(wire_d43_36),.data_out(wire_d43_37),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4404338(.data_in(wire_d43_37),.data_out(wire_d43_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404339(.data_in(wire_d43_38),.data_out(wire_d43_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404340(.data_in(wire_d43_39),.data_out(wire_d43_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4404341(.data_in(wire_d43_40),.data_out(wire_d43_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4404342(.data_in(wire_d43_41),.data_out(wire_d43_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404343(.data_in(wire_d43_42),.data_out(wire_d43_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404344(.data_in(wire_d43_43),.data_out(wire_d43_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404345(.data_in(wire_d43_44),.data_out(wire_d43_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4404346(.data_in(wire_d43_45),.data_out(wire_d43_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404347(.data_in(wire_d43_46),.data_out(wire_d43_47),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4404348(.data_in(wire_d43_47),.data_out(wire_d43_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404349(.data_in(wire_d43_48),.data_out(wire_d43_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4404350(.data_in(wire_d43_49),.data_out(wire_d43_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404351(.data_in(wire_d43_50),.data_out(wire_d43_51),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4404352(.data_in(wire_d43_51),.data_out(wire_d43_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404353(.data_in(wire_d43_52),.data_out(wire_d43_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4404354(.data_in(wire_d43_53),.data_out(wire_d43_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4404355(.data_in(wire_d43_54),.data_out(wire_d43_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4404356(.data_in(wire_d43_55),.data_out(wire_d43_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4404357(.data_in(wire_d43_56),.data_out(wire_d43_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404358(.data_in(wire_d43_57),.data_out(wire_d43_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404359(.data_in(wire_d43_58),.data_out(wire_d43_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4404360(.data_in(wire_d43_59),.data_out(wire_d43_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404361(.data_in(wire_d43_60),.data_out(wire_d43_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404362(.data_in(wire_d43_61),.data_out(wire_d43_62),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404363(.data_in(wire_d43_62),.data_out(wire_d43_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404364(.data_in(wire_d43_63),.data_out(wire_d43_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4404365(.data_in(wire_d43_64),.data_out(wire_d43_65),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4404366(.data_in(wire_d43_65),.data_out(wire_d43_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4404367(.data_in(wire_d43_66),.data_out(wire_d43_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404368(.data_in(wire_d43_67),.data_out(wire_d43_68),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404369(.data_in(wire_d43_68),.data_out(wire_d43_69),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404370(.data_in(wire_d43_69),.data_out(wire_d43_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404371(.data_in(wire_d43_70),.data_out(wire_d43_71),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404372(.data_in(wire_d43_71),.data_out(wire_d43_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404373(.data_in(wire_d43_72),.data_out(wire_d43_73),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404374(.data_in(wire_d43_73),.data_out(wire_d43_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4404375(.data_in(wire_d43_74),.data_out(wire_d43_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404376(.data_in(wire_d43_75),.data_out(wire_d43_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404377(.data_in(wire_d43_76),.data_out(wire_d43_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4404378(.data_in(wire_d43_77),.data_out(wire_d43_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4404379(.data_in(wire_d43_78),.data_out(wire_d43_79),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404380(.data_in(wire_d43_79),.data_out(wire_d43_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4404381(.data_in(wire_d43_80),.data_out(wire_d43_81),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404382(.data_in(wire_d43_81),.data_out(wire_d43_82),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404383(.data_in(wire_d43_82),.data_out(wire_d43_83),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404384(.data_in(wire_d43_83),.data_out(wire_d43_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404385(.data_in(wire_d43_84),.data_out(wire_d43_85),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404386(.data_in(wire_d43_85),.data_out(wire_d43_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4404387(.data_in(wire_d43_86),.data_out(wire_d43_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404388(.data_in(wire_d43_87),.data_out(wire_d43_88),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404389(.data_in(wire_d43_88),.data_out(wire_d43_89),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404390(.data_in(wire_d43_89),.data_out(wire_d43_90),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404391(.data_in(wire_d43_90),.data_out(wire_d43_91),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4404392(.data_in(wire_d43_91),.data_out(wire_d43_92),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4404393(.data_in(wire_d43_92),.data_out(wire_d43_93),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404394(.data_in(wire_d43_93),.data_out(wire_d43_94),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404395(.data_in(wire_d43_94),.data_out(wire_d43_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404396(.data_in(wire_d43_95),.data_out(wire_d43_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404397(.data_in(wire_d43_96),.data_out(wire_d43_97),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404398(.data_in(wire_d43_97),.data_out(wire_d43_98),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404399(.data_in(wire_d43_98),.data_out(wire_d43_99),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance44043100(.data_in(wire_d43_99),.data_out(wire_d43_100),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance44043101(.data_in(wire_d43_100),.data_out(wire_d43_101),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance44043102(.data_in(wire_d43_101),.data_out(wire_d43_102),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance44043103(.data_in(wire_d43_102),.data_out(wire_d43_103),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance44043104(.data_in(wire_d43_103),.data_out(wire_d43_104),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance44043105(.data_in(wire_d43_104),.data_out(wire_d43_105),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance44043106(.data_in(wire_d43_105),.data_out(wire_d43_106),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance44043107(.data_in(wire_d43_106),.data_out(wire_d43_107),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance44043108(.data_in(wire_d43_107),.data_out(wire_d43_108),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance44043109(.data_in(wire_d43_108),.data_out(wire_d43_109),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance44043110(.data_in(wire_d43_109),.data_out(wire_d43_110),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance44043111(.data_in(wire_d43_110),.data_out(wire_d43_111),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance44043112(.data_in(wire_d43_111),.data_out(wire_d43_112),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance44043113(.data_in(wire_d43_112),.data_out(wire_d43_113),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance44043114(.data_in(wire_d43_113),.data_out(wire_d43_114),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance44043115(.data_in(wire_d43_114),.data_out(wire_d43_115),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance44043116(.data_in(wire_d43_115),.data_out(wire_d43_116),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance44043117(.data_in(wire_d43_116),.data_out(wire_d43_117),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance44043118(.data_in(wire_d43_117),.data_out(wire_d43_118),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance44043119(.data_in(wire_d43_118),.data_out(d_out43),.clk(clk),.rst(rst));

	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance450440(.data_in(d_in44),.data_out(wire_d44_0),.clk(clk),.rst(rst));            //channel 45
	encoder #(.WIDTH(WIDTH)) encoder_instance450441(.data_in(wire_d44_0),.data_out(wire_d44_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance450442(.data_in(wire_d44_1),.data_out(wire_d44_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance450443(.data_in(wire_d44_2),.data_out(wire_d44_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance450444(.data_in(wire_d44_3),.data_out(wire_d44_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance450445(.data_in(wire_d44_4),.data_out(wire_d44_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance450446(.data_in(wire_d44_5),.data_out(wire_d44_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance450447(.data_in(wire_d44_6),.data_out(wire_d44_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance450448(.data_in(wire_d44_7),.data_out(wire_d44_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance450449(.data_in(wire_d44_8),.data_out(wire_d44_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504410(.data_in(wire_d44_9),.data_out(wire_d44_10),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4504411(.data_in(wire_d44_10),.data_out(wire_d44_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4504412(.data_in(wire_d44_11),.data_out(wire_d44_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504413(.data_in(wire_d44_12),.data_out(wire_d44_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4504414(.data_in(wire_d44_13),.data_out(wire_d44_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504415(.data_in(wire_d44_14),.data_out(wire_d44_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504416(.data_in(wire_d44_15),.data_out(wire_d44_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504417(.data_in(wire_d44_16),.data_out(wire_d44_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504418(.data_in(wire_d44_17),.data_out(wire_d44_18),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4504419(.data_in(wire_d44_18),.data_out(wire_d44_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504420(.data_in(wire_d44_19),.data_out(wire_d44_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4504421(.data_in(wire_d44_20),.data_out(wire_d44_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4504422(.data_in(wire_d44_21),.data_out(wire_d44_22),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4504423(.data_in(wire_d44_22),.data_out(wire_d44_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4504424(.data_in(wire_d44_23),.data_out(wire_d44_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504425(.data_in(wire_d44_24),.data_out(wire_d44_25),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4504426(.data_in(wire_d44_25),.data_out(wire_d44_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4504427(.data_in(wire_d44_26),.data_out(wire_d44_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504428(.data_in(wire_d44_27),.data_out(wire_d44_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504429(.data_in(wire_d44_28),.data_out(wire_d44_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504430(.data_in(wire_d44_29),.data_out(wire_d44_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4504431(.data_in(wire_d44_30),.data_out(wire_d44_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504432(.data_in(wire_d44_31),.data_out(wire_d44_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4504433(.data_in(wire_d44_32),.data_out(wire_d44_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504434(.data_in(wire_d44_33),.data_out(wire_d44_34),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4504435(.data_in(wire_d44_34),.data_out(wire_d44_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504436(.data_in(wire_d44_35),.data_out(wire_d44_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4504437(.data_in(wire_d44_36),.data_out(wire_d44_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504438(.data_in(wire_d44_37),.data_out(wire_d44_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4504439(.data_in(wire_d44_38),.data_out(wire_d44_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504440(.data_in(wire_d44_39),.data_out(wire_d44_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504441(.data_in(wire_d44_40),.data_out(wire_d44_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504442(.data_in(wire_d44_41),.data_out(wire_d44_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4504443(.data_in(wire_d44_42),.data_out(wire_d44_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4504444(.data_in(wire_d44_43),.data_out(wire_d44_44),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504445(.data_in(wire_d44_44),.data_out(wire_d44_45),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504446(.data_in(wire_d44_45),.data_out(wire_d44_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4504447(.data_in(wire_d44_46),.data_out(wire_d44_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4504448(.data_in(wire_d44_47),.data_out(wire_d44_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504449(.data_in(wire_d44_48),.data_out(wire_d44_49),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504450(.data_in(wire_d44_49),.data_out(wire_d44_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504451(.data_in(wire_d44_50),.data_out(wire_d44_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504452(.data_in(wire_d44_51),.data_out(wire_d44_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4504453(.data_in(wire_d44_52),.data_out(wire_d44_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4504454(.data_in(wire_d44_53),.data_out(wire_d44_54),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4504455(.data_in(wire_d44_54),.data_out(wire_d44_55),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504456(.data_in(wire_d44_55),.data_out(wire_d44_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504457(.data_in(wire_d44_56),.data_out(wire_d44_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4504458(.data_in(wire_d44_57),.data_out(wire_d44_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504459(.data_in(wire_d44_58),.data_out(wire_d44_59),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4504460(.data_in(wire_d44_59),.data_out(wire_d44_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4504461(.data_in(wire_d44_60),.data_out(wire_d44_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4504462(.data_in(wire_d44_61),.data_out(wire_d44_62),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504463(.data_in(wire_d44_62),.data_out(wire_d44_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504464(.data_in(wire_d44_63),.data_out(wire_d44_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504465(.data_in(wire_d44_64),.data_out(wire_d44_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504466(.data_in(wire_d44_65),.data_out(wire_d44_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4504467(.data_in(wire_d44_66),.data_out(wire_d44_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4504468(.data_in(wire_d44_67),.data_out(wire_d44_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4504469(.data_in(wire_d44_68),.data_out(wire_d44_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504470(.data_in(wire_d44_69),.data_out(wire_d44_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4504471(.data_in(wire_d44_70),.data_out(wire_d44_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504472(.data_in(wire_d44_71),.data_out(wire_d44_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504473(.data_in(wire_d44_72),.data_out(wire_d44_73),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504474(.data_in(wire_d44_73),.data_out(wire_d44_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504475(.data_in(wire_d44_74),.data_out(wire_d44_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4504476(.data_in(wire_d44_75),.data_out(wire_d44_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504477(.data_in(wire_d44_76),.data_out(wire_d44_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4504478(.data_in(wire_d44_77),.data_out(wire_d44_78),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504479(.data_in(wire_d44_78),.data_out(wire_d44_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504480(.data_in(wire_d44_79),.data_out(wire_d44_80),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504481(.data_in(wire_d44_80),.data_out(wire_d44_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4504482(.data_in(wire_d44_81),.data_out(wire_d44_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4504483(.data_in(wire_d44_82),.data_out(wire_d44_83),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504484(.data_in(wire_d44_83),.data_out(wire_d44_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504485(.data_in(wire_d44_84),.data_out(wire_d44_85),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504486(.data_in(wire_d44_85),.data_out(wire_d44_86),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4504487(.data_in(wire_d44_86),.data_out(wire_d44_87),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504488(.data_in(wire_d44_87),.data_out(wire_d44_88),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4504489(.data_in(wire_d44_88),.data_out(wire_d44_89),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4504490(.data_in(wire_d44_89),.data_out(wire_d44_90),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504491(.data_in(wire_d44_90),.data_out(wire_d44_91),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4504492(.data_in(wire_d44_91),.data_out(wire_d44_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4504493(.data_in(wire_d44_92),.data_out(wire_d44_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4504494(.data_in(wire_d44_93),.data_out(wire_d44_94),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504495(.data_in(wire_d44_94),.data_out(wire_d44_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4504496(.data_in(wire_d44_95),.data_out(wire_d44_96),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504497(.data_in(wire_d44_96),.data_out(wire_d44_97),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504498(.data_in(wire_d44_97),.data_out(wire_d44_98),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504499(.data_in(wire_d44_98),.data_out(wire_d44_99),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance45044100(.data_in(wire_d44_99),.data_out(wire_d44_100),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance45044101(.data_in(wire_d44_100),.data_out(wire_d44_101),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance45044102(.data_in(wire_d44_101),.data_out(wire_d44_102),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance45044103(.data_in(wire_d44_102),.data_out(wire_d44_103),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance45044104(.data_in(wire_d44_103),.data_out(wire_d44_104),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance45044105(.data_in(wire_d44_104),.data_out(wire_d44_105),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance45044106(.data_in(wire_d44_105),.data_out(wire_d44_106),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance45044107(.data_in(wire_d44_106),.data_out(wire_d44_107),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance45044108(.data_in(wire_d44_107),.data_out(wire_d44_108),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance45044109(.data_in(wire_d44_108),.data_out(wire_d44_109),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance45044110(.data_in(wire_d44_109),.data_out(wire_d44_110),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance45044111(.data_in(wire_d44_110),.data_out(wire_d44_111),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance45044112(.data_in(wire_d44_111),.data_out(wire_d44_112),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance45044113(.data_in(wire_d44_112),.data_out(wire_d44_113),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance45044114(.data_in(wire_d44_113),.data_out(wire_d44_114),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance45044115(.data_in(wire_d44_114),.data_out(wire_d44_115),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance45044116(.data_in(wire_d44_115),.data_out(wire_d44_116),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance45044117(.data_in(wire_d44_116),.data_out(wire_d44_117),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance45044118(.data_in(wire_d44_117),.data_out(wire_d44_118),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance45044119(.data_in(wire_d44_118),.data_out(d_out44),.clk(clk),.rst(rst));

	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance460450(.data_in(d_in45),.data_out(wire_d45_0),.clk(clk),.rst(rst));            //channel 46
	large_mux #(.WIDTH(WIDTH)) large_mux_instance460451(.data_in(wire_d45_0),.data_out(wire_d45_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance460452(.data_in(wire_d45_1),.data_out(wire_d45_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance460453(.data_in(wire_d45_2),.data_out(wire_d45_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance460454(.data_in(wire_d45_3),.data_out(wire_d45_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance460455(.data_in(wire_d45_4),.data_out(wire_d45_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance460456(.data_in(wire_d45_5),.data_out(wire_d45_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance460457(.data_in(wire_d45_6),.data_out(wire_d45_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance460458(.data_in(wire_d45_7),.data_out(wire_d45_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance460459(.data_in(wire_d45_8),.data_out(wire_d45_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604510(.data_in(wire_d45_9),.data_out(wire_d45_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4604511(.data_in(wire_d45_10),.data_out(wire_d45_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604512(.data_in(wire_d45_11),.data_out(wire_d45_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604513(.data_in(wire_d45_12),.data_out(wire_d45_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4604514(.data_in(wire_d45_13),.data_out(wire_d45_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604515(.data_in(wire_d45_14),.data_out(wire_d45_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4604516(.data_in(wire_d45_15),.data_out(wire_d45_16),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4604517(.data_in(wire_d45_16),.data_out(wire_d45_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604518(.data_in(wire_d45_17),.data_out(wire_d45_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604519(.data_in(wire_d45_18),.data_out(wire_d45_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4604520(.data_in(wire_d45_19),.data_out(wire_d45_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4604521(.data_in(wire_d45_20),.data_out(wire_d45_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604522(.data_in(wire_d45_21),.data_out(wire_d45_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604523(.data_in(wire_d45_22),.data_out(wire_d45_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4604524(.data_in(wire_d45_23),.data_out(wire_d45_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604525(.data_in(wire_d45_24),.data_out(wire_d45_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604526(.data_in(wire_d45_25),.data_out(wire_d45_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604527(.data_in(wire_d45_26),.data_out(wire_d45_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604528(.data_in(wire_d45_27),.data_out(wire_d45_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4604529(.data_in(wire_d45_28),.data_out(wire_d45_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4604530(.data_in(wire_d45_29),.data_out(wire_d45_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4604531(.data_in(wire_d45_30),.data_out(wire_d45_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604532(.data_in(wire_d45_31),.data_out(wire_d45_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4604533(.data_in(wire_d45_32),.data_out(wire_d45_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4604534(.data_in(wire_d45_33),.data_out(wire_d45_34),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604535(.data_in(wire_d45_34),.data_out(wire_d45_35),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4604536(.data_in(wire_d45_35),.data_out(wire_d45_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4604537(.data_in(wire_d45_36),.data_out(wire_d45_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4604538(.data_in(wire_d45_37),.data_out(wire_d45_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4604539(.data_in(wire_d45_38),.data_out(wire_d45_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604540(.data_in(wire_d45_39),.data_out(wire_d45_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4604541(.data_in(wire_d45_40),.data_out(wire_d45_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604542(.data_in(wire_d45_41),.data_out(wire_d45_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4604543(.data_in(wire_d45_42),.data_out(wire_d45_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604544(.data_in(wire_d45_43),.data_out(wire_d45_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604545(.data_in(wire_d45_44),.data_out(wire_d45_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4604546(.data_in(wire_d45_45),.data_out(wire_d45_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4604547(.data_in(wire_d45_46),.data_out(wire_d45_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604548(.data_in(wire_d45_47),.data_out(wire_d45_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604549(.data_in(wire_d45_48),.data_out(wire_d45_49),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4604550(.data_in(wire_d45_49),.data_out(wire_d45_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4604551(.data_in(wire_d45_50),.data_out(wire_d45_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604552(.data_in(wire_d45_51),.data_out(wire_d45_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604553(.data_in(wire_d45_52),.data_out(wire_d45_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4604554(.data_in(wire_d45_53),.data_out(wire_d45_54),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4604555(.data_in(wire_d45_54),.data_out(wire_d45_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604556(.data_in(wire_d45_55),.data_out(wire_d45_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4604557(.data_in(wire_d45_56),.data_out(wire_d45_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4604558(.data_in(wire_d45_57),.data_out(wire_d45_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4604559(.data_in(wire_d45_58),.data_out(wire_d45_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4604560(.data_in(wire_d45_59),.data_out(wire_d45_60),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604561(.data_in(wire_d45_60),.data_out(wire_d45_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604562(.data_in(wire_d45_61),.data_out(wire_d45_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4604563(.data_in(wire_d45_62),.data_out(wire_d45_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604564(.data_in(wire_d45_63),.data_out(wire_d45_64),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604565(.data_in(wire_d45_64),.data_out(wire_d45_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4604566(.data_in(wire_d45_65),.data_out(wire_d45_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4604567(.data_in(wire_d45_66),.data_out(wire_d45_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4604568(.data_in(wire_d45_67),.data_out(wire_d45_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604569(.data_in(wire_d45_68),.data_out(wire_d45_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4604570(.data_in(wire_d45_69),.data_out(wire_d45_70),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4604571(.data_in(wire_d45_70),.data_out(wire_d45_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4604572(.data_in(wire_d45_71),.data_out(wire_d45_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604573(.data_in(wire_d45_72),.data_out(wire_d45_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604574(.data_in(wire_d45_73),.data_out(wire_d45_74),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4604575(.data_in(wire_d45_74),.data_out(wire_d45_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4604576(.data_in(wire_d45_75),.data_out(wire_d45_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4604577(.data_in(wire_d45_76),.data_out(wire_d45_77),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4604578(.data_in(wire_d45_77),.data_out(wire_d45_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604579(.data_in(wire_d45_78),.data_out(wire_d45_79),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604580(.data_in(wire_d45_79),.data_out(wire_d45_80),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4604581(.data_in(wire_d45_80),.data_out(wire_d45_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4604582(.data_in(wire_d45_81),.data_out(wire_d45_82),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4604583(.data_in(wire_d45_82),.data_out(wire_d45_83),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604584(.data_in(wire_d45_83),.data_out(wire_d45_84),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4604585(.data_in(wire_d45_84),.data_out(wire_d45_85),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604586(.data_in(wire_d45_85),.data_out(wire_d45_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4604587(.data_in(wire_d45_86),.data_out(wire_d45_87),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604588(.data_in(wire_d45_87),.data_out(wire_d45_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4604589(.data_in(wire_d45_88),.data_out(wire_d45_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4604590(.data_in(wire_d45_89),.data_out(wire_d45_90),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4604591(.data_in(wire_d45_90),.data_out(wire_d45_91),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604592(.data_in(wire_d45_91),.data_out(wire_d45_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4604593(.data_in(wire_d45_92),.data_out(wire_d45_93),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4604594(.data_in(wire_d45_93),.data_out(wire_d45_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4604595(.data_in(wire_d45_94),.data_out(wire_d45_95),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604596(.data_in(wire_d45_95),.data_out(wire_d45_96),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4604597(.data_in(wire_d45_96),.data_out(wire_d45_97),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604598(.data_in(wire_d45_97),.data_out(wire_d45_98),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604599(.data_in(wire_d45_98),.data_out(wire_d45_99),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance46045100(.data_in(wire_d45_99),.data_out(wire_d45_100),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance46045101(.data_in(wire_d45_100),.data_out(wire_d45_101),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance46045102(.data_in(wire_d45_101),.data_out(wire_d45_102),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance46045103(.data_in(wire_d45_102),.data_out(wire_d45_103),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance46045104(.data_in(wire_d45_103),.data_out(wire_d45_104),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance46045105(.data_in(wire_d45_104),.data_out(wire_d45_105),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance46045106(.data_in(wire_d45_105),.data_out(wire_d45_106),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance46045107(.data_in(wire_d45_106),.data_out(wire_d45_107),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance46045108(.data_in(wire_d45_107),.data_out(wire_d45_108),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance46045109(.data_in(wire_d45_108),.data_out(wire_d45_109),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance46045110(.data_in(wire_d45_109),.data_out(wire_d45_110),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance46045111(.data_in(wire_d45_110),.data_out(wire_d45_111),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance46045112(.data_in(wire_d45_111),.data_out(wire_d45_112),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance46045113(.data_in(wire_d45_112),.data_out(wire_d45_113),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance46045114(.data_in(wire_d45_113),.data_out(wire_d45_114),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance46045115(.data_in(wire_d45_114),.data_out(wire_d45_115),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance46045116(.data_in(wire_d45_115),.data_out(wire_d45_116),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance46045117(.data_in(wire_d45_116),.data_out(wire_d45_117),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance46045118(.data_in(wire_d45_117),.data_out(wire_d45_118),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance46045119(.data_in(wire_d45_118),.data_out(d_out45),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance470460(.data_in(d_in46),.data_out(wire_d46_0),.clk(clk),.rst(rst));            //channel 47
	register #(.WIDTH(WIDTH)) register_instance470461(.data_in(wire_d46_0),.data_out(wire_d46_1),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance470462(.data_in(wire_d46_1),.data_out(wire_d46_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance470463(.data_in(wire_d46_2),.data_out(wire_d46_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance470464(.data_in(wire_d46_3),.data_out(wire_d46_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance470465(.data_in(wire_d46_4),.data_out(wire_d46_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance470466(.data_in(wire_d46_5),.data_out(wire_d46_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance470467(.data_in(wire_d46_6),.data_out(wire_d46_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance470468(.data_in(wire_d46_7),.data_out(wire_d46_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance470469(.data_in(wire_d46_8),.data_out(wire_d46_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4704610(.data_in(wire_d46_9),.data_out(wire_d46_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704611(.data_in(wire_d46_10),.data_out(wire_d46_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4704612(.data_in(wire_d46_11),.data_out(wire_d46_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704613(.data_in(wire_d46_12),.data_out(wire_d46_13),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704614(.data_in(wire_d46_13),.data_out(wire_d46_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704615(.data_in(wire_d46_14),.data_out(wire_d46_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704616(.data_in(wire_d46_15),.data_out(wire_d46_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704617(.data_in(wire_d46_16),.data_out(wire_d46_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704618(.data_in(wire_d46_17),.data_out(wire_d46_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704619(.data_in(wire_d46_18),.data_out(wire_d46_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704620(.data_in(wire_d46_19),.data_out(wire_d46_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4704621(.data_in(wire_d46_20),.data_out(wire_d46_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4704622(.data_in(wire_d46_21),.data_out(wire_d46_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4704623(.data_in(wire_d46_22),.data_out(wire_d46_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4704624(.data_in(wire_d46_23),.data_out(wire_d46_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704625(.data_in(wire_d46_24),.data_out(wire_d46_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704626(.data_in(wire_d46_25),.data_out(wire_d46_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704627(.data_in(wire_d46_26),.data_out(wire_d46_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4704628(.data_in(wire_d46_27),.data_out(wire_d46_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704629(.data_in(wire_d46_28),.data_out(wire_d46_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704630(.data_in(wire_d46_29),.data_out(wire_d46_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704631(.data_in(wire_d46_30),.data_out(wire_d46_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4704632(.data_in(wire_d46_31),.data_out(wire_d46_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704633(.data_in(wire_d46_32),.data_out(wire_d46_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4704634(.data_in(wire_d46_33),.data_out(wire_d46_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4704635(.data_in(wire_d46_34),.data_out(wire_d46_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704636(.data_in(wire_d46_35),.data_out(wire_d46_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704637(.data_in(wire_d46_36),.data_out(wire_d46_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4704638(.data_in(wire_d46_37),.data_out(wire_d46_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704639(.data_in(wire_d46_38),.data_out(wire_d46_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4704640(.data_in(wire_d46_39),.data_out(wire_d46_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704641(.data_in(wire_d46_40),.data_out(wire_d46_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704642(.data_in(wire_d46_41),.data_out(wire_d46_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4704643(.data_in(wire_d46_42),.data_out(wire_d46_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4704644(.data_in(wire_d46_43),.data_out(wire_d46_44),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704645(.data_in(wire_d46_44),.data_out(wire_d46_45),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704646(.data_in(wire_d46_45),.data_out(wire_d46_46),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704647(.data_in(wire_d46_46),.data_out(wire_d46_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704648(.data_in(wire_d46_47),.data_out(wire_d46_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704649(.data_in(wire_d46_48),.data_out(wire_d46_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704650(.data_in(wire_d46_49),.data_out(wire_d46_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704651(.data_in(wire_d46_50),.data_out(wire_d46_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4704652(.data_in(wire_d46_51),.data_out(wire_d46_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704653(.data_in(wire_d46_52),.data_out(wire_d46_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4704654(.data_in(wire_d46_53),.data_out(wire_d46_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704655(.data_in(wire_d46_54),.data_out(wire_d46_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4704656(.data_in(wire_d46_55),.data_out(wire_d46_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704657(.data_in(wire_d46_56),.data_out(wire_d46_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704658(.data_in(wire_d46_57),.data_out(wire_d46_58),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4704659(.data_in(wire_d46_58),.data_out(wire_d46_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704660(.data_in(wire_d46_59),.data_out(wire_d46_60),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4704661(.data_in(wire_d46_60),.data_out(wire_d46_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704662(.data_in(wire_d46_61),.data_out(wire_d46_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704663(.data_in(wire_d46_62),.data_out(wire_d46_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704664(.data_in(wire_d46_63),.data_out(wire_d46_64),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704665(.data_in(wire_d46_64),.data_out(wire_d46_65),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4704666(.data_in(wire_d46_65),.data_out(wire_d46_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704667(.data_in(wire_d46_66),.data_out(wire_d46_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704668(.data_in(wire_d46_67),.data_out(wire_d46_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704669(.data_in(wire_d46_68),.data_out(wire_d46_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704670(.data_in(wire_d46_69),.data_out(wire_d46_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4704671(.data_in(wire_d46_70),.data_out(wire_d46_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4704672(.data_in(wire_d46_71),.data_out(wire_d46_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704673(.data_in(wire_d46_72),.data_out(wire_d46_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4704674(.data_in(wire_d46_73),.data_out(wire_d46_74),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4704675(.data_in(wire_d46_74),.data_out(wire_d46_75),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4704676(.data_in(wire_d46_75),.data_out(wire_d46_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4704677(.data_in(wire_d46_76),.data_out(wire_d46_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704678(.data_in(wire_d46_77),.data_out(wire_d46_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704679(.data_in(wire_d46_78),.data_out(wire_d46_79),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704680(.data_in(wire_d46_79),.data_out(wire_d46_80),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704681(.data_in(wire_d46_80),.data_out(wire_d46_81),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4704682(.data_in(wire_d46_81),.data_out(wire_d46_82),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704683(.data_in(wire_d46_82),.data_out(wire_d46_83),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4704684(.data_in(wire_d46_83),.data_out(wire_d46_84),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704685(.data_in(wire_d46_84),.data_out(wire_d46_85),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704686(.data_in(wire_d46_85),.data_out(wire_d46_86),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4704687(.data_in(wire_d46_86),.data_out(wire_d46_87),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704688(.data_in(wire_d46_87),.data_out(wire_d46_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4704689(.data_in(wire_d46_88),.data_out(wire_d46_89),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704690(.data_in(wire_d46_89),.data_out(wire_d46_90),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704691(.data_in(wire_d46_90),.data_out(wire_d46_91),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704692(.data_in(wire_d46_91),.data_out(wire_d46_92),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4704693(.data_in(wire_d46_92),.data_out(wire_d46_93),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704694(.data_in(wire_d46_93),.data_out(wire_d46_94),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4704695(.data_in(wire_d46_94),.data_out(wire_d46_95),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704696(.data_in(wire_d46_95),.data_out(wire_d46_96),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704697(.data_in(wire_d46_96),.data_out(wire_d46_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4704698(.data_in(wire_d46_97),.data_out(wire_d46_98),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4704699(.data_in(wire_d46_98),.data_out(wire_d46_99),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance47046100(.data_in(wire_d46_99),.data_out(wire_d46_100),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance47046101(.data_in(wire_d46_100),.data_out(wire_d46_101),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance47046102(.data_in(wire_d46_101),.data_out(wire_d46_102),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance47046103(.data_in(wire_d46_102),.data_out(wire_d46_103),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance47046104(.data_in(wire_d46_103),.data_out(wire_d46_104),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance47046105(.data_in(wire_d46_104),.data_out(wire_d46_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance47046106(.data_in(wire_d46_105),.data_out(wire_d46_106),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance47046107(.data_in(wire_d46_106),.data_out(wire_d46_107),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance47046108(.data_in(wire_d46_107),.data_out(wire_d46_108),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance47046109(.data_in(wire_d46_108),.data_out(wire_d46_109),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance47046110(.data_in(wire_d46_109),.data_out(wire_d46_110),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance47046111(.data_in(wire_d46_110),.data_out(wire_d46_111),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance47046112(.data_in(wire_d46_111),.data_out(wire_d46_112),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance47046113(.data_in(wire_d46_112),.data_out(wire_d46_113),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance47046114(.data_in(wire_d46_113),.data_out(wire_d46_114),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance47046115(.data_in(wire_d46_114),.data_out(wire_d46_115),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance47046116(.data_in(wire_d46_115),.data_out(wire_d46_116),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance47046117(.data_in(wire_d46_116),.data_out(wire_d46_117),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance47046118(.data_in(wire_d46_117),.data_out(wire_d46_118),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance47046119(.data_in(wire_d46_118),.data_out(d_out46),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance480470(.data_in(d_in47),.data_out(wire_d47_0),.clk(clk),.rst(rst));            //channel 48
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance480471(.data_in(wire_d47_0),.data_out(wire_d47_1),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance480472(.data_in(wire_d47_1),.data_out(wire_d47_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance480473(.data_in(wire_d47_2),.data_out(wire_d47_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance480474(.data_in(wire_d47_3),.data_out(wire_d47_4),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance480475(.data_in(wire_d47_4),.data_out(wire_d47_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance480476(.data_in(wire_d47_5),.data_out(wire_d47_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance480477(.data_in(wire_d47_6),.data_out(wire_d47_7),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance480478(.data_in(wire_d47_7),.data_out(wire_d47_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance480479(.data_in(wire_d47_8),.data_out(wire_d47_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804710(.data_in(wire_d47_9),.data_out(wire_d47_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4804711(.data_in(wire_d47_10),.data_out(wire_d47_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804712(.data_in(wire_d47_11),.data_out(wire_d47_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804713(.data_in(wire_d47_12),.data_out(wire_d47_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4804714(.data_in(wire_d47_13),.data_out(wire_d47_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804715(.data_in(wire_d47_14),.data_out(wire_d47_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4804716(.data_in(wire_d47_15),.data_out(wire_d47_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4804717(.data_in(wire_d47_16),.data_out(wire_d47_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4804718(.data_in(wire_d47_17),.data_out(wire_d47_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804719(.data_in(wire_d47_18),.data_out(wire_d47_19),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4804720(.data_in(wire_d47_19),.data_out(wire_d47_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4804721(.data_in(wire_d47_20),.data_out(wire_d47_21),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4804722(.data_in(wire_d47_21),.data_out(wire_d47_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804723(.data_in(wire_d47_22),.data_out(wire_d47_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4804724(.data_in(wire_d47_23),.data_out(wire_d47_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804725(.data_in(wire_d47_24),.data_out(wire_d47_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804726(.data_in(wire_d47_25),.data_out(wire_d47_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804727(.data_in(wire_d47_26),.data_out(wire_d47_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804728(.data_in(wire_d47_27),.data_out(wire_d47_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4804729(.data_in(wire_d47_28),.data_out(wire_d47_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804730(.data_in(wire_d47_29),.data_out(wire_d47_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4804731(.data_in(wire_d47_30),.data_out(wire_d47_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804732(.data_in(wire_d47_31),.data_out(wire_d47_32),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804733(.data_in(wire_d47_32),.data_out(wire_d47_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804734(.data_in(wire_d47_33),.data_out(wire_d47_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4804735(.data_in(wire_d47_34),.data_out(wire_d47_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4804736(.data_in(wire_d47_35),.data_out(wire_d47_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4804737(.data_in(wire_d47_36),.data_out(wire_d47_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4804738(.data_in(wire_d47_37),.data_out(wire_d47_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804739(.data_in(wire_d47_38),.data_out(wire_d47_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804740(.data_in(wire_d47_39),.data_out(wire_d47_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4804741(.data_in(wire_d47_40),.data_out(wire_d47_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804742(.data_in(wire_d47_41),.data_out(wire_d47_42),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804743(.data_in(wire_d47_42),.data_out(wire_d47_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804744(.data_in(wire_d47_43),.data_out(wire_d47_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804745(.data_in(wire_d47_44),.data_out(wire_d47_45),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804746(.data_in(wire_d47_45),.data_out(wire_d47_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804747(.data_in(wire_d47_46),.data_out(wire_d47_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804748(.data_in(wire_d47_47),.data_out(wire_d47_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4804749(.data_in(wire_d47_48),.data_out(wire_d47_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804750(.data_in(wire_d47_49),.data_out(wire_d47_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804751(.data_in(wire_d47_50),.data_out(wire_d47_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804752(.data_in(wire_d47_51),.data_out(wire_d47_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804753(.data_in(wire_d47_52),.data_out(wire_d47_53),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804754(.data_in(wire_d47_53),.data_out(wire_d47_54),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4804755(.data_in(wire_d47_54),.data_out(wire_d47_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804756(.data_in(wire_d47_55),.data_out(wire_d47_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804757(.data_in(wire_d47_56),.data_out(wire_d47_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4804758(.data_in(wire_d47_57),.data_out(wire_d47_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4804759(.data_in(wire_d47_58),.data_out(wire_d47_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804760(.data_in(wire_d47_59),.data_out(wire_d47_60),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804761(.data_in(wire_d47_60),.data_out(wire_d47_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4804762(.data_in(wire_d47_61),.data_out(wire_d47_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804763(.data_in(wire_d47_62),.data_out(wire_d47_63),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804764(.data_in(wire_d47_63),.data_out(wire_d47_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804765(.data_in(wire_d47_64),.data_out(wire_d47_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804766(.data_in(wire_d47_65),.data_out(wire_d47_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4804767(.data_in(wire_d47_66),.data_out(wire_d47_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4804768(.data_in(wire_d47_67),.data_out(wire_d47_68),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804769(.data_in(wire_d47_68),.data_out(wire_d47_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4804770(.data_in(wire_d47_69),.data_out(wire_d47_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4804771(.data_in(wire_d47_70),.data_out(wire_d47_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804772(.data_in(wire_d47_71),.data_out(wire_d47_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4804773(.data_in(wire_d47_72),.data_out(wire_d47_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804774(.data_in(wire_d47_73),.data_out(wire_d47_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804775(.data_in(wire_d47_74),.data_out(wire_d47_75),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804776(.data_in(wire_d47_75),.data_out(wire_d47_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804777(.data_in(wire_d47_76),.data_out(wire_d47_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804778(.data_in(wire_d47_77),.data_out(wire_d47_78),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804779(.data_in(wire_d47_78),.data_out(wire_d47_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4804780(.data_in(wire_d47_79),.data_out(wire_d47_80),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804781(.data_in(wire_d47_80),.data_out(wire_d47_81),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804782(.data_in(wire_d47_81),.data_out(wire_d47_82),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4804783(.data_in(wire_d47_82),.data_out(wire_d47_83),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4804784(.data_in(wire_d47_83),.data_out(wire_d47_84),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804785(.data_in(wire_d47_84),.data_out(wire_d47_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4804786(.data_in(wire_d47_85),.data_out(wire_d47_86),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4804787(.data_in(wire_d47_86),.data_out(wire_d47_87),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804788(.data_in(wire_d47_87),.data_out(wire_d47_88),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804789(.data_in(wire_d47_88),.data_out(wire_d47_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4804790(.data_in(wire_d47_89),.data_out(wire_d47_90),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804791(.data_in(wire_d47_90),.data_out(wire_d47_91),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804792(.data_in(wire_d47_91),.data_out(wire_d47_92),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804793(.data_in(wire_d47_92),.data_out(wire_d47_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804794(.data_in(wire_d47_93),.data_out(wire_d47_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804795(.data_in(wire_d47_94),.data_out(wire_d47_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804796(.data_in(wire_d47_95),.data_out(wire_d47_96),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804797(.data_in(wire_d47_96),.data_out(wire_d47_97),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804798(.data_in(wire_d47_97),.data_out(wire_d47_98),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804799(.data_in(wire_d47_98),.data_out(wire_d47_99),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance48047100(.data_in(wire_d47_99),.data_out(wire_d47_100),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance48047101(.data_in(wire_d47_100),.data_out(wire_d47_101),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance48047102(.data_in(wire_d47_101),.data_out(wire_d47_102),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance48047103(.data_in(wire_d47_102),.data_out(wire_d47_103),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance48047104(.data_in(wire_d47_103),.data_out(wire_d47_104),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance48047105(.data_in(wire_d47_104),.data_out(wire_d47_105),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance48047106(.data_in(wire_d47_105),.data_out(wire_d47_106),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance48047107(.data_in(wire_d47_106),.data_out(wire_d47_107),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance48047108(.data_in(wire_d47_107),.data_out(wire_d47_108),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance48047109(.data_in(wire_d47_108),.data_out(wire_d47_109),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance48047110(.data_in(wire_d47_109),.data_out(wire_d47_110),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance48047111(.data_in(wire_d47_110),.data_out(wire_d47_111),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance48047112(.data_in(wire_d47_111),.data_out(wire_d47_112),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance48047113(.data_in(wire_d47_112),.data_out(wire_d47_113),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance48047114(.data_in(wire_d47_113),.data_out(wire_d47_114),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance48047115(.data_in(wire_d47_114),.data_out(wire_d47_115),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance48047116(.data_in(wire_d47_115),.data_out(wire_d47_116),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance48047117(.data_in(wire_d47_116),.data_out(wire_d47_117),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance48047118(.data_in(wire_d47_117),.data_out(wire_d47_118),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance48047119(.data_in(wire_d47_118),.data_out(d_out47),.clk(clk),.rst(rst));

	large_adder #(.WIDTH(WIDTH)) large_adder_instance490480(.data_in(d_in48),.data_out(wire_d48_0),.clk(clk),.rst(rst));            //channel 49
	encoder #(.WIDTH(WIDTH)) encoder_instance490481(.data_in(wire_d48_0),.data_out(wire_d48_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance490482(.data_in(wire_d48_1),.data_out(wire_d48_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance490483(.data_in(wire_d48_2),.data_out(wire_d48_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance490484(.data_in(wire_d48_3),.data_out(wire_d48_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance490485(.data_in(wire_d48_4),.data_out(wire_d48_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance490486(.data_in(wire_d48_5),.data_out(wire_d48_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance490487(.data_in(wire_d48_6),.data_out(wire_d48_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance490488(.data_in(wire_d48_7),.data_out(wire_d48_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance490489(.data_in(wire_d48_8),.data_out(wire_d48_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904810(.data_in(wire_d48_9),.data_out(wire_d48_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904811(.data_in(wire_d48_10),.data_out(wire_d48_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904812(.data_in(wire_d48_11),.data_out(wire_d48_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904813(.data_in(wire_d48_12),.data_out(wire_d48_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4904814(.data_in(wire_d48_13),.data_out(wire_d48_14),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904815(.data_in(wire_d48_14),.data_out(wire_d48_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904816(.data_in(wire_d48_15),.data_out(wire_d48_16),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4904817(.data_in(wire_d48_16),.data_out(wire_d48_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904818(.data_in(wire_d48_17),.data_out(wire_d48_18),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4904819(.data_in(wire_d48_18),.data_out(wire_d48_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904820(.data_in(wire_d48_19),.data_out(wire_d48_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4904821(.data_in(wire_d48_20),.data_out(wire_d48_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904822(.data_in(wire_d48_21),.data_out(wire_d48_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4904823(.data_in(wire_d48_22),.data_out(wire_d48_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4904824(.data_in(wire_d48_23),.data_out(wire_d48_24),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904825(.data_in(wire_d48_24),.data_out(wire_d48_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4904826(.data_in(wire_d48_25),.data_out(wire_d48_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4904827(.data_in(wire_d48_26),.data_out(wire_d48_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904828(.data_in(wire_d48_27),.data_out(wire_d48_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904829(.data_in(wire_d48_28),.data_out(wire_d48_29),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904830(.data_in(wire_d48_29),.data_out(wire_d48_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4904831(.data_in(wire_d48_30),.data_out(wire_d48_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904832(.data_in(wire_d48_31),.data_out(wire_d48_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904833(.data_in(wire_d48_32),.data_out(wire_d48_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4904834(.data_in(wire_d48_33),.data_out(wire_d48_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904835(.data_in(wire_d48_34),.data_out(wire_d48_35),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4904836(.data_in(wire_d48_35),.data_out(wire_d48_36),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904837(.data_in(wire_d48_36),.data_out(wire_d48_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4904838(.data_in(wire_d48_37),.data_out(wire_d48_38),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4904839(.data_in(wire_d48_38),.data_out(wire_d48_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904840(.data_in(wire_d48_39),.data_out(wire_d48_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4904841(.data_in(wire_d48_40),.data_out(wire_d48_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904842(.data_in(wire_d48_41),.data_out(wire_d48_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4904843(.data_in(wire_d48_42),.data_out(wire_d48_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904844(.data_in(wire_d48_43),.data_out(wire_d48_44),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904845(.data_in(wire_d48_44),.data_out(wire_d48_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904846(.data_in(wire_d48_45),.data_out(wire_d48_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4904847(.data_in(wire_d48_46),.data_out(wire_d48_47),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4904848(.data_in(wire_d48_47),.data_out(wire_d48_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4904849(.data_in(wire_d48_48),.data_out(wire_d48_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904850(.data_in(wire_d48_49),.data_out(wire_d48_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4904851(.data_in(wire_d48_50),.data_out(wire_d48_51),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904852(.data_in(wire_d48_51),.data_out(wire_d48_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904853(.data_in(wire_d48_52),.data_out(wire_d48_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4904854(.data_in(wire_d48_53),.data_out(wire_d48_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904855(.data_in(wire_d48_54),.data_out(wire_d48_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904856(.data_in(wire_d48_55),.data_out(wire_d48_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904857(.data_in(wire_d48_56),.data_out(wire_d48_57),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4904858(.data_in(wire_d48_57),.data_out(wire_d48_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904859(.data_in(wire_d48_58),.data_out(wire_d48_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904860(.data_in(wire_d48_59),.data_out(wire_d48_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4904861(.data_in(wire_d48_60),.data_out(wire_d48_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904862(.data_in(wire_d48_61),.data_out(wire_d48_62),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4904863(.data_in(wire_d48_62),.data_out(wire_d48_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4904864(.data_in(wire_d48_63),.data_out(wire_d48_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904865(.data_in(wire_d48_64),.data_out(wire_d48_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4904866(.data_in(wire_d48_65),.data_out(wire_d48_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904867(.data_in(wire_d48_66),.data_out(wire_d48_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904868(.data_in(wire_d48_67),.data_out(wire_d48_68),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904869(.data_in(wire_d48_68),.data_out(wire_d48_69),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904870(.data_in(wire_d48_69),.data_out(wire_d48_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904871(.data_in(wire_d48_70),.data_out(wire_d48_71),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904872(.data_in(wire_d48_71),.data_out(wire_d48_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904873(.data_in(wire_d48_72),.data_out(wire_d48_73),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4904874(.data_in(wire_d48_73),.data_out(wire_d48_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904875(.data_in(wire_d48_74),.data_out(wire_d48_75),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904876(.data_in(wire_d48_75),.data_out(wire_d48_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4904877(.data_in(wire_d48_76),.data_out(wire_d48_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904878(.data_in(wire_d48_77),.data_out(wire_d48_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904879(.data_in(wire_d48_78),.data_out(wire_d48_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4904880(.data_in(wire_d48_79),.data_out(wire_d48_80),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904881(.data_in(wire_d48_80),.data_out(wire_d48_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4904882(.data_in(wire_d48_81),.data_out(wire_d48_82),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4904883(.data_in(wire_d48_82),.data_out(wire_d48_83),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904884(.data_in(wire_d48_83),.data_out(wire_d48_84),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4904885(.data_in(wire_d48_84),.data_out(wire_d48_85),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904886(.data_in(wire_d48_85),.data_out(wire_d48_86),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904887(.data_in(wire_d48_86),.data_out(wire_d48_87),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904888(.data_in(wire_d48_87),.data_out(wire_d48_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4904889(.data_in(wire_d48_88),.data_out(wire_d48_89),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904890(.data_in(wire_d48_89),.data_out(wire_d48_90),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904891(.data_in(wire_d48_90),.data_out(wire_d48_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4904892(.data_in(wire_d48_91),.data_out(wire_d48_92),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904893(.data_in(wire_d48_92),.data_out(wire_d48_93),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4904894(.data_in(wire_d48_93),.data_out(wire_d48_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904895(.data_in(wire_d48_94),.data_out(wire_d48_95),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904896(.data_in(wire_d48_95),.data_out(wire_d48_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4904897(.data_in(wire_d48_96),.data_out(wire_d48_97),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904898(.data_in(wire_d48_97),.data_out(wire_d48_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4904899(.data_in(wire_d48_98),.data_out(wire_d48_99),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance49048100(.data_in(wire_d48_99),.data_out(wire_d48_100),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance49048101(.data_in(wire_d48_100),.data_out(wire_d48_101),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance49048102(.data_in(wire_d48_101),.data_out(wire_d48_102),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance49048103(.data_in(wire_d48_102),.data_out(wire_d48_103),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance49048104(.data_in(wire_d48_103),.data_out(wire_d48_104),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance49048105(.data_in(wire_d48_104),.data_out(wire_d48_105),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance49048106(.data_in(wire_d48_105),.data_out(wire_d48_106),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance49048107(.data_in(wire_d48_106),.data_out(wire_d48_107),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance49048108(.data_in(wire_d48_107),.data_out(wire_d48_108),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance49048109(.data_in(wire_d48_108),.data_out(wire_d48_109),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance49048110(.data_in(wire_d48_109),.data_out(wire_d48_110),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance49048111(.data_in(wire_d48_110),.data_out(wire_d48_111),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance49048112(.data_in(wire_d48_111),.data_out(wire_d48_112),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance49048113(.data_in(wire_d48_112),.data_out(wire_d48_113),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance49048114(.data_in(wire_d48_113),.data_out(wire_d48_114),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance49048115(.data_in(wire_d48_114),.data_out(wire_d48_115),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance49048116(.data_in(wire_d48_115),.data_out(wire_d48_116),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance49048117(.data_in(wire_d48_116),.data_out(wire_d48_117),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance49048118(.data_in(wire_d48_117),.data_out(wire_d48_118),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance49048119(.data_in(wire_d48_118),.data_out(d_out48),.clk(clk),.rst(rst));

	large_adder #(.WIDTH(WIDTH)) large_adder_instance500490(.data_in(d_in49),.data_out(wire_d49_0),.clk(clk),.rst(rst));            //channel 50
	large_mux #(.WIDTH(WIDTH)) large_mux_instance500491(.data_in(wire_d49_0),.data_out(wire_d49_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance500492(.data_in(wire_d49_1),.data_out(wire_d49_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance500493(.data_in(wire_d49_2),.data_out(wire_d49_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance500494(.data_in(wire_d49_3),.data_out(wire_d49_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance500495(.data_in(wire_d49_4),.data_out(wire_d49_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance500496(.data_in(wire_d49_5),.data_out(wire_d49_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance500497(.data_in(wire_d49_6),.data_out(wire_d49_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance500498(.data_in(wire_d49_7),.data_out(wire_d49_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance500499(.data_in(wire_d49_8),.data_out(wire_d49_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5004910(.data_in(wire_d49_9),.data_out(wire_d49_10),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5004911(.data_in(wire_d49_10),.data_out(wire_d49_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004912(.data_in(wire_d49_11),.data_out(wire_d49_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004913(.data_in(wire_d49_12),.data_out(wire_d49_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004914(.data_in(wire_d49_13),.data_out(wire_d49_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004915(.data_in(wire_d49_14),.data_out(wire_d49_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004916(.data_in(wire_d49_15),.data_out(wire_d49_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004917(.data_in(wire_d49_16),.data_out(wire_d49_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004918(.data_in(wire_d49_17),.data_out(wire_d49_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5004919(.data_in(wire_d49_18),.data_out(wire_d49_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004920(.data_in(wire_d49_19),.data_out(wire_d49_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5004921(.data_in(wire_d49_20),.data_out(wire_d49_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004922(.data_in(wire_d49_21),.data_out(wire_d49_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004923(.data_in(wire_d49_22),.data_out(wire_d49_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5004924(.data_in(wire_d49_23),.data_out(wire_d49_24),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004925(.data_in(wire_d49_24),.data_out(wire_d49_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004926(.data_in(wire_d49_25),.data_out(wire_d49_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004927(.data_in(wire_d49_26),.data_out(wire_d49_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004928(.data_in(wire_d49_27),.data_out(wire_d49_28),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5004929(.data_in(wire_d49_28),.data_out(wire_d49_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5004930(.data_in(wire_d49_29),.data_out(wire_d49_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004931(.data_in(wire_d49_30),.data_out(wire_d49_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004932(.data_in(wire_d49_31),.data_out(wire_d49_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5004933(.data_in(wire_d49_32),.data_out(wire_d49_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004934(.data_in(wire_d49_33),.data_out(wire_d49_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004935(.data_in(wire_d49_34),.data_out(wire_d49_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004936(.data_in(wire_d49_35),.data_out(wire_d49_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5004937(.data_in(wire_d49_36),.data_out(wire_d49_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004938(.data_in(wire_d49_37),.data_out(wire_d49_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004939(.data_in(wire_d49_38),.data_out(wire_d49_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004940(.data_in(wire_d49_39),.data_out(wire_d49_40),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5004941(.data_in(wire_d49_40),.data_out(wire_d49_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5004942(.data_in(wire_d49_41),.data_out(wire_d49_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004943(.data_in(wire_d49_42),.data_out(wire_d49_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004944(.data_in(wire_d49_43),.data_out(wire_d49_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004945(.data_in(wire_d49_44),.data_out(wire_d49_45),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5004946(.data_in(wire_d49_45),.data_out(wire_d49_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004947(.data_in(wire_d49_46),.data_out(wire_d49_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5004948(.data_in(wire_d49_47),.data_out(wire_d49_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5004949(.data_in(wire_d49_48),.data_out(wire_d49_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004950(.data_in(wire_d49_49),.data_out(wire_d49_50),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5004951(.data_in(wire_d49_50),.data_out(wire_d49_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004952(.data_in(wire_d49_51),.data_out(wire_d49_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004953(.data_in(wire_d49_52),.data_out(wire_d49_53),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004954(.data_in(wire_d49_53),.data_out(wire_d49_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004955(.data_in(wire_d49_54),.data_out(wire_d49_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004956(.data_in(wire_d49_55),.data_out(wire_d49_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5004957(.data_in(wire_d49_56),.data_out(wire_d49_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5004958(.data_in(wire_d49_57),.data_out(wire_d49_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5004959(.data_in(wire_d49_58),.data_out(wire_d49_59),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5004960(.data_in(wire_d49_59),.data_out(wire_d49_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004961(.data_in(wire_d49_60),.data_out(wire_d49_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004962(.data_in(wire_d49_61),.data_out(wire_d49_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004963(.data_in(wire_d49_62),.data_out(wire_d49_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5004964(.data_in(wire_d49_63),.data_out(wire_d49_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004965(.data_in(wire_d49_64),.data_out(wire_d49_65),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5004966(.data_in(wire_d49_65),.data_out(wire_d49_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004967(.data_in(wire_d49_66),.data_out(wire_d49_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5004968(.data_in(wire_d49_67),.data_out(wire_d49_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004969(.data_in(wire_d49_68),.data_out(wire_d49_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5004970(.data_in(wire_d49_69),.data_out(wire_d49_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004971(.data_in(wire_d49_70),.data_out(wire_d49_71),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004972(.data_in(wire_d49_71),.data_out(wire_d49_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004973(.data_in(wire_d49_72),.data_out(wire_d49_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004974(.data_in(wire_d49_73),.data_out(wire_d49_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004975(.data_in(wire_d49_74),.data_out(wire_d49_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004976(.data_in(wire_d49_75),.data_out(wire_d49_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004977(.data_in(wire_d49_76),.data_out(wire_d49_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004978(.data_in(wire_d49_77),.data_out(wire_d49_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004979(.data_in(wire_d49_78),.data_out(wire_d49_79),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004980(.data_in(wire_d49_79),.data_out(wire_d49_80),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004981(.data_in(wire_d49_80),.data_out(wire_d49_81),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004982(.data_in(wire_d49_81),.data_out(wire_d49_82),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004983(.data_in(wire_d49_82),.data_out(wire_d49_83),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5004984(.data_in(wire_d49_83),.data_out(wire_d49_84),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004985(.data_in(wire_d49_84),.data_out(wire_d49_85),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004986(.data_in(wire_d49_85),.data_out(wire_d49_86),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004987(.data_in(wire_d49_86),.data_out(wire_d49_87),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004988(.data_in(wire_d49_87),.data_out(wire_d49_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004989(.data_in(wire_d49_88),.data_out(wire_d49_89),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004990(.data_in(wire_d49_89),.data_out(wire_d49_90),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5004991(.data_in(wire_d49_90),.data_out(wire_d49_91),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004992(.data_in(wire_d49_91),.data_out(wire_d49_92),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5004993(.data_in(wire_d49_92),.data_out(wire_d49_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5004994(.data_in(wire_d49_93),.data_out(wire_d49_94),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5004995(.data_in(wire_d49_94),.data_out(wire_d49_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5004996(.data_in(wire_d49_95),.data_out(wire_d49_96),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004997(.data_in(wire_d49_96),.data_out(wire_d49_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5004998(.data_in(wire_d49_97),.data_out(wire_d49_98),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004999(.data_in(wire_d49_98),.data_out(wire_d49_99),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance50049100(.data_in(wire_d49_99),.data_out(wire_d49_100),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance50049101(.data_in(wire_d49_100),.data_out(wire_d49_101),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance50049102(.data_in(wire_d49_101),.data_out(wire_d49_102),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance50049103(.data_in(wire_d49_102),.data_out(wire_d49_103),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance50049104(.data_in(wire_d49_103),.data_out(wire_d49_104),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance50049105(.data_in(wire_d49_104),.data_out(wire_d49_105),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance50049106(.data_in(wire_d49_105),.data_out(wire_d49_106),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance50049107(.data_in(wire_d49_106),.data_out(wire_d49_107),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance50049108(.data_in(wire_d49_107),.data_out(wire_d49_108),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance50049109(.data_in(wire_d49_108),.data_out(wire_d49_109),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance50049110(.data_in(wire_d49_109),.data_out(wire_d49_110),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance50049111(.data_in(wire_d49_110),.data_out(wire_d49_111),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance50049112(.data_in(wire_d49_111),.data_out(wire_d49_112),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance50049113(.data_in(wire_d49_112),.data_out(wire_d49_113),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance50049114(.data_in(wire_d49_113),.data_out(wire_d49_114),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance50049115(.data_in(wire_d49_114),.data_out(wire_d49_115),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance50049116(.data_in(wire_d49_115),.data_out(wire_d49_116),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance50049117(.data_in(wire_d49_116),.data_out(wire_d49_117),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance50049118(.data_in(wire_d49_117),.data_out(wire_d49_118),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance50049119(.data_in(wire_d49_118),.data_out(d_out49),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance510500(.data_in(d_in50),.data_out(wire_d50_0),.clk(clk),.rst(rst));            //channel 51
	encoder #(.WIDTH(WIDTH)) encoder_instance510501(.data_in(wire_d50_0),.data_out(wire_d50_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance510502(.data_in(wire_d50_1),.data_out(wire_d50_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance510503(.data_in(wire_d50_2),.data_out(wire_d50_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance510504(.data_in(wire_d50_3),.data_out(wire_d50_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance510505(.data_in(wire_d50_4),.data_out(wire_d50_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance510506(.data_in(wire_d50_5),.data_out(wire_d50_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance510507(.data_in(wire_d50_6),.data_out(wire_d50_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance510508(.data_in(wire_d50_7),.data_out(wire_d50_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance510509(.data_in(wire_d50_8),.data_out(wire_d50_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5105010(.data_in(wire_d50_9),.data_out(wire_d50_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5105011(.data_in(wire_d50_10),.data_out(wire_d50_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5105012(.data_in(wire_d50_11),.data_out(wire_d50_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5105013(.data_in(wire_d50_12),.data_out(wire_d50_13),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5105014(.data_in(wire_d50_13),.data_out(wire_d50_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5105015(.data_in(wire_d50_14),.data_out(wire_d50_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5105016(.data_in(wire_d50_15),.data_out(wire_d50_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105017(.data_in(wire_d50_16),.data_out(wire_d50_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5105018(.data_in(wire_d50_17),.data_out(wire_d50_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5105019(.data_in(wire_d50_18),.data_out(wire_d50_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105020(.data_in(wire_d50_19),.data_out(wire_d50_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105021(.data_in(wire_d50_20),.data_out(wire_d50_21),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105022(.data_in(wire_d50_21),.data_out(wire_d50_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5105023(.data_in(wire_d50_22),.data_out(wire_d50_23),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5105024(.data_in(wire_d50_23),.data_out(wire_d50_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105025(.data_in(wire_d50_24),.data_out(wire_d50_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5105026(.data_in(wire_d50_25),.data_out(wire_d50_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105027(.data_in(wire_d50_26),.data_out(wire_d50_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5105028(.data_in(wire_d50_27),.data_out(wire_d50_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5105029(.data_in(wire_d50_28),.data_out(wire_d50_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5105030(.data_in(wire_d50_29),.data_out(wire_d50_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5105031(.data_in(wire_d50_30),.data_out(wire_d50_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5105032(.data_in(wire_d50_31),.data_out(wire_d50_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105033(.data_in(wire_d50_32),.data_out(wire_d50_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105034(.data_in(wire_d50_33),.data_out(wire_d50_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105035(.data_in(wire_d50_34),.data_out(wire_d50_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105036(.data_in(wire_d50_35),.data_out(wire_d50_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105037(.data_in(wire_d50_36),.data_out(wire_d50_37),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105038(.data_in(wire_d50_37),.data_out(wire_d50_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5105039(.data_in(wire_d50_38),.data_out(wire_d50_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5105040(.data_in(wire_d50_39),.data_out(wire_d50_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5105041(.data_in(wire_d50_40),.data_out(wire_d50_41),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5105042(.data_in(wire_d50_41),.data_out(wire_d50_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5105043(.data_in(wire_d50_42),.data_out(wire_d50_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105044(.data_in(wire_d50_43),.data_out(wire_d50_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5105045(.data_in(wire_d50_44),.data_out(wire_d50_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5105046(.data_in(wire_d50_45),.data_out(wire_d50_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105047(.data_in(wire_d50_46),.data_out(wire_d50_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105048(.data_in(wire_d50_47),.data_out(wire_d50_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5105049(.data_in(wire_d50_48),.data_out(wire_d50_49),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5105050(.data_in(wire_d50_49),.data_out(wire_d50_50),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5105051(.data_in(wire_d50_50),.data_out(wire_d50_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5105052(.data_in(wire_d50_51),.data_out(wire_d50_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5105053(.data_in(wire_d50_52),.data_out(wire_d50_53),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105054(.data_in(wire_d50_53),.data_out(wire_d50_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105055(.data_in(wire_d50_54),.data_out(wire_d50_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105056(.data_in(wire_d50_55),.data_out(wire_d50_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5105057(.data_in(wire_d50_56),.data_out(wire_d50_57),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5105058(.data_in(wire_d50_57),.data_out(wire_d50_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5105059(.data_in(wire_d50_58),.data_out(wire_d50_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5105060(.data_in(wire_d50_59),.data_out(wire_d50_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5105061(.data_in(wire_d50_60),.data_out(wire_d50_61),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5105062(.data_in(wire_d50_61),.data_out(wire_d50_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5105063(.data_in(wire_d50_62),.data_out(wire_d50_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105064(.data_in(wire_d50_63),.data_out(wire_d50_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5105065(.data_in(wire_d50_64),.data_out(wire_d50_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105066(.data_in(wire_d50_65),.data_out(wire_d50_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5105067(.data_in(wire_d50_66),.data_out(wire_d50_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105068(.data_in(wire_d50_67),.data_out(wire_d50_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105069(.data_in(wire_d50_68),.data_out(wire_d50_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5105070(.data_in(wire_d50_69),.data_out(wire_d50_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5105071(.data_in(wire_d50_70),.data_out(wire_d50_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5105072(.data_in(wire_d50_71),.data_out(wire_d50_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105073(.data_in(wire_d50_72),.data_out(wire_d50_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105074(.data_in(wire_d50_73),.data_out(wire_d50_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105075(.data_in(wire_d50_74),.data_out(wire_d50_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105076(.data_in(wire_d50_75),.data_out(wire_d50_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5105077(.data_in(wire_d50_76),.data_out(wire_d50_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105078(.data_in(wire_d50_77),.data_out(wire_d50_78),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105079(.data_in(wire_d50_78),.data_out(wire_d50_79),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105080(.data_in(wire_d50_79),.data_out(wire_d50_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105081(.data_in(wire_d50_80),.data_out(wire_d50_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5105082(.data_in(wire_d50_81),.data_out(wire_d50_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105083(.data_in(wire_d50_82),.data_out(wire_d50_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105084(.data_in(wire_d50_83),.data_out(wire_d50_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5105085(.data_in(wire_d50_84),.data_out(wire_d50_85),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5105086(.data_in(wire_d50_85),.data_out(wire_d50_86),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5105087(.data_in(wire_d50_86),.data_out(wire_d50_87),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5105088(.data_in(wire_d50_87),.data_out(wire_d50_88),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105089(.data_in(wire_d50_88),.data_out(wire_d50_89),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105090(.data_in(wire_d50_89),.data_out(wire_d50_90),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105091(.data_in(wire_d50_90),.data_out(wire_d50_91),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105092(.data_in(wire_d50_91),.data_out(wire_d50_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105093(.data_in(wire_d50_92),.data_out(wire_d50_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5105094(.data_in(wire_d50_93),.data_out(wire_d50_94),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5105095(.data_in(wire_d50_94),.data_out(wire_d50_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5105096(.data_in(wire_d50_95),.data_out(wire_d50_96),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105097(.data_in(wire_d50_96),.data_out(wire_d50_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105098(.data_in(wire_d50_97),.data_out(wire_d50_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5105099(.data_in(wire_d50_98),.data_out(wire_d50_99),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance51050100(.data_in(wire_d50_99),.data_out(wire_d50_100),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance51050101(.data_in(wire_d50_100),.data_out(wire_d50_101),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance51050102(.data_in(wire_d50_101),.data_out(wire_d50_102),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance51050103(.data_in(wire_d50_102),.data_out(wire_d50_103),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance51050104(.data_in(wire_d50_103),.data_out(wire_d50_104),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance51050105(.data_in(wire_d50_104),.data_out(wire_d50_105),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance51050106(.data_in(wire_d50_105),.data_out(wire_d50_106),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance51050107(.data_in(wire_d50_106),.data_out(wire_d50_107),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance51050108(.data_in(wire_d50_107),.data_out(wire_d50_108),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance51050109(.data_in(wire_d50_108),.data_out(wire_d50_109),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance51050110(.data_in(wire_d50_109),.data_out(wire_d50_110),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance51050111(.data_in(wire_d50_110),.data_out(wire_d50_111),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance51050112(.data_in(wire_d50_111),.data_out(wire_d50_112),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance51050113(.data_in(wire_d50_112),.data_out(wire_d50_113),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance51050114(.data_in(wire_d50_113),.data_out(wire_d50_114),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance51050115(.data_in(wire_d50_114),.data_out(wire_d50_115),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance51050116(.data_in(wire_d50_115),.data_out(wire_d50_116),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance51050117(.data_in(wire_d50_116),.data_out(wire_d50_117),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance51050118(.data_in(wire_d50_117),.data_out(wire_d50_118),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance51050119(.data_in(wire_d50_118),.data_out(d_out50),.clk(clk),.rst(rst));

	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance520510(.data_in(d_in51),.data_out(wire_d51_0),.clk(clk),.rst(rst));            //channel 52
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance520511(.data_in(wire_d51_0),.data_out(wire_d51_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance520512(.data_in(wire_d51_1),.data_out(wire_d51_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance520513(.data_in(wire_d51_2),.data_out(wire_d51_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance520514(.data_in(wire_d51_3),.data_out(wire_d51_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance520515(.data_in(wire_d51_4),.data_out(wire_d51_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance520516(.data_in(wire_d51_5),.data_out(wire_d51_6),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance520517(.data_in(wire_d51_6),.data_out(wire_d51_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance520518(.data_in(wire_d51_7),.data_out(wire_d51_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance520519(.data_in(wire_d51_8),.data_out(wire_d51_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205110(.data_in(wire_d51_9),.data_out(wire_d51_10),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5205111(.data_in(wire_d51_10),.data_out(wire_d51_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205112(.data_in(wire_d51_11),.data_out(wire_d51_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205113(.data_in(wire_d51_12),.data_out(wire_d51_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205114(.data_in(wire_d51_13),.data_out(wire_d51_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205115(.data_in(wire_d51_14),.data_out(wire_d51_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205116(.data_in(wire_d51_15),.data_out(wire_d51_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205117(.data_in(wire_d51_16),.data_out(wire_d51_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5205118(.data_in(wire_d51_17),.data_out(wire_d51_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205119(.data_in(wire_d51_18),.data_out(wire_d51_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205120(.data_in(wire_d51_19),.data_out(wire_d51_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205121(.data_in(wire_d51_20),.data_out(wire_d51_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205122(.data_in(wire_d51_21),.data_out(wire_d51_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5205123(.data_in(wire_d51_22),.data_out(wire_d51_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205124(.data_in(wire_d51_23),.data_out(wire_d51_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5205125(.data_in(wire_d51_24),.data_out(wire_d51_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5205126(.data_in(wire_d51_25),.data_out(wire_d51_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205127(.data_in(wire_d51_26),.data_out(wire_d51_27),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5205128(.data_in(wire_d51_27),.data_out(wire_d51_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205129(.data_in(wire_d51_28),.data_out(wire_d51_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5205130(.data_in(wire_d51_29),.data_out(wire_d51_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205131(.data_in(wire_d51_30),.data_out(wire_d51_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205132(.data_in(wire_d51_31),.data_out(wire_d51_32),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205133(.data_in(wire_d51_32),.data_out(wire_d51_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5205134(.data_in(wire_d51_33),.data_out(wire_d51_34),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205135(.data_in(wire_d51_34),.data_out(wire_d51_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205136(.data_in(wire_d51_35),.data_out(wire_d51_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205137(.data_in(wire_d51_36),.data_out(wire_d51_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5205138(.data_in(wire_d51_37),.data_out(wire_d51_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5205139(.data_in(wire_d51_38),.data_out(wire_d51_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5205140(.data_in(wire_d51_39),.data_out(wire_d51_40),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5205141(.data_in(wire_d51_40),.data_out(wire_d51_41),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5205142(.data_in(wire_d51_41),.data_out(wire_d51_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5205143(.data_in(wire_d51_42),.data_out(wire_d51_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205144(.data_in(wire_d51_43),.data_out(wire_d51_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205145(.data_in(wire_d51_44),.data_out(wire_d51_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5205146(.data_in(wire_d51_45),.data_out(wire_d51_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5205147(.data_in(wire_d51_46),.data_out(wire_d51_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5205148(.data_in(wire_d51_47),.data_out(wire_d51_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205149(.data_in(wire_d51_48),.data_out(wire_d51_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5205150(.data_in(wire_d51_49),.data_out(wire_d51_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5205151(.data_in(wire_d51_50),.data_out(wire_d51_51),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5205152(.data_in(wire_d51_51),.data_out(wire_d51_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205153(.data_in(wire_d51_52),.data_out(wire_d51_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5205154(.data_in(wire_d51_53),.data_out(wire_d51_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5205155(.data_in(wire_d51_54),.data_out(wire_d51_55),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5205156(.data_in(wire_d51_55),.data_out(wire_d51_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5205157(.data_in(wire_d51_56),.data_out(wire_d51_57),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5205158(.data_in(wire_d51_57),.data_out(wire_d51_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205159(.data_in(wire_d51_58),.data_out(wire_d51_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5205160(.data_in(wire_d51_59),.data_out(wire_d51_60),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205161(.data_in(wire_d51_60),.data_out(wire_d51_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205162(.data_in(wire_d51_61),.data_out(wire_d51_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205163(.data_in(wire_d51_62),.data_out(wire_d51_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5205164(.data_in(wire_d51_63),.data_out(wire_d51_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205165(.data_in(wire_d51_64),.data_out(wire_d51_65),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205166(.data_in(wire_d51_65),.data_out(wire_d51_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205167(.data_in(wire_d51_66),.data_out(wire_d51_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5205168(.data_in(wire_d51_67),.data_out(wire_d51_68),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205169(.data_in(wire_d51_68),.data_out(wire_d51_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205170(.data_in(wire_d51_69),.data_out(wire_d51_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5205171(.data_in(wire_d51_70),.data_out(wire_d51_71),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5205172(.data_in(wire_d51_71),.data_out(wire_d51_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205173(.data_in(wire_d51_72),.data_out(wire_d51_73),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5205174(.data_in(wire_d51_73),.data_out(wire_d51_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5205175(.data_in(wire_d51_74),.data_out(wire_d51_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205176(.data_in(wire_d51_75),.data_out(wire_d51_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5205177(.data_in(wire_d51_76),.data_out(wire_d51_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205178(.data_in(wire_d51_77),.data_out(wire_d51_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205179(.data_in(wire_d51_78),.data_out(wire_d51_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5205180(.data_in(wire_d51_79),.data_out(wire_d51_80),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205181(.data_in(wire_d51_80),.data_out(wire_d51_81),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205182(.data_in(wire_d51_81),.data_out(wire_d51_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5205183(.data_in(wire_d51_82),.data_out(wire_d51_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205184(.data_in(wire_d51_83),.data_out(wire_d51_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5205185(.data_in(wire_d51_84),.data_out(wire_d51_85),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205186(.data_in(wire_d51_85),.data_out(wire_d51_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5205187(.data_in(wire_d51_86),.data_out(wire_d51_87),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205188(.data_in(wire_d51_87),.data_out(wire_d51_88),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205189(.data_in(wire_d51_88),.data_out(wire_d51_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205190(.data_in(wire_d51_89),.data_out(wire_d51_90),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205191(.data_in(wire_d51_90),.data_out(wire_d51_91),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205192(.data_in(wire_d51_91),.data_out(wire_d51_92),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205193(.data_in(wire_d51_92),.data_out(wire_d51_93),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5205194(.data_in(wire_d51_93),.data_out(wire_d51_94),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205195(.data_in(wire_d51_94),.data_out(wire_d51_95),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205196(.data_in(wire_d51_95),.data_out(wire_d51_96),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205197(.data_in(wire_d51_96),.data_out(wire_d51_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5205198(.data_in(wire_d51_97),.data_out(wire_d51_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5205199(.data_in(wire_d51_98),.data_out(wire_d51_99),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance52051100(.data_in(wire_d51_99),.data_out(wire_d51_100),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance52051101(.data_in(wire_d51_100),.data_out(wire_d51_101),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance52051102(.data_in(wire_d51_101),.data_out(wire_d51_102),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance52051103(.data_in(wire_d51_102),.data_out(wire_d51_103),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance52051104(.data_in(wire_d51_103),.data_out(wire_d51_104),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance52051105(.data_in(wire_d51_104),.data_out(wire_d51_105),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance52051106(.data_in(wire_d51_105),.data_out(wire_d51_106),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance52051107(.data_in(wire_d51_106),.data_out(wire_d51_107),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance52051108(.data_in(wire_d51_107),.data_out(wire_d51_108),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance52051109(.data_in(wire_d51_108),.data_out(wire_d51_109),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance52051110(.data_in(wire_d51_109),.data_out(wire_d51_110),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance52051111(.data_in(wire_d51_110),.data_out(wire_d51_111),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance52051112(.data_in(wire_d51_111),.data_out(wire_d51_112),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance52051113(.data_in(wire_d51_112),.data_out(wire_d51_113),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance52051114(.data_in(wire_d51_113),.data_out(wire_d51_114),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance52051115(.data_in(wire_d51_114),.data_out(wire_d51_115),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance52051116(.data_in(wire_d51_115),.data_out(wire_d51_116),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance52051117(.data_in(wire_d51_116),.data_out(wire_d51_117),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance52051118(.data_in(wire_d51_117),.data_out(wire_d51_118),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance52051119(.data_in(wire_d51_118),.data_out(d_out51),.clk(clk),.rst(rst));

	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance530520(.data_in(d_in52),.data_out(wire_d52_0),.clk(clk),.rst(rst));            //channel 53
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance530521(.data_in(wire_d52_0),.data_out(wire_d52_1),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance530522(.data_in(wire_d52_1),.data_out(wire_d52_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance530523(.data_in(wire_d52_2),.data_out(wire_d52_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance530524(.data_in(wire_d52_3),.data_out(wire_d52_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance530525(.data_in(wire_d52_4),.data_out(wire_d52_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance530526(.data_in(wire_d52_5),.data_out(wire_d52_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance530527(.data_in(wire_d52_6),.data_out(wire_d52_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance530528(.data_in(wire_d52_7),.data_out(wire_d52_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance530529(.data_in(wire_d52_8),.data_out(wire_d52_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5305210(.data_in(wire_d52_9),.data_out(wire_d52_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305211(.data_in(wire_d52_10),.data_out(wire_d52_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5305212(.data_in(wire_d52_11),.data_out(wire_d52_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305213(.data_in(wire_d52_12),.data_out(wire_d52_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5305214(.data_in(wire_d52_13),.data_out(wire_d52_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5305215(.data_in(wire_d52_14),.data_out(wire_d52_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5305216(.data_in(wire_d52_15),.data_out(wire_d52_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305217(.data_in(wire_d52_16),.data_out(wire_d52_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305218(.data_in(wire_d52_17),.data_out(wire_d52_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305219(.data_in(wire_d52_18),.data_out(wire_d52_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305220(.data_in(wire_d52_19),.data_out(wire_d52_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305221(.data_in(wire_d52_20),.data_out(wire_d52_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305222(.data_in(wire_d52_21),.data_out(wire_d52_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305223(.data_in(wire_d52_22),.data_out(wire_d52_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5305224(.data_in(wire_d52_23),.data_out(wire_d52_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305225(.data_in(wire_d52_24),.data_out(wire_d52_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5305226(.data_in(wire_d52_25),.data_out(wire_d52_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5305227(.data_in(wire_d52_26),.data_out(wire_d52_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305228(.data_in(wire_d52_27),.data_out(wire_d52_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5305229(.data_in(wire_d52_28),.data_out(wire_d52_29),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5305230(.data_in(wire_d52_29),.data_out(wire_d52_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305231(.data_in(wire_d52_30),.data_out(wire_d52_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305232(.data_in(wire_d52_31),.data_out(wire_d52_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5305233(.data_in(wire_d52_32),.data_out(wire_d52_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305234(.data_in(wire_d52_33),.data_out(wire_d52_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305235(.data_in(wire_d52_34),.data_out(wire_d52_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5305236(.data_in(wire_d52_35),.data_out(wire_d52_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305237(.data_in(wire_d52_36),.data_out(wire_d52_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5305238(.data_in(wire_d52_37),.data_out(wire_d52_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5305239(.data_in(wire_d52_38),.data_out(wire_d52_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5305240(.data_in(wire_d52_39),.data_out(wire_d52_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305241(.data_in(wire_d52_40),.data_out(wire_d52_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305242(.data_in(wire_d52_41),.data_out(wire_d52_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305243(.data_in(wire_d52_42),.data_out(wire_d52_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305244(.data_in(wire_d52_43),.data_out(wire_d52_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5305245(.data_in(wire_d52_44),.data_out(wire_d52_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305246(.data_in(wire_d52_45),.data_out(wire_d52_46),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305247(.data_in(wire_d52_46),.data_out(wire_d52_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5305248(.data_in(wire_d52_47),.data_out(wire_d52_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305249(.data_in(wire_d52_48),.data_out(wire_d52_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305250(.data_in(wire_d52_49),.data_out(wire_d52_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5305251(.data_in(wire_d52_50),.data_out(wire_d52_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5305252(.data_in(wire_d52_51),.data_out(wire_d52_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305253(.data_in(wire_d52_52),.data_out(wire_d52_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305254(.data_in(wire_d52_53),.data_out(wire_d52_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305255(.data_in(wire_d52_54),.data_out(wire_d52_55),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305256(.data_in(wire_d52_55),.data_out(wire_d52_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305257(.data_in(wire_d52_56),.data_out(wire_d52_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5305258(.data_in(wire_d52_57),.data_out(wire_d52_58),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305259(.data_in(wire_d52_58),.data_out(wire_d52_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305260(.data_in(wire_d52_59),.data_out(wire_d52_60),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305261(.data_in(wire_d52_60),.data_out(wire_d52_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305262(.data_in(wire_d52_61),.data_out(wire_d52_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5305263(.data_in(wire_d52_62),.data_out(wire_d52_63),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5305264(.data_in(wire_d52_63),.data_out(wire_d52_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305265(.data_in(wire_d52_64),.data_out(wire_d52_65),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305266(.data_in(wire_d52_65),.data_out(wire_d52_66),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305267(.data_in(wire_d52_66),.data_out(wire_d52_67),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5305268(.data_in(wire_d52_67),.data_out(wire_d52_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305269(.data_in(wire_d52_68),.data_out(wire_d52_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305270(.data_in(wire_d52_69),.data_out(wire_d52_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5305271(.data_in(wire_d52_70),.data_out(wire_d52_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305272(.data_in(wire_d52_71),.data_out(wire_d52_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305273(.data_in(wire_d52_72),.data_out(wire_d52_73),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305274(.data_in(wire_d52_73),.data_out(wire_d52_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305275(.data_in(wire_d52_74),.data_out(wire_d52_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305276(.data_in(wire_d52_75),.data_out(wire_d52_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5305277(.data_in(wire_d52_76),.data_out(wire_d52_77),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305278(.data_in(wire_d52_77),.data_out(wire_d52_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305279(.data_in(wire_d52_78),.data_out(wire_d52_79),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305280(.data_in(wire_d52_79),.data_out(wire_d52_80),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305281(.data_in(wire_d52_80),.data_out(wire_d52_81),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305282(.data_in(wire_d52_81),.data_out(wire_d52_82),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305283(.data_in(wire_d52_82),.data_out(wire_d52_83),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5305284(.data_in(wire_d52_83),.data_out(wire_d52_84),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5305285(.data_in(wire_d52_84),.data_out(wire_d52_85),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305286(.data_in(wire_d52_85),.data_out(wire_d52_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5305287(.data_in(wire_d52_86),.data_out(wire_d52_87),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5305288(.data_in(wire_d52_87),.data_out(wire_d52_88),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305289(.data_in(wire_d52_88),.data_out(wire_d52_89),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305290(.data_in(wire_d52_89),.data_out(wire_d52_90),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305291(.data_in(wire_d52_90),.data_out(wire_d52_91),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305292(.data_in(wire_d52_91),.data_out(wire_d52_92),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305293(.data_in(wire_d52_92),.data_out(wire_d52_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5305294(.data_in(wire_d52_93),.data_out(wire_d52_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5305295(.data_in(wire_d52_94),.data_out(wire_d52_95),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305296(.data_in(wire_d52_95),.data_out(wire_d52_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305297(.data_in(wire_d52_96),.data_out(wire_d52_97),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305298(.data_in(wire_d52_97),.data_out(wire_d52_98),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305299(.data_in(wire_d52_98),.data_out(wire_d52_99),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance53052100(.data_in(wire_d52_99),.data_out(wire_d52_100),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance53052101(.data_in(wire_d52_100),.data_out(wire_d52_101),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance53052102(.data_in(wire_d52_101),.data_out(wire_d52_102),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance53052103(.data_in(wire_d52_102),.data_out(wire_d52_103),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance53052104(.data_in(wire_d52_103),.data_out(wire_d52_104),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance53052105(.data_in(wire_d52_104),.data_out(wire_d52_105),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance53052106(.data_in(wire_d52_105),.data_out(wire_d52_106),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance53052107(.data_in(wire_d52_106),.data_out(wire_d52_107),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance53052108(.data_in(wire_d52_107),.data_out(wire_d52_108),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance53052109(.data_in(wire_d52_108),.data_out(wire_d52_109),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance53052110(.data_in(wire_d52_109),.data_out(wire_d52_110),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance53052111(.data_in(wire_d52_110),.data_out(wire_d52_111),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance53052112(.data_in(wire_d52_111),.data_out(wire_d52_112),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance53052113(.data_in(wire_d52_112),.data_out(wire_d52_113),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance53052114(.data_in(wire_d52_113),.data_out(wire_d52_114),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance53052115(.data_in(wire_d52_114),.data_out(wire_d52_115),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance53052116(.data_in(wire_d52_115),.data_out(wire_d52_116),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance53052117(.data_in(wire_d52_116),.data_out(wire_d52_117),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance53052118(.data_in(wire_d52_117),.data_out(wire_d52_118),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance53052119(.data_in(wire_d52_118),.data_out(d_out52),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance540530(.data_in(d_in53),.data_out(wire_d53_0),.clk(clk),.rst(rst));            //channel 54
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance540531(.data_in(wire_d53_0),.data_out(wire_d53_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance540532(.data_in(wire_d53_1),.data_out(wire_d53_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance540533(.data_in(wire_d53_2),.data_out(wire_d53_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance540534(.data_in(wire_d53_3),.data_out(wire_d53_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance540535(.data_in(wire_d53_4),.data_out(wire_d53_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance540536(.data_in(wire_d53_5),.data_out(wire_d53_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance540537(.data_in(wire_d53_6),.data_out(wire_d53_7),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance540538(.data_in(wire_d53_7),.data_out(wire_d53_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance540539(.data_in(wire_d53_8),.data_out(wire_d53_9),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405310(.data_in(wire_d53_9),.data_out(wire_d53_10),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5405311(.data_in(wire_d53_10),.data_out(wire_d53_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5405312(.data_in(wire_d53_11),.data_out(wire_d53_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405313(.data_in(wire_d53_12),.data_out(wire_d53_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405314(.data_in(wire_d53_13),.data_out(wire_d53_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405315(.data_in(wire_d53_14),.data_out(wire_d53_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405316(.data_in(wire_d53_15),.data_out(wire_d53_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405317(.data_in(wire_d53_16),.data_out(wire_d53_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405318(.data_in(wire_d53_17),.data_out(wire_d53_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405319(.data_in(wire_d53_18),.data_out(wire_d53_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5405320(.data_in(wire_d53_19),.data_out(wire_d53_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405321(.data_in(wire_d53_20),.data_out(wire_d53_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405322(.data_in(wire_d53_21),.data_out(wire_d53_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405323(.data_in(wire_d53_22),.data_out(wire_d53_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5405324(.data_in(wire_d53_23),.data_out(wire_d53_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5405325(.data_in(wire_d53_24),.data_out(wire_d53_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5405326(.data_in(wire_d53_25),.data_out(wire_d53_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405327(.data_in(wire_d53_26),.data_out(wire_d53_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405328(.data_in(wire_d53_27),.data_out(wire_d53_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405329(.data_in(wire_d53_28),.data_out(wire_d53_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405330(.data_in(wire_d53_29),.data_out(wire_d53_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405331(.data_in(wire_d53_30),.data_out(wire_d53_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405332(.data_in(wire_d53_31),.data_out(wire_d53_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5405333(.data_in(wire_d53_32),.data_out(wire_d53_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405334(.data_in(wire_d53_33),.data_out(wire_d53_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5405335(.data_in(wire_d53_34),.data_out(wire_d53_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405336(.data_in(wire_d53_35),.data_out(wire_d53_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5405337(.data_in(wire_d53_36),.data_out(wire_d53_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405338(.data_in(wire_d53_37),.data_out(wire_d53_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405339(.data_in(wire_d53_38),.data_out(wire_d53_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405340(.data_in(wire_d53_39),.data_out(wire_d53_40),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5405341(.data_in(wire_d53_40),.data_out(wire_d53_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5405342(.data_in(wire_d53_41),.data_out(wire_d53_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5405343(.data_in(wire_d53_42),.data_out(wire_d53_43),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5405344(.data_in(wire_d53_43),.data_out(wire_d53_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5405345(.data_in(wire_d53_44),.data_out(wire_d53_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5405346(.data_in(wire_d53_45),.data_out(wire_d53_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5405347(.data_in(wire_d53_46),.data_out(wire_d53_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405348(.data_in(wire_d53_47),.data_out(wire_d53_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405349(.data_in(wire_d53_48),.data_out(wire_d53_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405350(.data_in(wire_d53_49),.data_out(wire_d53_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405351(.data_in(wire_d53_50),.data_out(wire_d53_51),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5405352(.data_in(wire_d53_51),.data_out(wire_d53_52),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5405353(.data_in(wire_d53_52),.data_out(wire_d53_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405354(.data_in(wire_d53_53),.data_out(wire_d53_54),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5405355(.data_in(wire_d53_54),.data_out(wire_d53_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405356(.data_in(wire_d53_55),.data_out(wire_d53_56),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5405357(.data_in(wire_d53_56),.data_out(wire_d53_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405358(.data_in(wire_d53_57),.data_out(wire_d53_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5405359(.data_in(wire_d53_58),.data_out(wire_d53_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405360(.data_in(wire_d53_59),.data_out(wire_d53_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5405361(.data_in(wire_d53_60),.data_out(wire_d53_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5405362(.data_in(wire_d53_61),.data_out(wire_d53_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5405363(.data_in(wire_d53_62),.data_out(wire_d53_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405364(.data_in(wire_d53_63),.data_out(wire_d53_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405365(.data_in(wire_d53_64),.data_out(wire_d53_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5405366(.data_in(wire_d53_65),.data_out(wire_d53_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5405367(.data_in(wire_d53_66),.data_out(wire_d53_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405368(.data_in(wire_d53_67),.data_out(wire_d53_68),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405369(.data_in(wire_d53_68),.data_out(wire_d53_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5405370(.data_in(wire_d53_69),.data_out(wire_d53_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5405371(.data_in(wire_d53_70),.data_out(wire_d53_71),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5405372(.data_in(wire_d53_71),.data_out(wire_d53_72),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5405373(.data_in(wire_d53_72),.data_out(wire_d53_73),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405374(.data_in(wire_d53_73),.data_out(wire_d53_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405375(.data_in(wire_d53_74),.data_out(wire_d53_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5405376(.data_in(wire_d53_75),.data_out(wire_d53_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405377(.data_in(wire_d53_76),.data_out(wire_d53_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405378(.data_in(wire_d53_77),.data_out(wire_d53_78),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405379(.data_in(wire_d53_78),.data_out(wire_d53_79),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405380(.data_in(wire_d53_79),.data_out(wire_d53_80),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405381(.data_in(wire_d53_80),.data_out(wire_d53_81),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5405382(.data_in(wire_d53_81),.data_out(wire_d53_82),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405383(.data_in(wire_d53_82),.data_out(wire_d53_83),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405384(.data_in(wire_d53_83),.data_out(wire_d53_84),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405385(.data_in(wire_d53_84),.data_out(wire_d53_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5405386(.data_in(wire_d53_85),.data_out(wire_d53_86),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405387(.data_in(wire_d53_86),.data_out(wire_d53_87),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405388(.data_in(wire_d53_87),.data_out(wire_d53_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5405389(.data_in(wire_d53_88),.data_out(wire_d53_89),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405390(.data_in(wire_d53_89),.data_out(wire_d53_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405391(.data_in(wire_d53_90),.data_out(wire_d53_91),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5405392(.data_in(wire_d53_91),.data_out(wire_d53_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5405393(.data_in(wire_d53_92),.data_out(wire_d53_93),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405394(.data_in(wire_d53_93),.data_out(wire_d53_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405395(.data_in(wire_d53_94),.data_out(wire_d53_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5405396(.data_in(wire_d53_95),.data_out(wire_d53_96),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5405397(.data_in(wire_d53_96),.data_out(wire_d53_97),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405398(.data_in(wire_d53_97),.data_out(wire_d53_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5405399(.data_in(wire_d53_98),.data_out(wire_d53_99),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance54053100(.data_in(wire_d53_99),.data_out(wire_d53_100),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance54053101(.data_in(wire_d53_100),.data_out(wire_d53_101),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance54053102(.data_in(wire_d53_101),.data_out(wire_d53_102),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance54053103(.data_in(wire_d53_102),.data_out(wire_d53_103),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance54053104(.data_in(wire_d53_103),.data_out(wire_d53_104),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance54053105(.data_in(wire_d53_104),.data_out(wire_d53_105),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance54053106(.data_in(wire_d53_105),.data_out(wire_d53_106),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance54053107(.data_in(wire_d53_106),.data_out(wire_d53_107),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance54053108(.data_in(wire_d53_107),.data_out(wire_d53_108),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance54053109(.data_in(wire_d53_108),.data_out(wire_d53_109),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance54053110(.data_in(wire_d53_109),.data_out(wire_d53_110),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance54053111(.data_in(wire_d53_110),.data_out(wire_d53_111),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance54053112(.data_in(wire_d53_111),.data_out(wire_d53_112),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance54053113(.data_in(wire_d53_112),.data_out(wire_d53_113),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance54053114(.data_in(wire_d53_113),.data_out(wire_d53_114),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance54053115(.data_in(wire_d53_114),.data_out(wire_d53_115),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance54053116(.data_in(wire_d53_115),.data_out(wire_d53_116),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance54053117(.data_in(wire_d53_116),.data_out(wire_d53_117),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance54053118(.data_in(wire_d53_117),.data_out(wire_d53_118),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance54053119(.data_in(wire_d53_118),.data_out(d_out53),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance550540(.data_in(d_in54),.data_out(wire_d54_0),.clk(clk),.rst(rst));            //channel 55
	large_mux #(.WIDTH(WIDTH)) large_mux_instance550541(.data_in(wire_d54_0),.data_out(wire_d54_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance550542(.data_in(wire_d54_1),.data_out(wire_d54_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance550543(.data_in(wire_d54_2),.data_out(wire_d54_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance550544(.data_in(wire_d54_3),.data_out(wire_d54_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance550545(.data_in(wire_d54_4),.data_out(wire_d54_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance550546(.data_in(wire_d54_5),.data_out(wire_d54_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance550547(.data_in(wire_d54_6),.data_out(wire_d54_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance550548(.data_in(wire_d54_7),.data_out(wire_d54_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance550549(.data_in(wire_d54_8),.data_out(wire_d54_9),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5505410(.data_in(wire_d54_9),.data_out(wire_d54_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5505411(.data_in(wire_d54_10),.data_out(wire_d54_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5505412(.data_in(wire_d54_11),.data_out(wire_d54_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505413(.data_in(wire_d54_12),.data_out(wire_d54_13),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505414(.data_in(wire_d54_13),.data_out(wire_d54_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5505415(.data_in(wire_d54_14),.data_out(wire_d54_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505416(.data_in(wire_d54_15),.data_out(wire_d54_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505417(.data_in(wire_d54_16),.data_out(wire_d54_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5505418(.data_in(wire_d54_17),.data_out(wire_d54_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5505419(.data_in(wire_d54_18),.data_out(wire_d54_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5505420(.data_in(wire_d54_19),.data_out(wire_d54_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505421(.data_in(wire_d54_20),.data_out(wire_d54_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505422(.data_in(wire_d54_21),.data_out(wire_d54_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5505423(.data_in(wire_d54_22),.data_out(wire_d54_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5505424(.data_in(wire_d54_23),.data_out(wire_d54_24),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5505425(.data_in(wire_d54_24),.data_out(wire_d54_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505426(.data_in(wire_d54_25),.data_out(wire_d54_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5505427(.data_in(wire_d54_26),.data_out(wire_d54_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505428(.data_in(wire_d54_27),.data_out(wire_d54_28),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5505429(.data_in(wire_d54_28),.data_out(wire_d54_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5505430(.data_in(wire_d54_29),.data_out(wire_d54_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5505431(.data_in(wire_d54_30),.data_out(wire_d54_31),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5505432(.data_in(wire_d54_31),.data_out(wire_d54_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5505433(.data_in(wire_d54_32),.data_out(wire_d54_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505434(.data_in(wire_d54_33),.data_out(wire_d54_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505435(.data_in(wire_d54_34),.data_out(wire_d54_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505436(.data_in(wire_d54_35),.data_out(wire_d54_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5505437(.data_in(wire_d54_36),.data_out(wire_d54_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505438(.data_in(wire_d54_37),.data_out(wire_d54_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505439(.data_in(wire_d54_38),.data_out(wire_d54_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505440(.data_in(wire_d54_39),.data_out(wire_d54_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5505441(.data_in(wire_d54_40),.data_out(wire_d54_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505442(.data_in(wire_d54_41),.data_out(wire_d54_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505443(.data_in(wire_d54_42),.data_out(wire_d54_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505444(.data_in(wire_d54_43),.data_out(wire_d54_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505445(.data_in(wire_d54_44),.data_out(wire_d54_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505446(.data_in(wire_d54_45),.data_out(wire_d54_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505447(.data_in(wire_d54_46),.data_out(wire_d54_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5505448(.data_in(wire_d54_47),.data_out(wire_d54_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505449(.data_in(wire_d54_48),.data_out(wire_d54_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5505450(.data_in(wire_d54_49),.data_out(wire_d54_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5505451(.data_in(wire_d54_50),.data_out(wire_d54_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5505452(.data_in(wire_d54_51),.data_out(wire_d54_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505453(.data_in(wire_d54_52),.data_out(wire_d54_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5505454(.data_in(wire_d54_53),.data_out(wire_d54_54),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5505455(.data_in(wire_d54_54),.data_out(wire_d54_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5505456(.data_in(wire_d54_55),.data_out(wire_d54_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505457(.data_in(wire_d54_56),.data_out(wire_d54_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505458(.data_in(wire_d54_57),.data_out(wire_d54_58),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5505459(.data_in(wire_d54_58),.data_out(wire_d54_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505460(.data_in(wire_d54_59),.data_out(wire_d54_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5505461(.data_in(wire_d54_60),.data_out(wire_d54_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505462(.data_in(wire_d54_61),.data_out(wire_d54_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505463(.data_in(wire_d54_62),.data_out(wire_d54_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505464(.data_in(wire_d54_63),.data_out(wire_d54_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505465(.data_in(wire_d54_64),.data_out(wire_d54_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505466(.data_in(wire_d54_65),.data_out(wire_d54_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5505467(.data_in(wire_d54_66),.data_out(wire_d54_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505468(.data_in(wire_d54_67),.data_out(wire_d54_68),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505469(.data_in(wire_d54_68),.data_out(wire_d54_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5505470(.data_in(wire_d54_69),.data_out(wire_d54_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505471(.data_in(wire_d54_70),.data_out(wire_d54_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5505472(.data_in(wire_d54_71),.data_out(wire_d54_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505473(.data_in(wire_d54_72),.data_out(wire_d54_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5505474(.data_in(wire_d54_73),.data_out(wire_d54_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505475(.data_in(wire_d54_74),.data_out(wire_d54_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505476(.data_in(wire_d54_75),.data_out(wire_d54_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505477(.data_in(wire_d54_76),.data_out(wire_d54_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5505478(.data_in(wire_d54_77),.data_out(wire_d54_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505479(.data_in(wire_d54_78),.data_out(wire_d54_79),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505480(.data_in(wire_d54_79),.data_out(wire_d54_80),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505481(.data_in(wire_d54_80),.data_out(wire_d54_81),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5505482(.data_in(wire_d54_81),.data_out(wire_d54_82),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505483(.data_in(wire_d54_82),.data_out(wire_d54_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505484(.data_in(wire_d54_83),.data_out(wire_d54_84),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505485(.data_in(wire_d54_84),.data_out(wire_d54_85),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5505486(.data_in(wire_d54_85),.data_out(wire_d54_86),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505487(.data_in(wire_d54_86),.data_out(wire_d54_87),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505488(.data_in(wire_d54_87),.data_out(wire_d54_88),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505489(.data_in(wire_d54_88),.data_out(wire_d54_89),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5505490(.data_in(wire_d54_89),.data_out(wire_d54_90),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505491(.data_in(wire_d54_90),.data_out(wire_d54_91),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505492(.data_in(wire_d54_91),.data_out(wire_d54_92),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5505493(.data_in(wire_d54_92),.data_out(wire_d54_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505494(.data_in(wire_d54_93),.data_out(wire_d54_94),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505495(.data_in(wire_d54_94),.data_out(wire_d54_95),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505496(.data_in(wire_d54_95),.data_out(wire_d54_96),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5505497(.data_in(wire_d54_96),.data_out(wire_d54_97),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5505498(.data_in(wire_d54_97),.data_out(wire_d54_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505499(.data_in(wire_d54_98),.data_out(wire_d54_99),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance55054100(.data_in(wire_d54_99),.data_out(wire_d54_100),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance55054101(.data_in(wire_d54_100),.data_out(wire_d54_101),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance55054102(.data_in(wire_d54_101),.data_out(wire_d54_102),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance55054103(.data_in(wire_d54_102),.data_out(wire_d54_103),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance55054104(.data_in(wire_d54_103),.data_out(wire_d54_104),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance55054105(.data_in(wire_d54_104),.data_out(wire_d54_105),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance55054106(.data_in(wire_d54_105),.data_out(wire_d54_106),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance55054107(.data_in(wire_d54_106),.data_out(wire_d54_107),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance55054108(.data_in(wire_d54_107),.data_out(wire_d54_108),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance55054109(.data_in(wire_d54_108),.data_out(wire_d54_109),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance55054110(.data_in(wire_d54_109),.data_out(wire_d54_110),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance55054111(.data_in(wire_d54_110),.data_out(wire_d54_111),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance55054112(.data_in(wire_d54_111),.data_out(wire_d54_112),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance55054113(.data_in(wire_d54_112),.data_out(wire_d54_113),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance55054114(.data_in(wire_d54_113),.data_out(wire_d54_114),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance55054115(.data_in(wire_d54_114),.data_out(wire_d54_115),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance55054116(.data_in(wire_d54_115),.data_out(wire_d54_116),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance55054117(.data_in(wire_d54_116),.data_out(wire_d54_117),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance55054118(.data_in(wire_d54_117),.data_out(wire_d54_118),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance55054119(.data_in(wire_d54_118),.data_out(d_out54),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance560550(.data_in(d_in55),.data_out(wire_d55_0),.clk(clk),.rst(rst));            //channel 56
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance560551(.data_in(wire_d55_0),.data_out(wire_d55_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance560552(.data_in(wire_d55_1),.data_out(wire_d55_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance560553(.data_in(wire_d55_2),.data_out(wire_d55_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance560554(.data_in(wire_d55_3),.data_out(wire_d55_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance560555(.data_in(wire_d55_4),.data_out(wire_d55_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance560556(.data_in(wire_d55_5),.data_out(wire_d55_6),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance560557(.data_in(wire_d55_6),.data_out(wire_d55_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance560558(.data_in(wire_d55_7),.data_out(wire_d55_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance560559(.data_in(wire_d55_8),.data_out(wire_d55_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605510(.data_in(wire_d55_9),.data_out(wire_d55_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5605511(.data_in(wire_d55_10),.data_out(wire_d55_11),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5605512(.data_in(wire_d55_11),.data_out(wire_d55_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605513(.data_in(wire_d55_12),.data_out(wire_d55_13),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605514(.data_in(wire_d55_13),.data_out(wire_d55_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5605515(.data_in(wire_d55_14),.data_out(wire_d55_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605516(.data_in(wire_d55_15),.data_out(wire_d55_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5605517(.data_in(wire_d55_16),.data_out(wire_d55_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5605518(.data_in(wire_d55_17),.data_out(wire_d55_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5605519(.data_in(wire_d55_18),.data_out(wire_d55_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5605520(.data_in(wire_d55_19),.data_out(wire_d55_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5605521(.data_in(wire_d55_20),.data_out(wire_d55_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5605522(.data_in(wire_d55_21),.data_out(wire_d55_22),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5605523(.data_in(wire_d55_22),.data_out(wire_d55_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605524(.data_in(wire_d55_23),.data_out(wire_d55_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5605525(.data_in(wire_d55_24),.data_out(wire_d55_25),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5605526(.data_in(wire_d55_25),.data_out(wire_d55_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5605527(.data_in(wire_d55_26),.data_out(wire_d55_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5605528(.data_in(wire_d55_27),.data_out(wire_d55_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5605529(.data_in(wire_d55_28),.data_out(wire_d55_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605530(.data_in(wire_d55_29),.data_out(wire_d55_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5605531(.data_in(wire_d55_30),.data_out(wire_d55_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5605532(.data_in(wire_d55_31),.data_out(wire_d55_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5605533(.data_in(wire_d55_32),.data_out(wire_d55_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605534(.data_in(wire_d55_33),.data_out(wire_d55_34),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5605535(.data_in(wire_d55_34),.data_out(wire_d55_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5605536(.data_in(wire_d55_35),.data_out(wire_d55_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5605537(.data_in(wire_d55_36),.data_out(wire_d55_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5605538(.data_in(wire_d55_37),.data_out(wire_d55_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605539(.data_in(wire_d55_38),.data_out(wire_d55_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605540(.data_in(wire_d55_39),.data_out(wire_d55_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605541(.data_in(wire_d55_40),.data_out(wire_d55_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5605542(.data_in(wire_d55_41),.data_out(wire_d55_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605543(.data_in(wire_d55_42),.data_out(wire_d55_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605544(.data_in(wire_d55_43),.data_out(wire_d55_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5605545(.data_in(wire_d55_44),.data_out(wire_d55_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5605546(.data_in(wire_d55_45),.data_out(wire_d55_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5605547(.data_in(wire_d55_46),.data_out(wire_d55_47),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5605548(.data_in(wire_d55_47),.data_out(wire_d55_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5605549(.data_in(wire_d55_48),.data_out(wire_d55_49),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605550(.data_in(wire_d55_49),.data_out(wire_d55_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5605551(.data_in(wire_d55_50),.data_out(wire_d55_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5605552(.data_in(wire_d55_51),.data_out(wire_d55_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5605553(.data_in(wire_d55_52),.data_out(wire_d55_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605554(.data_in(wire_d55_53),.data_out(wire_d55_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605555(.data_in(wire_d55_54),.data_out(wire_d55_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5605556(.data_in(wire_d55_55),.data_out(wire_d55_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5605557(.data_in(wire_d55_56),.data_out(wire_d55_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5605558(.data_in(wire_d55_57),.data_out(wire_d55_58),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5605559(.data_in(wire_d55_58),.data_out(wire_d55_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5605560(.data_in(wire_d55_59),.data_out(wire_d55_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605561(.data_in(wire_d55_60),.data_out(wire_d55_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5605562(.data_in(wire_d55_61),.data_out(wire_d55_62),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5605563(.data_in(wire_d55_62),.data_out(wire_d55_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5605564(.data_in(wire_d55_63),.data_out(wire_d55_64),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5605565(.data_in(wire_d55_64),.data_out(wire_d55_65),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5605566(.data_in(wire_d55_65),.data_out(wire_d55_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605567(.data_in(wire_d55_66),.data_out(wire_d55_67),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5605568(.data_in(wire_d55_67),.data_out(wire_d55_68),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5605569(.data_in(wire_d55_68),.data_out(wire_d55_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605570(.data_in(wire_d55_69),.data_out(wire_d55_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5605571(.data_in(wire_d55_70),.data_out(wire_d55_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5605572(.data_in(wire_d55_71),.data_out(wire_d55_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5605573(.data_in(wire_d55_72),.data_out(wire_d55_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5605574(.data_in(wire_d55_73),.data_out(wire_d55_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605575(.data_in(wire_d55_74),.data_out(wire_d55_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5605576(.data_in(wire_d55_75),.data_out(wire_d55_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5605577(.data_in(wire_d55_76),.data_out(wire_d55_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5605578(.data_in(wire_d55_77),.data_out(wire_d55_78),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5605579(.data_in(wire_d55_78),.data_out(wire_d55_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605580(.data_in(wire_d55_79),.data_out(wire_d55_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5605581(.data_in(wire_d55_80),.data_out(wire_d55_81),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5605582(.data_in(wire_d55_81),.data_out(wire_d55_82),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5605583(.data_in(wire_d55_82),.data_out(wire_d55_83),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5605584(.data_in(wire_d55_83),.data_out(wire_d55_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5605585(.data_in(wire_d55_84),.data_out(wire_d55_85),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5605586(.data_in(wire_d55_85),.data_out(wire_d55_86),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5605587(.data_in(wire_d55_86),.data_out(wire_d55_87),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5605588(.data_in(wire_d55_87),.data_out(wire_d55_88),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5605589(.data_in(wire_d55_88),.data_out(wire_d55_89),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5605590(.data_in(wire_d55_89),.data_out(wire_d55_90),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5605591(.data_in(wire_d55_90),.data_out(wire_d55_91),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5605592(.data_in(wire_d55_91),.data_out(wire_d55_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5605593(.data_in(wire_d55_92),.data_out(wire_d55_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5605594(.data_in(wire_d55_93),.data_out(wire_d55_94),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605595(.data_in(wire_d55_94),.data_out(wire_d55_95),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5605596(.data_in(wire_d55_95),.data_out(wire_d55_96),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5605597(.data_in(wire_d55_96),.data_out(wire_d55_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5605598(.data_in(wire_d55_97),.data_out(wire_d55_98),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5605599(.data_in(wire_d55_98),.data_out(wire_d55_99),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance56055100(.data_in(wire_d55_99),.data_out(wire_d55_100),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance56055101(.data_in(wire_d55_100),.data_out(wire_d55_101),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance56055102(.data_in(wire_d55_101),.data_out(wire_d55_102),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance56055103(.data_in(wire_d55_102),.data_out(wire_d55_103),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance56055104(.data_in(wire_d55_103),.data_out(wire_d55_104),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance56055105(.data_in(wire_d55_104),.data_out(wire_d55_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance56055106(.data_in(wire_d55_105),.data_out(wire_d55_106),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance56055107(.data_in(wire_d55_106),.data_out(wire_d55_107),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance56055108(.data_in(wire_d55_107),.data_out(wire_d55_108),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance56055109(.data_in(wire_d55_108),.data_out(wire_d55_109),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance56055110(.data_in(wire_d55_109),.data_out(wire_d55_110),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance56055111(.data_in(wire_d55_110),.data_out(wire_d55_111),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance56055112(.data_in(wire_d55_111),.data_out(wire_d55_112),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance56055113(.data_in(wire_d55_112),.data_out(wire_d55_113),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance56055114(.data_in(wire_d55_113),.data_out(wire_d55_114),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance56055115(.data_in(wire_d55_114),.data_out(wire_d55_115),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance56055116(.data_in(wire_d55_115),.data_out(wire_d55_116),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance56055117(.data_in(wire_d55_116),.data_out(wire_d55_117),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance56055118(.data_in(wire_d55_117),.data_out(wire_d55_118),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance56055119(.data_in(wire_d55_118),.data_out(d_out55),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance570560(.data_in(d_in56),.data_out(wire_d56_0),.clk(clk),.rst(rst));            //channel 57
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance570561(.data_in(wire_d56_0),.data_out(wire_d56_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance570562(.data_in(wire_d56_1),.data_out(wire_d56_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance570563(.data_in(wire_d56_2),.data_out(wire_d56_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance570564(.data_in(wire_d56_3),.data_out(wire_d56_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance570565(.data_in(wire_d56_4),.data_out(wire_d56_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance570566(.data_in(wire_d56_5),.data_out(wire_d56_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance570567(.data_in(wire_d56_6),.data_out(wire_d56_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance570568(.data_in(wire_d56_7),.data_out(wire_d56_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance570569(.data_in(wire_d56_8),.data_out(wire_d56_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5705610(.data_in(wire_d56_9),.data_out(wire_d56_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705611(.data_in(wire_d56_10),.data_out(wire_d56_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5705612(.data_in(wire_d56_11),.data_out(wire_d56_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5705613(.data_in(wire_d56_12),.data_out(wire_d56_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5705614(.data_in(wire_d56_13),.data_out(wire_d56_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705615(.data_in(wire_d56_14),.data_out(wire_d56_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5705616(.data_in(wire_d56_15),.data_out(wire_d56_16),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5705617(.data_in(wire_d56_16),.data_out(wire_d56_17),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5705618(.data_in(wire_d56_17),.data_out(wire_d56_18),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705619(.data_in(wire_d56_18),.data_out(wire_d56_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705620(.data_in(wire_d56_19),.data_out(wire_d56_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705621(.data_in(wire_d56_20),.data_out(wire_d56_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5705622(.data_in(wire_d56_21),.data_out(wire_d56_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705623(.data_in(wire_d56_22),.data_out(wire_d56_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5705624(.data_in(wire_d56_23),.data_out(wire_d56_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5705625(.data_in(wire_d56_24),.data_out(wire_d56_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5705626(.data_in(wire_d56_25),.data_out(wire_d56_26),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5705627(.data_in(wire_d56_26),.data_out(wire_d56_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705628(.data_in(wire_d56_27),.data_out(wire_d56_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5705629(.data_in(wire_d56_28),.data_out(wire_d56_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5705630(.data_in(wire_d56_29),.data_out(wire_d56_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5705631(.data_in(wire_d56_30),.data_out(wire_d56_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705632(.data_in(wire_d56_31),.data_out(wire_d56_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705633(.data_in(wire_d56_32),.data_out(wire_d56_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5705634(.data_in(wire_d56_33),.data_out(wire_d56_34),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5705635(.data_in(wire_d56_34),.data_out(wire_d56_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5705636(.data_in(wire_d56_35),.data_out(wire_d56_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5705637(.data_in(wire_d56_36),.data_out(wire_d56_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705638(.data_in(wire_d56_37),.data_out(wire_d56_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705639(.data_in(wire_d56_38),.data_out(wire_d56_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5705640(.data_in(wire_d56_39),.data_out(wire_d56_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5705641(.data_in(wire_d56_40),.data_out(wire_d56_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5705642(.data_in(wire_d56_41),.data_out(wire_d56_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705643(.data_in(wire_d56_42),.data_out(wire_d56_43),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705644(.data_in(wire_d56_43),.data_out(wire_d56_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705645(.data_in(wire_d56_44),.data_out(wire_d56_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5705646(.data_in(wire_d56_45),.data_out(wire_d56_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5705647(.data_in(wire_d56_46),.data_out(wire_d56_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5705648(.data_in(wire_d56_47),.data_out(wire_d56_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5705649(.data_in(wire_d56_48),.data_out(wire_d56_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705650(.data_in(wire_d56_49),.data_out(wire_d56_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5705651(.data_in(wire_d56_50),.data_out(wire_d56_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5705652(.data_in(wire_d56_51),.data_out(wire_d56_52),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5705653(.data_in(wire_d56_52),.data_out(wire_d56_53),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5705654(.data_in(wire_d56_53),.data_out(wire_d56_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5705655(.data_in(wire_d56_54),.data_out(wire_d56_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5705656(.data_in(wire_d56_55),.data_out(wire_d56_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5705657(.data_in(wire_d56_56),.data_out(wire_d56_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5705658(.data_in(wire_d56_57),.data_out(wire_d56_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5705659(.data_in(wire_d56_58),.data_out(wire_d56_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705660(.data_in(wire_d56_59),.data_out(wire_d56_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5705661(.data_in(wire_d56_60),.data_out(wire_d56_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5705662(.data_in(wire_d56_61),.data_out(wire_d56_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5705663(.data_in(wire_d56_62),.data_out(wire_d56_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705664(.data_in(wire_d56_63),.data_out(wire_d56_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5705665(.data_in(wire_d56_64),.data_out(wire_d56_65),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5705666(.data_in(wire_d56_65),.data_out(wire_d56_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705667(.data_in(wire_d56_66),.data_out(wire_d56_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5705668(.data_in(wire_d56_67),.data_out(wire_d56_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5705669(.data_in(wire_d56_68),.data_out(wire_d56_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705670(.data_in(wire_d56_69),.data_out(wire_d56_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5705671(.data_in(wire_d56_70),.data_out(wire_d56_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5705672(.data_in(wire_d56_71),.data_out(wire_d56_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705673(.data_in(wire_d56_72),.data_out(wire_d56_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5705674(.data_in(wire_d56_73),.data_out(wire_d56_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5705675(.data_in(wire_d56_74),.data_out(wire_d56_75),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5705676(.data_in(wire_d56_75),.data_out(wire_d56_76),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5705677(.data_in(wire_d56_76),.data_out(wire_d56_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5705678(.data_in(wire_d56_77),.data_out(wire_d56_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5705679(.data_in(wire_d56_78),.data_out(wire_d56_79),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5705680(.data_in(wire_d56_79),.data_out(wire_d56_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5705681(.data_in(wire_d56_80),.data_out(wire_d56_81),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705682(.data_in(wire_d56_81),.data_out(wire_d56_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5705683(.data_in(wire_d56_82),.data_out(wire_d56_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5705684(.data_in(wire_d56_83),.data_out(wire_d56_84),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705685(.data_in(wire_d56_84),.data_out(wire_d56_85),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5705686(.data_in(wire_d56_85),.data_out(wire_d56_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5705687(.data_in(wire_d56_86),.data_out(wire_d56_87),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5705688(.data_in(wire_d56_87),.data_out(wire_d56_88),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5705689(.data_in(wire_d56_88),.data_out(wire_d56_89),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705690(.data_in(wire_d56_89),.data_out(wire_d56_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5705691(.data_in(wire_d56_90),.data_out(wire_d56_91),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705692(.data_in(wire_d56_91),.data_out(wire_d56_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5705693(.data_in(wire_d56_92),.data_out(wire_d56_93),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5705694(.data_in(wire_d56_93),.data_out(wire_d56_94),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5705695(.data_in(wire_d56_94),.data_out(wire_d56_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5705696(.data_in(wire_d56_95),.data_out(wire_d56_96),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5705697(.data_in(wire_d56_96),.data_out(wire_d56_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5705698(.data_in(wire_d56_97),.data_out(wire_d56_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5705699(.data_in(wire_d56_98),.data_out(wire_d56_99),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance57056100(.data_in(wire_d56_99),.data_out(wire_d56_100),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance57056101(.data_in(wire_d56_100),.data_out(wire_d56_101),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance57056102(.data_in(wire_d56_101),.data_out(wire_d56_102),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance57056103(.data_in(wire_d56_102),.data_out(wire_d56_103),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance57056104(.data_in(wire_d56_103),.data_out(wire_d56_104),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance57056105(.data_in(wire_d56_104),.data_out(wire_d56_105),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance57056106(.data_in(wire_d56_105),.data_out(wire_d56_106),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance57056107(.data_in(wire_d56_106),.data_out(wire_d56_107),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance57056108(.data_in(wire_d56_107),.data_out(wire_d56_108),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance57056109(.data_in(wire_d56_108),.data_out(wire_d56_109),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance57056110(.data_in(wire_d56_109),.data_out(wire_d56_110),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance57056111(.data_in(wire_d56_110),.data_out(wire_d56_111),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance57056112(.data_in(wire_d56_111),.data_out(wire_d56_112),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance57056113(.data_in(wire_d56_112),.data_out(wire_d56_113),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance57056114(.data_in(wire_d56_113),.data_out(wire_d56_114),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance57056115(.data_in(wire_d56_114),.data_out(wire_d56_115),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance57056116(.data_in(wire_d56_115),.data_out(wire_d56_116),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance57056117(.data_in(wire_d56_116),.data_out(wire_d56_117),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance57056118(.data_in(wire_d56_117),.data_out(wire_d56_118),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance57056119(.data_in(wire_d56_118),.data_out(d_out56),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance580570(.data_in(d_in57),.data_out(wire_d57_0),.clk(clk),.rst(rst));            //channel 58
	register #(.WIDTH(WIDTH)) register_instance580571(.data_in(wire_d57_0),.data_out(wire_d57_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance580572(.data_in(wire_d57_1),.data_out(wire_d57_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance580573(.data_in(wire_d57_2),.data_out(wire_d57_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance580574(.data_in(wire_d57_3),.data_out(wire_d57_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance580575(.data_in(wire_d57_4),.data_out(wire_d57_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance580576(.data_in(wire_d57_5),.data_out(wire_d57_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance580577(.data_in(wire_d57_6),.data_out(wire_d57_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance580578(.data_in(wire_d57_7),.data_out(wire_d57_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance580579(.data_in(wire_d57_8),.data_out(wire_d57_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5805710(.data_in(wire_d57_9),.data_out(wire_d57_10),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805711(.data_in(wire_d57_10),.data_out(wire_d57_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805712(.data_in(wire_d57_11),.data_out(wire_d57_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805713(.data_in(wire_d57_12),.data_out(wire_d57_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5805714(.data_in(wire_d57_13),.data_out(wire_d57_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805715(.data_in(wire_d57_14),.data_out(wire_d57_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5805716(.data_in(wire_d57_15),.data_out(wire_d57_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5805717(.data_in(wire_d57_16),.data_out(wire_d57_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5805718(.data_in(wire_d57_17),.data_out(wire_d57_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5805719(.data_in(wire_d57_18),.data_out(wire_d57_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5805720(.data_in(wire_d57_19),.data_out(wire_d57_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805721(.data_in(wire_d57_20),.data_out(wire_d57_21),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5805722(.data_in(wire_d57_21),.data_out(wire_d57_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805723(.data_in(wire_d57_22),.data_out(wire_d57_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5805724(.data_in(wire_d57_23),.data_out(wire_d57_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5805725(.data_in(wire_d57_24),.data_out(wire_d57_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5805726(.data_in(wire_d57_25),.data_out(wire_d57_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5805727(.data_in(wire_d57_26),.data_out(wire_d57_27),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5805728(.data_in(wire_d57_27),.data_out(wire_d57_28),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5805729(.data_in(wire_d57_28),.data_out(wire_d57_29),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805730(.data_in(wire_d57_29),.data_out(wire_d57_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5805731(.data_in(wire_d57_30),.data_out(wire_d57_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5805732(.data_in(wire_d57_31),.data_out(wire_d57_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805733(.data_in(wire_d57_32),.data_out(wire_d57_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5805734(.data_in(wire_d57_33),.data_out(wire_d57_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5805735(.data_in(wire_d57_34),.data_out(wire_d57_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5805736(.data_in(wire_d57_35),.data_out(wire_d57_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5805737(.data_in(wire_d57_36),.data_out(wire_d57_37),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5805738(.data_in(wire_d57_37),.data_out(wire_d57_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5805739(.data_in(wire_d57_38),.data_out(wire_d57_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805740(.data_in(wire_d57_39),.data_out(wire_d57_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5805741(.data_in(wire_d57_40),.data_out(wire_d57_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5805742(.data_in(wire_d57_41),.data_out(wire_d57_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805743(.data_in(wire_d57_42),.data_out(wire_d57_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5805744(.data_in(wire_d57_43),.data_out(wire_d57_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5805745(.data_in(wire_d57_44),.data_out(wire_d57_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805746(.data_in(wire_d57_45),.data_out(wire_d57_46),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5805747(.data_in(wire_d57_46),.data_out(wire_d57_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5805748(.data_in(wire_d57_47),.data_out(wire_d57_48),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5805749(.data_in(wire_d57_48),.data_out(wire_d57_49),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5805750(.data_in(wire_d57_49),.data_out(wire_d57_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805751(.data_in(wire_d57_50),.data_out(wire_d57_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5805752(.data_in(wire_d57_51),.data_out(wire_d57_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5805753(.data_in(wire_d57_52),.data_out(wire_d57_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805754(.data_in(wire_d57_53),.data_out(wire_d57_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5805755(.data_in(wire_d57_54),.data_out(wire_d57_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805756(.data_in(wire_d57_55),.data_out(wire_d57_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5805757(.data_in(wire_d57_56),.data_out(wire_d57_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805758(.data_in(wire_d57_57),.data_out(wire_d57_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5805759(.data_in(wire_d57_58),.data_out(wire_d57_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5805760(.data_in(wire_d57_59),.data_out(wire_d57_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5805761(.data_in(wire_d57_60),.data_out(wire_d57_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5805762(.data_in(wire_d57_61),.data_out(wire_d57_62),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805763(.data_in(wire_d57_62),.data_out(wire_d57_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5805764(.data_in(wire_d57_63),.data_out(wire_d57_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805765(.data_in(wire_d57_64),.data_out(wire_d57_65),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5805766(.data_in(wire_d57_65),.data_out(wire_d57_66),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5805767(.data_in(wire_d57_66),.data_out(wire_d57_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805768(.data_in(wire_d57_67),.data_out(wire_d57_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805769(.data_in(wire_d57_68),.data_out(wire_d57_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5805770(.data_in(wire_d57_69),.data_out(wire_d57_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5805771(.data_in(wire_d57_70),.data_out(wire_d57_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5805772(.data_in(wire_d57_71),.data_out(wire_d57_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805773(.data_in(wire_d57_72),.data_out(wire_d57_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805774(.data_in(wire_d57_73),.data_out(wire_d57_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5805775(.data_in(wire_d57_74),.data_out(wire_d57_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5805776(.data_in(wire_d57_75),.data_out(wire_d57_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5805777(.data_in(wire_d57_76),.data_out(wire_d57_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5805778(.data_in(wire_d57_77),.data_out(wire_d57_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5805779(.data_in(wire_d57_78),.data_out(wire_d57_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5805780(.data_in(wire_d57_79),.data_out(wire_d57_80),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805781(.data_in(wire_d57_80),.data_out(wire_d57_81),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805782(.data_in(wire_d57_81),.data_out(wire_d57_82),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805783(.data_in(wire_d57_82),.data_out(wire_d57_83),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805784(.data_in(wire_d57_83),.data_out(wire_d57_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5805785(.data_in(wire_d57_84),.data_out(wire_d57_85),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5805786(.data_in(wire_d57_85),.data_out(wire_d57_86),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5805787(.data_in(wire_d57_86),.data_out(wire_d57_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5805788(.data_in(wire_d57_87),.data_out(wire_d57_88),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805789(.data_in(wire_d57_88),.data_out(wire_d57_89),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805790(.data_in(wire_d57_89),.data_out(wire_d57_90),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805791(.data_in(wire_d57_90),.data_out(wire_d57_91),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5805792(.data_in(wire_d57_91),.data_out(wire_d57_92),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805793(.data_in(wire_d57_92),.data_out(wire_d57_93),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5805794(.data_in(wire_d57_93),.data_out(wire_d57_94),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805795(.data_in(wire_d57_94),.data_out(wire_d57_95),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5805796(.data_in(wire_d57_95),.data_out(wire_d57_96),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5805797(.data_in(wire_d57_96),.data_out(wire_d57_97),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5805798(.data_in(wire_d57_97),.data_out(wire_d57_98),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5805799(.data_in(wire_d57_98),.data_out(wire_d57_99),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance58057100(.data_in(wire_d57_99),.data_out(wire_d57_100),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance58057101(.data_in(wire_d57_100),.data_out(wire_d57_101),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance58057102(.data_in(wire_d57_101),.data_out(wire_d57_102),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance58057103(.data_in(wire_d57_102),.data_out(wire_d57_103),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance58057104(.data_in(wire_d57_103),.data_out(wire_d57_104),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance58057105(.data_in(wire_d57_104),.data_out(wire_d57_105),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance58057106(.data_in(wire_d57_105),.data_out(wire_d57_106),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance58057107(.data_in(wire_d57_106),.data_out(wire_d57_107),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance58057108(.data_in(wire_d57_107),.data_out(wire_d57_108),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance58057109(.data_in(wire_d57_108),.data_out(wire_d57_109),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance58057110(.data_in(wire_d57_109),.data_out(wire_d57_110),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance58057111(.data_in(wire_d57_110),.data_out(wire_d57_111),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance58057112(.data_in(wire_d57_111),.data_out(wire_d57_112),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance58057113(.data_in(wire_d57_112),.data_out(wire_d57_113),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance58057114(.data_in(wire_d57_113),.data_out(wire_d57_114),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance58057115(.data_in(wire_d57_114),.data_out(wire_d57_115),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance58057116(.data_in(wire_d57_115),.data_out(wire_d57_116),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance58057117(.data_in(wire_d57_116),.data_out(wire_d57_117),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance58057118(.data_in(wire_d57_117),.data_out(wire_d57_118),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance58057119(.data_in(wire_d57_118),.data_out(d_out57),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance590580(.data_in(d_in58),.data_out(wire_d58_0),.clk(clk),.rst(rst));            //channel 59
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance590581(.data_in(wire_d58_0),.data_out(wire_d58_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance590582(.data_in(wire_d58_1),.data_out(wire_d58_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance590583(.data_in(wire_d58_2),.data_out(wire_d58_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance590584(.data_in(wire_d58_3),.data_out(wire_d58_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance590585(.data_in(wire_d58_4),.data_out(wire_d58_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance590586(.data_in(wire_d58_5),.data_out(wire_d58_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance590587(.data_in(wire_d58_6),.data_out(wire_d58_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance590588(.data_in(wire_d58_7),.data_out(wire_d58_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance590589(.data_in(wire_d58_8),.data_out(wire_d58_9),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5905810(.data_in(wire_d58_9),.data_out(wire_d58_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5905811(.data_in(wire_d58_10),.data_out(wire_d58_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905812(.data_in(wire_d58_11),.data_out(wire_d58_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5905813(.data_in(wire_d58_12),.data_out(wire_d58_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905814(.data_in(wire_d58_13),.data_out(wire_d58_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5905815(.data_in(wire_d58_14),.data_out(wire_d58_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5905816(.data_in(wire_d58_15),.data_out(wire_d58_16),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5905817(.data_in(wire_d58_16),.data_out(wire_d58_17),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905818(.data_in(wire_d58_17),.data_out(wire_d58_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5905819(.data_in(wire_d58_18),.data_out(wire_d58_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5905820(.data_in(wire_d58_19),.data_out(wire_d58_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5905821(.data_in(wire_d58_20),.data_out(wire_d58_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5905822(.data_in(wire_d58_21),.data_out(wire_d58_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905823(.data_in(wire_d58_22),.data_out(wire_d58_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5905824(.data_in(wire_d58_23),.data_out(wire_d58_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5905825(.data_in(wire_d58_24),.data_out(wire_d58_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5905826(.data_in(wire_d58_25),.data_out(wire_d58_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5905827(.data_in(wire_d58_26),.data_out(wire_d58_27),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5905828(.data_in(wire_d58_27),.data_out(wire_d58_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905829(.data_in(wire_d58_28),.data_out(wire_d58_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5905830(.data_in(wire_d58_29),.data_out(wire_d58_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5905831(.data_in(wire_d58_30),.data_out(wire_d58_31),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5905832(.data_in(wire_d58_31),.data_out(wire_d58_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5905833(.data_in(wire_d58_32),.data_out(wire_d58_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5905834(.data_in(wire_d58_33),.data_out(wire_d58_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5905835(.data_in(wire_d58_34),.data_out(wire_d58_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5905836(.data_in(wire_d58_35),.data_out(wire_d58_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5905837(.data_in(wire_d58_36),.data_out(wire_d58_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5905838(.data_in(wire_d58_37),.data_out(wire_d58_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905839(.data_in(wire_d58_38),.data_out(wire_d58_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5905840(.data_in(wire_d58_39),.data_out(wire_d58_40),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5905841(.data_in(wire_d58_40),.data_out(wire_d58_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905842(.data_in(wire_d58_41),.data_out(wire_d58_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5905843(.data_in(wire_d58_42),.data_out(wire_d58_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5905844(.data_in(wire_d58_43),.data_out(wire_d58_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5905845(.data_in(wire_d58_44),.data_out(wire_d58_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905846(.data_in(wire_d58_45),.data_out(wire_d58_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905847(.data_in(wire_d58_46),.data_out(wire_d58_47),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905848(.data_in(wire_d58_47),.data_out(wire_d58_48),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5905849(.data_in(wire_d58_48),.data_out(wire_d58_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5905850(.data_in(wire_d58_49),.data_out(wire_d58_50),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5905851(.data_in(wire_d58_50),.data_out(wire_d58_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5905852(.data_in(wire_d58_51),.data_out(wire_d58_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5905853(.data_in(wire_d58_52),.data_out(wire_d58_53),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5905854(.data_in(wire_d58_53),.data_out(wire_d58_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5905855(.data_in(wire_d58_54),.data_out(wire_d58_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5905856(.data_in(wire_d58_55),.data_out(wire_d58_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5905857(.data_in(wire_d58_56),.data_out(wire_d58_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5905858(.data_in(wire_d58_57),.data_out(wire_d58_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5905859(.data_in(wire_d58_58),.data_out(wire_d58_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905860(.data_in(wire_d58_59),.data_out(wire_d58_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5905861(.data_in(wire_d58_60),.data_out(wire_d58_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905862(.data_in(wire_d58_61),.data_out(wire_d58_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5905863(.data_in(wire_d58_62),.data_out(wire_d58_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5905864(.data_in(wire_d58_63),.data_out(wire_d58_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5905865(.data_in(wire_d58_64),.data_out(wire_d58_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5905866(.data_in(wire_d58_65),.data_out(wire_d58_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5905867(.data_in(wire_d58_66),.data_out(wire_d58_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5905868(.data_in(wire_d58_67),.data_out(wire_d58_68),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5905869(.data_in(wire_d58_68),.data_out(wire_d58_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5905870(.data_in(wire_d58_69),.data_out(wire_d58_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5905871(.data_in(wire_d58_70),.data_out(wire_d58_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905872(.data_in(wire_d58_71),.data_out(wire_d58_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905873(.data_in(wire_d58_72),.data_out(wire_d58_73),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5905874(.data_in(wire_d58_73),.data_out(wire_d58_74),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5905875(.data_in(wire_d58_74),.data_out(wire_d58_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5905876(.data_in(wire_d58_75),.data_out(wire_d58_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5905877(.data_in(wire_d58_76),.data_out(wire_d58_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5905878(.data_in(wire_d58_77),.data_out(wire_d58_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5905879(.data_in(wire_d58_78),.data_out(wire_d58_79),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5905880(.data_in(wire_d58_79),.data_out(wire_d58_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5905881(.data_in(wire_d58_80),.data_out(wire_d58_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5905882(.data_in(wire_d58_81),.data_out(wire_d58_82),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905883(.data_in(wire_d58_82),.data_out(wire_d58_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5905884(.data_in(wire_d58_83),.data_out(wire_d58_84),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5905885(.data_in(wire_d58_84),.data_out(wire_d58_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5905886(.data_in(wire_d58_85),.data_out(wire_d58_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5905887(.data_in(wire_d58_86),.data_out(wire_d58_87),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5905888(.data_in(wire_d58_87),.data_out(wire_d58_88),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5905889(.data_in(wire_d58_88),.data_out(wire_d58_89),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905890(.data_in(wire_d58_89),.data_out(wire_d58_90),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5905891(.data_in(wire_d58_90),.data_out(wire_d58_91),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5905892(.data_in(wire_d58_91),.data_out(wire_d58_92),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5905893(.data_in(wire_d58_92),.data_out(wire_d58_93),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5905894(.data_in(wire_d58_93),.data_out(wire_d58_94),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905895(.data_in(wire_d58_94),.data_out(wire_d58_95),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5905896(.data_in(wire_d58_95),.data_out(wire_d58_96),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5905897(.data_in(wire_d58_96),.data_out(wire_d58_97),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5905898(.data_in(wire_d58_97),.data_out(wire_d58_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5905899(.data_in(wire_d58_98),.data_out(wire_d58_99),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance59058100(.data_in(wire_d58_99),.data_out(wire_d58_100),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance59058101(.data_in(wire_d58_100),.data_out(wire_d58_101),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance59058102(.data_in(wire_d58_101),.data_out(wire_d58_102),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance59058103(.data_in(wire_d58_102),.data_out(wire_d58_103),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance59058104(.data_in(wire_d58_103),.data_out(wire_d58_104),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance59058105(.data_in(wire_d58_104),.data_out(wire_d58_105),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance59058106(.data_in(wire_d58_105),.data_out(wire_d58_106),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance59058107(.data_in(wire_d58_106),.data_out(wire_d58_107),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance59058108(.data_in(wire_d58_107),.data_out(wire_d58_108),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance59058109(.data_in(wire_d58_108),.data_out(wire_d58_109),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance59058110(.data_in(wire_d58_109),.data_out(wire_d58_110),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance59058111(.data_in(wire_d58_110),.data_out(wire_d58_111),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance59058112(.data_in(wire_d58_111),.data_out(wire_d58_112),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance59058113(.data_in(wire_d58_112),.data_out(wire_d58_113),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance59058114(.data_in(wire_d58_113),.data_out(wire_d58_114),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance59058115(.data_in(wire_d58_114),.data_out(wire_d58_115),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance59058116(.data_in(wire_d58_115),.data_out(wire_d58_116),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance59058117(.data_in(wire_d58_116),.data_out(wire_d58_117),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance59058118(.data_in(wire_d58_117),.data_out(wire_d58_118),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance59058119(.data_in(wire_d58_118),.data_out(d_out58),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance600590(.data_in(d_in59),.data_out(wire_d59_0),.clk(clk),.rst(rst));            //channel 60
	large_mux #(.WIDTH(WIDTH)) large_mux_instance600591(.data_in(wire_d59_0),.data_out(wire_d59_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance600592(.data_in(wire_d59_1),.data_out(wire_d59_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance600593(.data_in(wire_d59_2),.data_out(wire_d59_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance600594(.data_in(wire_d59_3),.data_out(wire_d59_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance600595(.data_in(wire_d59_4),.data_out(wire_d59_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance600596(.data_in(wire_d59_5),.data_out(wire_d59_6),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance600597(.data_in(wire_d59_6),.data_out(wire_d59_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance600598(.data_in(wire_d59_7),.data_out(wire_d59_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance600599(.data_in(wire_d59_8),.data_out(wire_d59_9),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005910(.data_in(wire_d59_9),.data_out(wire_d59_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6005911(.data_in(wire_d59_10),.data_out(wire_d59_11),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6005912(.data_in(wire_d59_11),.data_out(wire_d59_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6005913(.data_in(wire_d59_12),.data_out(wire_d59_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005914(.data_in(wire_d59_13),.data_out(wire_d59_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6005915(.data_in(wire_d59_14),.data_out(wire_d59_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6005916(.data_in(wire_d59_15),.data_out(wire_d59_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6005917(.data_in(wire_d59_16),.data_out(wire_d59_17),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6005918(.data_in(wire_d59_17),.data_out(wire_d59_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005919(.data_in(wire_d59_18),.data_out(wire_d59_19),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6005920(.data_in(wire_d59_19),.data_out(wire_d59_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6005921(.data_in(wire_d59_20),.data_out(wire_d59_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6005922(.data_in(wire_d59_21),.data_out(wire_d59_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6005923(.data_in(wire_d59_22),.data_out(wire_d59_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005924(.data_in(wire_d59_23),.data_out(wire_d59_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005925(.data_in(wire_d59_24),.data_out(wire_d59_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005926(.data_in(wire_d59_25),.data_out(wire_d59_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005927(.data_in(wire_d59_26),.data_out(wire_d59_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005928(.data_in(wire_d59_27),.data_out(wire_d59_28),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6005929(.data_in(wire_d59_28),.data_out(wire_d59_29),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6005930(.data_in(wire_d59_29),.data_out(wire_d59_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005931(.data_in(wire_d59_30),.data_out(wire_d59_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6005932(.data_in(wire_d59_31),.data_out(wire_d59_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6005933(.data_in(wire_d59_32),.data_out(wire_d59_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005934(.data_in(wire_d59_33),.data_out(wire_d59_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6005935(.data_in(wire_d59_34),.data_out(wire_d59_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6005936(.data_in(wire_d59_35),.data_out(wire_d59_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6005937(.data_in(wire_d59_36),.data_out(wire_d59_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6005938(.data_in(wire_d59_37),.data_out(wire_d59_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005939(.data_in(wire_d59_38),.data_out(wire_d59_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005940(.data_in(wire_d59_39),.data_out(wire_d59_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6005941(.data_in(wire_d59_40),.data_out(wire_d59_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6005942(.data_in(wire_d59_41),.data_out(wire_d59_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6005943(.data_in(wire_d59_42),.data_out(wire_d59_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6005944(.data_in(wire_d59_43),.data_out(wire_d59_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6005945(.data_in(wire_d59_44),.data_out(wire_d59_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6005946(.data_in(wire_d59_45),.data_out(wire_d59_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6005947(.data_in(wire_d59_46),.data_out(wire_d59_47),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005948(.data_in(wire_d59_47),.data_out(wire_d59_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005949(.data_in(wire_d59_48),.data_out(wire_d59_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6005950(.data_in(wire_d59_49),.data_out(wire_d59_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6005951(.data_in(wire_d59_50),.data_out(wire_d59_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005952(.data_in(wire_d59_51),.data_out(wire_d59_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6005953(.data_in(wire_d59_52),.data_out(wire_d59_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005954(.data_in(wire_d59_53),.data_out(wire_d59_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005955(.data_in(wire_d59_54),.data_out(wire_d59_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6005956(.data_in(wire_d59_55),.data_out(wire_d59_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6005957(.data_in(wire_d59_56),.data_out(wire_d59_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6005958(.data_in(wire_d59_57),.data_out(wire_d59_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6005959(.data_in(wire_d59_58),.data_out(wire_d59_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005960(.data_in(wire_d59_59),.data_out(wire_d59_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6005961(.data_in(wire_d59_60),.data_out(wire_d59_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6005962(.data_in(wire_d59_61),.data_out(wire_d59_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6005963(.data_in(wire_d59_62),.data_out(wire_d59_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005964(.data_in(wire_d59_63),.data_out(wire_d59_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005965(.data_in(wire_d59_64),.data_out(wire_d59_65),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6005966(.data_in(wire_d59_65),.data_out(wire_d59_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6005967(.data_in(wire_d59_66),.data_out(wire_d59_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6005968(.data_in(wire_d59_67),.data_out(wire_d59_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6005969(.data_in(wire_d59_68),.data_out(wire_d59_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005970(.data_in(wire_d59_69),.data_out(wire_d59_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6005971(.data_in(wire_d59_70),.data_out(wire_d59_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6005972(.data_in(wire_d59_71),.data_out(wire_d59_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005973(.data_in(wire_d59_72),.data_out(wire_d59_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005974(.data_in(wire_d59_73),.data_out(wire_d59_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6005975(.data_in(wire_d59_74),.data_out(wire_d59_75),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005976(.data_in(wire_d59_75),.data_out(wire_d59_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6005977(.data_in(wire_d59_76),.data_out(wire_d59_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6005978(.data_in(wire_d59_77),.data_out(wire_d59_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6005979(.data_in(wire_d59_78),.data_out(wire_d59_79),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005980(.data_in(wire_d59_79),.data_out(wire_d59_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6005981(.data_in(wire_d59_80),.data_out(wire_d59_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6005982(.data_in(wire_d59_81),.data_out(wire_d59_82),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005983(.data_in(wire_d59_82),.data_out(wire_d59_83),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005984(.data_in(wire_d59_83),.data_out(wire_d59_84),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005985(.data_in(wire_d59_84),.data_out(wire_d59_85),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005986(.data_in(wire_d59_85),.data_out(wire_d59_86),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005987(.data_in(wire_d59_86),.data_out(wire_d59_87),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6005988(.data_in(wire_d59_87),.data_out(wire_d59_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6005989(.data_in(wire_d59_88),.data_out(wire_d59_89),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6005990(.data_in(wire_d59_89),.data_out(wire_d59_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6005991(.data_in(wire_d59_90),.data_out(wire_d59_91),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6005992(.data_in(wire_d59_91),.data_out(wire_d59_92),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6005993(.data_in(wire_d59_92),.data_out(wire_d59_93),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6005994(.data_in(wire_d59_93),.data_out(wire_d59_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6005995(.data_in(wire_d59_94),.data_out(wire_d59_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6005996(.data_in(wire_d59_95),.data_out(wire_d59_96),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6005997(.data_in(wire_d59_96),.data_out(wire_d59_97),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6005998(.data_in(wire_d59_97),.data_out(wire_d59_98),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6005999(.data_in(wire_d59_98),.data_out(wire_d59_99),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance60059100(.data_in(wire_d59_99),.data_out(wire_d59_100),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance60059101(.data_in(wire_d59_100),.data_out(wire_d59_101),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance60059102(.data_in(wire_d59_101),.data_out(wire_d59_102),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance60059103(.data_in(wire_d59_102),.data_out(wire_d59_103),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance60059104(.data_in(wire_d59_103),.data_out(wire_d59_104),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance60059105(.data_in(wire_d59_104),.data_out(wire_d59_105),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance60059106(.data_in(wire_d59_105),.data_out(wire_d59_106),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance60059107(.data_in(wire_d59_106),.data_out(wire_d59_107),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance60059108(.data_in(wire_d59_107),.data_out(wire_d59_108),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance60059109(.data_in(wire_d59_108),.data_out(wire_d59_109),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance60059110(.data_in(wire_d59_109),.data_out(wire_d59_110),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance60059111(.data_in(wire_d59_110),.data_out(wire_d59_111),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance60059112(.data_in(wire_d59_111),.data_out(wire_d59_112),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance60059113(.data_in(wire_d59_112),.data_out(wire_d59_113),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance60059114(.data_in(wire_d59_113),.data_out(wire_d59_114),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance60059115(.data_in(wire_d59_114),.data_out(wire_d59_115),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance60059116(.data_in(wire_d59_115),.data_out(wire_d59_116),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance60059117(.data_in(wire_d59_116),.data_out(wire_d59_117),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance60059118(.data_in(wire_d59_117),.data_out(wire_d59_118),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance60059119(.data_in(wire_d59_118),.data_out(d_out59),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance610600(.data_in(d_in60),.data_out(wire_d60_0),.clk(clk),.rst(rst));            //channel 61
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance610601(.data_in(wire_d60_0),.data_out(wire_d60_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance610602(.data_in(wire_d60_1),.data_out(wire_d60_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance610603(.data_in(wire_d60_2),.data_out(wire_d60_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance610604(.data_in(wire_d60_3),.data_out(wire_d60_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance610605(.data_in(wire_d60_4),.data_out(wire_d60_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance610606(.data_in(wire_d60_5),.data_out(wire_d60_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance610607(.data_in(wire_d60_6),.data_out(wire_d60_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance610608(.data_in(wire_d60_7),.data_out(wire_d60_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance610609(.data_in(wire_d60_8),.data_out(wire_d60_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6106010(.data_in(wire_d60_9),.data_out(wire_d60_10),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6106011(.data_in(wire_d60_10),.data_out(wire_d60_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6106012(.data_in(wire_d60_11),.data_out(wire_d60_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6106013(.data_in(wire_d60_12),.data_out(wire_d60_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6106014(.data_in(wire_d60_13),.data_out(wire_d60_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6106015(.data_in(wire_d60_14),.data_out(wire_d60_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6106016(.data_in(wire_d60_15),.data_out(wire_d60_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6106017(.data_in(wire_d60_16),.data_out(wire_d60_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6106018(.data_in(wire_d60_17),.data_out(wire_d60_18),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6106019(.data_in(wire_d60_18),.data_out(wire_d60_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6106020(.data_in(wire_d60_19),.data_out(wire_d60_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6106021(.data_in(wire_d60_20),.data_out(wire_d60_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6106022(.data_in(wire_d60_21),.data_out(wire_d60_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6106023(.data_in(wire_d60_22),.data_out(wire_d60_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6106024(.data_in(wire_d60_23),.data_out(wire_d60_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6106025(.data_in(wire_d60_24),.data_out(wire_d60_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6106026(.data_in(wire_d60_25),.data_out(wire_d60_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6106027(.data_in(wire_d60_26),.data_out(wire_d60_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6106028(.data_in(wire_d60_27),.data_out(wire_d60_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6106029(.data_in(wire_d60_28),.data_out(wire_d60_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6106030(.data_in(wire_d60_29),.data_out(wire_d60_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6106031(.data_in(wire_d60_30),.data_out(wire_d60_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6106032(.data_in(wire_d60_31),.data_out(wire_d60_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6106033(.data_in(wire_d60_32),.data_out(wire_d60_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6106034(.data_in(wire_d60_33),.data_out(wire_d60_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6106035(.data_in(wire_d60_34),.data_out(wire_d60_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6106036(.data_in(wire_d60_35),.data_out(wire_d60_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6106037(.data_in(wire_d60_36),.data_out(wire_d60_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6106038(.data_in(wire_d60_37),.data_out(wire_d60_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6106039(.data_in(wire_d60_38),.data_out(wire_d60_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6106040(.data_in(wire_d60_39),.data_out(wire_d60_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6106041(.data_in(wire_d60_40),.data_out(wire_d60_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6106042(.data_in(wire_d60_41),.data_out(wire_d60_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6106043(.data_in(wire_d60_42),.data_out(wire_d60_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6106044(.data_in(wire_d60_43),.data_out(wire_d60_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6106045(.data_in(wire_d60_44),.data_out(wire_d60_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6106046(.data_in(wire_d60_45),.data_out(wire_d60_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6106047(.data_in(wire_d60_46),.data_out(wire_d60_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6106048(.data_in(wire_d60_47),.data_out(wire_d60_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6106049(.data_in(wire_d60_48),.data_out(wire_d60_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6106050(.data_in(wire_d60_49),.data_out(wire_d60_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6106051(.data_in(wire_d60_50),.data_out(wire_d60_51),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6106052(.data_in(wire_d60_51),.data_out(wire_d60_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6106053(.data_in(wire_d60_52),.data_out(wire_d60_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6106054(.data_in(wire_d60_53),.data_out(wire_d60_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6106055(.data_in(wire_d60_54),.data_out(wire_d60_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6106056(.data_in(wire_d60_55),.data_out(wire_d60_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6106057(.data_in(wire_d60_56),.data_out(wire_d60_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6106058(.data_in(wire_d60_57),.data_out(wire_d60_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6106059(.data_in(wire_d60_58),.data_out(wire_d60_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6106060(.data_in(wire_d60_59),.data_out(wire_d60_60),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6106061(.data_in(wire_d60_60),.data_out(wire_d60_61),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6106062(.data_in(wire_d60_61),.data_out(wire_d60_62),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6106063(.data_in(wire_d60_62),.data_out(wire_d60_63),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6106064(.data_in(wire_d60_63),.data_out(wire_d60_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6106065(.data_in(wire_d60_64),.data_out(wire_d60_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6106066(.data_in(wire_d60_65),.data_out(wire_d60_66),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6106067(.data_in(wire_d60_66),.data_out(wire_d60_67),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6106068(.data_in(wire_d60_67),.data_out(wire_d60_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6106069(.data_in(wire_d60_68),.data_out(wire_d60_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6106070(.data_in(wire_d60_69),.data_out(wire_d60_70),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6106071(.data_in(wire_d60_70),.data_out(wire_d60_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6106072(.data_in(wire_d60_71),.data_out(wire_d60_72),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6106073(.data_in(wire_d60_72),.data_out(wire_d60_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6106074(.data_in(wire_d60_73),.data_out(wire_d60_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6106075(.data_in(wire_d60_74),.data_out(wire_d60_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6106076(.data_in(wire_d60_75),.data_out(wire_d60_76),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6106077(.data_in(wire_d60_76),.data_out(wire_d60_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6106078(.data_in(wire_d60_77),.data_out(wire_d60_78),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6106079(.data_in(wire_d60_78),.data_out(wire_d60_79),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6106080(.data_in(wire_d60_79),.data_out(wire_d60_80),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6106081(.data_in(wire_d60_80),.data_out(wire_d60_81),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6106082(.data_in(wire_d60_81),.data_out(wire_d60_82),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6106083(.data_in(wire_d60_82),.data_out(wire_d60_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6106084(.data_in(wire_d60_83),.data_out(wire_d60_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6106085(.data_in(wire_d60_84),.data_out(wire_d60_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6106086(.data_in(wire_d60_85),.data_out(wire_d60_86),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6106087(.data_in(wire_d60_86),.data_out(wire_d60_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6106088(.data_in(wire_d60_87),.data_out(wire_d60_88),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6106089(.data_in(wire_d60_88),.data_out(wire_d60_89),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6106090(.data_in(wire_d60_89),.data_out(wire_d60_90),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6106091(.data_in(wire_d60_90),.data_out(wire_d60_91),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6106092(.data_in(wire_d60_91),.data_out(wire_d60_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6106093(.data_in(wire_d60_92),.data_out(wire_d60_93),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6106094(.data_in(wire_d60_93),.data_out(wire_d60_94),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6106095(.data_in(wire_d60_94),.data_out(wire_d60_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6106096(.data_in(wire_d60_95),.data_out(wire_d60_96),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6106097(.data_in(wire_d60_96),.data_out(wire_d60_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6106098(.data_in(wire_d60_97),.data_out(wire_d60_98),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6106099(.data_in(wire_d60_98),.data_out(wire_d60_99),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance61060100(.data_in(wire_d60_99),.data_out(wire_d60_100),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance61060101(.data_in(wire_d60_100),.data_out(wire_d60_101),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance61060102(.data_in(wire_d60_101),.data_out(wire_d60_102),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance61060103(.data_in(wire_d60_102),.data_out(wire_d60_103),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance61060104(.data_in(wire_d60_103),.data_out(wire_d60_104),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance61060105(.data_in(wire_d60_104),.data_out(wire_d60_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance61060106(.data_in(wire_d60_105),.data_out(wire_d60_106),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance61060107(.data_in(wire_d60_106),.data_out(wire_d60_107),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance61060108(.data_in(wire_d60_107),.data_out(wire_d60_108),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance61060109(.data_in(wire_d60_108),.data_out(wire_d60_109),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance61060110(.data_in(wire_d60_109),.data_out(wire_d60_110),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance61060111(.data_in(wire_d60_110),.data_out(wire_d60_111),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance61060112(.data_in(wire_d60_111),.data_out(wire_d60_112),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance61060113(.data_in(wire_d60_112),.data_out(wire_d60_113),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance61060114(.data_in(wire_d60_113),.data_out(wire_d60_114),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance61060115(.data_in(wire_d60_114),.data_out(wire_d60_115),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance61060116(.data_in(wire_d60_115),.data_out(wire_d60_116),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance61060117(.data_in(wire_d60_116),.data_out(wire_d60_117),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance61060118(.data_in(wire_d60_117),.data_out(wire_d60_118),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance61060119(.data_in(wire_d60_118),.data_out(d_out60),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance620610(.data_in(d_in61),.data_out(wire_d61_0),.clk(clk),.rst(rst));            //channel 62
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance620611(.data_in(wire_d61_0),.data_out(wire_d61_1),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance620612(.data_in(wire_d61_1),.data_out(wire_d61_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance620613(.data_in(wire_d61_2),.data_out(wire_d61_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance620614(.data_in(wire_d61_3),.data_out(wire_d61_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance620615(.data_in(wire_d61_4),.data_out(wire_d61_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance620616(.data_in(wire_d61_5),.data_out(wire_d61_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance620617(.data_in(wire_d61_6),.data_out(wire_d61_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance620618(.data_in(wire_d61_7),.data_out(wire_d61_8),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance620619(.data_in(wire_d61_8),.data_out(wire_d61_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6206110(.data_in(wire_d61_9),.data_out(wire_d61_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6206111(.data_in(wire_d61_10),.data_out(wire_d61_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6206112(.data_in(wire_d61_11),.data_out(wire_d61_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6206113(.data_in(wire_d61_12),.data_out(wire_d61_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6206114(.data_in(wire_d61_13),.data_out(wire_d61_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6206115(.data_in(wire_d61_14),.data_out(wire_d61_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6206116(.data_in(wire_d61_15),.data_out(wire_d61_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6206117(.data_in(wire_d61_16),.data_out(wire_d61_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6206118(.data_in(wire_d61_17),.data_out(wire_d61_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6206119(.data_in(wire_d61_18),.data_out(wire_d61_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6206120(.data_in(wire_d61_19),.data_out(wire_d61_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6206121(.data_in(wire_d61_20),.data_out(wire_d61_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6206122(.data_in(wire_d61_21),.data_out(wire_d61_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6206123(.data_in(wire_d61_22),.data_out(wire_d61_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6206124(.data_in(wire_d61_23),.data_out(wire_d61_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6206125(.data_in(wire_d61_24),.data_out(wire_d61_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6206126(.data_in(wire_d61_25),.data_out(wire_d61_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6206127(.data_in(wire_d61_26),.data_out(wire_d61_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6206128(.data_in(wire_d61_27),.data_out(wire_d61_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6206129(.data_in(wire_d61_28),.data_out(wire_d61_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6206130(.data_in(wire_d61_29),.data_out(wire_d61_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6206131(.data_in(wire_d61_30),.data_out(wire_d61_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6206132(.data_in(wire_d61_31),.data_out(wire_d61_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6206133(.data_in(wire_d61_32),.data_out(wire_d61_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6206134(.data_in(wire_d61_33),.data_out(wire_d61_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6206135(.data_in(wire_d61_34),.data_out(wire_d61_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6206136(.data_in(wire_d61_35),.data_out(wire_d61_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6206137(.data_in(wire_d61_36),.data_out(wire_d61_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6206138(.data_in(wire_d61_37),.data_out(wire_d61_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6206139(.data_in(wire_d61_38),.data_out(wire_d61_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6206140(.data_in(wire_d61_39),.data_out(wire_d61_40),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6206141(.data_in(wire_d61_40),.data_out(wire_d61_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6206142(.data_in(wire_d61_41),.data_out(wire_d61_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6206143(.data_in(wire_d61_42),.data_out(wire_d61_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6206144(.data_in(wire_d61_43),.data_out(wire_d61_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6206145(.data_in(wire_d61_44),.data_out(wire_d61_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6206146(.data_in(wire_d61_45),.data_out(wire_d61_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6206147(.data_in(wire_d61_46),.data_out(wire_d61_47),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6206148(.data_in(wire_d61_47),.data_out(wire_d61_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6206149(.data_in(wire_d61_48),.data_out(wire_d61_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6206150(.data_in(wire_d61_49),.data_out(wire_d61_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6206151(.data_in(wire_d61_50),.data_out(wire_d61_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6206152(.data_in(wire_d61_51),.data_out(wire_d61_52),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6206153(.data_in(wire_d61_52),.data_out(wire_d61_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6206154(.data_in(wire_d61_53),.data_out(wire_d61_54),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6206155(.data_in(wire_d61_54),.data_out(wire_d61_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6206156(.data_in(wire_d61_55),.data_out(wire_d61_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6206157(.data_in(wire_d61_56),.data_out(wire_d61_57),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6206158(.data_in(wire_d61_57),.data_out(wire_d61_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6206159(.data_in(wire_d61_58),.data_out(wire_d61_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6206160(.data_in(wire_d61_59),.data_out(wire_d61_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6206161(.data_in(wire_d61_60),.data_out(wire_d61_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6206162(.data_in(wire_d61_61),.data_out(wire_d61_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6206163(.data_in(wire_d61_62),.data_out(wire_d61_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6206164(.data_in(wire_d61_63),.data_out(wire_d61_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6206165(.data_in(wire_d61_64),.data_out(wire_d61_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6206166(.data_in(wire_d61_65),.data_out(wire_d61_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6206167(.data_in(wire_d61_66),.data_out(wire_d61_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6206168(.data_in(wire_d61_67),.data_out(wire_d61_68),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6206169(.data_in(wire_d61_68),.data_out(wire_d61_69),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6206170(.data_in(wire_d61_69),.data_out(wire_d61_70),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6206171(.data_in(wire_d61_70),.data_out(wire_d61_71),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6206172(.data_in(wire_d61_71),.data_out(wire_d61_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6206173(.data_in(wire_d61_72),.data_out(wire_d61_73),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6206174(.data_in(wire_d61_73),.data_out(wire_d61_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6206175(.data_in(wire_d61_74),.data_out(wire_d61_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6206176(.data_in(wire_d61_75),.data_out(wire_d61_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6206177(.data_in(wire_d61_76),.data_out(wire_d61_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6206178(.data_in(wire_d61_77),.data_out(wire_d61_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6206179(.data_in(wire_d61_78),.data_out(wire_d61_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6206180(.data_in(wire_d61_79),.data_out(wire_d61_80),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6206181(.data_in(wire_d61_80),.data_out(wire_d61_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6206182(.data_in(wire_d61_81),.data_out(wire_d61_82),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6206183(.data_in(wire_d61_82),.data_out(wire_d61_83),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6206184(.data_in(wire_d61_83),.data_out(wire_d61_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6206185(.data_in(wire_d61_84),.data_out(wire_d61_85),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6206186(.data_in(wire_d61_85),.data_out(wire_d61_86),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6206187(.data_in(wire_d61_86),.data_out(wire_d61_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6206188(.data_in(wire_d61_87),.data_out(wire_d61_88),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6206189(.data_in(wire_d61_88),.data_out(wire_d61_89),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6206190(.data_in(wire_d61_89),.data_out(wire_d61_90),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6206191(.data_in(wire_d61_90),.data_out(wire_d61_91),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6206192(.data_in(wire_d61_91),.data_out(wire_d61_92),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6206193(.data_in(wire_d61_92),.data_out(wire_d61_93),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6206194(.data_in(wire_d61_93),.data_out(wire_d61_94),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6206195(.data_in(wire_d61_94),.data_out(wire_d61_95),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6206196(.data_in(wire_d61_95),.data_out(wire_d61_96),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6206197(.data_in(wire_d61_96),.data_out(wire_d61_97),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6206198(.data_in(wire_d61_97),.data_out(wire_d61_98),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6206199(.data_in(wire_d61_98),.data_out(wire_d61_99),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance62061100(.data_in(wire_d61_99),.data_out(wire_d61_100),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance62061101(.data_in(wire_d61_100),.data_out(wire_d61_101),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance62061102(.data_in(wire_d61_101),.data_out(wire_d61_102),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance62061103(.data_in(wire_d61_102),.data_out(wire_d61_103),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance62061104(.data_in(wire_d61_103),.data_out(wire_d61_104),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance62061105(.data_in(wire_d61_104),.data_out(wire_d61_105),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance62061106(.data_in(wire_d61_105),.data_out(wire_d61_106),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance62061107(.data_in(wire_d61_106),.data_out(wire_d61_107),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance62061108(.data_in(wire_d61_107),.data_out(wire_d61_108),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance62061109(.data_in(wire_d61_108),.data_out(wire_d61_109),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance62061110(.data_in(wire_d61_109),.data_out(wire_d61_110),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance62061111(.data_in(wire_d61_110),.data_out(wire_d61_111),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance62061112(.data_in(wire_d61_111),.data_out(wire_d61_112),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance62061113(.data_in(wire_d61_112),.data_out(wire_d61_113),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance62061114(.data_in(wire_d61_113),.data_out(wire_d61_114),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance62061115(.data_in(wire_d61_114),.data_out(wire_d61_115),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance62061116(.data_in(wire_d61_115),.data_out(wire_d61_116),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance62061117(.data_in(wire_d61_116),.data_out(wire_d61_117),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance62061118(.data_in(wire_d61_117),.data_out(wire_d61_118),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance62061119(.data_in(wire_d61_118),.data_out(d_out61),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance630620(.data_in(d_in62),.data_out(wire_d62_0),.clk(clk),.rst(rst));            //channel 63
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance630621(.data_in(wire_d62_0),.data_out(wire_d62_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance630622(.data_in(wire_d62_1),.data_out(wire_d62_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance630623(.data_in(wire_d62_2),.data_out(wire_d62_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance630624(.data_in(wire_d62_3),.data_out(wire_d62_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance630625(.data_in(wire_d62_4),.data_out(wire_d62_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance630626(.data_in(wire_d62_5),.data_out(wire_d62_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance630627(.data_in(wire_d62_6),.data_out(wire_d62_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance630628(.data_in(wire_d62_7),.data_out(wire_d62_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance630629(.data_in(wire_d62_8),.data_out(wire_d62_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6306210(.data_in(wire_d62_9),.data_out(wire_d62_10),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6306211(.data_in(wire_d62_10),.data_out(wire_d62_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6306212(.data_in(wire_d62_11),.data_out(wire_d62_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6306213(.data_in(wire_d62_12),.data_out(wire_d62_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6306214(.data_in(wire_d62_13),.data_out(wire_d62_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6306215(.data_in(wire_d62_14),.data_out(wire_d62_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6306216(.data_in(wire_d62_15),.data_out(wire_d62_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6306217(.data_in(wire_d62_16),.data_out(wire_d62_17),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6306218(.data_in(wire_d62_17),.data_out(wire_d62_18),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6306219(.data_in(wire_d62_18),.data_out(wire_d62_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6306220(.data_in(wire_d62_19),.data_out(wire_d62_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6306221(.data_in(wire_d62_20),.data_out(wire_d62_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6306222(.data_in(wire_d62_21),.data_out(wire_d62_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6306223(.data_in(wire_d62_22),.data_out(wire_d62_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6306224(.data_in(wire_d62_23),.data_out(wire_d62_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6306225(.data_in(wire_d62_24),.data_out(wire_d62_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6306226(.data_in(wire_d62_25),.data_out(wire_d62_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6306227(.data_in(wire_d62_26),.data_out(wire_d62_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6306228(.data_in(wire_d62_27),.data_out(wire_d62_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6306229(.data_in(wire_d62_28),.data_out(wire_d62_29),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6306230(.data_in(wire_d62_29),.data_out(wire_d62_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6306231(.data_in(wire_d62_30),.data_out(wire_d62_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6306232(.data_in(wire_d62_31),.data_out(wire_d62_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6306233(.data_in(wire_d62_32),.data_out(wire_d62_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6306234(.data_in(wire_d62_33),.data_out(wire_d62_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6306235(.data_in(wire_d62_34),.data_out(wire_d62_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6306236(.data_in(wire_d62_35),.data_out(wire_d62_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6306237(.data_in(wire_d62_36),.data_out(wire_d62_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6306238(.data_in(wire_d62_37),.data_out(wire_d62_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6306239(.data_in(wire_d62_38),.data_out(wire_d62_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6306240(.data_in(wire_d62_39),.data_out(wire_d62_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6306241(.data_in(wire_d62_40),.data_out(wire_d62_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6306242(.data_in(wire_d62_41),.data_out(wire_d62_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6306243(.data_in(wire_d62_42),.data_out(wire_d62_43),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6306244(.data_in(wire_d62_43),.data_out(wire_d62_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6306245(.data_in(wire_d62_44),.data_out(wire_d62_45),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6306246(.data_in(wire_d62_45),.data_out(wire_d62_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6306247(.data_in(wire_d62_46),.data_out(wire_d62_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6306248(.data_in(wire_d62_47),.data_out(wire_d62_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6306249(.data_in(wire_d62_48),.data_out(wire_d62_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6306250(.data_in(wire_d62_49),.data_out(wire_d62_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6306251(.data_in(wire_d62_50),.data_out(wire_d62_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6306252(.data_in(wire_d62_51),.data_out(wire_d62_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6306253(.data_in(wire_d62_52),.data_out(wire_d62_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6306254(.data_in(wire_d62_53),.data_out(wire_d62_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6306255(.data_in(wire_d62_54),.data_out(wire_d62_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6306256(.data_in(wire_d62_55),.data_out(wire_d62_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6306257(.data_in(wire_d62_56),.data_out(wire_d62_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6306258(.data_in(wire_d62_57),.data_out(wire_d62_58),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6306259(.data_in(wire_d62_58),.data_out(wire_d62_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6306260(.data_in(wire_d62_59),.data_out(wire_d62_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6306261(.data_in(wire_d62_60),.data_out(wire_d62_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6306262(.data_in(wire_d62_61),.data_out(wire_d62_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6306263(.data_in(wire_d62_62),.data_out(wire_d62_63),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6306264(.data_in(wire_d62_63),.data_out(wire_d62_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6306265(.data_in(wire_d62_64),.data_out(wire_d62_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6306266(.data_in(wire_d62_65),.data_out(wire_d62_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6306267(.data_in(wire_d62_66),.data_out(wire_d62_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6306268(.data_in(wire_d62_67),.data_out(wire_d62_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6306269(.data_in(wire_d62_68),.data_out(wire_d62_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6306270(.data_in(wire_d62_69),.data_out(wire_d62_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6306271(.data_in(wire_d62_70),.data_out(wire_d62_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6306272(.data_in(wire_d62_71),.data_out(wire_d62_72),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6306273(.data_in(wire_d62_72),.data_out(wire_d62_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6306274(.data_in(wire_d62_73),.data_out(wire_d62_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6306275(.data_in(wire_d62_74),.data_out(wire_d62_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6306276(.data_in(wire_d62_75),.data_out(wire_d62_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6306277(.data_in(wire_d62_76),.data_out(wire_d62_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6306278(.data_in(wire_d62_77),.data_out(wire_d62_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6306279(.data_in(wire_d62_78),.data_out(wire_d62_79),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6306280(.data_in(wire_d62_79),.data_out(wire_d62_80),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6306281(.data_in(wire_d62_80),.data_out(wire_d62_81),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6306282(.data_in(wire_d62_81),.data_out(wire_d62_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6306283(.data_in(wire_d62_82),.data_out(wire_d62_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6306284(.data_in(wire_d62_83),.data_out(wire_d62_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6306285(.data_in(wire_d62_84),.data_out(wire_d62_85),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6306286(.data_in(wire_d62_85),.data_out(wire_d62_86),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6306287(.data_in(wire_d62_86),.data_out(wire_d62_87),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6306288(.data_in(wire_d62_87),.data_out(wire_d62_88),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6306289(.data_in(wire_d62_88),.data_out(wire_d62_89),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6306290(.data_in(wire_d62_89),.data_out(wire_d62_90),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6306291(.data_in(wire_d62_90),.data_out(wire_d62_91),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6306292(.data_in(wire_d62_91),.data_out(wire_d62_92),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6306293(.data_in(wire_d62_92),.data_out(wire_d62_93),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6306294(.data_in(wire_d62_93),.data_out(wire_d62_94),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6306295(.data_in(wire_d62_94),.data_out(wire_d62_95),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6306296(.data_in(wire_d62_95),.data_out(wire_d62_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6306297(.data_in(wire_d62_96),.data_out(wire_d62_97),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6306298(.data_in(wire_d62_97),.data_out(wire_d62_98),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6306299(.data_in(wire_d62_98),.data_out(wire_d62_99),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance63062100(.data_in(wire_d62_99),.data_out(wire_d62_100),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance63062101(.data_in(wire_d62_100),.data_out(wire_d62_101),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance63062102(.data_in(wire_d62_101),.data_out(wire_d62_102),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance63062103(.data_in(wire_d62_102),.data_out(wire_d62_103),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance63062104(.data_in(wire_d62_103),.data_out(wire_d62_104),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance63062105(.data_in(wire_d62_104),.data_out(wire_d62_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance63062106(.data_in(wire_d62_105),.data_out(wire_d62_106),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance63062107(.data_in(wire_d62_106),.data_out(wire_d62_107),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance63062108(.data_in(wire_d62_107),.data_out(wire_d62_108),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance63062109(.data_in(wire_d62_108),.data_out(wire_d62_109),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance63062110(.data_in(wire_d62_109),.data_out(wire_d62_110),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance63062111(.data_in(wire_d62_110),.data_out(wire_d62_111),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance63062112(.data_in(wire_d62_111),.data_out(wire_d62_112),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance63062113(.data_in(wire_d62_112),.data_out(wire_d62_113),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance63062114(.data_in(wire_d62_113),.data_out(wire_d62_114),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance63062115(.data_in(wire_d62_114),.data_out(wire_d62_115),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance63062116(.data_in(wire_d62_115),.data_out(wire_d62_116),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance63062117(.data_in(wire_d62_116),.data_out(wire_d62_117),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance63062118(.data_in(wire_d62_117),.data_out(wire_d62_118),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance63062119(.data_in(wire_d62_118),.data_out(d_out62),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance640630(.data_in(d_in63),.data_out(wire_d63_0),.clk(clk),.rst(rst));            //channel 64
	decoder_top #(.WIDTH(WIDTH)) decoder_instance640631(.data_in(wire_d63_0),.data_out(wire_d63_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance640632(.data_in(wire_d63_1),.data_out(wire_d63_2),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance640633(.data_in(wire_d63_2),.data_out(wire_d63_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance640634(.data_in(wire_d63_3),.data_out(wire_d63_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance640635(.data_in(wire_d63_4),.data_out(wire_d63_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance640636(.data_in(wire_d63_5),.data_out(wire_d63_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance640637(.data_in(wire_d63_6),.data_out(wire_d63_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance640638(.data_in(wire_d63_7),.data_out(wire_d63_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance640639(.data_in(wire_d63_8),.data_out(wire_d63_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6406310(.data_in(wire_d63_9),.data_out(wire_d63_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6406311(.data_in(wire_d63_10),.data_out(wire_d63_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6406312(.data_in(wire_d63_11),.data_out(wire_d63_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6406313(.data_in(wire_d63_12),.data_out(wire_d63_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6406314(.data_in(wire_d63_13),.data_out(wire_d63_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6406315(.data_in(wire_d63_14),.data_out(wire_d63_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6406316(.data_in(wire_d63_15),.data_out(wire_d63_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6406317(.data_in(wire_d63_16),.data_out(wire_d63_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6406318(.data_in(wire_d63_17),.data_out(wire_d63_18),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6406319(.data_in(wire_d63_18),.data_out(wire_d63_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6406320(.data_in(wire_d63_19),.data_out(wire_d63_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6406321(.data_in(wire_d63_20),.data_out(wire_d63_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6406322(.data_in(wire_d63_21),.data_out(wire_d63_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6406323(.data_in(wire_d63_22),.data_out(wire_d63_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6406324(.data_in(wire_d63_23),.data_out(wire_d63_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6406325(.data_in(wire_d63_24),.data_out(wire_d63_25),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6406326(.data_in(wire_d63_25),.data_out(wire_d63_26),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6406327(.data_in(wire_d63_26),.data_out(wire_d63_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6406328(.data_in(wire_d63_27),.data_out(wire_d63_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6406329(.data_in(wire_d63_28),.data_out(wire_d63_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6406330(.data_in(wire_d63_29),.data_out(wire_d63_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6406331(.data_in(wire_d63_30),.data_out(wire_d63_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6406332(.data_in(wire_d63_31),.data_out(wire_d63_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6406333(.data_in(wire_d63_32),.data_out(wire_d63_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6406334(.data_in(wire_d63_33),.data_out(wire_d63_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6406335(.data_in(wire_d63_34),.data_out(wire_d63_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6406336(.data_in(wire_d63_35),.data_out(wire_d63_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6406337(.data_in(wire_d63_36),.data_out(wire_d63_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6406338(.data_in(wire_d63_37),.data_out(wire_d63_38),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6406339(.data_in(wire_d63_38),.data_out(wire_d63_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6406340(.data_in(wire_d63_39),.data_out(wire_d63_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6406341(.data_in(wire_d63_40),.data_out(wire_d63_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6406342(.data_in(wire_d63_41),.data_out(wire_d63_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6406343(.data_in(wire_d63_42),.data_out(wire_d63_43),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6406344(.data_in(wire_d63_43),.data_out(wire_d63_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6406345(.data_in(wire_d63_44),.data_out(wire_d63_45),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6406346(.data_in(wire_d63_45),.data_out(wire_d63_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6406347(.data_in(wire_d63_46),.data_out(wire_d63_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6406348(.data_in(wire_d63_47),.data_out(wire_d63_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6406349(.data_in(wire_d63_48),.data_out(wire_d63_49),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6406350(.data_in(wire_d63_49),.data_out(wire_d63_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6406351(.data_in(wire_d63_50),.data_out(wire_d63_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6406352(.data_in(wire_d63_51),.data_out(wire_d63_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6406353(.data_in(wire_d63_52),.data_out(wire_d63_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6406354(.data_in(wire_d63_53),.data_out(wire_d63_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6406355(.data_in(wire_d63_54),.data_out(wire_d63_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6406356(.data_in(wire_d63_55),.data_out(wire_d63_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6406357(.data_in(wire_d63_56),.data_out(wire_d63_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6406358(.data_in(wire_d63_57),.data_out(wire_d63_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6406359(.data_in(wire_d63_58),.data_out(wire_d63_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6406360(.data_in(wire_d63_59),.data_out(wire_d63_60),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6406361(.data_in(wire_d63_60),.data_out(wire_d63_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6406362(.data_in(wire_d63_61),.data_out(wire_d63_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6406363(.data_in(wire_d63_62),.data_out(wire_d63_63),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6406364(.data_in(wire_d63_63),.data_out(wire_d63_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6406365(.data_in(wire_d63_64),.data_out(wire_d63_65),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6406366(.data_in(wire_d63_65),.data_out(wire_d63_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6406367(.data_in(wire_d63_66),.data_out(wire_d63_67),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6406368(.data_in(wire_d63_67),.data_out(wire_d63_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6406369(.data_in(wire_d63_68),.data_out(wire_d63_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6406370(.data_in(wire_d63_69),.data_out(wire_d63_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6406371(.data_in(wire_d63_70),.data_out(wire_d63_71),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6406372(.data_in(wire_d63_71),.data_out(wire_d63_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6406373(.data_in(wire_d63_72),.data_out(wire_d63_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6406374(.data_in(wire_d63_73),.data_out(wire_d63_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6406375(.data_in(wire_d63_74),.data_out(wire_d63_75),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6406376(.data_in(wire_d63_75),.data_out(wire_d63_76),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6406377(.data_in(wire_d63_76),.data_out(wire_d63_77),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6406378(.data_in(wire_d63_77),.data_out(wire_d63_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6406379(.data_in(wire_d63_78),.data_out(wire_d63_79),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6406380(.data_in(wire_d63_79),.data_out(wire_d63_80),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6406381(.data_in(wire_d63_80),.data_out(wire_d63_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6406382(.data_in(wire_d63_81),.data_out(wire_d63_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6406383(.data_in(wire_d63_82),.data_out(wire_d63_83),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6406384(.data_in(wire_d63_83),.data_out(wire_d63_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6406385(.data_in(wire_d63_84),.data_out(wire_d63_85),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6406386(.data_in(wire_d63_85),.data_out(wire_d63_86),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6406387(.data_in(wire_d63_86),.data_out(wire_d63_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6406388(.data_in(wire_d63_87),.data_out(wire_d63_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6406389(.data_in(wire_d63_88),.data_out(wire_d63_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6406390(.data_in(wire_d63_89),.data_out(wire_d63_90),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6406391(.data_in(wire_d63_90),.data_out(wire_d63_91),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6406392(.data_in(wire_d63_91),.data_out(wire_d63_92),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6406393(.data_in(wire_d63_92),.data_out(wire_d63_93),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6406394(.data_in(wire_d63_93),.data_out(wire_d63_94),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6406395(.data_in(wire_d63_94),.data_out(wire_d63_95),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6406396(.data_in(wire_d63_95),.data_out(wire_d63_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6406397(.data_in(wire_d63_96),.data_out(wire_d63_97),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6406398(.data_in(wire_d63_97),.data_out(wire_d63_98),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6406399(.data_in(wire_d63_98),.data_out(wire_d63_99),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance64063100(.data_in(wire_d63_99),.data_out(wire_d63_100),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance64063101(.data_in(wire_d63_100),.data_out(wire_d63_101),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance64063102(.data_in(wire_d63_101),.data_out(wire_d63_102),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance64063103(.data_in(wire_d63_102),.data_out(wire_d63_103),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance64063104(.data_in(wire_d63_103),.data_out(wire_d63_104),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance64063105(.data_in(wire_d63_104),.data_out(wire_d63_105),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance64063106(.data_in(wire_d63_105),.data_out(wire_d63_106),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance64063107(.data_in(wire_d63_106),.data_out(wire_d63_107),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance64063108(.data_in(wire_d63_107),.data_out(wire_d63_108),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance64063109(.data_in(wire_d63_108),.data_out(wire_d63_109),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance64063110(.data_in(wire_d63_109),.data_out(wire_d63_110),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance64063111(.data_in(wire_d63_110),.data_out(wire_d63_111),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance64063112(.data_in(wire_d63_111),.data_out(wire_d63_112),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance64063113(.data_in(wire_d63_112),.data_out(wire_d63_113),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance64063114(.data_in(wire_d63_113),.data_out(wire_d63_114),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance64063115(.data_in(wire_d63_114),.data_out(wire_d63_115),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance64063116(.data_in(wire_d63_115),.data_out(wire_d63_116),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance64063117(.data_in(wire_d63_116),.data_out(wire_d63_117),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance64063118(.data_in(wire_d63_117),.data_out(wire_d63_118),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance64063119(.data_in(wire_d63_118),.data_out(d_out63),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance650640(.data_in(d_in64),.data_out(wire_d64_0),.clk(clk),.rst(rst));            //channel 65
	invertion #(.WIDTH(WIDTH)) invertion_instance650641(.data_in(wire_d64_0),.data_out(wire_d64_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance650642(.data_in(wire_d64_1),.data_out(wire_d64_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance650643(.data_in(wire_d64_2),.data_out(wire_d64_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance650644(.data_in(wire_d64_3),.data_out(wire_d64_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance650645(.data_in(wire_d64_4),.data_out(wire_d64_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance650646(.data_in(wire_d64_5),.data_out(wire_d64_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance650647(.data_in(wire_d64_6),.data_out(wire_d64_7),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance650648(.data_in(wire_d64_7),.data_out(wire_d64_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance650649(.data_in(wire_d64_8),.data_out(wire_d64_9),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6506410(.data_in(wire_d64_9),.data_out(wire_d64_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6506411(.data_in(wire_d64_10),.data_out(wire_d64_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6506412(.data_in(wire_d64_11),.data_out(wire_d64_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6506413(.data_in(wire_d64_12),.data_out(wire_d64_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6506414(.data_in(wire_d64_13),.data_out(wire_d64_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6506415(.data_in(wire_d64_14),.data_out(wire_d64_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6506416(.data_in(wire_d64_15),.data_out(wire_d64_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6506417(.data_in(wire_d64_16),.data_out(wire_d64_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6506418(.data_in(wire_d64_17),.data_out(wire_d64_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6506419(.data_in(wire_d64_18),.data_out(wire_d64_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6506420(.data_in(wire_d64_19),.data_out(wire_d64_20),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6506421(.data_in(wire_d64_20),.data_out(wire_d64_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6506422(.data_in(wire_d64_21),.data_out(wire_d64_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6506423(.data_in(wire_d64_22),.data_out(wire_d64_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6506424(.data_in(wire_d64_23),.data_out(wire_d64_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6506425(.data_in(wire_d64_24),.data_out(wire_d64_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6506426(.data_in(wire_d64_25),.data_out(wire_d64_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6506427(.data_in(wire_d64_26),.data_out(wire_d64_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6506428(.data_in(wire_d64_27),.data_out(wire_d64_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6506429(.data_in(wire_d64_28),.data_out(wire_d64_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6506430(.data_in(wire_d64_29),.data_out(wire_d64_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6506431(.data_in(wire_d64_30),.data_out(wire_d64_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6506432(.data_in(wire_d64_31),.data_out(wire_d64_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6506433(.data_in(wire_d64_32),.data_out(wire_d64_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6506434(.data_in(wire_d64_33),.data_out(wire_d64_34),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6506435(.data_in(wire_d64_34),.data_out(wire_d64_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6506436(.data_in(wire_d64_35),.data_out(wire_d64_36),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6506437(.data_in(wire_d64_36),.data_out(wire_d64_37),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6506438(.data_in(wire_d64_37),.data_out(wire_d64_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6506439(.data_in(wire_d64_38),.data_out(wire_d64_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6506440(.data_in(wire_d64_39),.data_out(wire_d64_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6506441(.data_in(wire_d64_40),.data_out(wire_d64_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6506442(.data_in(wire_d64_41),.data_out(wire_d64_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6506443(.data_in(wire_d64_42),.data_out(wire_d64_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6506444(.data_in(wire_d64_43),.data_out(wire_d64_44),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6506445(.data_in(wire_d64_44),.data_out(wire_d64_45),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6506446(.data_in(wire_d64_45),.data_out(wire_d64_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6506447(.data_in(wire_d64_46),.data_out(wire_d64_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6506448(.data_in(wire_d64_47),.data_out(wire_d64_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6506449(.data_in(wire_d64_48),.data_out(wire_d64_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6506450(.data_in(wire_d64_49),.data_out(wire_d64_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6506451(.data_in(wire_d64_50),.data_out(wire_d64_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6506452(.data_in(wire_d64_51),.data_out(wire_d64_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6506453(.data_in(wire_d64_52),.data_out(wire_d64_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6506454(.data_in(wire_d64_53),.data_out(wire_d64_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6506455(.data_in(wire_d64_54),.data_out(wire_d64_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6506456(.data_in(wire_d64_55),.data_out(wire_d64_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6506457(.data_in(wire_d64_56),.data_out(wire_d64_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6506458(.data_in(wire_d64_57),.data_out(wire_d64_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6506459(.data_in(wire_d64_58),.data_out(wire_d64_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6506460(.data_in(wire_d64_59),.data_out(wire_d64_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6506461(.data_in(wire_d64_60),.data_out(wire_d64_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6506462(.data_in(wire_d64_61),.data_out(wire_d64_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6506463(.data_in(wire_d64_62),.data_out(wire_d64_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6506464(.data_in(wire_d64_63),.data_out(wire_d64_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6506465(.data_in(wire_d64_64),.data_out(wire_d64_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6506466(.data_in(wire_d64_65),.data_out(wire_d64_66),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6506467(.data_in(wire_d64_66),.data_out(wire_d64_67),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6506468(.data_in(wire_d64_67),.data_out(wire_d64_68),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6506469(.data_in(wire_d64_68),.data_out(wire_d64_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6506470(.data_in(wire_d64_69),.data_out(wire_d64_70),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6506471(.data_in(wire_d64_70),.data_out(wire_d64_71),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6506472(.data_in(wire_d64_71),.data_out(wire_d64_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6506473(.data_in(wire_d64_72),.data_out(wire_d64_73),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6506474(.data_in(wire_d64_73),.data_out(wire_d64_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6506475(.data_in(wire_d64_74),.data_out(wire_d64_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6506476(.data_in(wire_d64_75),.data_out(wire_d64_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6506477(.data_in(wire_d64_76),.data_out(wire_d64_77),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6506478(.data_in(wire_d64_77),.data_out(wire_d64_78),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6506479(.data_in(wire_d64_78),.data_out(wire_d64_79),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6506480(.data_in(wire_d64_79),.data_out(wire_d64_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6506481(.data_in(wire_d64_80),.data_out(wire_d64_81),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6506482(.data_in(wire_d64_81),.data_out(wire_d64_82),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6506483(.data_in(wire_d64_82),.data_out(wire_d64_83),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6506484(.data_in(wire_d64_83),.data_out(wire_d64_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6506485(.data_in(wire_d64_84),.data_out(wire_d64_85),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6506486(.data_in(wire_d64_85),.data_out(wire_d64_86),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6506487(.data_in(wire_d64_86),.data_out(wire_d64_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6506488(.data_in(wire_d64_87),.data_out(wire_d64_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6506489(.data_in(wire_d64_88),.data_out(wire_d64_89),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6506490(.data_in(wire_d64_89),.data_out(wire_d64_90),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6506491(.data_in(wire_d64_90),.data_out(wire_d64_91),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6506492(.data_in(wire_d64_91),.data_out(wire_d64_92),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6506493(.data_in(wire_d64_92),.data_out(wire_d64_93),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6506494(.data_in(wire_d64_93),.data_out(wire_d64_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6506495(.data_in(wire_d64_94),.data_out(wire_d64_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6506496(.data_in(wire_d64_95),.data_out(wire_d64_96),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6506497(.data_in(wire_d64_96),.data_out(wire_d64_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6506498(.data_in(wire_d64_97),.data_out(wire_d64_98),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6506499(.data_in(wire_d64_98),.data_out(wire_d64_99),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65064100(.data_in(wire_d64_99),.data_out(wire_d64_100),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance65064101(.data_in(wire_d64_100),.data_out(wire_d64_101),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance65064102(.data_in(wire_d64_101),.data_out(wire_d64_102),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance65064103(.data_in(wire_d64_102),.data_out(wire_d64_103),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance65064104(.data_in(wire_d64_103),.data_out(wire_d64_104),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance65064105(.data_in(wire_d64_104),.data_out(wire_d64_105),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance65064106(.data_in(wire_d64_105),.data_out(wire_d64_106),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance65064107(.data_in(wire_d64_106),.data_out(wire_d64_107),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance65064108(.data_in(wire_d64_107),.data_out(wire_d64_108),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance65064109(.data_in(wire_d64_108),.data_out(wire_d64_109),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance65064110(.data_in(wire_d64_109),.data_out(wire_d64_110),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance65064111(.data_in(wire_d64_110),.data_out(wire_d64_111),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance65064112(.data_in(wire_d64_111),.data_out(wire_d64_112),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance65064113(.data_in(wire_d64_112),.data_out(wire_d64_113),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance65064114(.data_in(wire_d64_113),.data_out(wire_d64_114),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance65064115(.data_in(wire_d64_114),.data_out(wire_d64_115),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance65064116(.data_in(wire_d64_115),.data_out(wire_d64_116),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance65064117(.data_in(wire_d64_116),.data_out(wire_d64_117),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance65064118(.data_in(wire_d64_117),.data_out(wire_d64_118),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance65064119(.data_in(wire_d64_118),.data_out(d_out64),.clk(clk),.rst(rst));

	large_adder #(.WIDTH(WIDTH)) large_adder_instance660650(.data_in(d_in65),.data_out(wire_d65_0),.clk(clk),.rst(rst));            //channel 66
	register #(.WIDTH(WIDTH)) register_instance660651(.data_in(wire_d65_0),.data_out(wire_d65_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance660652(.data_in(wire_d65_1),.data_out(wire_d65_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance660653(.data_in(wire_d65_2),.data_out(wire_d65_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance660654(.data_in(wire_d65_3),.data_out(wire_d65_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance660655(.data_in(wire_d65_4),.data_out(wire_d65_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance660656(.data_in(wire_d65_5),.data_out(wire_d65_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance660657(.data_in(wire_d65_6),.data_out(wire_d65_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance660658(.data_in(wire_d65_7),.data_out(wire_d65_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance660659(.data_in(wire_d65_8),.data_out(wire_d65_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6606510(.data_in(wire_d65_9),.data_out(wire_d65_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6606511(.data_in(wire_d65_10),.data_out(wire_d65_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6606512(.data_in(wire_d65_11),.data_out(wire_d65_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6606513(.data_in(wire_d65_12),.data_out(wire_d65_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6606514(.data_in(wire_d65_13),.data_out(wire_d65_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6606515(.data_in(wire_d65_14),.data_out(wire_d65_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6606516(.data_in(wire_d65_15),.data_out(wire_d65_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6606517(.data_in(wire_d65_16),.data_out(wire_d65_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6606518(.data_in(wire_d65_17),.data_out(wire_d65_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6606519(.data_in(wire_d65_18),.data_out(wire_d65_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6606520(.data_in(wire_d65_19),.data_out(wire_d65_20),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6606521(.data_in(wire_d65_20),.data_out(wire_d65_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6606522(.data_in(wire_d65_21),.data_out(wire_d65_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6606523(.data_in(wire_d65_22),.data_out(wire_d65_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6606524(.data_in(wire_d65_23),.data_out(wire_d65_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6606525(.data_in(wire_d65_24),.data_out(wire_d65_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6606526(.data_in(wire_d65_25),.data_out(wire_d65_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6606527(.data_in(wire_d65_26),.data_out(wire_d65_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6606528(.data_in(wire_d65_27),.data_out(wire_d65_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6606529(.data_in(wire_d65_28),.data_out(wire_d65_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6606530(.data_in(wire_d65_29),.data_out(wire_d65_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6606531(.data_in(wire_d65_30),.data_out(wire_d65_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6606532(.data_in(wire_d65_31),.data_out(wire_d65_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6606533(.data_in(wire_d65_32),.data_out(wire_d65_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6606534(.data_in(wire_d65_33),.data_out(wire_d65_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6606535(.data_in(wire_d65_34),.data_out(wire_d65_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6606536(.data_in(wire_d65_35),.data_out(wire_d65_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6606537(.data_in(wire_d65_36),.data_out(wire_d65_37),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6606538(.data_in(wire_d65_37),.data_out(wire_d65_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6606539(.data_in(wire_d65_38),.data_out(wire_d65_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6606540(.data_in(wire_d65_39),.data_out(wire_d65_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6606541(.data_in(wire_d65_40),.data_out(wire_d65_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6606542(.data_in(wire_d65_41),.data_out(wire_d65_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6606543(.data_in(wire_d65_42),.data_out(wire_d65_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6606544(.data_in(wire_d65_43),.data_out(wire_d65_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6606545(.data_in(wire_d65_44),.data_out(wire_d65_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6606546(.data_in(wire_d65_45),.data_out(wire_d65_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6606547(.data_in(wire_d65_46),.data_out(wire_d65_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6606548(.data_in(wire_d65_47),.data_out(wire_d65_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6606549(.data_in(wire_d65_48),.data_out(wire_d65_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6606550(.data_in(wire_d65_49),.data_out(wire_d65_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6606551(.data_in(wire_d65_50),.data_out(wire_d65_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6606552(.data_in(wire_d65_51),.data_out(wire_d65_52),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6606553(.data_in(wire_d65_52),.data_out(wire_d65_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6606554(.data_in(wire_d65_53),.data_out(wire_d65_54),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6606555(.data_in(wire_d65_54),.data_out(wire_d65_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6606556(.data_in(wire_d65_55),.data_out(wire_d65_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6606557(.data_in(wire_d65_56),.data_out(wire_d65_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6606558(.data_in(wire_d65_57),.data_out(wire_d65_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6606559(.data_in(wire_d65_58),.data_out(wire_d65_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6606560(.data_in(wire_d65_59),.data_out(wire_d65_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6606561(.data_in(wire_d65_60),.data_out(wire_d65_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6606562(.data_in(wire_d65_61),.data_out(wire_d65_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6606563(.data_in(wire_d65_62),.data_out(wire_d65_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6606564(.data_in(wire_d65_63),.data_out(wire_d65_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6606565(.data_in(wire_d65_64),.data_out(wire_d65_65),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6606566(.data_in(wire_d65_65),.data_out(wire_d65_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6606567(.data_in(wire_d65_66),.data_out(wire_d65_67),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6606568(.data_in(wire_d65_67),.data_out(wire_d65_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6606569(.data_in(wire_d65_68),.data_out(wire_d65_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6606570(.data_in(wire_d65_69),.data_out(wire_d65_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6606571(.data_in(wire_d65_70),.data_out(wire_d65_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6606572(.data_in(wire_d65_71),.data_out(wire_d65_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6606573(.data_in(wire_d65_72),.data_out(wire_d65_73),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6606574(.data_in(wire_d65_73),.data_out(wire_d65_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6606575(.data_in(wire_d65_74),.data_out(wire_d65_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6606576(.data_in(wire_d65_75),.data_out(wire_d65_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6606577(.data_in(wire_d65_76),.data_out(wire_d65_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6606578(.data_in(wire_d65_77),.data_out(wire_d65_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6606579(.data_in(wire_d65_78),.data_out(wire_d65_79),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6606580(.data_in(wire_d65_79),.data_out(wire_d65_80),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6606581(.data_in(wire_d65_80),.data_out(wire_d65_81),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6606582(.data_in(wire_d65_81),.data_out(wire_d65_82),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6606583(.data_in(wire_d65_82),.data_out(wire_d65_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6606584(.data_in(wire_d65_83),.data_out(wire_d65_84),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6606585(.data_in(wire_d65_84),.data_out(wire_d65_85),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6606586(.data_in(wire_d65_85),.data_out(wire_d65_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6606587(.data_in(wire_d65_86),.data_out(wire_d65_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6606588(.data_in(wire_d65_87),.data_out(wire_d65_88),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6606589(.data_in(wire_d65_88),.data_out(wire_d65_89),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6606590(.data_in(wire_d65_89),.data_out(wire_d65_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6606591(.data_in(wire_d65_90),.data_out(wire_d65_91),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6606592(.data_in(wire_d65_91),.data_out(wire_d65_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6606593(.data_in(wire_d65_92),.data_out(wire_d65_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6606594(.data_in(wire_d65_93),.data_out(wire_d65_94),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6606595(.data_in(wire_d65_94),.data_out(wire_d65_95),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6606596(.data_in(wire_d65_95),.data_out(wire_d65_96),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6606597(.data_in(wire_d65_96),.data_out(wire_d65_97),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6606598(.data_in(wire_d65_97),.data_out(wire_d65_98),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6606599(.data_in(wire_d65_98),.data_out(wire_d65_99),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance66065100(.data_in(wire_d65_99),.data_out(wire_d65_100),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance66065101(.data_in(wire_d65_100),.data_out(wire_d65_101),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance66065102(.data_in(wire_d65_101),.data_out(wire_d65_102),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance66065103(.data_in(wire_d65_102),.data_out(wire_d65_103),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance66065104(.data_in(wire_d65_103),.data_out(wire_d65_104),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance66065105(.data_in(wire_d65_104),.data_out(wire_d65_105),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance66065106(.data_in(wire_d65_105),.data_out(wire_d65_106),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance66065107(.data_in(wire_d65_106),.data_out(wire_d65_107),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance66065108(.data_in(wire_d65_107),.data_out(wire_d65_108),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance66065109(.data_in(wire_d65_108),.data_out(wire_d65_109),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance66065110(.data_in(wire_d65_109),.data_out(wire_d65_110),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance66065111(.data_in(wire_d65_110),.data_out(wire_d65_111),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance66065112(.data_in(wire_d65_111),.data_out(wire_d65_112),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance66065113(.data_in(wire_d65_112),.data_out(wire_d65_113),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance66065114(.data_in(wire_d65_113),.data_out(wire_d65_114),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance66065115(.data_in(wire_d65_114),.data_out(wire_d65_115),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance66065116(.data_in(wire_d65_115),.data_out(wire_d65_116),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance66065117(.data_in(wire_d65_116),.data_out(wire_d65_117),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance66065118(.data_in(wire_d65_117),.data_out(wire_d65_118),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance66065119(.data_in(wire_d65_118),.data_out(d_out65),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance670660(.data_in(d_in66),.data_out(wire_d66_0),.clk(clk),.rst(rst));            //channel 67
	decoder_top #(.WIDTH(WIDTH)) decoder_instance670661(.data_in(wire_d66_0),.data_out(wire_d66_1),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance670662(.data_in(wire_d66_1),.data_out(wire_d66_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance670663(.data_in(wire_d66_2),.data_out(wire_d66_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance670664(.data_in(wire_d66_3),.data_out(wire_d66_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance670665(.data_in(wire_d66_4),.data_out(wire_d66_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance670666(.data_in(wire_d66_5),.data_out(wire_d66_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance670667(.data_in(wire_d66_6),.data_out(wire_d66_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance670668(.data_in(wire_d66_7),.data_out(wire_d66_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance670669(.data_in(wire_d66_8),.data_out(wire_d66_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6706610(.data_in(wire_d66_9),.data_out(wire_d66_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6706611(.data_in(wire_d66_10),.data_out(wire_d66_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6706612(.data_in(wire_d66_11),.data_out(wire_d66_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6706613(.data_in(wire_d66_12),.data_out(wire_d66_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6706614(.data_in(wire_d66_13),.data_out(wire_d66_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6706615(.data_in(wire_d66_14),.data_out(wire_d66_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6706616(.data_in(wire_d66_15),.data_out(wire_d66_16),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6706617(.data_in(wire_d66_16),.data_out(wire_d66_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6706618(.data_in(wire_d66_17),.data_out(wire_d66_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6706619(.data_in(wire_d66_18),.data_out(wire_d66_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6706620(.data_in(wire_d66_19),.data_out(wire_d66_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6706621(.data_in(wire_d66_20),.data_out(wire_d66_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6706622(.data_in(wire_d66_21),.data_out(wire_d66_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6706623(.data_in(wire_d66_22),.data_out(wire_d66_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6706624(.data_in(wire_d66_23),.data_out(wire_d66_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6706625(.data_in(wire_d66_24),.data_out(wire_d66_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6706626(.data_in(wire_d66_25),.data_out(wire_d66_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6706627(.data_in(wire_d66_26),.data_out(wire_d66_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6706628(.data_in(wire_d66_27),.data_out(wire_d66_28),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6706629(.data_in(wire_d66_28),.data_out(wire_d66_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6706630(.data_in(wire_d66_29),.data_out(wire_d66_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6706631(.data_in(wire_d66_30),.data_out(wire_d66_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6706632(.data_in(wire_d66_31),.data_out(wire_d66_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6706633(.data_in(wire_d66_32),.data_out(wire_d66_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6706634(.data_in(wire_d66_33),.data_out(wire_d66_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6706635(.data_in(wire_d66_34),.data_out(wire_d66_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6706636(.data_in(wire_d66_35),.data_out(wire_d66_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6706637(.data_in(wire_d66_36),.data_out(wire_d66_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6706638(.data_in(wire_d66_37),.data_out(wire_d66_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6706639(.data_in(wire_d66_38),.data_out(wire_d66_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6706640(.data_in(wire_d66_39),.data_out(wire_d66_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6706641(.data_in(wire_d66_40),.data_out(wire_d66_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6706642(.data_in(wire_d66_41),.data_out(wire_d66_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6706643(.data_in(wire_d66_42),.data_out(wire_d66_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6706644(.data_in(wire_d66_43),.data_out(wire_d66_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6706645(.data_in(wire_d66_44),.data_out(wire_d66_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6706646(.data_in(wire_d66_45),.data_out(wire_d66_46),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6706647(.data_in(wire_d66_46),.data_out(wire_d66_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6706648(.data_in(wire_d66_47),.data_out(wire_d66_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6706649(.data_in(wire_d66_48),.data_out(wire_d66_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6706650(.data_in(wire_d66_49),.data_out(wire_d66_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6706651(.data_in(wire_d66_50),.data_out(wire_d66_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6706652(.data_in(wire_d66_51),.data_out(wire_d66_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6706653(.data_in(wire_d66_52),.data_out(wire_d66_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6706654(.data_in(wire_d66_53),.data_out(wire_d66_54),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6706655(.data_in(wire_d66_54),.data_out(wire_d66_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6706656(.data_in(wire_d66_55),.data_out(wire_d66_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6706657(.data_in(wire_d66_56),.data_out(wire_d66_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6706658(.data_in(wire_d66_57),.data_out(wire_d66_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6706659(.data_in(wire_d66_58),.data_out(wire_d66_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6706660(.data_in(wire_d66_59),.data_out(wire_d66_60),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6706661(.data_in(wire_d66_60),.data_out(wire_d66_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6706662(.data_in(wire_d66_61),.data_out(wire_d66_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6706663(.data_in(wire_d66_62),.data_out(wire_d66_63),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6706664(.data_in(wire_d66_63),.data_out(wire_d66_64),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6706665(.data_in(wire_d66_64),.data_out(wire_d66_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6706666(.data_in(wire_d66_65),.data_out(wire_d66_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6706667(.data_in(wire_d66_66),.data_out(wire_d66_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6706668(.data_in(wire_d66_67),.data_out(wire_d66_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6706669(.data_in(wire_d66_68),.data_out(wire_d66_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6706670(.data_in(wire_d66_69),.data_out(wire_d66_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6706671(.data_in(wire_d66_70),.data_out(wire_d66_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6706672(.data_in(wire_d66_71),.data_out(wire_d66_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6706673(.data_in(wire_d66_72),.data_out(wire_d66_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6706674(.data_in(wire_d66_73),.data_out(wire_d66_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6706675(.data_in(wire_d66_74),.data_out(wire_d66_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6706676(.data_in(wire_d66_75),.data_out(wire_d66_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6706677(.data_in(wire_d66_76),.data_out(wire_d66_77),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6706678(.data_in(wire_d66_77),.data_out(wire_d66_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6706679(.data_in(wire_d66_78),.data_out(wire_d66_79),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6706680(.data_in(wire_d66_79),.data_out(wire_d66_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6706681(.data_in(wire_d66_80),.data_out(wire_d66_81),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6706682(.data_in(wire_d66_81),.data_out(wire_d66_82),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6706683(.data_in(wire_d66_82),.data_out(wire_d66_83),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6706684(.data_in(wire_d66_83),.data_out(wire_d66_84),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6706685(.data_in(wire_d66_84),.data_out(wire_d66_85),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6706686(.data_in(wire_d66_85),.data_out(wire_d66_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6706687(.data_in(wire_d66_86),.data_out(wire_d66_87),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6706688(.data_in(wire_d66_87),.data_out(wire_d66_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6706689(.data_in(wire_d66_88),.data_out(wire_d66_89),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6706690(.data_in(wire_d66_89),.data_out(wire_d66_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6706691(.data_in(wire_d66_90),.data_out(wire_d66_91),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6706692(.data_in(wire_d66_91),.data_out(wire_d66_92),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6706693(.data_in(wire_d66_92),.data_out(wire_d66_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6706694(.data_in(wire_d66_93),.data_out(wire_d66_94),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6706695(.data_in(wire_d66_94),.data_out(wire_d66_95),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6706696(.data_in(wire_d66_95),.data_out(wire_d66_96),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6706697(.data_in(wire_d66_96),.data_out(wire_d66_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6706698(.data_in(wire_d66_97),.data_out(wire_d66_98),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6706699(.data_in(wire_d66_98),.data_out(wire_d66_99),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance67066100(.data_in(wire_d66_99),.data_out(wire_d66_100),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance67066101(.data_in(wire_d66_100),.data_out(wire_d66_101),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance67066102(.data_in(wire_d66_101),.data_out(wire_d66_102),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance67066103(.data_in(wire_d66_102),.data_out(wire_d66_103),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance67066104(.data_in(wire_d66_103),.data_out(wire_d66_104),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance67066105(.data_in(wire_d66_104),.data_out(wire_d66_105),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance67066106(.data_in(wire_d66_105),.data_out(wire_d66_106),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance67066107(.data_in(wire_d66_106),.data_out(wire_d66_107),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance67066108(.data_in(wire_d66_107),.data_out(wire_d66_108),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance67066109(.data_in(wire_d66_108),.data_out(wire_d66_109),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance67066110(.data_in(wire_d66_109),.data_out(wire_d66_110),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance67066111(.data_in(wire_d66_110),.data_out(wire_d66_111),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance67066112(.data_in(wire_d66_111),.data_out(wire_d66_112),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance67066113(.data_in(wire_d66_112),.data_out(wire_d66_113),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance67066114(.data_in(wire_d66_113),.data_out(wire_d66_114),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance67066115(.data_in(wire_d66_114),.data_out(wire_d66_115),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance67066116(.data_in(wire_d66_115),.data_out(wire_d66_116),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance67066117(.data_in(wire_d66_116),.data_out(wire_d66_117),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance67066118(.data_in(wire_d66_117),.data_out(wire_d66_118),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance67066119(.data_in(wire_d66_118),.data_out(d_out66),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance680670(.data_in(d_in67),.data_out(wire_d67_0),.clk(clk),.rst(rst));            //channel 68
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance680671(.data_in(wire_d67_0),.data_out(wire_d67_1),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance680672(.data_in(wire_d67_1),.data_out(wire_d67_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance680673(.data_in(wire_d67_2),.data_out(wire_d67_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance680674(.data_in(wire_d67_3),.data_out(wire_d67_4),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance680675(.data_in(wire_d67_4),.data_out(wire_d67_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance680676(.data_in(wire_d67_5),.data_out(wire_d67_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance680677(.data_in(wire_d67_6),.data_out(wire_d67_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance680678(.data_in(wire_d67_7),.data_out(wire_d67_8),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance680679(.data_in(wire_d67_8),.data_out(wire_d67_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6806710(.data_in(wire_d67_9),.data_out(wire_d67_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6806711(.data_in(wire_d67_10),.data_out(wire_d67_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6806712(.data_in(wire_d67_11),.data_out(wire_d67_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6806713(.data_in(wire_d67_12),.data_out(wire_d67_13),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6806714(.data_in(wire_d67_13),.data_out(wire_d67_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6806715(.data_in(wire_d67_14),.data_out(wire_d67_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6806716(.data_in(wire_d67_15),.data_out(wire_d67_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6806717(.data_in(wire_d67_16),.data_out(wire_d67_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6806718(.data_in(wire_d67_17),.data_out(wire_d67_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6806719(.data_in(wire_d67_18),.data_out(wire_d67_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6806720(.data_in(wire_d67_19),.data_out(wire_d67_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6806721(.data_in(wire_d67_20),.data_out(wire_d67_21),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6806722(.data_in(wire_d67_21),.data_out(wire_d67_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6806723(.data_in(wire_d67_22),.data_out(wire_d67_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6806724(.data_in(wire_d67_23),.data_out(wire_d67_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6806725(.data_in(wire_d67_24),.data_out(wire_d67_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6806726(.data_in(wire_d67_25),.data_out(wire_d67_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6806727(.data_in(wire_d67_26),.data_out(wire_d67_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6806728(.data_in(wire_d67_27),.data_out(wire_d67_28),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6806729(.data_in(wire_d67_28),.data_out(wire_d67_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6806730(.data_in(wire_d67_29),.data_out(wire_d67_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6806731(.data_in(wire_d67_30),.data_out(wire_d67_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6806732(.data_in(wire_d67_31),.data_out(wire_d67_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6806733(.data_in(wire_d67_32),.data_out(wire_d67_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6806734(.data_in(wire_d67_33),.data_out(wire_d67_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6806735(.data_in(wire_d67_34),.data_out(wire_d67_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6806736(.data_in(wire_d67_35),.data_out(wire_d67_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6806737(.data_in(wire_d67_36),.data_out(wire_d67_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6806738(.data_in(wire_d67_37),.data_out(wire_d67_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6806739(.data_in(wire_d67_38),.data_out(wire_d67_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6806740(.data_in(wire_d67_39),.data_out(wire_d67_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6806741(.data_in(wire_d67_40),.data_out(wire_d67_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6806742(.data_in(wire_d67_41),.data_out(wire_d67_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6806743(.data_in(wire_d67_42),.data_out(wire_d67_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6806744(.data_in(wire_d67_43),.data_out(wire_d67_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6806745(.data_in(wire_d67_44),.data_out(wire_d67_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6806746(.data_in(wire_d67_45),.data_out(wire_d67_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6806747(.data_in(wire_d67_46),.data_out(wire_d67_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6806748(.data_in(wire_d67_47),.data_out(wire_d67_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6806749(.data_in(wire_d67_48),.data_out(wire_d67_49),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6806750(.data_in(wire_d67_49),.data_out(wire_d67_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6806751(.data_in(wire_d67_50),.data_out(wire_d67_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6806752(.data_in(wire_d67_51),.data_out(wire_d67_52),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6806753(.data_in(wire_d67_52),.data_out(wire_d67_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6806754(.data_in(wire_d67_53),.data_out(wire_d67_54),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6806755(.data_in(wire_d67_54),.data_out(wire_d67_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6806756(.data_in(wire_d67_55),.data_out(wire_d67_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6806757(.data_in(wire_d67_56),.data_out(wire_d67_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6806758(.data_in(wire_d67_57),.data_out(wire_d67_58),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6806759(.data_in(wire_d67_58),.data_out(wire_d67_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6806760(.data_in(wire_d67_59),.data_out(wire_d67_60),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6806761(.data_in(wire_d67_60),.data_out(wire_d67_61),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6806762(.data_in(wire_d67_61),.data_out(wire_d67_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6806763(.data_in(wire_d67_62),.data_out(wire_d67_63),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6806764(.data_in(wire_d67_63),.data_out(wire_d67_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6806765(.data_in(wire_d67_64),.data_out(wire_d67_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6806766(.data_in(wire_d67_65),.data_out(wire_d67_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6806767(.data_in(wire_d67_66),.data_out(wire_d67_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6806768(.data_in(wire_d67_67),.data_out(wire_d67_68),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6806769(.data_in(wire_d67_68),.data_out(wire_d67_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6806770(.data_in(wire_d67_69),.data_out(wire_d67_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6806771(.data_in(wire_d67_70),.data_out(wire_d67_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6806772(.data_in(wire_d67_71),.data_out(wire_d67_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6806773(.data_in(wire_d67_72),.data_out(wire_d67_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6806774(.data_in(wire_d67_73),.data_out(wire_d67_74),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6806775(.data_in(wire_d67_74),.data_out(wire_d67_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6806776(.data_in(wire_d67_75),.data_out(wire_d67_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6806777(.data_in(wire_d67_76),.data_out(wire_d67_77),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6806778(.data_in(wire_d67_77),.data_out(wire_d67_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6806779(.data_in(wire_d67_78),.data_out(wire_d67_79),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6806780(.data_in(wire_d67_79),.data_out(wire_d67_80),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6806781(.data_in(wire_d67_80),.data_out(wire_d67_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6806782(.data_in(wire_d67_81),.data_out(wire_d67_82),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6806783(.data_in(wire_d67_82),.data_out(wire_d67_83),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6806784(.data_in(wire_d67_83),.data_out(wire_d67_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6806785(.data_in(wire_d67_84),.data_out(wire_d67_85),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6806786(.data_in(wire_d67_85),.data_out(wire_d67_86),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6806787(.data_in(wire_d67_86),.data_out(wire_d67_87),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6806788(.data_in(wire_d67_87),.data_out(wire_d67_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6806789(.data_in(wire_d67_88),.data_out(wire_d67_89),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6806790(.data_in(wire_d67_89),.data_out(wire_d67_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6806791(.data_in(wire_d67_90),.data_out(wire_d67_91),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6806792(.data_in(wire_d67_91),.data_out(wire_d67_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6806793(.data_in(wire_d67_92),.data_out(wire_d67_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6806794(.data_in(wire_d67_93),.data_out(wire_d67_94),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6806795(.data_in(wire_d67_94),.data_out(wire_d67_95),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6806796(.data_in(wire_d67_95),.data_out(wire_d67_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6806797(.data_in(wire_d67_96),.data_out(wire_d67_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6806798(.data_in(wire_d67_97),.data_out(wire_d67_98),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6806799(.data_in(wire_d67_98),.data_out(wire_d67_99),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance68067100(.data_in(wire_d67_99),.data_out(wire_d67_100),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance68067101(.data_in(wire_d67_100),.data_out(wire_d67_101),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance68067102(.data_in(wire_d67_101),.data_out(wire_d67_102),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance68067103(.data_in(wire_d67_102),.data_out(wire_d67_103),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance68067104(.data_in(wire_d67_103),.data_out(wire_d67_104),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance68067105(.data_in(wire_d67_104),.data_out(wire_d67_105),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance68067106(.data_in(wire_d67_105),.data_out(wire_d67_106),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance68067107(.data_in(wire_d67_106),.data_out(wire_d67_107),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance68067108(.data_in(wire_d67_107),.data_out(wire_d67_108),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance68067109(.data_in(wire_d67_108),.data_out(wire_d67_109),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance68067110(.data_in(wire_d67_109),.data_out(wire_d67_110),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance68067111(.data_in(wire_d67_110),.data_out(wire_d67_111),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance68067112(.data_in(wire_d67_111),.data_out(wire_d67_112),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance68067113(.data_in(wire_d67_112),.data_out(wire_d67_113),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance68067114(.data_in(wire_d67_113),.data_out(wire_d67_114),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance68067115(.data_in(wire_d67_114),.data_out(wire_d67_115),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance68067116(.data_in(wire_d67_115),.data_out(wire_d67_116),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance68067117(.data_in(wire_d67_116),.data_out(wire_d67_117),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance68067118(.data_in(wire_d67_117),.data_out(wire_d67_118),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance68067119(.data_in(wire_d67_118),.data_out(d_out67),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance690680(.data_in(d_in68),.data_out(wire_d68_0),.clk(clk),.rst(rst));            //channel 69
	decoder_top #(.WIDTH(WIDTH)) decoder_instance690681(.data_in(wire_d68_0),.data_out(wire_d68_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance690682(.data_in(wire_d68_1),.data_out(wire_d68_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance690683(.data_in(wire_d68_2),.data_out(wire_d68_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance690684(.data_in(wire_d68_3),.data_out(wire_d68_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance690685(.data_in(wire_d68_4),.data_out(wire_d68_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance690686(.data_in(wire_d68_5),.data_out(wire_d68_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance690687(.data_in(wire_d68_6),.data_out(wire_d68_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance690688(.data_in(wire_d68_7),.data_out(wire_d68_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance690689(.data_in(wire_d68_8),.data_out(wire_d68_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6906810(.data_in(wire_d68_9),.data_out(wire_d68_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6906811(.data_in(wire_d68_10),.data_out(wire_d68_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6906812(.data_in(wire_d68_11),.data_out(wire_d68_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6906813(.data_in(wire_d68_12),.data_out(wire_d68_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6906814(.data_in(wire_d68_13),.data_out(wire_d68_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6906815(.data_in(wire_d68_14),.data_out(wire_d68_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6906816(.data_in(wire_d68_15),.data_out(wire_d68_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6906817(.data_in(wire_d68_16),.data_out(wire_d68_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6906818(.data_in(wire_d68_17),.data_out(wire_d68_18),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6906819(.data_in(wire_d68_18),.data_out(wire_d68_19),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6906820(.data_in(wire_d68_19),.data_out(wire_d68_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6906821(.data_in(wire_d68_20),.data_out(wire_d68_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6906822(.data_in(wire_d68_21),.data_out(wire_d68_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6906823(.data_in(wire_d68_22),.data_out(wire_d68_23),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6906824(.data_in(wire_d68_23),.data_out(wire_d68_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6906825(.data_in(wire_d68_24),.data_out(wire_d68_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6906826(.data_in(wire_d68_25),.data_out(wire_d68_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6906827(.data_in(wire_d68_26),.data_out(wire_d68_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6906828(.data_in(wire_d68_27),.data_out(wire_d68_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6906829(.data_in(wire_d68_28),.data_out(wire_d68_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6906830(.data_in(wire_d68_29),.data_out(wire_d68_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6906831(.data_in(wire_d68_30),.data_out(wire_d68_31),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6906832(.data_in(wire_d68_31),.data_out(wire_d68_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6906833(.data_in(wire_d68_32),.data_out(wire_d68_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6906834(.data_in(wire_d68_33),.data_out(wire_d68_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6906835(.data_in(wire_d68_34),.data_out(wire_d68_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6906836(.data_in(wire_d68_35),.data_out(wire_d68_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6906837(.data_in(wire_d68_36),.data_out(wire_d68_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6906838(.data_in(wire_d68_37),.data_out(wire_d68_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6906839(.data_in(wire_d68_38),.data_out(wire_d68_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6906840(.data_in(wire_d68_39),.data_out(wire_d68_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6906841(.data_in(wire_d68_40),.data_out(wire_d68_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6906842(.data_in(wire_d68_41),.data_out(wire_d68_42),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6906843(.data_in(wire_d68_42),.data_out(wire_d68_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6906844(.data_in(wire_d68_43),.data_out(wire_d68_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6906845(.data_in(wire_d68_44),.data_out(wire_d68_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6906846(.data_in(wire_d68_45),.data_out(wire_d68_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6906847(.data_in(wire_d68_46),.data_out(wire_d68_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6906848(.data_in(wire_d68_47),.data_out(wire_d68_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6906849(.data_in(wire_d68_48),.data_out(wire_d68_49),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6906850(.data_in(wire_d68_49),.data_out(wire_d68_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6906851(.data_in(wire_d68_50),.data_out(wire_d68_51),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6906852(.data_in(wire_d68_51),.data_out(wire_d68_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6906853(.data_in(wire_d68_52),.data_out(wire_d68_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6906854(.data_in(wire_d68_53),.data_out(wire_d68_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6906855(.data_in(wire_d68_54),.data_out(wire_d68_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6906856(.data_in(wire_d68_55),.data_out(wire_d68_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6906857(.data_in(wire_d68_56),.data_out(wire_d68_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6906858(.data_in(wire_d68_57),.data_out(wire_d68_58),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6906859(.data_in(wire_d68_58),.data_out(wire_d68_59),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6906860(.data_in(wire_d68_59),.data_out(wire_d68_60),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6906861(.data_in(wire_d68_60),.data_out(wire_d68_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6906862(.data_in(wire_d68_61),.data_out(wire_d68_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6906863(.data_in(wire_d68_62),.data_out(wire_d68_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6906864(.data_in(wire_d68_63),.data_out(wire_d68_64),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6906865(.data_in(wire_d68_64),.data_out(wire_d68_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6906866(.data_in(wire_d68_65),.data_out(wire_d68_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6906867(.data_in(wire_d68_66),.data_out(wire_d68_67),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6906868(.data_in(wire_d68_67),.data_out(wire_d68_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6906869(.data_in(wire_d68_68),.data_out(wire_d68_69),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6906870(.data_in(wire_d68_69),.data_out(wire_d68_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6906871(.data_in(wire_d68_70),.data_out(wire_d68_71),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6906872(.data_in(wire_d68_71),.data_out(wire_d68_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6906873(.data_in(wire_d68_72),.data_out(wire_d68_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6906874(.data_in(wire_d68_73),.data_out(wire_d68_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6906875(.data_in(wire_d68_74),.data_out(wire_d68_75),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6906876(.data_in(wire_d68_75),.data_out(wire_d68_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6906877(.data_in(wire_d68_76),.data_out(wire_d68_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6906878(.data_in(wire_d68_77),.data_out(wire_d68_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6906879(.data_in(wire_d68_78),.data_out(wire_d68_79),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6906880(.data_in(wire_d68_79),.data_out(wire_d68_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6906881(.data_in(wire_d68_80),.data_out(wire_d68_81),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6906882(.data_in(wire_d68_81),.data_out(wire_d68_82),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6906883(.data_in(wire_d68_82),.data_out(wire_d68_83),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6906884(.data_in(wire_d68_83),.data_out(wire_d68_84),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6906885(.data_in(wire_d68_84),.data_out(wire_d68_85),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6906886(.data_in(wire_d68_85),.data_out(wire_d68_86),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6906887(.data_in(wire_d68_86),.data_out(wire_d68_87),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6906888(.data_in(wire_d68_87),.data_out(wire_d68_88),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6906889(.data_in(wire_d68_88),.data_out(wire_d68_89),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6906890(.data_in(wire_d68_89),.data_out(wire_d68_90),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6906891(.data_in(wire_d68_90),.data_out(wire_d68_91),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6906892(.data_in(wire_d68_91),.data_out(wire_d68_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6906893(.data_in(wire_d68_92),.data_out(wire_d68_93),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6906894(.data_in(wire_d68_93),.data_out(wire_d68_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6906895(.data_in(wire_d68_94),.data_out(wire_d68_95),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6906896(.data_in(wire_d68_95),.data_out(wire_d68_96),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6906897(.data_in(wire_d68_96),.data_out(wire_d68_97),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6906898(.data_in(wire_d68_97),.data_out(wire_d68_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6906899(.data_in(wire_d68_98),.data_out(wire_d68_99),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance69068100(.data_in(wire_d68_99),.data_out(wire_d68_100),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance69068101(.data_in(wire_d68_100),.data_out(wire_d68_101),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance69068102(.data_in(wire_d68_101),.data_out(wire_d68_102),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance69068103(.data_in(wire_d68_102),.data_out(wire_d68_103),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance69068104(.data_in(wire_d68_103),.data_out(wire_d68_104),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance69068105(.data_in(wire_d68_104),.data_out(wire_d68_105),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance69068106(.data_in(wire_d68_105),.data_out(wire_d68_106),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance69068107(.data_in(wire_d68_106),.data_out(wire_d68_107),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance69068108(.data_in(wire_d68_107),.data_out(wire_d68_108),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance69068109(.data_in(wire_d68_108),.data_out(wire_d68_109),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance69068110(.data_in(wire_d68_109),.data_out(wire_d68_110),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance69068111(.data_in(wire_d68_110),.data_out(wire_d68_111),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance69068112(.data_in(wire_d68_111),.data_out(wire_d68_112),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance69068113(.data_in(wire_d68_112),.data_out(wire_d68_113),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance69068114(.data_in(wire_d68_113),.data_out(wire_d68_114),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance69068115(.data_in(wire_d68_114),.data_out(wire_d68_115),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance69068116(.data_in(wire_d68_115),.data_out(wire_d68_116),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance69068117(.data_in(wire_d68_116),.data_out(wire_d68_117),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance69068118(.data_in(wire_d68_117),.data_out(wire_d68_118),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance69068119(.data_in(wire_d68_118),.data_out(d_out68),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance700690(.data_in(d_in69),.data_out(wire_d69_0),.clk(clk),.rst(rst));            //channel 70
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance700691(.data_in(wire_d69_0),.data_out(wire_d69_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance700692(.data_in(wire_d69_1),.data_out(wire_d69_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance700693(.data_in(wire_d69_2),.data_out(wire_d69_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance700694(.data_in(wire_d69_3),.data_out(wire_d69_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance700695(.data_in(wire_d69_4),.data_out(wire_d69_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance700696(.data_in(wire_d69_5),.data_out(wire_d69_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance700697(.data_in(wire_d69_6),.data_out(wire_d69_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance700698(.data_in(wire_d69_7),.data_out(wire_d69_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance700699(.data_in(wire_d69_8),.data_out(wire_d69_9),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7006910(.data_in(wire_d69_9),.data_out(wire_d69_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7006911(.data_in(wire_d69_10),.data_out(wire_d69_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7006912(.data_in(wire_d69_11),.data_out(wire_d69_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7006913(.data_in(wire_d69_12),.data_out(wire_d69_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7006914(.data_in(wire_d69_13),.data_out(wire_d69_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7006915(.data_in(wire_d69_14),.data_out(wire_d69_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7006916(.data_in(wire_d69_15),.data_out(wire_d69_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7006917(.data_in(wire_d69_16),.data_out(wire_d69_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7006918(.data_in(wire_d69_17),.data_out(wire_d69_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7006919(.data_in(wire_d69_18),.data_out(wire_d69_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7006920(.data_in(wire_d69_19),.data_out(wire_d69_20),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7006921(.data_in(wire_d69_20),.data_out(wire_d69_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7006922(.data_in(wire_d69_21),.data_out(wire_d69_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7006923(.data_in(wire_d69_22),.data_out(wire_d69_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7006924(.data_in(wire_d69_23),.data_out(wire_d69_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7006925(.data_in(wire_d69_24),.data_out(wire_d69_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7006926(.data_in(wire_d69_25),.data_out(wire_d69_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7006927(.data_in(wire_d69_26),.data_out(wire_d69_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7006928(.data_in(wire_d69_27),.data_out(wire_d69_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7006929(.data_in(wire_d69_28),.data_out(wire_d69_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7006930(.data_in(wire_d69_29),.data_out(wire_d69_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7006931(.data_in(wire_d69_30),.data_out(wire_d69_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7006932(.data_in(wire_d69_31),.data_out(wire_d69_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7006933(.data_in(wire_d69_32),.data_out(wire_d69_33),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7006934(.data_in(wire_d69_33),.data_out(wire_d69_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7006935(.data_in(wire_d69_34),.data_out(wire_d69_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7006936(.data_in(wire_d69_35),.data_out(wire_d69_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7006937(.data_in(wire_d69_36),.data_out(wire_d69_37),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7006938(.data_in(wire_d69_37),.data_out(wire_d69_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7006939(.data_in(wire_d69_38),.data_out(wire_d69_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7006940(.data_in(wire_d69_39),.data_out(wire_d69_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7006941(.data_in(wire_d69_40),.data_out(wire_d69_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7006942(.data_in(wire_d69_41),.data_out(wire_d69_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7006943(.data_in(wire_d69_42),.data_out(wire_d69_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7006944(.data_in(wire_d69_43),.data_out(wire_d69_44),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7006945(.data_in(wire_d69_44),.data_out(wire_d69_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7006946(.data_in(wire_d69_45),.data_out(wire_d69_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7006947(.data_in(wire_d69_46),.data_out(wire_d69_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7006948(.data_in(wire_d69_47),.data_out(wire_d69_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7006949(.data_in(wire_d69_48),.data_out(wire_d69_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7006950(.data_in(wire_d69_49),.data_out(wire_d69_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7006951(.data_in(wire_d69_50),.data_out(wire_d69_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7006952(.data_in(wire_d69_51),.data_out(wire_d69_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7006953(.data_in(wire_d69_52),.data_out(wire_d69_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7006954(.data_in(wire_d69_53),.data_out(wire_d69_54),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7006955(.data_in(wire_d69_54),.data_out(wire_d69_55),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7006956(.data_in(wire_d69_55),.data_out(wire_d69_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7006957(.data_in(wire_d69_56),.data_out(wire_d69_57),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7006958(.data_in(wire_d69_57),.data_out(wire_d69_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7006959(.data_in(wire_d69_58),.data_out(wire_d69_59),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7006960(.data_in(wire_d69_59),.data_out(wire_d69_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7006961(.data_in(wire_d69_60),.data_out(wire_d69_61),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7006962(.data_in(wire_d69_61),.data_out(wire_d69_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7006963(.data_in(wire_d69_62),.data_out(wire_d69_63),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7006964(.data_in(wire_d69_63),.data_out(wire_d69_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7006965(.data_in(wire_d69_64),.data_out(wire_d69_65),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7006966(.data_in(wire_d69_65),.data_out(wire_d69_66),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7006967(.data_in(wire_d69_66),.data_out(wire_d69_67),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7006968(.data_in(wire_d69_67),.data_out(wire_d69_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7006969(.data_in(wire_d69_68),.data_out(wire_d69_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7006970(.data_in(wire_d69_69),.data_out(wire_d69_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7006971(.data_in(wire_d69_70),.data_out(wire_d69_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7006972(.data_in(wire_d69_71),.data_out(wire_d69_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7006973(.data_in(wire_d69_72),.data_out(wire_d69_73),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7006974(.data_in(wire_d69_73),.data_out(wire_d69_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7006975(.data_in(wire_d69_74),.data_out(wire_d69_75),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7006976(.data_in(wire_d69_75),.data_out(wire_d69_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7006977(.data_in(wire_d69_76),.data_out(wire_d69_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7006978(.data_in(wire_d69_77),.data_out(wire_d69_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7006979(.data_in(wire_d69_78),.data_out(wire_d69_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7006980(.data_in(wire_d69_79),.data_out(wire_d69_80),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7006981(.data_in(wire_d69_80),.data_out(wire_d69_81),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7006982(.data_in(wire_d69_81),.data_out(wire_d69_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7006983(.data_in(wire_d69_82),.data_out(wire_d69_83),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7006984(.data_in(wire_d69_83),.data_out(wire_d69_84),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7006985(.data_in(wire_d69_84),.data_out(wire_d69_85),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7006986(.data_in(wire_d69_85),.data_out(wire_d69_86),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7006987(.data_in(wire_d69_86),.data_out(wire_d69_87),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7006988(.data_in(wire_d69_87),.data_out(wire_d69_88),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7006989(.data_in(wire_d69_88),.data_out(wire_d69_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7006990(.data_in(wire_d69_89),.data_out(wire_d69_90),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7006991(.data_in(wire_d69_90),.data_out(wire_d69_91),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7006992(.data_in(wire_d69_91),.data_out(wire_d69_92),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7006993(.data_in(wire_d69_92),.data_out(wire_d69_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7006994(.data_in(wire_d69_93),.data_out(wire_d69_94),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7006995(.data_in(wire_d69_94),.data_out(wire_d69_95),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7006996(.data_in(wire_d69_95),.data_out(wire_d69_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7006997(.data_in(wire_d69_96),.data_out(wire_d69_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7006998(.data_in(wire_d69_97),.data_out(wire_d69_98),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7006999(.data_in(wire_d69_98),.data_out(wire_d69_99),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance70069100(.data_in(wire_d69_99),.data_out(wire_d69_100),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance70069101(.data_in(wire_d69_100),.data_out(wire_d69_101),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance70069102(.data_in(wire_d69_101),.data_out(wire_d69_102),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance70069103(.data_in(wire_d69_102),.data_out(wire_d69_103),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance70069104(.data_in(wire_d69_103),.data_out(wire_d69_104),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance70069105(.data_in(wire_d69_104),.data_out(wire_d69_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance70069106(.data_in(wire_d69_105),.data_out(wire_d69_106),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance70069107(.data_in(wire_d69_106),.data_out(wire_d69_107),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance70069108(.data_in(wire_d69_107),.data_out(wire_d69_108),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance70069109(.data_in(wire_d69_108),.data_out(wire_d69_109),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance70069110(.data_in(wire_d69_109),.data_out(wire_d69_110),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance70069111(.data_in(wire_d69_110),.data_out(wire_d69_111),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance70069112(.data_in(wire_d69_111),.data_out(wire_d69_112),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance70069113(.data_in(wire_d69_112),.data_out(wire_d69_113),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance70069114(.data_in(wire_d69_113),.data_out(wire_d69_114),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance70069115(.data_in(wire_d69_114),.data_out(wire_d69_115),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance70069116(.data_in(wire_d69_115),.data_out(wire_d69_116),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance70069117(.data_in(wire_d69_116),.data_out(wire_d69_117),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance70069118(.data_in(wire_d69_117),.data_out(wire_d69_118),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance70069119(.data_in(wire_d69_118),.data_out(d_out69),.clk(clk),.rst(rst));

	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance710700(.data_in(d_in70),.data_out(wire_d70_0),.clk(clk),.rst(rst));            //channel 71
	decoder_top #(.WIDTH(WIDTH)) decoder_instance710701(.data_in(wire_d70_0),.data_out(wire_d70_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance710702(.data_in(wire_d70_1),.data_out(wire_d70_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance710703(.data_in(wire_d70_2),.data_out(wire_d70_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance710704(.data_in(wire_d70_3),.data_out(wire_d70_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance710705(.data_in(wire_d70_4),.data_out(wire_d70_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance710706(.data_in(wire_d70_5),.data_out(wire_d70_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance710707(.data_in(wire_d70_6),.data_out(wire_d70_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance710708(.data_in(wire_d70_7),.data_out(wire_d70_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance710709(.data_in(wire_d70_8),.data_out(wire_d70_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7107010(.data_in(wire_d70_9),.data_out(wire_d70_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7107011(.data_in(wire_d70_10),.data_out(wire_d70_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7107012(.data_in(wire_d70_11),.data_out(wire_d70_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7107013(.data_in(wire_d70_12),.data_out(wire_d70_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7107014(.data_in(wire_d70_13),.data_out(wire_d70_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7107015(.data_in(wire_d70_14),.data_out(wire_d70_15),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7107016(.data_in(wire_d70_15),.data_out(wire_d70_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7107017(.data_in(wire_d70_16),.data_out(wire_d70_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7107018(.data_in(wire_d70_17),.data_out(wire_d70_18),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7107019(.data_in(wire_d70_18),.data_out(wire_d70_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7107020(.data_in(wire_d70_19),.data_out(wire_d70_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7107021(.data_in(wire_d70_20),.data_out(wire_d70_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7107022(.data_in(wire_d70_21),.data_out(wire_d70_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7107023(.data_in(wire_d70_22),.data_out(wire_d70_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7107024(.data_in(wire_d70_23),.data_out(wire_d70_24),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7107025(.data_in(wire_d70_24),.data_out(wire_d70_25),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7107026(.data_in(wire_d70_25),.data_out(wire_d70_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7107027(.data_in(wire_d70_26),.data_out(wire_d70_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7107028(.data_in(wire_d70_27),.data_out(wire_d70_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7107029(.data_in(wire_d70_28),.data_out(wire_d70_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7107030(.data_in(wire_d70_29),.data_out(wire_d70_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7107031(.data_in(wire_d70_30),.data_out(wire_d70_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7107032(.data_in(wire_d70_31),.data_out(wire_d70_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7107033(.data_in(wire_d70_32),.data_out(wire_d70_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7107034(.data_in(wire_d70_33),.data_out(wire_d70_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7107035(.data_in(wire_d70_34),.data_out(wire_d70_35),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7107036(.data_in(wire_d70_35),.data_out(wire_d70_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7107037(.data_in(wire_d70_36),.data_out(wire_d70_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7107038(.data_in(wire_d70_37),.data_out(wire_d70_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7107039(.data_in(wire_d70_38),.data_out(wire_d70_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7107040(.data_in(wire_d70_39),.data_out(wire_d70_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7107041(.data_in(wire_d70_40),.data_out(wire_d70_41),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7107042(.data_in(wire_d70_41),.data_out(wire_d70_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7107043(.data_in(wire_d70_42),.data_out(wire_d70_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7107044(.data_in(wire_d70_43),.data_out(wire_d70_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7107045(.data_in(wire_d70_44),.data_out(wire_d70_45),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7107046(.data_in(wire_d70_45),.data_out(wire_d70_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7107047(.data_in(wire_d70_46),.data_out(wire_d70_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7107048(.data_in(wire_d70_47),.data_out(wire_d70_48),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7107049(.data_in(wire_d70_48),.data_out(wire_d70_49),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7107050(.data_in(wire_d70_49),.data_out(wire_d70_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7107051(.data_in(wire_d70_50),.data_out(wire_d70_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7107052(.data_in(wire_d70_51),.data_out(wire_d70_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7107053(.data_in(wire_d70_52),.data_out(wire_d70_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7107054(.data_in(wire_d70_53),.data_out(wire_d70_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7107055(.data_in(wire_d70_54),.data_out(wire_d70_55),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7107056(.data_in(wire_d70_55),.data_out(wire_d70_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7107057(.data_in(wire_d70_56),.data_out(wire_d70_57),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7107058(.data_in(wire_d70_57),.data_out(wire_d70_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7107059(.data_in(wire_d70_58),.data_out(wire_d70_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7107060(.data_in(wire_d70_59),.data_out(wire_d70_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7107061(.data_in(wire_d70_60),.data_out(wire_d70_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7107062(.data_in(wire_d70_61),.data_out(wire_d70_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7107063(.data_in(wire_d70_62),.data_out(wire_d70_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7107064(.data_in(wire_d70_63),.data_out(wire_d70_64),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7107065(.data_in(wire_d70_64),.data_out(wire_d70_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7107066(.data_in(wire_d70_65),.data_out(wire_d70_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7107067(.data_in(wire_d70_66),.data_out(wire_d70_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7107068(.data_in(wire_d70_67),.data_out(wire_d70_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7107069(.data_in(wire_d70_68),.data_out(wire_d70_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7107070(.data_in(wire_d70_69),.data_out(wire_d70_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7107071(.data_in(wire_d70_70),.data_out(wire_d70_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7107072(.data_in(wire_d70_71),.data_out(wire_d70_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7107073(.data_in(wire_d70_72),.data_out(wire_d70_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7107074(.data_in(wire_d70_73),.data_out(wire_d70_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7107075(.data_in(wire_d70_74),.data_out(wire_d70_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7107076(.data_in(wire_d70_75),.data_out(wire_d70_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7107077(.data_in(wire_d70_76),.data_out(wire_d70_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7107078(.data_in(wire_d70_77),.data_out(wire_d70_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7107079(.data_in(wire_d70_78),.data_out(wire_d70_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7107080(.data_in(wire_d70_79),.data_out(wire_d70_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7107081(.data_in(wire_d70_80),.data_out(wire_d70_81),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7107082(.data_in(wire_d70_81),.data_out(wire_d70_82),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7107083(.data_in(wire_d70_82),.data_out(wire_d70_83),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7107084(.data_in(wire_d70_83),.data_out(wire_d70_84),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7107085(.data_in(wire_d70_84),.data_out(wire_d70_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7107086(.data_in(wire_d70_85),.data_out(wire_d70_86),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7107087(.data_in(wire_d70_86),.data_out(wire_d70_87),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7107088(.data_in(wire_d70_87),.data_out(wire_d70_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7107089(.data_in(wire_d70_88),.data_out(wire_d70_89),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7107090(.data_in(wire_d70_89),.data_out(wire_d70_90),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7107091(.data_in(wire_d70_90),.data_out(wire_d70_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7107092(.data_in(wire_d70_91),.data_out(wire_d70_92),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7107093(.data_in(wire_d70_92),.data_out(wire_d70_93),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7107094(.data_in(wire_d70_93),.data_out(wire_d70_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7107095(.data_in(wire_d70_94),.data_out(wire_d70_95),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7107096(.data_in(wire_d70_95),.data_out(wire_d70_96),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7107097(.data_in(wire_d70_96),.data_out(wire_d70_97),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7107098(.data_in(wire_d70_97),.data_out(wire_d70_98),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7107099(.data_in(wire_d70_98),.data_out(wire_d70_99),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance71070100(.data_in(wire_d70_99),.data_out(wire_d70_100),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance71070101(.data_in(wire_d70_100),.data_out(wire_d70_101),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance71070102(.data_in(wire_d70_101),.data_out(wire_d70_102),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance71070103(.data_in(wire_d70_102),.data_out(wire_d70_103),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance71070104(.data_in(wire_d70_103),.data_out(wire_d70_104),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance71070105(.data_in(wire_d70_104),.data_out(wire_d70_105),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance71070106(.data_in(wire_d70_105),.data_out(wire_d70_106),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance71070107(.data_in(wire_d70_106),.data_out(wire_d70_107),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance71070108(.data_in(wire_d70_107),.data_out(wire_d70_108),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance71070109(.data_in(wire_d70_108),.data_out(wire_d70_109),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance71070110(.data_in(wire_d70_109),.data_out(wire_d70_110),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance71070111(.data_in(wire_d70_110),.data_out(wire_d70_111),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance71070112(.data_in(wire_d70_111),.data_out(wire_d70_112),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance71070113(.data_in(wire_d70_112),.data_out(wire_d70_113),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance71070114(.data_in(wire_d70_113),.data_out(wire_d70_114),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance71070115(.data_in(wire_d70_114),.data_out(wire_d70_115),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance71070116(.data_in(wire_d70_115),.data_out(wire_d70_116),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance71070117(.data_in(wire_d70_116),.data_out(wire_d70_117),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance71070118(.data_in(wire_d70_117),.data_out(wire_d70_118),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance71070119(.data_in(wire_d70_118),.data_out(d_out70),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance720710(.data_in(d_in71),.data_out(wire_d71_0),.clk(clk),.rst(rst));            //channel 72
	large_mux #(.WIDTH(WIDTH)) large_mux_instance720711(.data_in(wire_d71_0),.data_out(wire_d71_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance720712(.data_in(wire_d71_1),.data_out(wire_d71_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance720713(.data_in(wire_d71_2),.data_out(wire_d71_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance720714(.data_in(wire_d71_3),.data_out(wire_d71_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance720715(.data_in(wire_d71_4),.data_out(wire_d71_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance720716(.data_in(wire_d71_5),.data_out(wire_d71_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance720717(.data_in(wire_d71_6),.data_out(wire_d71_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance720718(.data_in(wire_d71_7),.data_out(wire_d71_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance720719(.data_in(wire_d71_8),.data_out(wire_d71_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7207110(.data_in(wire_d71_9),.data_out(wire_d71_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7207111(.data_in(wire_d71_10),.data_out(wire_d71_11),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7207112(.data_in(wire_d71_11),.data_out(wire_d71_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7207113(.data_in(wire_d71_12),.data_out(wire_d71_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7207114(.data_in(wire_d71_13),.data_out(wire_d71_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7207115(.data_in(wire_d71_14),.data_out(wire_d71_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7207116(.data_in(wire_d71_15),.data_out(wire_d71_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7207117(.data_in(wire_d71_16),.data_out(wire_d71_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7207118(.data_in(wire_d71_17),.data_out(wire_d71_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7207119(.data_in(wire_d71_18),.data_out(wire_d71_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7207120(.data_in(wire_d71_19),.data_out(wire_d71_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7207121(.data_in(wire_d71_20),.data_out(wire_d71_21),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7207122(.data_in(wire_d71_21),.data_out(wire_d71_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7207123(.data_in(wire_d71_22),.data_out(wire_d71_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7207124(.data_in(wire_d71_23),.data_out(wire_d71_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7207125(.data_in(wire_d71_24),.data_out(wire_d71_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7207126(.data_in(wire_d71_25),.data_out(wire_d71_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7207127(.data_in(wire_d71_26),.data_out(wire_d71_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7207128(.data_in(wire_d71_27),.data_out(wire_d71_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7207129(.data_in(wire_d71_28),.data_out(wire_d71_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7207130(.data_in(wire_d71_29),.data_out(wire_d71_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7207131(.data_in(wire_d71_30),.data_out(wire_d71_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7207132(.data_in(wire_d71_31),.data_out(wire_d71_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7207133(.data_in(wire_d71_32),.data_out(wire_d71_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7207134(.data_in(wire_d71_33),.data_out(wire_d71_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7207135(.data_in(wire_d71_34),.data_out(wire_d71_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7207136(.data_in(wire_d71_35),.data_out(wire_d71_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7207137(.data_in(wire_d71_36),.data_out(wire_d71_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7207138(.data_in(wire_d71_37),.data_out(wire_d71_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7207139(.data_in(wire_d71_38),.data_out(wire_d71_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7207140(.data_in(wire_d71_39),.data_out(wire_d71_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7207141(.data_in(wire_d71_40),.data_out(wire_d71_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7207142(.data_in(wire_d71_41),.data_out(wire_d71_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7207143(.data_in(wire_d71_42),.data_out(wire_d71_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7207144(.data_in(wire_d71_43),.data_out(wire_d71_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7207145(.data_in(wire_d71_44),.data_out(wire_d71_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7207146(.data_in(wire_d71_45),.data_out(wire_d71_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7207147(.data_in(wire_d71_46),.data_out(wire_d71_47),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7207148(.data_in(wire_d71_47),.data_out(wire_d71_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7207149(.data_in(wire_d71_48),.data_out(wire_d71_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7207150(.data_in(wire_d71_49),.data_out(wire_d71_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7207151(.data_in(wire_d71_50),.data_out(wire_d71_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7207152(.data_in(wire_d71_51),.data_out(wire_d71_52),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7207153(.data_in(wire_d71_52),.data_out(wire_d71_53),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7207154(.data_in(wire_d71_53),.data_out(wire_d71_54),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7207155(.data_in(wire_d71_54),.data_out(wire_d71_55),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7207156(.data_in(wire_d71_55),.data_out(wire_d71_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7207157(.data_in(wire_d71_56),.data_out(wire_d71_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7207158(.data_in(wire_d71_57),.data_out(wire_d71_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7207159(.data_in(wire_d71_58),.data_out(wire_d71_59),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7207160(.data_in(wire_d71_59),.data_out(wire_d71_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7207161(.data_in(wire_d71_60),.data_out(wire_d71_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7207162(.data_in(wire_d71_61),.data_out(wire_d71_62),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7207163(.data_in(wire_d71_62),.data_out(wire_d71_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7207164(.data_in(wire_d71_63),.data_out(wire_d71_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7207165(.data_in(wire_d71_64),.data_out(wire_d71_65),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7207166(.data_in(wire_d71_65),.data_out(wire_d71_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7207167(.data_in(wire_d71_66),.data_out(wire_d71_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7207168(.data_in(wire_d71_67),.data_out(wire_d71_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7207169(.data_in(wire_d71_68),.data_out(wire_d71_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7207170(.data_in(wire_d71_69),.data_out(wire_d71_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7207171(.data_in(wire_d71_70),.data_out(wire_d71_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7207172(.data_in(wire_d71_71),.data_out(wire_d71_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7207173(.data_in(wire_d71_72),.data_out(wire_d71_73),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7207174(.data_in(wire_d71_73),.data_out(wire_d71_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7207175(.data_in(wire_d71_74),.data_out(wire_d71_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7207176(.data_in(wire_d71_75),.data_out(wire_d71_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7207177(.data_in(wire_d71_76),.data_out(wire_d71_77),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7207178(.data_in(wire_d71_77),.data_out(wire_d71_78),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7207179(.data_in(wire_d71_78),.data_out(wire_d71_79),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7207180(.data_in(wire_d71_79),.data_out(wire_d71_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7207181(.data_in(wire_d71_80),.data_out(wire_d71_81),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7207182(.data_in(wire_d71_81),.data_out(wire_d71_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7207183(.data_in(wire_d71_82),.data_out(wire_d71_83),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7207184(.data_in(wire_d71_83),.data_out(wire_d71_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7207185(.data_in(wire_d71_84),.data_out(wire_d71_85),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7207186(.data_in(wire_d71_85),.data_out(wire_d71_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7207187(.data_in(wire_d71_86),.data_out(wire_d71_87),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7207188(.data_in(wire_d71_87),.data_out(wire_d71_88),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7207189(.data_in(wire_d71_88),.data_out(wire_d71_89),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7207190(.data_in(wire_d71_89),.data_out(wire_d71_90),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7207191(.data_in(wire_d71_90),.data_out(wire_d71_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7207192(.data_in(wire_d71_91),.data_out(wire_d71_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7207193(.data_in(wire_d71_92),.data_out(wire_d71_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7207194(.data_in(wire_d71_93),.data_out(wire_d71_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7207195(.data_in(wire_d71_94),.data_out(wire_d71_95),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7207196(.data_in(wire_d71_95),.data_out(wire_d71_96),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7207197(.data_in(wire_d71_96),.data_out(wire_d71_97),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7207198(.data_in(wire_d71_97),.data_out(wire_d71_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7207199(.data_in(wire_d71_98),.data_out(wire_d71_99),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance72071100(.data_in(wire_d71_99),.data_out(wire_d71_100),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance72071101(.data_in(wire_d71_100),.data_out(wire_d71_101),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance72071102(.data_in(wire_d71_101),.data_out(wire_d71_102),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance72071103(.data_in(wire_d71_102),.data_out(wire_d71_103),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance72071104(.data_in(wire_d71_103),.data_out(wire_d71_104),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance72071105(.data_in(wire_d71_104),.data_out(wire_d71_105),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance72071106(.data_in(wire_d71_105),.data_out(wire_d71_106),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance72071107(.data_in(wire_d71_106),.data_out(wire_d71_107),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance72071108(.data_in(wire_d71_107),.data_out(wire_d71_108),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance72071109(.data_in(wire_d71_108),.data_out(wire_d71_109),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance72071110(.data_in(wire_d71_109),.data_out(wire_d71_110),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance72071111(.data_in(wire_d71_110),.data_out(wire_d71_111),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance72071112(.data_in(wire_d71_111),.data_out(wire_d71_112),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance72071113(.data_in(wire_d71_112),.data_out(wire_d71_113),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance72071114(.data_in(wire_d71_113),.data_out(wire_d71_114),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance72071115(.data_in(wire_d71_114),.data_out(wire_d71_115),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance72071116(.data_in(wire_d71_115),.data_out(wire_d71_116),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance72071117(.data_in(wire_d71_116),.data_out(wire_d71_117),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance72071118(.data_in(wire_d71_117),.data_out(wire_d71_118),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance72071119(.data_in(wire_d71_118),.data_out(d_out71),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance730720(.data_in(d_in72),.data_out(wire_d72_0),.clk(clk),.rst(rst));            //channel 73
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance730721(.data_in(wire_d72_0),.data_out(wire_d72_1),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance730722(.data_in(wire_d72_1),.data_out(wire_d72_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance730723(.data_in(wire_d72_2),.data_out(wire_d72_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance730724(.data_in(wire_d72_3),.data_out(wire_d72_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance730725(.data_in(wire_d72_4),.data_out(wire_d72_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance730726(.data_in(wire_d72_5),.data_out(wire_d72_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance730727(.data_in(wire_d72_6),.data_out(wire_d72_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance730728(.data_in(wire_d72_7),.data_out(wire_d72_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance730729(.data_in(wire_d72_8),.data_out(wire_d72_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7307210(.data_in(wire_d72_9),.data_out(wire_d72_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7307211(.data_in(wire_d72_10),.data_out(wire_d72_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7307212(.data_in(wire_d72_11),.data_out(wire_d72_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7307213(.data_in(wire_d72_12),.data_out(wire_d72_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7307214(.data_in(wire_d72_13),.data_out(wire_d72_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7307215(.data_in(wire_d72_14),.data_out(wire_d72_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7307216(.data_in(wire_d72_15),.data_out(wire_d72_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7307217(.data_in(wire_d72_16),.data_out(wire_d72_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7307218(.data_in(wire_d72_17),.data_out(wire_d72_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7307219(.data_in(wire_d72_18),.data_out(wire_d72_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7307220(.data_in(wire_d72_19),.data_out(wire_d72_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7307221(.data_in(wire_d72_20),.data_out(wire_d72_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7307222(.data_in(wire_d72_21),.data_out(wire_d72_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7307223(.data_in(wire_d72_22),.data_out(wire_d72_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7307224(.data_in(wire_d72_23),.data_out(wire_d72_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7307225(.data_in(wire_d72_24),.data_out(wire_d72_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7307226(.data_in(wire_d72_25),.data_out(wire_d72_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7307227(.data_in(wire_d72_26),.data_out(wire_d72_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7307228(.data_in(wire_d72_27),.data_out(wire_d72_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7307229(.data_in(wire_d72_28),.data_out(wire_d72_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7307230(.data_in(wire_d72_29),.data_out(wire_d72_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7307231(.data_in(wire_d72_30),.data_out(wire_d72_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7307232(.data_in(wire_d72_31),.data_out(wire_d72_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7307233(.data_in(wire_d72_32),.data_out(wire_d72_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7307234(.data_in(wire_d72_33),.data_out(wire_d72_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7307235(.data_in(wire_d72_34),.data_out(wire_d72_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7307236(.data_in(wire_d72_35),.data_out(wire_d72_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7307237(.data_in(wire_d72_36),.data_out(wire_d72_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7307238(.data_in(wire_d72_37),.data_out(wire_d72_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7307239(.data_in(wire_d72_38),.data_out(wire_d72_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7307240(.data_in(wire_d72_39),.data_out(wire_d72_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7307241(.data_in(wire_d72_40),.data_out(wire_d72_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7307242(.data_in(wire_d72_41),.data_out(wire_d72_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7307243(.data_in(wire_d72_42),.data_out(wire_d72_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7307244(.data_in(wire_d72_43),.data_out(wire_d72_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7307245(.data_in(wire_d72_44),.data_out(wire_d72_45),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7307246(.data_in(wire_d72_45),.data_out(wire_d72_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7307247(.data_in(wire_d72_46),.data_out(wire_d72_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7307248(.data_in(wire_d72_47),.data_out(wire_d72_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7307249(.data_in(wire_d72_48),.data_out(wire_d72_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7307250(.data_in(wire_d72_49),.data_out(wire_d72_50),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7307251(.data_in(wire_d72_50),.data_out(wire_d72_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7307252(.data_in(wire_d72_51),.data_out(wire_d72_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7307253(.data_in(wire_d72_52),.data_out(wire_d72_53),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7307254(.data_in(wire_d72_53),.data_out(wire_d72_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7307255(.data_in(wire_d72_54),.data_out(wire_d72_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7307256(.data_in(wire_d72_55),.data_out(wire_d72_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7307257(.data_in(wire_d72_56),.data_out(wire_d72_57),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7307258(.data_in(wire_d72_57),.data_out(wire_d72_58),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7307259(.data_in(wire_d72_58),.data_out(wire_d72_59),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7307260(.data_in(wire_d72_59),.data_out(wire_d72_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7307261(.data_in(wire_d72_60),.data_out(wire_d72_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7307262(.data_in(wire_d72_61),.data_out(wire_d72_62),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7307263(.data_in(wire_d72_62),.data_out(wire_d72_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7307264(.data_in(wire_d72_63),.data_out(wire_d72_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7307265(.data_in(wire_d72_64),.data_out(wire_d72_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7307266(.data_in(wire_d72_65),.data_out(wire_d72_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7307267(.data_in(wire_d72_66),.data_out(wire_d72_67),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7307268(.data_in(wire_d72_67),.data_out(wire_d72_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7307269(.data_in(wire_d72_68),.data_out(wire_d72_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7307270(.data_in(wire_d72_69),.data_out(wire_d72_70),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7307271(.data_in(wire_d72_70),.data_out(wire_d72_71),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7307272(.data_in(wire_d72_71),.data_out(wire_d72_72),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7307273(.data_in(wire_d72_72),.data_out(wire_d72_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7307274(.data_in(wire_d72_73),.data_out(wire_d72_74),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7307275(.data_in(wire_d72_74),.data_out(wire_d72_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7307276(.data_in(wire_d72_75),.data_out(wire_d72_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7307277(.data_in(wire_d72_76),.data_out(wire_d72_77),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7307278(.data_in(wire_d72_77),.data_out(wire_d72_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7307279(.data_in(wire_d72_78),.data_out(wire_d72_79),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7307280(.data_in(wire_d72_79),.data_out(wire_d72_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7307281(.data_in(wire_d72_80),.data_out(wire_d72_81),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7307282(.data_in(wire_d72_81),.data_out(wire_d72_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7307283(.data_in(wire_d72_82),.data_out(wire_d72_83),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7307284(.data_in(wire_d72_83),.data_out(wire_d72_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7307285(.data_in(wire_d72_84),.data_out(wire_d72_85),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7307286(.data_in(wire_d72_85),.data_out(wire_d72_86),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7307287(.data_in(wire_d72_86),.data_out(wire_d72_87),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7307288(.data_in(wire_d72_87),.data_out(wire_d72_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7307289(.data_in(wire_d72_88),.data_out(wire_d72_89),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7307290(.data_in(wire_d72_89),.data_out(wire_d72_90),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7307291(.data_in(wire_d72_90),.data_out(wire_d72_91),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7307292(.data_in(wire_d72_91),.data_out(wire_d72_92),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7307293(.data_in(wire_d72_92),.data_out(wire_d72_93),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7307294(.data_in(wire_d72_93),.data_out(wire_d72_94),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7307295(.data_in(wire_d72_94),.data_out(wire_d72_95),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7307296(.data_in(wire_d72_95),.data_out(wire_d72_96),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7307297(.data_in(wire_d72_96),.data_out(wire_d72_97),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7307298(.data_in(wire_d72_97),.data_out(wire_d72_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7307299(.data_in(wire_d72_98),.data_out(wire_d72_99),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance73072100(.data_in(wire_d72_99),.data_out(wire_d72_100),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance73072101(.data_in(wire_d72_100),.data_out(wire_d72_101),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance73072102(.data_in(wire_d72_101),.data_out(wire_d72_102),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance73072103(.data_in(wire_d72_102),.data_out(wire_d72_103),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance73072104(.data_in(wire_d72_103),.data_out(wire_d72_104),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance73072105(.data_in(wire_d72_104),.data_out(wire_d72_105),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance73072106(.data_in(wire_d72_105),.data_out(wire_d72_106),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance73072107(.data_in(wire_d72_106),.data_out(wire_d72_107),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance73072108(.data_in(wire_d72_107),.data_out(wire_d72_108),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance73072109(.data_in(wire_d72_108),.data_out(wire_d72_109),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance73072110(.data_in(wire_d72_109),.data_out(wire_d72_110),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance73072111(.data_in(wire_d72_110),.data_out(wire_d72_111),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance73072112(.data_in(wire_d72_111),.data_out(wire_d72_112),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance73072113(.data_in(wire_d72_112),.data_out(wire_d72_113),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance73072114(.data_in(wire_d72_113),.data_out(wire_d72_114),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance73072115(.data_in(wire_d72_114),.data_out(wire_d72_115),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance73072116(.data_in(wire_d72_115),.data_out(wire_d72_116),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance73072117(.data_in(wire_d72_116),.data_out(wire_d72_117),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance73072118(.data_in(wire_d72_117),.data_out(wire_d72_118),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance73072119(.data_in(wire_d72_118),.data_out(d_out72),.clk(clk),.rst(rst));

	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance740730(.data_in(d_in73),.data_out(wire_d73_0),.clk(clk),.rst(rst));            //channel 74
	register #(.WIDTH(WIDTH)) register_instance740731(.data_in(wire_d73_0),.data_out(wire_d73_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance740732(.data_in(wire_d73_1),.data_out(wire_d73_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance740733(.data_in(wire_d73_2),.data_out(wire_d73_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance740734(.data_in(wire_d73_3),.data_out(wire_d73_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance740735(.data_in(wire_d73_4),.data_out(wire_d73_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance740736(.data_in(wire_d73_5),.data_out(wire_d73_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance740737(.data_in(wire_d73_6),.data_out(wire_d73_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance740738(.data_in(wire_d73_7),.data_out(wire_d73_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance740739(.data_in(wire_d73_8),.data_out(wire_d73_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7407310(.data_in(wire_d73_9),.data_out(wire_d73_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7407311(.data_in(wire_d73_10),.data_out(wire_d73_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7407312(.data_in(wire_d73_11),.data_out(wire_d73_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7407313(.data_in(wire_d73_12),.data_out(wire_d73_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7407314(.data_in(wire_d73_13),.data_out(wire_d73_14),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7407315(.data_in(wire_d73_14),.data_out(wire_d73_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7407316(.data_in(wire_d73_15),.data_out(wire_d73_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7407317(.data_in(wire_d73_16),.data_out(wire_d73_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7407318(.data_in(wire_d73_17),.data_out(wire_d73_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7407319(.data_in(wire_d73_18),.data_out(wire_d73_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7407320(.data_in(wire_d73_19),.data_out(wire_d73_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7407321(.data_in(wire_d73_20),.data_out(wire_d73_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7407322(.data_in(wire_d73_21),.data_out(wire_d73_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7407323(.data_in(wire_d73_22),.data_out(wire_d73_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7407324(.data_in(wire_d73_23),.data_out(wire_d73_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7407325(.data_in(wire_d73_24),.data_out(wire_d73_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7407326(.data_in(wire_d73_25),.data_out(wire_d73_26),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7407327(.data_in(wire_d73_26),.data_out(wire_d73_27),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7407328(.data_in(wire_d73_27),.data_out(wire_d73_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7407329(.data_in(wire_d73_28),.data_out(wire_d73_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7407330(.data_in(wire_d73_29),.data_out(wire_d73_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7407331(.data_in(wire_d73_30),.data_out(wire_d73_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7407332(.data_in(wire_d73_31),.data_out(wire_d73_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7407333(.data_in(wire_d73_32),.data_out(wire_d73_33),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7407334(.data_in(wire_d73_33),.data_out(wire_d73_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7407335(.data_in(wire_d73_34),.data_out(wire_d73_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7407336(.data_in(wire_d73_35),.data_out(wire_d73_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7407337(.data_in(wire_d73_36),.data_out(wire_d73_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7407338(.data_in(wire_d73_37),.data_out(wire_d73_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7407339(.data_in(wire_d73_38),.data_out(wire_d73_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7407340(.data_in(wire_d73_39),.data_out(wire_d73_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7407341(.data_in(wire_d73_40),.data_out(wire_d73_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7407342(.data_in(wire_d73_41),.data_out(wire_d73_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7407343(.data_in(wire_d73_42),.data_out(wire_d73_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7407344(.data_in(wire_d73_43),.data_out(wire_d73_44),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7407345(.data_in(wire_d73_44),.data_out(wire_d73_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7407346(.data_in(wire_d73_45),.data_out(wire_d73_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7407347(.data_in(wire_d73_46),.data_out(wire_d73_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7407348(.data_in(wire_d73_47),.data_out(wire_d73_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7407349(.data_in(wire_d73_48),.data_out(wire_d73_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7407350(.data_in(wire_d73_49),.data_out(wire_d73_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7407351(.data_in(wire_d73_50),.data_out(wire_d73_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7407352(.data_in(wire_d73_51),.data_out(wire_d73_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7407353(.data_in(wire_d73_52),.data_out(wire_d73_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7407354(.data_in(wire_d73_53),.data_out(wire_d73_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7407355(.data_in(wire_d73_54),.data_out(wire_d73_55),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7407356(.data_in(wire_d73_55),.data_out(wire_d73_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7407357(.data_in(wire_d73_56),.data_out(wire_d73_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7407358(.data_in(wire_d73_57),.data_out(wire_d73_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7407359(.data_in(wire_d73_58),.data_out(wire_d73_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7407360(.data_in(wire_d73_59),.data_out(wire_d73_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7407361(.data_in(wire_d73_60),.data_out(wire_d73_61),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7407362(.data_in(wire_d73_61),.data_out(wire_d73_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7407363(.data_in(wire_d73_62),.data_out(wire_d73_63),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7407364(.data_in(wire_d73_63),.data_out(wire_d73_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7407365(.data_in(wire_d73_64),.data_out(wire_d73_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7407366(.data_in(wire_d73_65),.data_out(wire_d73_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7407367(.data_in(wire_d73_66),.data_out(wire_d73_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7407368(.data_in(wire_d73_67),.data_out(wire_d73_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7407369(.data_in(wire_d73_68),.data_out(wire_d73_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7407370(.data_in(wire_d73_69),.data_out(wire_d73_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7407371(.data_in(wire_d73_70),.data_out(wire_d73_71),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7407372(.data_in(wire_d73_71),.data_out(wire_d73_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7407373(.data_in(wire_d73_72),.data_out(wire_d73_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7407374(.data_in(wire_d73_73),.data_out(wire_d73_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7407375(.data_in(wire_d73_74),.data_out(wire_d73_75),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7407376(.data_in(wire_d73_75),.data_out(wire_d73_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7407377(.data_in(wire_d73_76),.data_out(wire_d73_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7407378(.data_in(wire_d73_77),.data_out(wire_d73_78),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7407379(.data_in(wire_d73_78),.data_out(wire_d73_79),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7407380(.data_in(wire_d73_79),.data_out(wire_d73_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7407381(.data_in(wire_d73_80),.data_out(wire_d73_81),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7407382(.data_in(wire_d73_81),.data_out(wire_d73_82),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7407383(.data_in(wire_d73_82),.data_out(wire_d73_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7407384(.data_in(wire_d73_83),.data_out(wire_d73_84),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7407385(.data_in(wire_d73_84),.data_out(wire_d73_85),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7407386(.data_in(wire_d73_85),.data_out(wire_d73_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7407387(.data_in(wire_d73_86),.data_out(wire_d73_87),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7407388(.data_in(wire_d73_87),.data_out(wire_d73_88),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7407389(.data_in(wire_d73_88),.data_out(wire_d73_89),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7407390(.data_in(wire_d73_89),.data_out(wire_d73_90),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7407391(.data_in(wire_d73_90),.data_out(wire_d73_91),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7407392(.data_in(wire_d73_91),.data_out(wire_d73_92),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7407393(.data_in(wire_d73_92),.data_out(wire_d73_93),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7407394(.data_in(wire_d73_93),.data_out(wire_d73_94),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7407395(.data_in(wire_d73_94),.data_out(wire_d73_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7407396(.data_in(wire_d73_95),.data_out(wire_d73_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7407397(.data_in(wire_d73_96),.data_out(wire_d73_97),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7407398(.data_in(wire_d73_97),.data_out(wire_d73_98),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7407399(.data_in(wire_d73_98),.data_out(wire_d73_99),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance74073100(.data_in(wire_d73_99),.data_out(wire_d73_100),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance74073101(.data_in(wire_d73_100),.data_out(wire_d73_101),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance74073102(.data_in(wire_d73_101),.data_out(wire_d73_102),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance74073103(.data_in(wire_d73_102),.data_out(wire_d73_103),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance74073104(.data_in(wire_d73_103),.data_out(wire_d73_104),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance74073105(.data_in(wire_d73_104),.data_out(wire_d73_105),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance74073106(.data_in(wire_d73_105),.data_out(wire_d73_106),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance74073107(.data_in(wire_d73_106),.data_out(wire_d73_107),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance74073108(.data_in(wire_d73_107),.data_out(wire_d73_108),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance74073109(.data_in(wire_d73_108),.data_out(wire_d73_109),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance74073110(.data_in(wire_d73_109),.data_out(wire_d73_110),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance74073111(.data_in(wire_d73_110),.data_out(wire_d73_111),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance74073112(.data_in(wire_d73_111),.data_out(wire_d73_112),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance74073113(.data_in(wire_d73_112),.data_out(wire_d73_113),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance74073114(.data_in(wire_d73_113),.data_out(wire_d73_114),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance74073115(.data_in(wire_d73_114),.data_out(wire_d73_115),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance74073116(.data_in(wire_d73_115),.data_out(wire_d73_116),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance74073117(.data_in(wire_d73_116),.data_out(wire_d73_117),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance74073118(.data_in(wire_d73_117),.data_out(wire_d73_118),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance74073119(.data_in(wire_d73_118),.data_out(d_out73),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance750740(.data_in(d_in74),.data_out(wire_d74_0),.clk(clk),.rst(rst));            //channel 75
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance750741(.data_in(wire_d74_0),.data_out(wire_d74_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance750742(.data_in(wire_d74_1),.data_out(wire_d74_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance750743(.data_in(wire_d74_2),.data_out(wire_d74_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance750744(.data_in(wire_d74_3),.data_out(wire_d74_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance750745(.data_in(wire_d74_4),.data_out(wire_d74_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance750746(.data_in(wire_d74_5),.data_out(wire_d74_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance750747(.data_in(wire_d74_6),.data_out(wire_d74_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance750748(.data_in(wire_d74_7),.data_out(wire_d74_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance750749(.data_in(wire_d74_8),.data_out(wire_d74_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7507410(.data_in(wire_d74_9),.data_out(wire_d74_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7507411(.data_in(wire_d74_10),.data_out(wire_d74_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7507412(.data_in(wire_d74_11),.data_out(wire_d74_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7507413(.data_in(wire_d74_12),.data_out(wire_d74_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7507414(.data_in(wire_d74_13),.data_out(wire_d74_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7507415(.data_in(wire_d74_14),.data_out(wire_d74_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7507416(.data_in(wire_d74_15),.data_out(wire_d74_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7507417(.data_in(wire_d74_16),.data_out(wire_d74_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7507418(.data_in(wire_d74_17),.data_out(wire_d74_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7507419(.data_in(wire_d74_18),.data_out(wire_d74_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7507420(.data_in(wire_d74_19),.data_out(wire_d74_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7507421(.data_in(wire_d74_20),.data_out(wire_d74_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7507422(.data_in(wire_d74_21),.data_out(wire_d74_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7507423(.data_in(wire_d74_22),.data_out(wire_d74_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7507424(.data_in(wire_d74_23),.data_out(wire_d74_24),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7507425(.data_in(wire_d74_24),.data_out(wire_d74_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7507426(.data_in(wire_d74_25),.data_out(wire_d74_26),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7507427(.data_in(wire_d74_26),.data_out(wire_d74_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7507428(.data_in(wire_d74_27),.data_out(wire_d74_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7507429(.data_in(wire_d74_28),.data_out(wire_d74_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7507430(.data_in(wire_d74_29),.data_out(wire_d74_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7507431(.data_in(wire_d74_30),.data_out(wire_d74_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7507432(.data_in(wire_d74_31),.data_out(wire_d74_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7507433(.data_in(wire_d74_32),.data_out(wire_d74_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7507434(.data_in(wire_d74_33),.data_out(wire_d74_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7507435(.data_in(wire_d74_34),.data_out(wire_d74_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7507436(.data_in(wire_d74_35),.data_out(wire_d74_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7507437(.data_in(wire_d74_36),.data_out(wire_d74_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7507438(.data_in(wire_d74_37),.data_out(wire_d74_38),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7507439(.data_in(wire_d74_38),.data_out(wire_d74_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7507440(.data_in(wire_d74_39),.data_out(wire_d74_40),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7507441(.data_in(wire_d74_40),.data_out(wire_d74_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7507442(.data_in(wire_d74_41),.data_out(wire_d74_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7507443(.data_in(wire_d74_42),.data_out(wire_d74_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7507444(.data_in(wire_d74_43),.data_out(wire_d74_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7507445(.data_in(wire_d74_44),.data_out(wire_d74_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7507446(.data_in(wire_d74_45),.data_out(wire_d74_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7507447(.data_in(wire_d74_46),.data_out(wire_d74_47),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7507448(.data_in(wire_d74_47),.data_out(wire_d74_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7507449(.data_in(wire_d74_48),.data_out(wire_d74_49),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7507450(.data_in(wire_d74_49),.data_out(wire_d74_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7507451(.data_in(wire_d74_50),.data_out(wire_d74_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7507452(.data_in(wire_d74_51),.data_out(wire_d74_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7507453(.data_in(wire_d74_52),.data_out(wire_d74_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7507454(.data_in(wire_d74_53),.data_out(wire_d74_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7507455(.data_in(wire_d74_54),.data_out(wire_d74_55),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7507456(.data_in(wire_d74_55),.data_out(wire_d74_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7507457(.data_in(wire_d74_56),.data_out(wire_d74_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7507458(.data_in(wire_d74_57),.data_out(wire_d74_58),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7507459(.data_in(wire_d74_58),.data_out(wire_d74_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7507460(.data_in(wire_d74_59),.data_out(wire_d74_60),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7507461(.data_in(wire_d74_60),.data_out(wire_d74_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7507462(.data_in(wire_d74_61),.data_out(wire_d74_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7507463(.data_in(wire_d74_62),.data_out(wire_d74_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7507464(.data_in(wire_d74_63),.data_out(wire_d74_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7507465(.data_in(wire_d74_64),.data_out(wire_d74_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7507466(.data_in(wire_d74_65),.data_out(wire_d74_66),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7507467(.data_in(wire_d74_66),.data_out(wire_d74_67),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7507468(.data_in(wire_d74_67),.data_out(wire_d74_68),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7507469(.data_in(wire_d74_68),.data_out(wire_d74_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7507470(.data_in(wire_d74_69),.data_out(wire_d74_70),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7507471(.data_in(wire_d74_70),.data_out(wire_d74_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7507472(.data_in(wire_d74_71),.data_out(wire_d74_72),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7507473(.data_in(wire_d74_72),.data_out(wire_d74_73),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7507474(.data_in(wire_d74_73),.data_out(wire_d74_74),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7507475(.data_in(wire_d74_74),.data_out(wire_d74_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7507476(.data_in(wire_d74_75),.data_out(wire_d74_76),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7507477(.data_in(wire_d74_76),.data_out(wire_d74_77),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7507478(.data_in(wire_d74_77),.data_out(wire_d74_78),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7507479(.data_in(wire_d74_78),.data_out(wire_d74_79),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7507480(.data_in(wire_d74_79),.data_out(wire_d74_80),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7507481(.data_in(wire_d74_80),.data_out(wire_d74_81),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7507482(.data_in(wire_d74_81),.data_out(wire_d74_82),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7507483(.data_in(wire_d74_82),.data_out(wire_d74_83),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7507484(.data_in(wire_d74_83),.data_out(wire_d74_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7507485(.data_in(wire_d74_84),.data_out(wire_d74_85),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7507486(.data_in(wire_d74_85),.data_out(wire_d74_86),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7507487(.data_in(wire_d74_86),.data_out(wire_d74_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7507488(.data_in(wire_d74_87),.data_out(wire_d74_88),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7507489(.data_in(wire_d74_88),.data_out(wire_d74_89),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7507490(.data_in(wire_d74_89),.data_out(wire_d74_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7507491(.data_in(wire_d74_90),.data_out(wire_d74_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7507492(.data_in(wire_d74_91),.data_out(wire_d74_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7507493(.data_in(wire_d74_92),.data_out(wire_d74_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7507494(.data_in(wire_d74_93),.data_out(wire_d74_94),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7507495(.data_in(wire_d74_94),.data_out(wire_d74_95),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7507496(.data_in(wire_d74_95),.data_out(wire_d74_96),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7507497(.data_in(wire_d74_96),.data_out(wire_d74_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7507498(.data_in(wire_d74_97),.data_out(wire_d74_98),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7507499(.data_in(wire_d74_98),.data_out(wire_d74_99),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance75074100(.data_in(wire_d74_99),.data_out(wire_d74_100),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance75074101(.data_in(wire_d74_100),.data_out(wire_d74_101),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance75074102(.data_in(wire_d74_101),.data_out(wire_d74_102),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance75074103(.data_in(wire_d74_102),.data_out(wire_d74_103),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance75074104(.data_in(wire_d74_103),.data_out(wire_d74_104),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance75074105(.data_in(wire_d74_104),.data_out(wire_d74_105),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance75074106(.data_in(wire_d74_105),.data_out(wire_d74_106),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance75074107(.data_in(wire_d74_106),.data_out(wire_d74_107),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance75074108(.data_in(wire_d74_107),.data_out(wire_d74_108),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance75074109(.data_in(wire_d74_108),.data_out(wire_d74_109),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance75074110(.data_in(wire_d74_109),.data_out(wire_d74_110),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance75074111(.data_in(wire_d74_110),.data_out(wire_d74_111),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance75074112(.data_in(wire_d74_111),.data_out(wire_d74_112),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance75074113(.data_in(wire_d74_112),.data_out(wire_d74_113),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance75074114(.data_in(wire_d74_113),.data_out(wire_d74_114),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance75074115(.data_in(wire_d74_114),.data_out(wire_d74_115),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance75074116(.data_in(wire_d74_115),.data_out(wire_d74_116),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance75074117(.data_in(wire_d74_116),.data_out(wire_d74_117),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance75074118(.data_in(wire_d74_117),.data_out(wire_d74_118),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance75074119(.data_in(wire_d74_118),.data_out(d_out74),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance760750(.data_in(d_in75),.data_out(wire_d75_0),.clk(clk),.rst(rst));            //channel 76
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance760751(.data_in(wire_d75_0),.data_out(wire_d75_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance760752(.data_in(wire_d75_1),.data_out(wire_d75_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance760753(.data_in(wire_d75_2),.data_out(wire_d75_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance760754(.data_in(wire_d75_3),.data_out(wire_d75_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance760755(.data_in(wire_d75_4),.data_out(wire_d75_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance760756(.data_in(wire_d75_5),.data_out(wire_d75_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance760757(.data_in(wire_d75_6),.data_out(wire_d75_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance760758(.data_in(wire_d75_7),.data_out(wire_d75_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance760759(.data_in(wire_d75_8),.data_out(wire_d75_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7607510(.data_in(wire_d75_9),.data_out(wire_d75_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7607511(.data_in(wire_d75_10),.data_out(wire_d75_11),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7607512(.data_in(wire_d75_11),.data_out(wire_d75_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7607513(.data_in(wire_d75_12),.data_out(wire_d75_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7607514(.data_in(wire_d75_13),.data_out(wire_d75_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7607515(.data_in(wire_d75_14),.data_out(wire_d75_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7607516(.data_in(wire_d75_15),.data_out(wire_d75_16),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7607517(.data_in(wire_d75_16),.data_out(wire_d75_17),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7607518(.data_in(wire_d75_17),.data_out(wire_d75_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7607519(.data_in(wire_d75_18),.data_out(wire_d75_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7607520(.data_in(wire_d75_19),.data_out(wire_d75_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7607521(.data_in(wire_d75_20),.data_out(wire_d75_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7607522(.data_in(wire_d75_21),.data_out(wire_d75_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7607523(.data_in(wire_d75_22),.data_out(wire_d75_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7607524(.data_in(wire_d75_23),.data_out(wire_d75_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7607525(.data_in(wire_d75_24),.data_out(wire_d75_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7607526(.data_in(wire_d75_25),.data_out(wire_d75_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7607527(.data_in(wire_d75_26),.data_out(wire_d75_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7607528(.data_in(wire_d75_27),.data_out(wire_d75_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7607529(.data_in(wire_d75_28),.data_out(wire_d75_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7607530(.data_in(wire_d75_29),.data_out(wire_d75_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7607531(.data_in(wire_d75_30),.data_out(wire_d75_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7607532(.data_in(wire_d75_31),.data_out(wire_d75_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7607533(.data_in(wire_d75_32),.data_out(wire_d75_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7607534(.data_in(wire_d75_33),.data_out(wire_d75_34),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7607535(.data_in(wire_d75_34),.data_out(wire_d75_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7607536(.data_in(wire_d75_35),.data_out(wire_d75_36),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7607537(.data_in(wire_d75_36),.data_out(wire_d75_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7607538(.data_in(wire_d75_37),.data_out(wire_d75_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7607539(.data_in(wire_d75_38),.data_out(wire_d75_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7607540(.data_in(wire_d75_39),.data_out(wire_d75_40),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7607541(.data_in(wire_d75_40),.data_out(wire_d75_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7607542(.data_in(wire_d75_41),.data_out(wire_d75_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7607543(.data_in(wire_d75_42),.data_out(wire_d75_43),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7607544(.data_in(wire_d75_43),.data_out(wire_d75_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7607545(.data_in(wire_d75_44),.data_out(wire_d75_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7607546(.data_in(wire_d75_45),.data_out(wire_d75_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7607547(.data_in(wire_d75_46),.data_out(wire_d75_47),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7607548(.data_in(wire_d75_47),.data_out(wire_d75_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7607549(.data_in(wire_d75_48),.data_out(wire_d75_49),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7607550(.data_in(wire_d75_49),.data_out(wire_d75_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7607551(.data_in(wire_d75_50),.data_out(wire_d75_51),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7607552(.data_in(wire_d75_51),.data_out(wire_d75_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7607553(.data_in(wire_d75_52),.data_out(wire_d75_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7607554(.data_in(wire_d75_53),.data_out(wire_d75_54),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7607555(.data_in(wire_d75_54),.data_out(wire_d75_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7607556(.data_in(wire_d75_55),.data_out(wire_d75_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7607557(.data_in(wire_d75_56),.data_out(wire_d75_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7607558(.data_in(wire_d75_57),.data_out(wire_d75_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7607559(.data_in(wire_d75_58),.data_out(wire_d75_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7607560(.data_in(wire_d75_59),.data_out(wire_d75_60),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7607561(.data_in(wire_d75_60),.data_out(wire_d75_61),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7607562(.data_in(wire_d75_61),.data_out(wire_d75_62),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7607563(.data_in(wire_d75_62),.data_out(wire_d75_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7607564(.data_in(wire_d75_63),.data_out(wire_d75_64),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7607565(.data_in(wire_d75_64),.data_out(wire_d75_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7607566(.data_in(wire_d75_65),.data_out(wire_d75_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7607567(.data_in(wire_d75_66),.data_out(wire_d75_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7607568(.data_in(wire_d75_67),.data_out(wire_d75_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7607569(.data_in(wire_d75_68),.data_out(wire_d75_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7607570(.data_in(wire_d75_69),.data_out(wire_d75_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7607571(.data_in(wire_d75_70),.data_out(wire_d75_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7607572(.data_in(wire_d75_71),.data_out(wire_d75_72),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7607573(.data_in(wire_d75_72),.data_out(wire_d75_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7607574(.data_in(wire_d75_73),.data_out(wire_d75_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7607575(.data_in(wire_d75_74),.data_out(wire_d75_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7607576(.data_in(wire_d75_75),.data_out(wire_d75_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7607577(.data_in(wire_d75_76),.data_out(wire_d75_77),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7607578(.data_in(wire_d75_77),.data_out(wire_d75_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7607579(.data_in(wire_d75_78),.data_out(wire_d75_79),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7607580(.data_in(wire_d75_79),.data_out(wire_d75_80),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7607581(.data_in(wire_d75_80),.data_out(wire_d75_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7607582(.data_in(wire_d75_81),.data_out(wire_d75_82),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7607583(.data_in(wire_d75_82),.data_out(wire_d75_83),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7607584(.data_in(wire_d75_83),.data_out(wire_d75_84),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7607585(.data_in(wire_d75_84),.data_out(wire_d75_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7607586(.data_in(wire_d75_85),.data_out(wire_d75_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7607587(.data_in(wire_d75_86),.data_out(wire_d75_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7607588(.data_in(wire_d75_87),.data_out(wire_d75_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7607589(.data_in(wire_d75_88),.data_out(wire_d75_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7607590(.data_in(wire_d75_89),.data_out(wire_d75_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7607591(.data_in(wire_d75_90),.data_out(wire_d75_91),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7607592(.data_in(wire_d75_91),.data_out(wire_d75_92),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7607593(.data_in(wire_d75_92),.data_out(wire_d75_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7607594(.data_in(wire_d75_93),.data_out(wire_d75_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7607595(.data_in(wire_d75_94),.data_out(wire_d75_95),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7607596(.data_in(wire_d75_95),.data_out(wire_d75_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7607597(.data_in(wire_d75_96),.data_out(wire_d75_97),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7607598(.data_in(wire_d75_97),.data_out(wire_d75_98),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7607599(.data_in(wire_d75_98),.data_out(wire_d75_99),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance76075100(.data_in(wire_d75_99),.data_out(wire_d75_100),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance76075101(.data_in(wire_d75_100),.data_out(wire_d75_101),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance76075102(.data_in(wire_d75_101),.data_out(wire_d75_102),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance76075103(.data_in(wire_d75_102),.data_out(wire_d75_103),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance76075104(.data_in(wire_d75_103),.data_out(wire_d75_104),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance76075105(.data_in(wire_d75_104),.data_out(wire_d75_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76075106(.data_in(wire_d75_105),.data_out(wire_d75_106),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance76075107(.data_in(wire_d75_106),.data_out(wire_d75_107),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance76075108(.data_in(wire_d75_107),.data_out(wire_d75_108),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance76075109(.data_in(wire_d75_108),.data_out(wire_d75_109),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance76075110(.data_in(wire_d75_109),.data_out(wire_d75_110),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance76075111(.data_in(wire_d75_110),.data_out(wire_d75_111),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance76075112(.data_in(wire_d75_111),.data_out(wire_d75_112),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance76075113(.data_in(wire_d75_112),.data_out(wire_d75_113),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance76075114(.data_in(wire_d75_113),.data_out(wire_d75_114),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance76075115(.data_in(wire_d75_114),.data_out(wire_d75_115),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance76075116(.data_in(wire_d75_115),.data_out(wire_d75_116),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76075117(.data_in(wire_d75_116),.data_out(wire_d75_117),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance76075118(.data_in(wire_d75_117),.data_out(wire_d75_118),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance76075119(.data_in(wire_d75_118),.data_out(d_out75),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance770760(.data_in(d_in76),.data_out(wire_d76_0),.clk(clk),.rst(rst));            //channel 77
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance770761(.data_in(wire_d76_0),.data_out(wire_d76_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance770762(.data_in(wire_d76_1),.data_out(wire_d76_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance770763(.data_in(wire_d76_2),.data_out(wire_d76_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance770764(.data_in(wire_d76_3),.data_out(wire_d76_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance770765(.data_in(wire_d76_4),.data_out(wire_d76_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance770766(.data_in(wire_d76_5),.data_out(wire_d76_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance770767(.data_in(wire_d76_6),.data_out(wire_d76_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance770768(.data_in(wire_d76_7),.data_out(wire_d76_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance770769(.data_in(wire_d76_8),.data_out(wire_d76_9),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7707610(.data_in(wire_d76_9),.data_out(wire_d76_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7707611(.data_in(wire_d76_10),.data_out(wire_d76_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7707612(.data_in(wire_d76_11),.data_out(wire_d76_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7707613(.data_in(wire_d76_12),.data_out(wire_d76_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7707614(.data_in(wire_d76_13),.data_out(wire_d76_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7707615(.data_in(wire_d76_14),.data_out(wire_d76_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7707616(.data_in(wire_d76_15),.data_out(wire_d76_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7707617(.data_in(wire_d76_16),.data_out(wire_d76_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7707618(.data_in(wire_d76_17),.data_out(wire_d76_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7707619(.data_in(wire_d76_18),.data_out(wire_d76_19),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7707620(.data_in(wire_d76_19),.data_out(wire_d76_20),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7707621(.data_in(wire_d76_20),.data_out(wire_d76_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7707622(.data_in(wire_d76_21),.data_out(wire_d76_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7707623(.data_in(wire_d76_22),.data_out(wire_d76_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7707624(.data_in(wire_d76_23),.data_out(wire_d76_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7707625(.data_in(wire_d76_24),.data_out(wire_d76_25),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7707626(.data_in(wire_d76_25),.data_out(wire_d76_26),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7707627(.data_in(wire_d76_26),.data_out(wire_d76_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7707628(.data_in(wire_d76_27),.data_out(wire_d76_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7707629(.data_in(wire_d76_28),.data_out(wire_d76_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7707630(.data_in(wire_d76_29),.data_out(wire_d76_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7707631(.data_in(wire_d76_30),.data_out(wire_d76_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7707632(.data_in(wire_d76_31),.data_out(wire_d76_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7707633(.data_in(wire_d76_32),.data_out(wire_d76_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7707634(.data_in(wire_d76_33),.data_out(wire_d76_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7707635(.data_in(wire_d76_34),.data_out(wire_d76_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7707636(.data_in(wire_d76_35),.data_out(wire_d76_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7707637(.data_in(wire_d76_36),.data_out(wire_d76_37),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7707638(.data_in(wire_d76_37),.data_out(wire_d76_38),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7707639(.data_in(wire_d76_38),.data_out(wire_d76_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7707640(.data_in(wire_d76_39),.data_out(wire_d76_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7707641(.data_in(wire_d76_40),.data_out(wire_d76_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7707642(.data_in(wire_d76_41),.data_out(wire_d76_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7707643(.data_in(wire_d76_42),.data_out(wire_d76_43),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7707644(.data_in(wire_d76_43),.data_out(wire_d76_44),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7707645(.data_in(wire_d76_44),.data_out(wire_d76_45),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7707646(.data_in(wire_d76_45),.data_out(wire_d76_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7707647(.data_in(wire_d76_46),.data_out(wire_d76_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7707648(.data_in(wire_d76_47),.data_out(wire_d76_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7707649(.data_in(wire_d76_48),.data_out(wire_d76_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7707650(.data_in(wire_d76_49),.data_out(wire_d76_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7707651(.data_in(wire_d76_50),.data_out(wire_d76_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7707652(.data_in(wire_d76_51),.data_out(wire_d76_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7707653(.data_in(wire_d76_52),.data_out(wire_d76_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7707654(.data_in(wire_d76_53),.data_out(wire_d76_54),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7707655(.data_in(wire_d76_54),.data_out(wire_d76_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7707656(.data_in(wire_d76_55),.data_out(wire_d76_56),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7707657(.data_in(wire_d76_56),.data_out(wire_d76_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7707658(.data_in(wire_d76_57),.data_out(wire_d76_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7707659(.data_in(wire_d76_58),.data_out(wire_d76_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7707660(.data_in(wire_d76_59),.data_out(wire_d76_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7707661(.data_in(wire_d76_60),.data_out(wire_d76_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7707662(.data_in(wire_d76_61),.data_out(wire_d76_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7707663(.data_in(wire_d76_62),.data_out(wire_d76_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7707664(.data_in(wire_d76_63),.data_out(wire_d76_64),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7707665(.data_in(wire_d76_64),.data_out(wire_d76_65),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7707666(.data_in(wire_d76_65),.data_out(wire_d76_66),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7707667(.data_in(wire_d76_66),.data_out(wire_d76_67),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7707668(.data_in(wire_d76_67),.data_out(wire_d76_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7707669(.data_in(wire_d76_68),.data_out(wire_d76_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7707670(.data_in(wire_d76_69),.data_out(wire_d76_70),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7707671(.data_in(wire_d76_70),.data_out(wire_d76_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7707672(.data_in(wire_d76_71),.data_out(wire_d76_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7707673(.data_in(wire_d76_72),.data_out(wire_d76_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7707674(.data_in(wire_d76_73),.data_out(wire_d76_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7707675(.data_in(wire_d76_74),.data_out(wire_d76_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7707676(.data_in(wire_d76_75),.data_out(wire_d76_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7707677(.data_in(wire_d76_76),.data_out(wire_d76_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7707678(.data_in(wire_d76_77),.data_out(wire_d76_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7707679(.data_in(wire_d76_78),.data_out(wire_d76_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7707680(.data_in(wire_d76_79),.data_out(wire_d76_80),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7707681(.data_in(wire_d76_80),.data_out(wire_d76_81),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7707682(.data_in(wire_d76_81),.data_out(wire_d76_82),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7707683(.data_in(wire_d76_82),.data_out(wire_d76_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7707684(.data_in(wire_d76_83),.data_out(wire_d76_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7707685(.data_in(wire_d76_84),.data_out(wire_d76_85),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7707686(.data_in(wire_d76_85),.data_out(wire_d76_86),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7707687(.data_in(wire_d76_86),.data_out(wire_d76_87),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7707688(.data_in(wire_d76_87),.data_out(wire_d76_88),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7707689(.data_in(wire_d76_88),.data_out(wire_d76_89),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7707690(.data_in(wire_d76_89),.data_out(wire_d76_90),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7707691(.data_in(wire_d76_90),.data_out(wire_d76_91),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7707692(.data_in(wire_d76_91),.data_out(wire_d76_92),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7707693(.data_in(wire_d76_92),.data_out(wire_d76_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7707694(.data_in(wire_d76_93),.data_out(wire_d76_94),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7707695(.data_in(wire_d76_94),.data_out(wire_d76_95),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7707696(.data_in(wire_d76_95),.data_out(wire_d76_96),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7707697(.data_in(wire_d76_96),.data_out(wire_d76_97),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7707698(.data_in(wire_d76_97),.data_out(wire_d76_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7707699(.data_in(wire_d76_98),.data_out(wire_d76_99),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance77076100(.data_in(wire_d76_99),.data_out(wire_d76_100),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance77076101(.data_in(wire_d76_100),.data_out(wire_d76_101),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance77076102(.data_in(wire_d76_101),.data_out(wire_d76_102),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance77076103(.data_in(wire_d76_102),.data_out(wire_d76_103),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance77076104(.data_in(wire_d76_103),.data_out(wire_d76_104),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance77076105(.data_in(wire_d76_104),.data_out(wire_d76_105),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance77076106(.data_in(wire_d76_105),.data_out(wire_d76_106),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance77076107(.data_in(wire_d76_106),.data_out(wire_d76_107),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance77076108(.data_in(wire_d76_107),.data_out(wire_d76_108),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance77076109(.data_in(wire_d76_108),.data_out(wire_d76_109),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance77076110(.data_in(wire_d76_109),.data_out(wire_d76_110),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance77076111(.data_in(wire_d76_110),.data_out(wire_d76_111),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance77076112(.data_in(wire_d76_111),.data_out(wire_d76_112),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance77076113(.data_in(wire_d76_112),.data_out(wire_d76_113),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance77076114(.data_in(wire_d76_113),.data_out(wire_d76_114),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance77076115(.data_in(wire_d76_114),.data_out(wire_d76_115),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance77076116(.data_in(wire_d76_115),.data_out(wire_d76_116),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance77076117(.data_in(wire_d76_116),.data_out(wire_d76_117),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance77076118(.data_in(wire_d76_117),.data_out(wire_d76_118),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance77076119(.data_in(wire_d76_118),.data_out(d_out76),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance780770(.data_in(d_in77),.data_out(wire_d77_0),.clk(clk),.rst(rst));            //channel 78
	encoder #(.WIDTH(WIDTH)) encoder_instance780771(.data_in(wire_d77_0),.data_out(wire_d77_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance780772(.data_in(wire_d77_1),.data_out(wire_d77_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance780773(.data_in(wire_d77_2),.data_out(wire_d77_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance780774(.data_in(wire_d77_3),.data_out(wire_d77_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance780775(.data_in(wire_d77_4),.data_out(wire_d77_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance780776(.data_in(wire_d77_5),.data_out(wire_d77_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance780777(.data_in(wire_d77_6),.data_out(wire_d77_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance780778(.data_in(wire_d77_7),.data_out(wire_d77_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance780779(.data_in(wire_d77_8),.data_out(wire_d77_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7807710(.data_in(wire_d77_9),.data_out(wire_d77_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7807711(.data_in(wire_d77_10),.data_out(wire_d77_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7807712(.data_in(wire_d77_11),.data_out(wire_d77_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7807713(.data_in(wire_d77_12),.data_out(wire_d77_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7807714(.data_in(wire_d77_13),.data_out(wire_d77_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7807715(.data_in(wire_d77_14),.data_out(wire_d77_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7807716(.data_in(wire_d77_15),.data_out(wire_d77_16),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7807717(.data_in(wire_d77_16),.data_out(wire_d77_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7807718(.data_in(wire_d77_17),.data_out(wire_d77_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7807719(.data_in(wire_d77_18),.data_out(wire_d77_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7807720(.data_in(wire_d77_19),.data_out(wire_d77_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7807721(.data_in(wire_d77_20),.data_out(wire_d77_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7807722(.data_in(wire_d77_21),.data_out(wire_d77_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7807723(.data_in(wire_d77_22),.data_out(wire_d77_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7807724(.data_in(wire_d77_23),.data_out(wire_d77_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7807725(.data_in(wire_d77_24),.data_out(wire_d77_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7807726(.data_in(wire_d77_25),.data_out(wire_d77_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7807727(.data_in(wire_d77_26),.data_out(wire_d77_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7807728(.data_in(wire_d77_27),.data_out(wire_d77_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7807729(.data_in(wire_d77_28),.data_out(wire_d77_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7807730(.data_in(wire_d77_29),.data_out(wire_d77_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7807731(.data_in(wire_d77_30),.data_out(wire_d77_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7807732(.data_in(wire_d77_31),.data_out(wire_d77_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7807733(.data_in(wire_d77_32),.data_out(wire_d77_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7807734(.data_in(wire_d77_33),.data_out(wire_d77_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7807735(.data_in(wire_d77_34),.data_out(wire_d77_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7807736(.data_in(wire_d77_35),.data_out(wire_d77_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7807737(.data_in(wire_d77_36),.data_out(wire_d77_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7807738(.data_in(wire_d77_37),.data_out(wire_d77_38),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7807739(.data_in(wire_d77_38),.data_out(wire_d77_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7807740(.data_in(wire_d77_39),.data_out(wire_d77_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7807741(.data_in(wire_d77_40),.data_out(wire_d77_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7807742(.data_in(wire_d77_41),.data_out(wire_d77_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7807743(.data_in(wire_d77_42),.data_out(wire_d77_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7807744(.data_in(wire_d77_43),.data_out(wire_d77_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7807745(.data_in(wire_d77_44),.data_out(wire_d77_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7807746(.data_in(wire_d77_45),.data_out(wire_d77_46),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7807747(.data_in(wire_d77_46),.data_out(wire_d77_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7807748(.data_in(wire_d77_47),.data_out(wire_d77_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7807749(.data_in(wire_d77_48),.data_out(wire_d77_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7807750(.data_in(wire_d77_49),.data_out(wire_d77_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7807751(.data_in(wire_d77_50),.data_out(wire_d77_51),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7807752(.data_in(wire_d77_51),.data_out(wire_d77_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7807753(.data_in(wire_d77_52),.data_out(wire_d77_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7807754(.data_in(wire_d77_53),.data_out(wire_d77_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7807755(.data_in(wire_d77_54),.data_out(wire_d77_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7807756(.data_in(wire_d77_55),.data_out(wire_d77_56),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7807757(.data_in(wire_d77_56),.data_out(wire_d77_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7807758(.data_in(wire_d77_57),.data_out(wire_d77_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7807759(.data_in(wire_d77_58),.data_out(wire_d77_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7807760(.data_in(wire_d77_59),.data_out(wire_d77_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7807761(.data_in(wire_d77_60),.data_out(wire_d77_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7807762(.data_in(wire_d77_61),.data_out(wire_d77_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7807763(.data_in(wire_d77_62),.data_out(wire_d77_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7807764(.data_in(wire_d77_63),.data_out(wire_d77_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7807765(.data_in(wire_d77_64),.data_out(wire_d77_65),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7807766(.data_in(wire_d77_65),.data_out(wire_d77_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7807767(.data_in(wire_d77_66),.data_out(wire_d77_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7807768(.data_in(wire_d77_67),.data_out(wire_d77_68),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7807769(.data_in(wire_d77_68),.data_out(wire_d77_69),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7807770(.data_in(wire_d77_69),.data_out(wire_d77_70),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7807771(.data_in(wire_d77_70),.data_out(wire_d77_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7807772(.data_in(wire_d77_71),.data_out(wire_d77_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7807773(.data_in(wire_d77_72),.data_out(wire_d77_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7807774(.data_in(wire_d77_73),.data_out(wire_d77_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7807775(.data_in(wire_d77_74),.data_out(wire_d77_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7807776(.data_in(wire_d77_75),.data_out(wire_d77_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7807777(.data_in(wire_d77_76),.data_out(wire_d77_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7807778(.data_in(wire_d77_77),.data_out(wire_d77_78),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7807779(.data_in(wire_d77_78),.data_out(wire_d77_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7807780(.data_in(wire_d77_79),.data_out(wire_d77_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7807781(.data_in(wire_d77_80),.data_out(wire_d77_81),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7807782(.data_in(wire_d77_81),.data_out(wire_d77_82),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7807783(.data_in(wire_d77_82),.data_out(wire_d77_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7807784(.data_in(wire_d77_83),.data_out(wire_d77_84),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7807785(.data_in(wire_d77_84),.data_out(wire_d77_85),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7807786(.data_in(wire_d77_85),.data_out(wire_d77_86),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7807787(.data_in(wire_d77_86),.data_out(wire_d77_87),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7807788(.data_in(wire_d77_87),.data_out(wire_d77_88),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7807789(.data_in(wire_d77_88),.data_out(wire_d77_89),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7807790(.data_in(wire_d77_89),.data_out(wire_d77_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7807791(.data_in(wire_d77_90),.data_out(wire_d77_91),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7807792(.data_in(wire_d77_91),.data_out(wire_d77_92),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7807793(.data_in(wire_d77_92),.data_out(wire_d77_93),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7807794(.data_in(wire_d77_93),.data_out(wire_d77_94),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7807795(.data_in(wire_d77_94),.data_out(wire_d77_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7807796(.data_in(wire_d77_95),.data_out(wire_d77_96),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7807797(.data_in(wire_d77_96),.data_out(wire_d77_97),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7807798(.data_in(wire_d77_97),.data_out(wire_d77_98),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7807799(.data_in(wire_d77_98),.data_out(wire_d77_99),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance78077100(.data_in(wire_d77_99),.data_out(wire_d77_100),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance78077101(.data_in(wire_d77_100),.data_out(wire_d77_101),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance78077102(.data_in(wire_d77_101),.data_out(wire_d77_102),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance78077103(.data_in(wire_d77_102),.data_out(wire_d77_103),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance78077104(.data_in(wire_d77_103),.data_out(wire_d77_104),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance78077105(.data_in(wire_d77_104),.data_out(wire_d77_105),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance78077106(.data_in(wire_d77_105),.data_out(wire_d77_106),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance78077107(.data_in(wire_d77_106),.data_out(wire_d77_107),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance78077108(.data_in(wire_d77_107),.data_out(wire_d77_108),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance78077109(.data_in(wire_d77_108),.data_out(wire_d77_109),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance78077110(.data_in(wire_d77_109),.data_out(wire_d77_110),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance78077111(.data_in(wire_d77_110),.data_out(wire_d77_111),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance78077112(.data_in(wire_d77_111),.data_out(wire_d77_112),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance78077113(.data_in(wire_d77_112),.data_out(wire_d77_113),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance78077114(.data_in(wire_d77_113),.data_out(wire_d77_114),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance78077115(.data_in(wire_d77_114),.data_out(wire_d77_115),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance78077116(.data_in(wire_d77_115),.data_out(wire_d77_116),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance78077117(.data_in(wire_d77_116),.data_out(wire_d77_117),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance78077118(.data_in(wire_d77_117),.data_out(wire_d77_118),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance78077119(.data_in(wire_d77_118),.data_out(d_out77),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance790780(.data_in(d_in78),.data_out(wire_d78_0),.clk(clk),.rst(rst));            //channel 79
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance790781(.data_in(wire_d78_0),.data_out(wire_d78_1),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance790782(.data_in(wire_d78_1),.data_out(wire_d78_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance790783(.data_in(wire_d78_2),.data_out(wire_d78_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance790784(.data_in(wire_d78_3),.data_out(wire_d78_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance790785(.data_in(wire_d78_4),.data_out(wire_d78_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance790786(.data_in(wire_d78_5),.data_out(wire_d78_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance790787(.data_in(wire_d78_6),.data_out(wire_d78_7),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance790788(.data_in(wire_d78_7),.data_out(wire_d78_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance790789(.data_in(wire_d78_8),.data_out(wire_d78_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7907810(.data_in(wire_d78_9),.data_out(wire_d78_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7907811(.data_in(wire_d78_10),.data_out(wire_d78_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7907812(.data_in(wire_d78_11),.data_out(wire_d78_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7907813(.data_in(wire_d78_12),.data_out(wire_d78_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7907814(.data_in(wire_d78_13),.data_out(wire_d78_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7907815(.data_in(wire_d78_14),.data_out(wire_d78_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7907816(.data_in(wire_d78_15),.data_out(wire_d78_16),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7907817(.data_in(wire_d78_16),.data_out(wire_d78_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7907818(.data_in(wire_d78_17),.data_out(wire_d78_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7907819(.data_in(wire_d78_18),.data_out(wire_d78_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7907820(.data_in(wire_d78_19),.data_out(wire_d78_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7907821(.data_in(wire_d78_20),.data_out(wire_d78_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7907822(.data_in(wire_d78_21),.data_out(wire_d78_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7907823(.data_in(wire_d78_22),.data_out(wire_d78_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7907824(.data_in(wire_d78_23),.data_out(wire_d78_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7907825(.data_in(wire_d78_24),.data_out(wire_d78_25),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7907826(.data_in(wire_d78_25),.data_out(wire_d78_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7907827(.data_in(wire_d78_26),.data_out(wire_d78_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7907828(.data_in(wire_d78_27),.data_out(wire_d78_28),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7907829(.data_in(wire_d78_28),.data_out(wire_d78_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7907830(.data_in(wire_d78_29),.data_out(wire_d78_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7907831(.data_in(wire_d78_30),.data_out(wire_d78_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7907832(.data_in(wire_d78_31),.data_out(wire_d78_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7907833(.data_in(wire_d78_32),.data_out(wire_d78_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7907834(.data_in(wire_d78_33),.data_out(wire_d78_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7907835(.data_in(wire_d78_34),.data_out(wire_d78_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7907836(.data_in(wire_d78_35),.data_out(wire_d78_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7907837(.data_in(wire_d78_36),.data_out(wire_d78_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7907838(.data_in(wire_d78_37),.data_out(wire_d78_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7907839(.data_in(wire_d78_38),.data_out(wire_d78_39),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7907840(.data_in(wire_d78_39),.data_out(wire_d78_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7907841(.data_in(wire_d78_40),.data_out(wire_d78_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7907842(.data_in(wire_d78_41),.data_out(wire_d78_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7907843(.data_in(wire_d78_42),.data_out(wire_d78_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7907844(.data_in(wire_d78_43),.data_out(wire_d78_44),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7907845(.data_in(wire_d78_44),.data_out(wire_d78_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7907846(.data_in(wire_d78_45),.data_out(wire_d78_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7907847(.data_in(wire_d78_46),.data_out(wire_d78_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7907848(.data_in(wire_d78_47),.data_out(wire_d78_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7907849(.data_in(wire_d78_48),.data_out(wire_d78_49),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7907850(.data_in(wire_d78_49),.data_out(wire_d78_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7907851(.data_in(wire_d78_50),.data_out(wire_d78_51),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7907852(.data_in(wire_d78_51),.data_out(wire_d78_52),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7907853(.data_in(wire_d78_52),.data_out(wire_d78_53),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7907854(.data_in(wire_d78_53),.data_out(wire_d78_54),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7907855(.data_in(wire_d78_54),.data_out(wire_d78_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7907856(.data_in(wire_d78_55),.data_out(wire_d78_56),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7907857(.data_in(wire_d78_56),.data_out(wire_d78_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7907858(.data_in(wire_d78_57),.data_out(wire_d78_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7907859(.data_in(wire_d78_58),.data_out(wire_d78_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7907860(.data_in(wire_d78_59),.data_out(wire_d78_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7907861(.data_in(wire_d78_60),.data_out(wire_d78_61),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7907862(.data_in(wire_d78_61),.data_out(wire_d78_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7907863(.data_in(wire_d78_62),.data_out(wire_d78_63),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7907864(.data_in(wire_d78_63),.data_out(wire_d78_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7907865(.data_in(wire_d78_64),.data_out(wire_d78_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7907866(.data_in(wire_d78_65),.data_out(wire_d78_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7907867(.data_in(wire_d78_66),.data_out(wire_d78_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7907868(.data_in(wire_d78_67),.data_out(wire_d78_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7907869(.data_in(wire_d78_68),.data_out(wire_d78_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7907870(.data_in(wire_d78_69),.data_out(wire_d78_70),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7907871(.data_in(wire_d78_70),.data_out(wire_d78_71),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7907872(.data_in(wire_d78_71),.data_out(wire_d78_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7907873(.data_in(wire_d78_72),.data_out(wire_d78_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7907874(.data_in(wire_d78_73),.data_out(wire_d78_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7907875(.data_in(wire_d78_74),.data_out(wire_d78_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7907876(.data_in(wire_d78_75),.data_out(wire_d78_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7907877(.data_in(wire_d78_76),.data_out(wire_d78_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7907878(.data_in(wire_d78_77),.data_out(wire_d78_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7907879(.data_in(wire_d78_78),.data_out(wire_d78_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7907880(.data_in(wire_d78_79),.data_out(wire_d78_80),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7907881(.data_in(wire_d78_80),.data_out(wire_d78_81),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7907882(.data_in(wire_d78_81),.data_out(wire_d78_82),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7907883(.data_in(wire_d78_82),.data_out(wire_d78_83),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7907884(.data_in(wire_d78_83),.data_out(wire_d78_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7907885(.data_in(wire_d78_84),.data_out(wire_d78_85),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7907886(.data_in(wire_d78_85),.data_out(wire_d78_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7907887(.data_in(wire_d78_86),.data_out(wire_d78_87),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7907888(.data_in(wire_d78_87),.data_out(wire_d78_88),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7907889(.data_in(wire_d78_88),.data_out(wire_d78_89),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7907890(.data_in(wire_d78_89),.data_out(wire_d78_90),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7907891(.data_in(wire_d78_90),.data_out(wire_d78_91),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7907892(.data_in(wire_d78_91),.data_out(wire_d78_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7907893(.data_in(wire_d78_92),.data_out(wire_d78_93),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7907894(.data_in(wire_d78_93),.data_out(wire_d78_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7907895(.data_in(wire_d78_94),.data_out(wire_d78_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7907896(.data_in(wire_d78_95),.data_out(wire_d78_96),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7907897(.data_in(wire_d78_96),.data_out(wire_d78_97),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7907898(.data_in(wire_d78_97),.data_out(wire_d78_98),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7907899(.data_in(wire_d78_98),.data_out(wire_d78_99),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance79078100(.data_in(wire_d78_99),.data_out(wire_d78_100),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance79078101(.data_in(wire_d78_100),.data_out(wire_d78_101),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance79078102(.data_in(wire_d78_101),.data_out(wire_d78_102),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance79078103(.data_in(wire_d78_102),.data_out(wire_d78_103),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance79078104(.data_in(wire_d78_103),.data_out(wire_d78_104),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance79078105(.data_in(wire_d78_104),.data_out(wire_d78_105),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance79078106(.data_in(wire_d78_105),.data_out(wire_d78_106),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance79078107(.data_in(wire_d78_106),.data_out(wire_d78_107),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance79078108(.data_in(wire_d78_107),.data_out(wire_d78_108),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance79078109(.data_in(wire_d78_108),.data_out(wire_d78_109),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance79078110(.data_in(wire_d78_109),.data_out(wire_d78_110),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance79078111(.data_in(wire_d78_110),.data_out(wire_d78_111),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance79078112(.data_in(wire_d78_111),.data_out(wire_d78_112),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance79078113(.data_in(wire_d78_112),.data_out(wire_d78_113),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance79078114(.data_in(wire_d78_113),.data_out(wire_d78_114),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance79078115(.data_in(wire_d78_114),.data_out(wire_d78_115),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance79078116(.data_in(wire_d78_115),.data_out(wire_d78_116),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance79078117(.data_in(wire_d78_116),.data_out(wire_d78_117),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance79078118(.data_in(wire_d78_117),.data_out(wire_d78_118),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance79078119(.data_in(wire_d78_118),.data_out(d_out78),.clk(clk),.rst(rst));

	large_adder #(.WIDTH(WIDTH)) large_adder_instance800790(.data_in(d_in79),.data_out(wire_d79_0),.clk(clk),.rst(rst));            //channel 80
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance800791(.data_in(wire_d79_0),.data_out(wire_d79_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance800792(.data_in(wire_d79_1),.data_out(wire_d79_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance800793(.data_in(wire_d79_2),.data_out(wire_d79_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance800794(.data_in(wire_d79_3),.data_out(wire_d79_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance800795(.data_in(wire_d79_4),.data_out(wire_d79_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance800796(.data_in(wire_d79_5),.data_out(wire_d79_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance800797(.data_in(wire_d79_6),.data_out(wire_d79_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance800798(.data_in(wire_d79_7),.data_out(wire_d79_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance800799(.data_in(wire_d79_8),.data_out(wire_d79_9),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8007910(.data_in(wire_d79_9),.data_out(wire_d79_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8007911(.data_in(wire_d79_10),.data_out(wire_d79_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8007912(.data_in(wire_d79_11),.data_out(wire_d79_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8007913(.data_in(wire_d79_12),.data_out(wire_d79_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8007914(.data_in(wire_d79_13),.data_out(wire_d79_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8007915(.data_in(wire_d79_14),.data_out(wire_d79_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8007916(.data_in(wire_d79_15),.data_out(wire_d79_16),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8007917(.data_in(wire_d79_16),.data_out(wire_d79_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8007918(.data_in(wire_d79_17),.data_out(wire_d79_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8007919(.data_in(wire_d79_18),.data_out(wire_d79_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8007920(.data_in(wire_d79_19),.data_out(wire_d79_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8007921(.data_in(wire_d79_20),.data_out(wire_d79_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8007922(.data_in(wire_d79_21),.data_out(wire_d79_22),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8007923(.data_in(wire_d79_22),.data_out(wire_d79_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8007924(.data_in(wire_d79_23),.data_out(wire_d79_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8007925(.data_in(wire_d79_24),.data_out(wire_d79_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8007926(.data_in(wire_d79_25),.data_out(wire_d79_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8007927(.data_in(wire_d79_26),.data_out(wire_d79_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8007928(.data_in(wire_d79_27),.data_out(wire_d79_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8007929(.data_in(wire_d79_28),.data_out(wire_d79_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8007930(.data_in(wire_d79_29),.data_out(wire_d79_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8007931(.data_in(wire_d79_30),.data_out(wire_d79_31),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8007932(.data_in(wire_d79_31),.data_out(wire_d79_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8007933(.data_in(wire_d79_32),.data_out(wire_d79_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8007934(.data_in(wire_d79_33),.data_out(wire_d79_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8007935(.data_in(wire_d79_34),.data_out(wire_d79_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8007936(.data_in(wire_d79_35),.data_out(wire_d79_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8007937(.data_in(wire_d79_36),.data_out(wire_d79_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8007938(.data_in(wire_d79_37),.data_out(wire_d79_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8007939(.data_in(wire_d79_38),.data_out(wire_d79_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8007940(.data_in(wire_d79_39),.data_out(wire_d79_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8007941(.data_in(wire_d79_40),.data_out(wire_d79_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8007942(.data_in(wire_d79_41),.data_out(wire_d79_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8007943(.data_in(wire_d79_42),.data_out(wire_d79_43),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8007944(.data_in(wire_d79_43),.data_out(wire_d79_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8007945(.data_in(wire_d79_44),.data_out(wire_d79_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8007946(.data_in(wire_d79_45),.data_out(wire_d79_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8007947(.data_in(wire_d79_46),.data_out(wire_d79_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8007948(.data_in(wire_d79_47),.data_out(wire_d79_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8007949(.data_in(wire_d79_48),.data_out(wire_d79_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8007950(.data_in(wire_d79_49),.data_out(wire_d79_50),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8007951(.data_in(wire_d79_50),.data_out(wire_d79_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8007952(.data_in(wire_d79_51),.data_out(wire_d79_52),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8007953(.data_in(wire_d79_52),.data_out(wire_d79_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8007954(.data_in(wire_d79_53),.data_out(wire_d79_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8007955(.data_in(wire_d79_54),.data_out(wire_d79_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8007956(.data_in(wire_d79_55),.data_out(wire_d79_56),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8007957(.data_in(wire_d79_56),.data_out(wire_d79_57),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8007958(.data_in(wire_d79_57),.data_out(wire_d79_58),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8007959(.data_in(wire_d79_58),.data_out(wire_d79_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8007960(.data_in(wire_d79_59),.data_out(wire_d79_60),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8007961(.data_in(wire_d79_60),.data_out(wire_d79_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8007962(.data_in(wire_d79_61),.data_out(wire_d79_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8007963(.data_in(wire_d79_62),.data_out(wire_d79_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8007964(.data_in(wire_d79_63),.data_out(wire_d79_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8007965(.data_in(wire_d79_64),.data_out(wire_d79_65),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8007966(.data_in(wire_d79_65),.data_out(wire_d79_66),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8007967(.data_in(wire_d79_66),.data_out(wire_d79_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8007968(.data_in(wire_d79_67),.data_out(wire_d79_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8007969(.data_in(wire_d79_68),.data_out(wire_d79_69),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8007970(.data_in(wire_d79_69),.data_out(wire_d79_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8007971(.data_in(wire_d79_70),.data_out(wire_d79_71),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8007972(.data_in(wire_d79_71),.data_out(wire_d79_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8007973(.data_in(wire_d79_72),.data_out(wire_d79_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8007974(.data_in(wire_d79_73),.data_out(wire_d79_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8007975(.data_in(wire_d79_74),.data_out(wire_d79_75),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8007976(.data_in(wire_d79_75),.data_out(wire_d79_76),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8007977(.data_in(wire_d79_76),.data_out(wire_d79_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8007978(.data_in(wire_d79_77),.data_out(wire_d79_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8007979(.data_in(wire_d79_78),.data_out(wire_d79_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8007980(.data_in(wire_d79_79),.data_out(wire_d79_80),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8007981(.data_in(wire_d79_80),.data_out(wire_d79_81),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8007982(.data_in(wire_d79_81),.data_out(wire_d79_82),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8007983(.data_in(wire_d79_82),.data_out(wire_d79_83),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8007984(.data_in(wire_d79_83),.data_out(wire_d79_84),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8007985(.data_in(wire_d79_84),.data_out(wire_d79_85),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8007986(.data_in(wire_d79_85),.data_out(wire_d79_86),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8007987(.data_in(wire_d79_86),.data_out(wire_d79_87),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8007988(.data_in(wire_d79_87),.data_out(wire_d79_88),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8007989(.data_in(wire_d79_88),.data_out(wire_d79_89),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8007990(.data_in(wire_d79_89),.data_out(wire_d79_90),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8007991(.data_in(wire_d79_90),.data_out(wire_d79_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8007992(.data_in(wire_d79_91),.data_out(wire_d79_92),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8007993(.data_in(wire_d79_92),.data_out(wire_d79_93),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8007994(.data_in(wire_d79_93),.data_out(wire_d79_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8007995(.data_in(wire_d79_94),.data_out(wire_d79_95),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8007996(.data_in(wire_d79_95),.data_out(wire_d79_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8007997(.data_in(wire_d79_96),.data_out(wire_d79_97),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8007998(.data_in(wire_d79_97),.data_out(wire_d79_98),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8007999(.data_in(wire_d79_98),.data_out(wire_d79_99),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance80079100(.data_in(wire_d79_99),.data_out(wire_d79_100),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance80079101(.data_in(wire_d79_100),.data_out(wire_d79_101),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance80079102(.data_in(wire_d79_101),.data_out(wire_d79_102),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance80079103(.data_in(wire_d79_102),.data_out(wire_d79_103),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance80079104(.data_in(wire_d79_103),.data_out(wire_d79_104),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance80079105(.data_in(wire_d79_104),.data_out(wire_d79_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance80079106(.data_in(wire_d79_105),.data_out(wire_d79_106),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance80079107(.data_in(wire_d79_106),.data_out(wire_d79_107),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance80079108(.data_in(wire_d79_107),.data_out(wire_d79_108),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance80079109(.data_in(wire_d79_108),.data_out(wire_d79_109),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance80079110(.data_in(wire_d79_109),.data_out(wire_d79_110),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance80079111(.data_in(wire_d79_110),.data_out(wire_d79_111),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance80079112(.data_in(wire_d79_111),.data_out(wire_d79_112),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance80079113(.data_in(wire_d79_112),.data_out(wire_d79_113),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance80079114(.data_in(wire_d79_113),.data_out(wire_d79_114),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance80079115(.data_in(wire_d79_114),.data_out(wire_d79_115),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance80079116(.data_in(wire_d79_115),.data_out(wire_d79_116),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance80079117(.data_in(wire_d79_116),.data_out(wire_d79_117),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance80079118(.data_in(wire_d79_117),.data_out(wire_d79_118),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance80079119(.data_in(wire_d79_118),.data_out(d_out79),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance810800(.data_in(d_in80),.data_out(wire_d80_0),.clk(clk),.rst(rst));            //channel 81
	register #(.WIDTH(WIDTH)) register_instance810801(.data_in(wire_d80_0),.data_out(wire_d80_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance810802(.data_in(wire_d80_1),.data_out(wire_d80_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance810803(.data_in(wire_d80_2),.data_out(wire_d80_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance810804(.data_in(wire_d80_3),.data_out(wire_d80_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance810805(.data_in(wire_d80_4),.data_out(wire_d80_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance810806(.data_in(wire_d80_5),.data_out(wire_d80_6),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance810807(.data_in(wire_d80_6),.data_out(wire_d80_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance810808(.data_in(wire_d80_7),.data_out(wire_d80_8),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance810809(.data_in(wire_d80_8),.data_out(wire_d80_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8108010(.data_in(wire_d80_9),.data_out(wire_d80_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8108011(.data_in(wire_d80_10),.data_out(wire_d80_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8108012(.data_in(wire_d80_11),.data_out(wire_d80_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8108013(.data_in(wire_d80_12),.data_out(wire_d80_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8108014(.data_in(wire_d80_13),.data_out(wire_d80_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8108015(.data_in(wire_d80_14),.data_out(wire_d80_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8108016(.data_in(wire_d80_15),.data_out(wire_d80_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8108017(.data_in(wire_d80_16),.data_out(wire_d80_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8108018(.data_in(wire_d80_17),.data_out(wire_d80_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8108019(.data_in(wire_d80_18),.data_out(wire_d80_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8108020(.data_in(wire_d80_19),.data_out(wire_d80_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8108021(.data_in(wire_d80_20),.data_out(wire_d80_21),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8108022(.data_in(wire_d80_21),.data_out(wire_d80_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8108023(.data_in(wire_d80_22),.data_out(wire_d80_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8108024(.data_in(wire_d80_23),.data_out(wire_d80_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8108025(.data_in(wire_d80_24),.data_out(wire_d80_25),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8108026(.data_in(wire_d80_25),.data_out(wire_d80_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8108027(.data_in(wire_d80_26),.data_out(wire_d80_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8108028(.data_in(wire_d80_27),.data_out(wire_d80_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8108029(.data_in(wire_d80_28),.data_out(wire_d80_29),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8108030(.data_in(wire_d80_29),.data_out(wire_d80_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8108031(.data_in(wire_d80_30),.data_out(wire_d80_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8108032(.data_in(wire_d80_31),.data_out(wire_d80_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8108033(.data_in(wire_d80_32),.data_out(wire_d80_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8108034(.data_in(wire_d80_33),.data_out(wire_d80_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8108035(.data_in(wire_d80_34),.data_out(wire_d80_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8108036(.data_in(wire_d80_35),.data_out(wire_d80_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8108037(.data_in(wire_d80_36),.data_out(wire_d80_37),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8108038(.data_in(wire_d80_37),.data_out(wire_d80_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8108039(.data_in(wire_d80_38),.data_out(wire_d80_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8108040(.data_in(wire_d80_39),.data_out(wire_d80_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8108041(.data_in(wire_d80_40),.data_out(wire_d80_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8108042(.data_in(wire_d80_41),.data_out(wire_d80_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8108043(.data_in(wire_d80_42),.data_out(wire_d80_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8108044(.data_in(wire_d80_43),.data_out(wire_d80_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8108045(.data_in(wire_d80_44),.data_out(wire_d80_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8108046(.data_in(wire_d80_45),.data_out(wire_d80_46),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8108047(.data_in(wire_d80_46),.data_out(wire_d80_47),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8108048(.data_in(wire_d80_47),.data_out(wire_d80_48),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8108049(.data_in(wire_d80_48),.data_out(wire_d80_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8108050(.data_in(wire_d80_49),.data_out(wire_d80_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8108051(.data_in(wire_d80_50),.data_out(wire_d80_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8108052(.data_in(wire_d80_51),.data_out(wire_d80_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8108053(.data_in(wire_d80_52),.data_out(wire_d80_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8108054(.data_in(wire_d80_53),.data_out(wire_d80_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8108055(.data_in(wire_d80_54),.data_out(wire_d80_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8108056(.data_in(wire_d80_55),.data_out(wire_d80_56),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8108057(.data_in(wire_d80_56),.data_out(wire_d80_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8108058(.data_in(wire_d80_57),.data_out(wire_d80_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8108059(.data_in(wire_d80_58),.data_out(wire_d80_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8108060(.data_in(wire_d80_59),.data_out(wire_d80_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8108061(.data_in(wire_d80_60),.data_out(wire_d80_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8108062(.data_in(wire_d80_61),.data_out(wire_d80_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8108063(.data_in(wire_d80_62),.data_out(wire_d80_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8108064(.data_in(wire_d80_63),.data_out(wire_d80_64),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8108065(.data_in(wire_d80_64),.data_out(wire_d80_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8108066(.data_in(wire_d80_65),.data_out(wire_d80_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8108067(.data_in(wire_d80_66),.data_out(wire_d80_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8108068(.data_in(wire_d80_67),.data_out(wire_d80_68),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8108069(.data_in(wire_d80_68),.data_out(wire_d80_69),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8108070(.data_in(wire_d80_69),.data_out(wire_d80_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8108071(.data_in(wire_d80_70),.data_out(wire_d80_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8108072(.data_in(wire_d80_71),.data_out(wire_d80_72),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8108073(.data_in(wire_d80_72),.data_out(wire_d80_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8108074(.data_in(wire_d80_73),.data_out(wire_d80_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8108075(.data_in(wire_d80_74),.data_out(wire_d80_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8108076(.data_in(wire_d80_75),.data_out(wire_d80_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8108077(.data_in(wire_d80_76),.data_out(wire_d80_77),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8108078(.data_in(wire_d80_77),.data_out(wire_d80_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8108079(.data_in(wire_d80_78),.data_out(wire_d80_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8108080(.data_in(wire_d80_79),.data_out(wire_d80_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8108081(.data_in(wire_d80_80),.data_out(wire_d80_81),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8108082(.data_in(wire_d80_81),.data_out(wire_d80_82),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8108083(.data_in(wire_d80_82),.data_out(wire_d80_83),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8108084(.data_in(wire_d80_83),.data_out(wire_d80_84),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8108085(.data_in(wire_d80_84),.data_out(wire_d80_85),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8108086(.data_in(wire_d80_85),.data_out(wire_d80_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8108087(.data_in(wire_d80_86),.data_out(wire_d80_87),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8108088(.data_in(wire_d80_87),.data_out(wire_d80_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8108089(.data_in(wire_d80_88),.data_out(wire_d80_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8108090(.data_in(wire_d80_89),.data_out(wire_d80_90),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8108091(.data_in(wire_d80_90),.data_out(wire_d80_91),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8108092(.data_in(wire_d80_91),.data_out(wire_d80_92),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8108093(.data_in(wire_d80_92),.data_out(wire_d80_93),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8108094(.data_in(wire_d80_93),.data_out(wire_d80_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8108095(.data_in(wire_d80_94),.data_out(wire_d80_95),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8108096(.data_in(wire_d80_95),.data_out(wire_d80_96),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8108097(.data_in(wire_d80_96),.data_out(wire_d80_97),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8108098(.data_in(wire_d80_97),.data_out(wire_d80_98),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8108099(.data_in(wire_d80_98),.data_out(wire_d80_99),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance81080100(.data_in(wire_d80_99),.data_out(wire_d80_100),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance81080101(.data_in(wire_d80_100),.data_out(wire_d80_101),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance81080102(.data_in(wire_d80_101),.data_out(wire_d80_102),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance81080103(.data_in(wire_d80_102),.data_out(wire_d80_103),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance81080104(.data_in(wire_d80_103),.data_out(wire_d80_104),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance81080105(.data_in(wire_d80_104),.data_out(wire_d80_105),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance81080106(.data_in(wire_d80_105),.data_out(wire_d80_106),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance81080107(.data_in(wire_d80_106),.data_out(wire_d80_107),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance81080108(.data_in(wire_d80_107),.data_out(wire_d80_108),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance81080109(.data_in(wire_d80_108),.data_out(wire_d80_109),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance81080110(.data_in(wire_d80_109),.data_out(wire_d80_110),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance81080111(.data_in(wire_d80_110),.data_out(wire_d80_111),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance81080112(.data_in(wire_d80_111),.data_out(wire_d80_112),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance81080113(.data_in(wire_d80_112),.data_out(wire_d80_113),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance81080114(.data_in(wire_d80_113),.data_out(wire_d80_114),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance81080115(.data_in(wire_d80_114),.data_out(wire_d80_115),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance81080116(.data_in(wire_d80_115),.data_out(wire_d80_116),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance81080117(.data_in(wire_d80_116),.data_out(wire_d80_117),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance81080118(.data_in(wire_d80_117),.data_out(wire_d80_118),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance81080119(.data_in(wire_d80_118),.data_out(d_out80),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance820810(.data_in(d_in81),.data_out(wire_d81_0),.clk(clk),.rst(rst));            //channel 82
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance820811(.data_in(wire_d81_0),.data_out(wire_d81_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance820812(.data_in(wire_d81_1),.data_out(wire_d81_2),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance820813(.data_in(wire_d81_2),.data_out(wire_d81_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance820814(.data_in(wire_d81_3),.data_out(wire_d81_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance820815(.data_in(wire_d81_4),.data_out(wire_d81_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance820816(.data_in(wire_d81_5),.data_out(wire_d81_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance820817(.data_in(wire_d81_6),.data_out(wire_d81_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance820818(.data_in(wire_d81_7),.data_out(wire_d81_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance820819(.data_in(wire_d81_8),.data_out(wire_d81_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8208110(.data_in(wire_d81_9),.data_out(wire_d81_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8208111(.data_in(wire_d81_10),.data_out(wire_d81_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8208112(.data_in(wire_d81_11),.data_out(wire_d81_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8208113(.data_in(wire_d81_12),.data_out(wire_d81_13),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8208114(.data_in(wire_d81_13),.data_out(wire_d81_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8208115(.data_in(wire_d81_14),.data_out(wire_d81_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8208116(.data_in(wire_d81_15),.data_out(wire_d81_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8208117(.data_in(wire_d81_16),.data_out(wire_d81_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8208118(.data_in(wire_d81_17),.data_out(wire_d81_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8208119(.data_in(wire_d81_18),.data_out(wire_d81_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8208120(.data_in(wire_d81_19),.data_out(wire_d81_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8208121(.data_in(wire_d81_20),.data_out(wire_d81_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8208122(.data_in(wire_d81_21),.data_out(wire_d81_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8208123(.data_in(wire_d81_22),.data_out(wire_d81_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8208124(.data_in(wire_d81_23),.data_out(wire_d81_24),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8208125(.data_in(wire_d81_24),.data_out(wire_d81_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8208126(.data_in(wire_d81_25),.data_out(wire_d81_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8208127(.data_in(wire_d81_26),.data_out(wire_d81_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8208128(.data_in(wire_d81_27),.data_out(wire_d81_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8208129(.data_in(wire_d81_28),.data_out(wire_d81_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8208130(.data_in(wire_d81_29),.data_out(wire_d81_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8208131(.data_in(wire_d81_30),.data_out(wire_d81_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8208132(.data_in(wire_d81_31),.data_out(wire_d81_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8208133(.data_in(wire_d81_32),.data_out(wire_d81_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8208134(.data_in(wire_d81_33),.data_out(wire_d81_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8208135(.data_in(wire_d81_34),.data_out(wire_d81_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8208136(.data_in(wire_d81_35),.data_out(wire_d81_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8208137(.data_in(wire_d81_36),.data_out(wire_d81_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8208138(.data_in(wire_d81_37),.data_out(wire_d81_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8208139(.data_in(wire_d81_38),.data_out(wire_d81_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8208140(.data_in(wire_d81_39),.data_out(wire_d81_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8208141(.data_in(wire_d81_40),.data_out(wire_d81_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8208142(.data_in(wire_d81_41),.data_out(wire_d81_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8208143(.data_in(wire_d81_42),.data_out(wire_d81_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8208144(.data_in(wire_d81_43),.data_out(wire_d81_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8208145(.data_in(wire_d81_44),.data_out(wire_d81_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8208146(.data_in(wire_d81_45),.data_out(wire_d81_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8208147(.data_in(wire_d81_46),.data_out(wire_d81_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8208148(.data_in(wire_d81_47),.data_out(wire_d81_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8208149(.data_in(wire_d81_48),.data_out(wire_d81_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8208150(.data_in(wire_d81_49),.data_out(wire_d81_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8208151(.data_in(wire_d81_50),.data_out(wire_d81_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8208152(.data_in(wire_d81_51),.data_out(wire_d81_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8208153(.data_in(wire_d81_52),.data_out(wire_d81_53),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8208154(.data_in(wire_d81_53),.data_out(wire_d81_54),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8208155(.data_in(wire_d81_54),.data_out(wire_d81_55),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8208156(.data_in(wire_d81_55),.data_out(wire_d81_56),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8208157(.data_in(wire_d81_56),.data_out(wire_d81_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8208158(.data_in(wire_d81_57),.data_out(wire_d81_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8208159(.data_in(wire_d81_58),.data_out(wire_d81_59),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8208160(.data_in(wire_d81_59),.data_out(wire_d81_60),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8208161(.data_in(wire_d81_60),.data_out(wire_d81_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8208162(.data_in(wire_d81_61),.data_out(wire_d81_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8208163(.data_in(wire_d81_62),.data_out(wire_d81_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8208164(.data_in(wire_d81_63),.data_out(wire_d81_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8208165(.data_in(wire_d81_64),.data_out(wire_d81_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8208166(.data_in(wire_d81_65),.data_out(wire_d81_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8208167(.data_in(wire_d81_66),.data_out(wire_d81_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8208168(.data_in(wire_d81_67),.data_out(wire_d81_68),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8208169(.data_in(wire_d81_68),.data_out(wire_d81_69),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8208170(.data_in(wire_d81_69),.data_out(wire_d81_70),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8208171(.data_in(wire_d81_70),.data_out(wire_d81_71),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8208172(.data_in(wire_d81_71),.data_out(wire_d81_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8208173(.data_in(wire_d81_72),.data_out(wire_d81_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8208174(.data_in(wire_d81_73),.data_out(wire_d81_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8208175(.data_in(wire_d81_74),.data_out(wire_d81_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8208176(.data_in(wire_d81_75),.data_out(wire_d81_76),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8208177(.data_in(wire_d81_76),.data_out(wire_d81_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8208178(.data_in(wire_d81_77),.data_out(wire_d81_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8208179(.data_in(wire_d81_78),.data_out(wire_d81_79),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8208180(.data_in(wire_d81_79),.data_out(wire_d81_80),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8208181(.data_in(wire_d81_80),.data_out(wire_d81_81),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8208182(.data_in(wire_d81_81),.data_out(wire_d81_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8208183(.data_in(wire_d81_82),.data_out(wire_d81_83),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8208184(.data_in(wire_d81_83),.data_out(wire_d81_84),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8208185(.data_in(wire_d81_84),.data_out(wire_d81_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8208186(.data_in(wire_d81_85),.data_out(wire_d81_86),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8208187(.data_in(wire_d81_86),.data_out(wire_d81_87),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8208188(.data_in(wire_d81_87),.data_out(wire_d81_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8208189(.data_in(wire_d81_88),.data_out(wire_d81_89),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8208190(.data_in(wire_d81_89),.data_out(wire_d81_90),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8208191(.data_in(wire_d81_90),.data_out(wire_d81_91),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8208192(.data_in(wire_d81_91),.data_out(wire_d81_92),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8208193(.data_in(wire_d81_92),.data_out(wire_d81_93),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8208194(.data_in(wire_d81_93),.data_out(wire_d81_94),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8208195(.data_in(wire_d81_94),.data_out(wire_d81_95),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8208196(.data_in(wire_d81_95),.data_out(wire_d81_96),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8208197(.data_in(wire_d81_96),.data_out(wire_d81_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8208198(.data_in(wire_d81_97),.data_out(wire_d81_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8208199(.data_in(wire_d81_98),.data_out(wire_d81_99),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance82081100(.data_in(wire_d81_99),.data_out(wire_d81_100),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance82081101(.data_in(wire_d81_100),.data_out(wire_d81_101),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance82081102(.data_in(wire_d81_101),.data_out(wire_d81_102),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance82081103(.data_in(wire_d81_102),.data_out(wire_d81_103),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance82081104(.data_in(wire_d81_103),.data_out(wire_d81_104),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance82081105(.data_in(wire_d81_104),.data_out(wire_d81_105),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance82081106(.data_in(wire_d81_105),.data_out(wire_d81_106),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance82081107(.data_in(wire_d81_106),.data_out(wire_d81_107),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance82081108(.data_in(wire_d81_107),.data_out(wire_d81_108),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance82081109(.data_in(wire_d81_108),.data_out(wire_d81_109),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance82081110(.data_in(wire_d81_109),.data_out(wire_d81_110),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance82081111(.data_in(wire_d81_110),.data_out(wire_d81_111),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance82081112(.data_in(wire_d81_111),.data_out(wire_d81_112),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance82081113(.data_in(wire_d81_112),.data_out(wire_d81_113),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance82081114(.data_in(wire_d81_113),.data_out(wire_d81_114),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance82081115(.data_in(wire_d81_114),.data_out(wire_d81_115),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance82081116(.data_in(wire_d81_115),.data_out(wire_d81_116),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance82081117(.data_in(wire_d81_116),.data_out(wire_d81_117),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance82081118(.data_in(wire_d81_117),.data_out(wire_d81_118),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance82081119(.data_in(wire_d81_118),.data_out(d_out81),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance830820(.data_in(d_in82),.data_out(wire_d82_0),.clk(clk),.rst(rst));            //channel 83
	register #(.WIDTH(WIDTH)) register_instance830821(.data_in(wire_d82_0),.data_out(wire_d82_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance830822(.data_in(wire_d82_1),.data_out(wire_d82_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance830823(.data_in(wire_d82_2),.data_out(wire_d82_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance830824(.data_in(wire_d82_3),.data_out(wire_d82_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance830825(.data_in(wire_d82_4),.data_out(wire_d82_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance830826(.data_in(wire_d82_5),.data_out(wire_d82_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance830827(.data_in(wire_d82_6),.data_out(wire_d82_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance830828(.data_in(wire_d82_7),.data_out(wire_d82_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance830829(.data_in(wire_d82_8),.data_out(wire_d82_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8308210(.data_in(wire_d82_9),.data_out(wire_d82_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8308211(.data_in(wire_d82_10),.data_out(wire_d82_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8308212(.data_in(wire_d82_11),.data_out(wire_d82_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8308213(.data_in(wire_d82_12),.data_out(wire_d82_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8308214(.data_in(wire_d82_13),.data_out(wire_d82_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8308215(.data_in(wire_d82_14),.data_out(wire_d82_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8308216(.data_in(wire_d82_15),.data_out(wire_d82_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8308217(.data_in(wire_d82_16),.data_out(wire_d82_17),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8308218(.data_in(wire_d82_17),.data_out(wire_d82_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8308219(.data_in(wire_d82_18),.data_out(wire_d82_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8308220(.data_in(wire_d82_19),.data_out(wire_d82_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8308221(.data_in(wire_d82_20),.data_out(wire_d82_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8308222(.data_in(wire_d82_21),.data_out(wire_d82_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8308223(.data_in(wire_d82_22),.data_out(wire_d82_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8308224(.data_in(wire_d82_23),.data_out(wire_d82_24),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8308225(.data_in(wire_d82_24),.data_out(wire_d82_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8308226(.data_in(wire_d82_25),.data_out(wire_d82_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8308227(.data_in(wire_d82_26),.data_out(wire_d82_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8308228(.data_in(wire_d82_27),.data_out(wire_d82_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8308229(.data_in(wire_d82_28),.data_out(wire_d82_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8308230(.data_in(wire_d82_29),.data_out(wire_d82_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8308231(.data_in(wire_d82_30),.data_out(wire_d82_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8308232(.data_in(wire_d82_31),.data_out(wire_d82_32),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8308233(.data_in(wire_d82_32),.data_out(wire_d82_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8308234(.data_in(wire_d82_33),.data_out(wire_d82_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8308235(.data_in(wire_d82_34),.data_out(wire_d82_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8308236(.data_in(wire_d82_35),.data_out(wire_d82_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8308237(.data_in(wire_d82_36),.data_out(wire_d82_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8308238(.data_in(wire_d82_37),.data_out(wire_d82_38),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8308239(.data_in(wire_d82_38),.data_out(wire_d82_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8308240(.data_in(wire_d82_39),.data_out(wire_d82_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8308241(.data_in(wire_d82_40),.data_out(wire_d82_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8308242(.data_in(wire_d82_41),.data_out(wire_d82_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8308243(.data_in(wire_d82_42),.data_out(wire_d82_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8308244(.data_in(wire_d82_43),.data_out(wire_d82_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8308245(.data_in(wire_d82_44),.data_out(wire_d82_45),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8308246(.data_in(wire_d82_45),.data_out(wire_d82_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8308247(.data_in(wire_d82_46),.data_out(wire_d82_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8308248(.data_in(wire_d82_47),.data_out(wire_d82_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8308249(.data_in(wire_d82_48),.data_out(wire_d82_49),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8308250(.data_in(wire_d82_49),.data_out(wire_d82_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8308251(.data_in(wire_d82_50),.data_out(wire_d82_51),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8308252(.data_in(wire_d82_51),.data_out(wire_d82_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8308253(.data_in(wire_d82_52),.data_out(wire_d82_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8308254(.data_in(wire_d82_53),.data_out(wire_d82_54),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8308255(.data_in(wire_d82_54),.data_out(wire_d82_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8308256(.data_in(wire_d82_55),.data_out(wire_d82_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8308257(.data_in(wire_d82_56),.data_out(wire_d82_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8308258(.data_in(wire_d82_57),.data_out(wire_d82_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8308259(.data_in(wire_d82_58),.data_out(wire_d82_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8308260(.data_in(wire_d82_59),.data_out(wire_d82_60),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8308261(.data_in(wire_d82_60),.data_out(wire_d82_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8308262(.data_in(wire_d82_61),.data_out(wire_d82_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8308263(.data_in(wire_d82_62),.data_out(wire_d82_63),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8308264(.data_in(wire_d82_63),.data_out(wire_d82_64),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8308265(.data_in(wire_d82_64),.data_out(wire_d82_65),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8308266(.data_in(wire_d82_65),.data_out(wire_d82_66),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8308267(.data_in(wire_d82_66),.data_out(wire_d82_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8308268(.data_in(wire_d82_67),.data_out(wire_d82_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8308269(.data_in(wire_d82_68),.data_out(wire_d82_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8308270(.data_in(wire_d82_69),.data_out(wire_d82_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8308271(.data_in(wire_d82_70),.data_out(wire_d82_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8308272(.data_in(wire_d82_71),.data_out(wire_d82_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8308273(.data_in(wire_d82_72),.data_out(wire_d82_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8308274(.data_in(wire_d82_73),.data_out(wire_d82_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8308275(.data_in(wire_d82_74),.data_out(wire_d82_75),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8308276(.data_in(wire_d82_75),.data_out(wire_d82_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8308277(.data_in(wire_d82_76),.data_out(wire_d82_77),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8308278(.data_in(wire_d82_77),.data_out(wire_d82_78),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8308279(.data_in(wire_d82_78),.data_out(wire_d82_79),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8308280(.data_in(wire_d82_79),.data_out(wire_d82_80),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8308281(.data_in(wire_d82_80),.data_out(wire_d82_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8308282(.data_in(wire_d82_81),.data_out(wire_d82_82),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8308283(.data_in(wire_d82_82),.data_out(wire_d82_83),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8308284(.data_in(wire_d82_83),.data_out(wire_d82_84),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8308285(.data_in(wire_d82_84),.data_out(wire_d82_85),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8308286(.data_in(wire_d82_85),.data_out(wire_d82_86),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8308287(.data_in(wire_d82_86),.data_out(wire_d82_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8308288(.data_in(wire_d82_87),.data_out(wire_d82_88),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8308289(.data_in(wire_d82_88),.data_out(wire_d82_89),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8308290(.data_in(wire_d82_89),.data_out(wire_d82_90),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8308291(.data_in(wire_d82_90),.data_out(wire_d82_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8308292(.data_in(wire_d82_91),.data_out(wire_d82_92),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8308293(.data_in(wire_d82_92),.data_out(wire_d82_93),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8308294(.data_in(wire_d82_93),.data_out(wire_d82_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8308295(.data_in(wire_d82_94),.data_out(wire_d82_95),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8308296(.data_in(wire_d82_95),.data_out(wire_d82_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8308297(.data_in(wire_d82_96),.data_out(wire_d82_97),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8308298(.data_in(wire_d82_97),.data_out(wire_d82_98),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8308299(.data_in(wire_d82_98),.data_out(wire_d82_99),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance83082100(.data_in(wire_d82_99),.data_out(wire_d82_100),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance83082101(.data_in(wire_d82_100),.data_out(wire_d82_101),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance83082102(.data_in(wire_d82_101),.data_out(wire_d82_102),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance83082103(.data_in(wire_d82_102),.data_out(wire_d82_103),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance83082104(.data_in(wire_d82_103),.data_out(wire_d82_104),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance83082105(.data_in(wire_d82_104),.data_out(wire_d82_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance83082106(.data_in(wire_d82_105),.data_out(wire_d82_106),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance83082107(.data_in(wire_d82_106),.data_out(wire_d82_107),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance83082108(.data_in(wire_d82_107),.data_out(wire_d82_108),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance83082109(.data_in(wire_d82_108),.data_out(wire_d82_109),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance83082110(.data_in(wire_d82_109),.data_out(wire_d82_110),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance83082111(.data_in(wire_d82_110),.data_out(wire_d82_111),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance83082112(.data_in(wire_d82_111),.data_out(wire_d82_112),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance83082113(.data_in(wire_d82_112),.data_out(wire_d82_113),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance83082114(.data_in(wire_d82_113),.data_out(wire_d82_114),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance83082115(.data_in(wire_d82_114),.data_out(wire_d82_115),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance83082116(.data_in(wire_d82_115),.data_out(wire_d82_116),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance83082117(.data_in(wire_d82_116),.data_out(wire_d82_117),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance83082118(.data_in(wire_d82_117),.data_out(wire_d82_118),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance83082119(.data_in(wire_d82_118),.data_out(d_out82),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance840830(.data_in(d_in83),.data_out(wire_d83_0),.clk(clk),.rst(rst));            //channel 84
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance840831(.data_in(wire_d83_0),.data_out(wire_d83_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance840832(.data_in(wire_d83_1),.data_out(wire_d83_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance840833(.data_in(wire_d83_2),.data_out(wire_d83_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance840834(.data_in(wire_d83_3),.data_out(wire_d83_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance840835(.data_in(wire_d83_4),.data_out(wire_d83_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance840836(.data_in(wire_d83_5),.data_out(wire_d83_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance840837(.data_in(wire_d83_6),.data_out(wire_d83_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance840838(.data_in(wire_d83_7),.data_out(wire_d83_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance840839(.data_in(wire_d83_8),.data_out(wire_d83_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8408310(.data_in(wire_d83_9),.data_out(wire_d83_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8408311(.data_in(wire_d83_10),.data_out(wire_d83_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8408312(.data_in(wire_d83_11),.data_out(wire_d83_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8408313(.data_in(wire_d83_12),.data_out(wire_d83_13),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8408314(.data_in(wire_d83_13),.data_out(wire_d83_14),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8408315(.data_in(wire_d83_14),.data_out(wire_d83_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8408316(.data_in(wire_d83_15),.data_out(wire_d83_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8408317(.data_in(wire_d83_16),.data_out(wire_d83_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8408318(.data_in(wire_d83_17),.data_out(wire_d83_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8408319(.data_in(wire_d83_18),.data_out(wire_d83_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8408320(.data_in(wire_d83_19),.data_out(wire_d83_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8408321(.data_in(wire_d83_20),.data_out(wire_d83_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8408322(.data_in(wire_d83_21),.data_out(wire_d83_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8408323(.data_in(wire_d83_22),.data_out(wire_d83_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8408324(.data_in(wire_d83_23),.data_out(wire_d83_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8408325(.data_in(wire_d83_24),.data_out(wire_d83_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8408326(.data_in(wire_d83_25),.data_out(wire_d83_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8408327(.data_in(wire_d83_26),.data_out(wire_d83_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8408328(.data_in(wire_d83_27),.data_out(wire_d83_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8408329(.data_in(wire_d83_28),.data_out(wire_d83_29),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8408330(.data_in(wire_d83_29),.data_out(wire_d83_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8408331(.data_in(wire_d83_30),.data_out(wire_d83_31),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8408332(.data_in(wire_d83_31),.data_out(wire_d83_32),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8408333(.data_in(wire_d83_32),.data_out(wire_d83_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8408334(.data_in(wire_d83_33),.data_out(wire_d83_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8408335(.data_in(wire_d83_34),.data_out(wire_d83_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8408336(.data_in(wire_d83_35),.data_out(wire_d83_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8408337(.data_in(wire_d83_36),.data_out(wire_d83_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8408338(.data_in(wire_d83_37),.data_out(wire_d83_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8408339(.data_in(wire_d83_38),.data_out(wire_d83_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8408340(.data_in(wire_d83_39),.data_out(wire_d83_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8408341(.data_in(wire_d83_40),.data_out(wire_d83_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8408342(.data_in(wire_d83_41),.data_out(wire_d83_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8408343(.data_in(wire_d83_42),.data_out(wire_d83_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8408344(.data_in(wire_d83_43),.data_out(wire_d83_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8408345(.data_in(wire_d83_44),.data_out(wire_d83_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8408346(.data_in(wire_d83_45),.data_out(wire_d83_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8408347(.data_in(wire_d83_46),.data_out(wire_d83_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8408348(.data_in(wire_d83_47),.data_out(wire_d83_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8408349(.data_in(wire_d83_48),.data_out(wire_d83_49),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8408350(.data_in(wire_d83_49),.data_out(wire_d83_50),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8408351(.data_in(wire_d83_50),.data_out(wire_d83_51),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8408352(.data_in(wire_d83_51),.data_out(wire_d83_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8408353(.data_in(wire_d83_52),.data_out(wire_d83_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8408354(.data_in(wire_d83_53),.data_out(wire_d83_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8408355(.data_in(wire_d83_54),.data_out(wire_d83_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8408356(.data_in(wire_d83_55),.data_out(wire_d83_56),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8408357(.data_in(wire_d83_56),.data_out(wire_d83_57),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8408358(.data_in(wire_d83_57),.data_out(wire_d83_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8408359(.data_in(wire_d83_58),.data_out(wire_d83_59),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8408360(.data_in(wire_d83_59),.data_out(wire_d83_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8408361(.data_in(wire_d83_60),.data_out(wire_d83_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8408362(.data_in(wire_d83_61),.data_out(wire_d83_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8408363(.data_in(wire_d83_62),.data_out(wire_d83_63),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8408364(.data_in(wire_d83_63),.data_out(wire_d83_64),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8408365(.data_in(wire_d83_64),.data_out(wire_d83_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8408366(.data_in(wire_d83_65),.data_out(wire_d83_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8408367(.data_in(wire_d83_66),.data_out(wire_d83_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8408368(.data_in(wire_d83_67),.data_out(wire_d83_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8408369(.data_in(wire_d83_68),.data_out(wire_d83_69),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8408370(.data_in(wire_d83_69),.data_out(wire_d83_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8408371(.data_in(wire_d83_70),.data_out(wire_d83_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8408372(.data_in(wire_d83_71),.data_out(wire_d83_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8408373(.data_in(wire_d83_72),.data_out(wire_d83_73),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8408374(.data_in(wire_d83_73),.data_out(wire_d83_74),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8408375(.data_in(wire_d83_74),.data_out(wire_d83_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8408376(.data_in(wire_d83_75),.data_out(wire_d83_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8408377(.data_in(wire_d83_76),.data_out(wire_d83_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8408378(.data_in(wire_d83_77),.data_out(wire_d83_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8408379(.data_in(wire_d83_78),.data_out(wire_d83_79),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8408380(.data_in(wire_d83_79),.data_out(wire_d83_80),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8408381(.data_in(wire_d83_80),.data_out(wire_d83_81),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8408382(.data_in(wire_d83_81),.data_out(wire_d83_82),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8408383(.data_in(wire_d83_82),.data_out(wire_d83_83),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8408384(.data_in(wire_d83_83),.data_out(wire_d83_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8408385(.data_in(wire_d83_84),.data_out(wire_d83_85),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8408386(.data_in(wire_d83_85),.data_out(wire_d83_86),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8408387(.data_in(wire_d83_86),.data_out(wire_d83_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8408388(.data_in(wire_d83_87),.data_out(wire_d83_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8408389(.data_in(wire_d83_88),.data_out(wire_d83_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8408390(.data_in(wire_d83_89),.data_out(wire_d83_90),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8408391(.data_in(wire_d83_90),.data_out(wire_d83_91),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8408392(.data_in(wire_d83_91),.data_out(wire_d83_92),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8408393(.data_in(wire_d83_92),.data_out(wire_d83_93),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8408394(.data_in(wire_d83_93),.data_out(wire_d83_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8408395(.data_in(wire_d83_94),.data_out(wire_d83_95),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8408396(.data_in(wire_d83_95),.data_out(wire_d83_96),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8408397(.data_in(wire_d83_96),.data_out(wire_d83_97),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8408398(.data_in(wire_d83_97),.data_out(wire_d83_98),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8408399(.data_in(wire_d83_98),.data_out(wire_d83_99),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance84083100(.data_in(wire_d83_99),.data_out(wire_d83_100),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance84083101(.data_in(wire_d83_100),.data_out(wire_d83_101),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance84083102(.data_in(wire_d83_101),.data_out(wire_d83_102),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance84083103(.data_in(wire_d83_102),.data_out(wire_d83_103),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance84083104(.data_in(wire_d83_103),.data_out(wire_d83_104),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance84083105(.data_in(wire_d83_104),.data_out(wire_d83_105),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance84083106(.data_in(wire_d83_105),.data_out(wire_d83_106),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance84083107(.data_in(wire_d83_106),.data_out(wire_d83_107),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance84083108(.data_in(wire_d83_107),.data_out(wire_d83_108),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance84083109(.data_in(wire_d83_108),.data_out(wire_d83_109),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance84083110(.data_in(wire_d83_109),.data_out(wire_d83_110),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance84083111(.data_in(wire_d83_110),.data_out(wire_d83_111),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance84083112(.data_in(wire_d83_111),.data_out(wire_d83_112),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance84083113(.data_in(wire_d83_112),.data_out(wire_d83_113),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance84083114(.data_in(wire_d83_113),.data_out(wire_d83_114),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance84083115(.data_in(wire_d83_114),.data_out(wire_d83_115),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance84083116(.data_in(wire_d83_115),.data_out(wire_d83_116),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance84083117(.data_in(wire_d83_116),.data_out(wire_d83_117),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance84083118(.data_in(wire_d83_117),.data_out(wire_d83_118),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance84083119(.data_in(wire_d83_118),.data_out(d_out83),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance850840(.data_in(d_in84),.data_out(wire_d84_0),.clk(clk),.rst(rst));            //channel 85
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance850841(.data_in(wire_d84_0),.data_out(wire_d84_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance850842(.data_in(wire_d84_1),.data_out(wire_d84_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance850843(.data_in(wire_d84_2),.data_out(wire_d84_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance850844(.data_in(wire_d84_3),.data_out(wire_d84_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance850845(.data_in(wire_d84_4),.data_out(wire_d84_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance850846(.data_in(wire_d84_5),.data_out(wire_d84_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance850847(.data_in(wire_d84_6),.data_out(wire_d84_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance850848(.data_in(wire_d84_7),.data_out(wire_d84_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance850849(.data_in(wire_d84_8),.data_out(wire_d84_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8508410(.data_in(wire_d84_9),.data_out(wire_d84_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8508411(.data_in(wire_d84_10),.data_out(wire_d84_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8508412(.data_in(wire_d84_11),.data_out(wire_d84_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8508413(.data_in(wire_d84_12),.data_out(wire_d84_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8508414(.data_in(wire_d84_13),.data_out(wire_d84_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8508415(.data_in(wire_d84_14),.data_out(wire_d84_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8508416(.data_in(wire_d84_15),.data_out(wire_d84_16),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8508417(.data_in(wire_d84_16),.data_out(wire_d84_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8508418(.data_in(wire_d84_17),.data_out(wire_d84_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8508419(.data_in(wire_d84_18),.data_out(wire_d84_19),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8508420(.data_in(wire_d84_19),.data_out(wire_d84_20),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8508421(.data_in(wire_d84_20),.data_out(wire_d84_21),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8508422(.data_in(wire_d84_21),.data_out(wire_d84_22),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8508423(.data_in(wire_d84_22),.data_out(wire_d84_23),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8508424(.data_in(wire_d84_23),.data_out(wire_d84_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8508425(.data_in(wire_d84_24),.data_out(wire_d84_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8508426(.data_in(wire_d84_25),.data_out(wire_d84_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8508427(.data_in(wire_d84_26),.data_out(wire_d84_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8508428(.data_in(wire_d84_27),.data_out(wire_d84_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8508429(.data_in(wire_d84_28),.data_out(wire_d84_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8508430(.data_in(wire_d84_29),.data_out(wire_d84_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8508431(.data_in(wire_d84_30),.data_out(wire_d84_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8508432(.data_in(wire_d84_31),.data_out(wire_d84_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8508433(.data_in(wire_d84_32),.data_out(wire_d84_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8508434(.data_in(wire_d84_33),.data_out(wire_d84_34),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8508435(.data_in(wire_d84_34),.data_out(wire_d84_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8508436(.data_in(wire_d84_35),.data_out(wire_d84_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8508437(.data_in(wire_d84_36),.data_out(wire_d84_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8508438(.data_in(wire_d84_37),.data_out(wire_d84_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8508439(.data_in(wire_d84_38),.data_out(wire_d84_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8508440(.data_in(wire_d84_39),.data_out(wire_d84_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8508441(.data_in(wire_d84_40),.data_out(wire_d84_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8508442(.data_in(wire_d84_41),.data_out(wire_d84_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8508443(.data_in(wire_d84_42),.data_out(wire_d84_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8508444(.data_in(wire_d84_43),.data_out(wire_d84_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8508445(.data_in(wire_d84_44),.data_out(wire_d84_45),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8508446(.data_in(wire_d84_45),.data_out(wire_d84_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8508447(.data_in(wire_d84_46),.data_out(wire_d84_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8508448(.data_in(wire_d84_47),.data_out(wire_d84_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8508449(.data_in(wire_d84_48),.data_out(wire_d84_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8508450(.data_in(wire_d84_49),.data_out(wire_d84_50),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8508451(.data_in(wire_d84_50),.data_out(wire_d84_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8508452(.data_in(wire_d84_51),.data_out(wire_d84_52),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8508453(.data_in(wire_d84_52),.data_out(wire_d84_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8508454(.data_in(wire_d84_53),.data_out(wire_d84_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8508455(.data_in(wire_d84_54),.data_out(wire_d84_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8508456(.data_in(wire_d84_55),.data_out(wire_d84_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8508457(.data_in(wire_d84_56),.data_out(wire_d84_57),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8508458(.data_in(wire_d84_57),.data_out(wire_d84_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8508459(.data_in(wire_d84_58),.data_out(wire_d84_59),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8508460(.data_in(wire_d84_59),.data_out(wire_d84_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8508461(.data_in(wire_d84_60),.data_out(wire_d84_61),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8508462(.data_in(wire_d84_61),.data_out(wire_d84_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8508463(.data_in(wire_d84_62),.data_out(wire_d84_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8508464(.data_in(wire_d84_63),.data_out(wire_d84_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8508465(.data_in(wire_d84_64),.data_out(wire_d84_65),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8508466(.data_in(wire_d84_65),.data_out(wire_d84_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8508467(.data_in(wire_d84_66),.data_out(wire_d84_67),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8508468(.data_in(wire_d84_67),.data_out(wire_d84_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8508469(.data_in(wire_d84_68),.data_out(wire_d84_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8508470(.data_in(wire_d84_69),.data_out(wire_d84_70),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8508471(.data_in(wire_d84_70),.data_out(wire_d84_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8508472(.data_in(wire_d84_71),.data_out(wire_d84_72),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8508473(.data_in(wire_d84_72),.data_out(wire_d84_73),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8508474(.data_in(wire_d84_73),.data_out(wire_d84_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8508475(.data_in(wire_d84_74),.data_out(wire_d84_75),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8508476(.data_in(wire_d84_75),.data_out(wire_d84_76),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8508477(.data_in(wire_d84_76),.data_out(wire_d84_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8508478(.data_in(wire_d84_77),.data_out(wire_d84_78),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8508479(.data_in(wire_d84_78),.data_out(wire_d84_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8508480(.data_in(wire_d84_79),.data_out(wire_d84_80),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8508481(.data_in(wire_d84_80),.data_out(wire_d84_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8508482(.data_in(wire_d84_81),.data_out(wire_d84_82),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8508483(.data_in(wire_d84_82),.data_out(wire_d84_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8508484(.data_in(wire_d84_83),.data_out(wire_d84_84),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8508485(.data_in(wire_d84_84),.data_out(wire_d84_85),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8508486(.data_in(wire_d84_85),.data_out(wire_d84_86),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8508487(.data_in(wire_d84_86),.data_out(wire_d84_87),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8508488(.data_in(wire_d84_87),.data_out(wire_d84_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8508489(.data_in(wire_d84_88),.data_out(wire_d84_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8508490(.data_in(wire_d84_89),.data_out(wire_d84_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8508491(.data_in(wire_d84_90),.data_out(wire_d84_91),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8508492(.data_in(wire_d84_91),.data_out(wire_d84_92),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8508493(.data_in(wire_d84_92),.data_out(wire_d84_93),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8508494(.data_in(wire_d84_93),.data_out(wire_d84_94),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8508495(.data_in(wire_d84_94),.data_out(wire_d84_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8508496(.data_in(wire_d84_95),.data_out(wire_d84_96),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8508497(.data_in(wire_d84_96),.data_out(wire_d84_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8508498(.data_in(wire_d84_97),.data_out(wire_d84_98),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8508499(.data_in(wire_d84_98),.data_out(wire_d84_99),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance85084100(.data_in(wire_d84_99),.data_out(wire_d84_100),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance85084101(.data_in(wire_d84_100),.data_out(wire_d84_101),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance85084102(.data_in(wire_d84_101),.data_out(wire_d84_102),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance85084103(.data_in(wire_d84_102),.data_out(wire_d84_103),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance85084104(.data_in(wire_d84_103),.data_out(wire_d84_104),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance85084105(.data_in(wire_d84_104),.data_out(wire_d84_105),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance85084106(.data_in(wire_d84_105),.data_out(wire_d84_106),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance85084107(.data_in(wire_d84_106),.data_out(wire_d84_107),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance85084108(.data_in(wire_d84_107),.data_out(wire_d84_108),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance85084109(.data_in(wire_d84_108),.data_out(wire_d84_109),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance85084110(.data_in(wire_d84_109),.data_out(wire_d84_110),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance85084111(.data_in(wire_d84_110),.data_out(wire_d84_111),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance85084112(.data_in(wire_d84_111),.data_out(wire_d84_112),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance85084113(.data_in(wire_d84_112),.data_out(wire_d84_113),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance85084114(.data_in(wire_d84_113),.data_out(wire_d84_114),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance85084115(.data_in(wire_d84_114),.data_out(wire_d84_115),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance85084116(.data_in(wire_d84_115),.data_out(wire_d84_116),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance85084117(.data_in(wire_d84_116),.data_out(wire_d84_117),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance85084118(.data_in(wire_d84_117),.data_out(wire_d84_118),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance85084119(.data_in(wire_d84_118),.data_out(d_out84),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance860850(.data_in(d_in85),.data_out(wire_d85_0),.clk(clk),.rst(rst));            //channel 86
	decoder_top #(.WIDTH(WIDTH)) decoder_instance860851(.data_in(wire_d85_0),.data_out(wire_d85_1),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance860852(.data_in(wire_d85_1),.data_out(wire_d85_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance860853(.data_in(wire_d85_2),.data_out(wire_d85_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance860854(.data_in(wire_d85_3),.data_out(wire_d85_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance860855(.data_in(wire_d85_4),.data_out(wire_d85_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance860856(.data_in(wire_d85_5),.data_out(wire_d85_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance860857(.data_in(wire_d85_6),.data_out(wire_d85_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance860858(.data_in(wire_d85_7),.data_out(wire_d85_8),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance860859(.data_in(wire_d85_8),.data_out(wire_d85_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8608510(.data_in(wire_d85_9),.data_out(wire_d85_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8608511(.data_in(wire_d85_10),.data_out(wire_d85_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8608512(.data_in(wire_d85_11),.data_out(wire_d85_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8608513(.data_in(wire_d85_12),.data_out(wire_d85_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8608514(.data_in(wire_d85_13),.data_out(wire_d85_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8608515(.data_in(wire_d85_14),.data_out(wire_d85_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8608516(.data_in(wire_d85_15),.data_out(wire_d85_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8608517(.data_in(wire_d85_16),.data_out(wire_d85_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8608518(.data_in(wire_d85_17),.data_out(wire_d85_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8608519(.data_in(wire_d85_18),.data_out(wire_d85_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8608520(.data_in(wire_d85_19),.data_out(wire_d85_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8608521(.data_in(wire_d85_20),.data_out(wire_d85_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8608522(.data_in(wire_d85_21),.data_out(wire_d85_22),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8608523(.data_in(wire_d85_22),.data_out(wire_d85_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8608524(.data_in(wire_d85_23),.data_out(wire_d85_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8608525(.data_in(wire_d85_24),.data_out(wire_d85_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8608526(.data_in(wire_d85_25),.data_out(wire_d85_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8608527(.data_in(wire_d85_26),.data_out(wire_d85_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8608528(.data_in(wire_d85_27),.data_out(wire_d85_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8608529(.data_in(wire_d85_28),.data_out(wire_d85_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8608530(.data_in(wire_d85_29),.data_out(wire_d85_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8608531(.data_in(wire_d85_30),.data_out(wire_d85_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8608532(.data_in(wire_d85_31),.data_out(wire_d85_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8608533(.data_in(wire_d85_32),.data_out(wire_d85_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8608534(.data_in(wire_d85_33),.data_out(wire_d85_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8608535(.data_in(wire_d85_34),.data_out(wire_d85_35),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8608536(.data_in(wire_d85_35),.data_out(wire_d85_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8608537(.data_in(wire_d85_36),.data_out(wire_d85_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8608538(.data_in(wire_d85_37),.data_out(wire_d85_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8608539(.data_in(wire_d85_38),.data_out(wire_d85_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8608540(.data_in(wire_d85_39),.data_out(wire_d85_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8608541(.data_in(wire_d85_40),.data_out(wire_d85_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8608542(.data_in(wire_d85_41),.data_out(wire_d85_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8608543(.data_in(wire_d85_42),.data_out(wire_d85_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8608544(.data_in(wire_d85_43),.data_out(wire_d85_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8608545(.data_in(wire_d85_44),.data_out(wire_d85_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8608546(.data_in(wire_d85_45),.data_out(wire_d85_46),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8608547(.data_in(wire_d85_46),.data_out(wire_d85_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8608548(.data_in(wire_d85_47),.data_out(wire_d85_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8608549(.data_in(wire_d85_48),.data_out(wire_d85_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8608550(.data_in(wire_d85_49),.data_out(wire_d85_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8608551(.data_in(wire_d85_50),.data_out(wire_d85_51),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8608552(.data_in(wire_d85_51),.data_out(wire_d85_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8608553(.data_in(wire_d85_52),.data_out(wire_d85_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8608554(.data_in(wire_d85_53),.data_out(wire_d85_54),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8608555(.data_in(wire_d85_54),.data_out(wire_d85_55),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8608556(.data_in(wire_d85_55),.data_out(wire_d85_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8608557(.data_in(wire_d85_56),.data_out(wire_d85_57),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8608558(.data_in(wire_d85_57),.data_out(wire_d85_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8608559(.data_in(wire_d85_58),.data_out(wire_d85_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8608560(.data_in(wire_d85_59),.data_out(wire_d85_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8608561(.data_in(wire_d85_60),.data_out(wire_d85_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8608562(.data_in(wire_d85_61),.data_out(wire_d85_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8608563(.data_in(wire_d85_62),.data_out(wire_d85_63),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8608564(.data_in(wire_d85_63),.data_out(wire_d85_64),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8608565(.data_in(wire_d85_64),.data_out(wire_d85_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8608566(.data_in(wire_d85_65),.data_out(wire_d85_66),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8608567(.data_in(wire_d85_66),.data_out(wire_d85_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8608568(.data_in(wire_d85_67),.data_out(wire_d85_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8608569(.data_in(wire_d85_68),.data_out(wire_d85_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8608570(.data_in(wire_d85_69),.data_out(wire_d85_70),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8608571(.data_in(wire_d85_70),.data_out(wire_d85_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8608572(.data_in(wire_d85_71),.data_out(wire_d85_72),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8608573(.data_in(wire_d85_72),.data_out(wire_d85_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8608574(.data_in(wire_d85_73),.data_out(wire_d85_74),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8608575(.data_in(wire_d85_74),.data_out(wire_d85_75),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8608576(.data_in(wire_d85_75),.data_out(wire_d85_76),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8608577(.data_in(wire_d85_76),.data_out(wire_d85_77),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8608578(.data_in(wire_d85_77),.data_out(wire_d85_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8608579(.data_in(wire_d85_78),.data_out(wire_d85_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8608580(.data_in(wire_d85_79),.data_out(wire_d85_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8608581(.data_in(wire_d85_80),.data_out(wire_d85_81),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8608582(.data_in(wire_d85_81),.data_out(wire_d85_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8608583(.data_in(wire_d85_82),.data_out(wire_d85_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8608584(.data_in(wire_d85_83),.data_out(wire_d85_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8608585(.data_in(wire_d85_84),.data_out(wire_d85_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8608586(.data_in(wire_d85_85),.data_out(wire_d85_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8608587(.data_in(wire_d85_86),.data_out(wire_d85_87),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8608588(.data_in(wire_d85_87),.data_out(wire_d85_88),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8608589(.data_in(wire_d85_88),.data_out(wire_d85_89),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8608590(.data_in(wire_d85_89),.data_out(wire_d85_90),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8608591(.data_in(wire_d85_90),.data_out(wire_d85_91),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8608592(.data_in(wire_d85_91),.data_out(wire_d85_92),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8608593(.data_in(wire_d85_92),.data_out(wire_d85_93),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8608594(.data_in(wire_d85_93),.data_out(wire_d85_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8608595(.data_in(wire_d85_94),.data_out(wire_d85_95),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8608596(.data_in(wire_d85_95),.data_out(wire_d85_96),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8608597(.data_in(wire_d85_96),.data_out(wire_d85_97),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8608598(.data_in(wire_d85_97),.data_out(wire_d85_98),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8608599(.data_in(wire_d85_98),.data_out(wire_d85_99),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance86085100(.data_in(wire_d85_99),.data_out(wire_d85_100),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance86085101(.data_in(wire_d85_100),.data_out(wire_d85_101),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance86085102(.data_in(wire_d85_101),.data_out(wire_d85_102),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance86085103(.data_in(wire_d85_102),.data_out(wire_d85_103),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance86085104(.data_in(wire_d85_103),.data_out(wire_d85_104),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance86085105(.data_in(wire_d85_104),.data_out(wire_d85_105),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance86085106(.data_in(wire_d85_105),.data_out(wire_d85_106),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance86085107(.data_in(wire_d85_106),.data_out(wire_d85_107),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance86085108(.data_in(wire_d85_107),.data_out(wire_d85_108),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance86085109(.data_in(wire_d85_108),.data_out(wire_d85_109),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance86085110(.data_in(wire_d85_109),.data_out(wire_d85_110),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance86085111(.data_in(wire_d85_110),.data_out(wire_d85_111),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance86085112(.data_in(wire_d85_111),.data_out(wire_d85_112),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance86085113(.data_in(wire_d85_112),.data_out(wire_d85_113),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance86085114(.data_in(wire_d85_113),.data_out(wire_d85_114),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance86085115(.data_in(wire_d85_114),.data_out(wire_d85_115),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance86085116(.data_in(wire_d85_115),.data_out(wire_d85_116),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance86085117(.data_in(wire_d85_116),.data_out(wire_d85_117),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance86085118(.data_in(wire_d85_117),.data_out(wire_d85_118),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance86085119(.data_in(wire_d85_118),.data_out(d_out85),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance870860(.data_in(d_in86),.data_out(wire_d86_0),.clk(clk),.rst(rst));            //channel 87
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance870861(.data_in(wire_d86_0),.data_out(wire_d86_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance870862(.data_in(wire_d86_1),.data_out(wire_d86_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance870863(.data_in(wire_d86_2),.data_out(wire_d86_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance870864(.data_in(wire_d86_3),.data_out(wire_d86_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance870865(.data_in(wire_d86_4),.data_out(wire_d86_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance870866(.data_in(wire_d86_5),.data_out(wire_d86_6),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance870867(.data_in(wire_d86_6),.data_out(wire_d86_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance870868(.data_in(wire_d86_7),.data_out(wire_d86_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance870869(.data_in(wire_d86_8),.data_out(wire_d86_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8708610(.data_in(wire_d86_9),.data_out(wire_d86_10),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8708611(.data_in(wire_d86_10),.data_out(wire_d86_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8708612(.data_in(wire_d86_11),.data_out(wire_d86_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8708613(.data_in(wire_d86_12),.data_out(wire_d86_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8708614(.data_in(wire_d86_13),.data_out(wire_d86_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8708615(.data_in(wire_d86_14),.data_out(wire_d86_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8708616(.data_in(wire_d86_15),.data_out(wire_d86_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8708617(.data_in(wire_d86_16),.data_out(wire_d86_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8708618(.data_in(wire_d86_17),.data_out(wire_d86_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8708619(.data_in(wire_d86_18),.data_out(wire_d86_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8708620(.data_in(wire_d86_19),.data_out(wire_d86_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8708621(.data_in(wire_d86_20),.data_out(wire_d86_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8708622(.data_in(wire_d86_21),.data_out(wire_d86_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8708623(.data_in(wire_d86_22),.data_out(wire_d86_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8708624(.data_in(wire_d86_23),.data_out(wire_d86_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8708625(.data_in(wire_d86_24),.data_out(wire_d86_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8708626(.data_in(wire_d86_25),.data_out(wire_d86_26),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8708627(.data_in(wire_d86_26),.data_out(wire_d86_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8708628(.data_in(wire_d86_27),.data_out(wire_d86_28),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8708629(.data_in(wire_d86_28),.data_out(wire_d86_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8708630(.data_in(wire_d86_29),.data_out(wire_d86_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8708631(.data_in(wire_d86_30),.data_out(wire_d86_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8708632(.data_in(wire_d86_31),.data_out(wire_d86_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8708633(.data_in(wire_d86_32),.data_out(wire_d86_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8708634(.data_in(wire_d86_33),.data_out(wire_d86_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8708635(.data_in(wire_d86_34),.data_out(wire_d86_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8708636(.data_in(wire_d86_35),.data_out(wire_d86_36),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8708637(.data_in(wire_d86_36),.data_out(wire_d86_37),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8708638(.data_in(wire_d86_37),.data_out(wire_d86_38),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8708639(.data_in(wire_d86_38),.data_out(wire_d86_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8708640(.data_in(wire_d86_39),.data_out(wire_d86_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8708641(.data_in(wire_d86_40),.data_out(wire_d86_41),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8708642(.data_in(wire_d86_41),.data_out(wire_d86_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8708643(.data_in(wire_d86_42),.data_out(wire_d86_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8708644(.data_in(wire_d86_43),.data_out(wire_d86_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8708645(.data_in(wire_d86_44),.data_out(wire_d86_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8708646(.data_in(wire_d86_45),.data_out(wire_d86_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8708647(.data_in(wire_d86_46),.data_out(wire_d86_47),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8708648(.data_in(wire_d86_47),.data_out(wire_d86_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8708649(.data_in(wire_d86_48),.data_out(wire_d86_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8708650(.data_in(wire_d86_49),.data_out(wire_d86_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8708651(.data_in(wire_d86_50),.data_out(wire_d86_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8708652(.data_in(wire_d86_51),.data_out(wire_d86_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8708653(.data_in(wire_d86_52),.data_out(wire_d86_53),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8708654(.data_in(wire_d86_53),.data_out(wire_d86_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8708655(.data_in(wire_d86_54),.data_out(wire_d86_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8708656(.data_in(wire_d86_55),.data_out(wire_d86_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8708657(.data_in(wire_d86_56),.data_out(wire_d86_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8708658(.data_in(wire_d86_57),.data_out(wire_d86_58),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8708659(.data_in(wire_d86_58),.data_out(wire_d86_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8708660(.data_in(wire_d86_59),.data_out(wire_d86_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8708661(.data_in(wire_d86_60),.data_out(wire_d86_61),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8708662(.data_in(wire_d86_61),.data_out(wire_d86_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8708663(.data_in(wire_d86_62),.data_out(wire_d86_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8708664(.data_in(wire_d86_63),.data_out(wire_d86_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8708665(.data_in(wire_d86_64),.data_out(wire_d86_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8708666(.data_in(wire_d86_65),.data_out(wire_d86_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8708667(.data_in(wire_d86_66),.data_out(wire_d86_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8708668(.data_in(wire_d86_67),.data_out(wire_d86_68),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8708669(.data_in(wire_d86_68),.data_out(wire_d86_69),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8708670(.data_in(wire_d86_69),.data_out(wire_d86_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8708671(.data_in(wire_d86_70),.data_out(wire_d86_71),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8708672(.data_in(wire_d86_71),.data_out(wire_d86_72),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8708673(.data_in(wire_d86_72),.data_out(wire_d86_73),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8708674(.data_in(wire_d86_73),.data_out(wire_d86_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8708675(.data_in(wire_d86_74),.data_out(wire_d86_75),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8708676(.data_in(wire_d86_75),.data_out(wire_d86_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8708677(.data_in(wire_d86_76),.data_out(wire_d86_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8708678(.data_in(wire_d86_77),.data_out(wire_d86_78),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8708679(.data_in(wire_d86_78),.data_out(wire_d86_79),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8708680(.data_in(wire_d86_79),.data_out(wire_d86_80),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8708681(.data_in(wire_d86_80),.data_out(wire_d86_81),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8708682(.data_in(wire_d86_81),.data_out(wire_d86_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8708683(.data_in(wire_d86_82),.data_out(wire_d86_83),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8708684(.data_in(wire_d86_83),.data_out(wire_d86_84),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8708685(.data_in(wire_d86_84),.data_out(wire_d86_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8708686(.data_in(wire_d86_85),.data_out(wire_d86_86),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8708687(.data_in(wire_d86_86),.data_out(wire_d86_87),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8708688(.data_in(wire_d86_87),.data_out(wire_d86_88),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8708689(.data_in(wire_d86_88),.data_out(wire_d86_89),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8708690(.data_in(wire_d86_89),.data_out(wire_d86_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8708691(.data_in(wire_d86_90),.data_out(wire_d86_91),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8708692(.data_in(wire_d86_91),.data_out(wire_d86_92),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8708693(.data_in(wire_d86_92),.data_out(wire_d86_93),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8708694(.data_in(wire_d86_93),.data_out(wire_d86_94),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8708695(.data_in(wire_d86_94),.data_out(wire_d86_95),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8708696(.data_in(wire_d86_95),.data_out(wire_d86_96),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8708697(.data_in(wire_d86_96),.data_out(wire_d86_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8708698(.data_in(wire_d86_97),.data_out(wire_d86_98),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8708699(.data_in(wire_d86_98),.data_out(wire_d86_99),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance87086100(.data_in(wire_d86_99),.data_out(wire_d86_100),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance87086101(.data_in(wire_d86_100),.data_out(wire_d86_101),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance87086102(.data_in(wire_d86_101),.data_out(wire_d86_102),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance87086103(.data_in(wire_d86_102),.data_out(wire_d86_103),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance87086104(.data_in(wire_d86_103),.data_out(wire_d86_104),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance87086105(.data_in(wire_d86_104),.data_out(wire_d86_105),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance87086106(.data_in(wire_d86_105),.data_out(wire_d86_106),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance87086107(.data_in(wire_d86_106),.data_out(wire_d86_107),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance87086108(.data_in(wire_d86_107),.data_out(wire_d86_108),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance87086109(.data_in(wire_d86_108),.data_out(wire_d86_109),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance87086110(.data_in(wire_d86_109),.data_out(wire_d86_110),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance87086111(.data_in(wire_d86_110),.data_out(wire_d86_111),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance87086112(.data_in(wire_d86_111),.data_out(wire_d86_112),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance87086113(.data_in(wire_d86_112),.data_out(wire_d86_113),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance87086114(.data_in(wire_d86_113),.data_out(wire_d86_114),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance87086115(.data_in(wire_d86_114),.data_out(wire_d86_115),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance87086116(.data_in(wire_d86_115),.data_out(wire_d86_116),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance87086117(.data_in(wire_d86_116),.data_out(wire_d86_117),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance87086118(.data_in(wire_d86_117),.data_out(wire_d86_118),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance87086119(.data_in(wire_d86_118),.data_out(d_out86),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance880870(.data_in(d_in87),.data_out(wire_d87_0),.clk(clk),.rst(rst));            //channel 88
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance880871(.data_in(wire_d87_0),.data_out(wire_d87_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance880872(.data_in(wire_d87_1),.data_out(wire_d87_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance880873(.data_in(wire_d87_2),.data_out(wire_d87_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance880874(.data_in(wire_d87_3),.data_out(wire_d87_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance880875(.data_in(wire_d87_4),.data_out(wire_d87_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance880876(.data_in(wire_d87_5),.data_out(wire_d87_6),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance880877(.data_in(wire_d87_6),.data_out(wire_d87_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance880878(.data_in(wire_d87_7),.data_out(wire_d87_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance880879(.data_in(wire_d87_8),.data_out(wire_d87_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8808710(.data_in(wire_d87_9),.data_out(wire_d87_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8808711(.data_in(wire_d87_10),.data_out(wire_d87_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8808712(.data_in(wire_d87_11),.data_out(wire_d87_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8808713(.data_in(wire_d87_12),.data_out(wire_d87_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8808714(.data_in(wire_d87_13),.data_out(wire_d87_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8808715(.data_in(wire_d87_14),.data_out(wire_d87_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8808716(.data_in(wire_d87_15),.data_out(wire_d87_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8808717(.data_in(wire_d87_16),.data_out(wire_d87_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8808718(.data_in(wire_d87_17),.data_out(wire_d87_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8808719(.data_in(wire_d87_18),.data_out(wire_d87_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8808720(.data_in(wire_d87_19),.data_out(wire_d87_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8808721(.data_in(wire_d87_20),.data_out(wire_d87_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8808722(.data_in(wire_d87_21),.data_out(wire_d87_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8808723(.data_in(wire_d87_22),.data_out(wire_d87_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8808724(.data_in(wire_d87_23),.data_out(wire_d87_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8808725(.data_in(wire_d87_24),.data_out(wire_d87_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8808726(.data_in(wire_d87_25),.data_out(wire_d87_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8808727(.data_in(wire_d87_26),.data_out(wire_d87_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8808728(.data_in(wire_d87_27),.data_out(wire_d87_28),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8808729(.data_in(wire_d87_28),.data_out(wire_d87_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8808730(.data_in(wire_d87_29),.data_out(wire_d87_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8808731(.data_in(wire_d87_30),.data_out(wire_d87_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8808732(.data_in(wire_d87_31),.data_out(wire_d87_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8808733(.data_in(wire_d87_32),.data_out(wire_d87_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8808734(.data_in(wire_d87_33),.data_out(wire_d87_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8808735(.data_in(wire_d87_34),.data_out(wire_d87_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8808736(.data_in(wire_d87_35),.data_out(wire_d87_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8808737(.data_in(wire_d87_36),.data_out(wire_d87_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8808738(.data_in(wire_d87_37),.data_out(wire_d87_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8808739(.data_in(wire_d87_38),.data_out(wire_d87_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8808740(.data_in(wire_d87_39),.data_out(wire_d87_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8808741(.data_in(wire_d87_40),.data_out(wire_d87_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8808742(.data_in(wire_d87_41),.data_out(wire_d87_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8808743(.data_in(wire_d87_42),.data_out(wire_d87_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8808744(.data_in(wire_d87_43),.data_out(wire_d87_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8808745(.data_in(wire_d87_44),.data_out(wire_d87_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8808746(.data_in(wire_d87_45),.data_out(wire_d87_46),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8808747(.data_in(wire_d87_46),.data_out(wire_d87_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8808748(.data_in(wire_d87_47),.data_out(wire_d87_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8808749(.data_in(wire_d87_48),.data_out(wire_d87_49),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8808750(.data_in(wire_d87_49),.data_out(wire_d87_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8808751(.data_in(wire_d87_50),.data_out(wire_d87_51),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8808752(.data_in(wire_d87_51),.data_out(wire_d87_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8808753(.data_in(wire_d87_52),.data_out(wire_d87_53),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8808754(.data_in(wire_d87_53),.data_out(wire_d87_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8808755(.data_in(wire_d87_54),.data_out(wire_d87_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8808756(.data_in(wire_d87_55),.data_out(wire_d87_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8808757(.data_in(wire_d87_56),.data_out(wire_d87_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8808758(.data_in(wire_d87_57),.data_out(wire_d87_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8808759(.data_in(wire_d87_58),.data_out(wire_d87_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8808760(.data_in(wire_d87_59),.data_out(wire_d87_60),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8808761(.data_in(wire_d87_60),.data_out(wire_d87_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8808762(.data_in(wire_d87_61),.data_out(wire_d87_62),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8808763(.data_in(wire_d87_62),.data_out(wire_d87_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8808764(.data_in(wire_d87_63),.data_out(wire_d87_64),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8808765(.data_in(wire_d87_64),.data_out(wire_d87_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8808766(.data_in(wire_d87_65),.data_out(wire_d87_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8808767(.data_in(wire_d87_66),.data_out(wire_d87_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8808768(.data_in(wire_d87_67),.data_out(wire_d87_68),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8808769(.data_in(wire_d87_68),.data_out(wire_d87_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8808770(.data_in(wire_d87_69),.data_out(wire_d87_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8808771(.data_in(wire_d87_70),.data_out(wire_d87_71),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8808772(.data_in(wire_d87_71),.data_out(wire_d87_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8808773(.data_in(wire_d87_72),.data_out(wire_d87_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8808774(.data_in(wire_d87_73),.data_out(wire_d87_74),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8808775(.data_in(wire_d87_74),.data_out(wire_d87_75),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8808776(.data_in(wire_d87_75),.data_out(wire_d87_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8808777(.data_in(wire_d87_76),.data_out(wire_d87_77),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8808778(.data_in(wire_d87_77),.data_out(wire_d87_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8808779(.data_in(wire_d87_78),.data_out(wire_d87_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8808780(.data_in(wire_d87_79),.data_out(wire_d87_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8808781(.data_in(wire_d87_80),.data_out(wire_d87_81),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8808782(.data_in(wire_d87_81),.data_out(wire_d87_82),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8808783(.data_in(wire_d87_82),.data_out(wire_d87_83),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8808784(.data_in(wire_d87_83),.data_out(wire_d87_84),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8808785(.data_in(wire_d87_84),.data_out(wire_d87_85),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8808786(.data_in(wire_d87_85),.data_out(wire_d87_86),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8808787(.data_in(wire_d87_86),.data_out(wire_d87_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8808788(.data_in(wire_d87_87),.data_out(wire_d87_88),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8808789(.data_in(wire_d87_88),.data_out(wire_d87_89),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8808790(.data_in(wire_d87_89),.data_out(wire_d87_90),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8808791(.data_in(wire_d87_90),.data_out(wire_d87_91),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8808792(.data_in(wire_d87_91),.data_out(wire_d87_92),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8808793(.data_in(wire_d87_92),.data_out(wire_d87_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8808794(.data_in(wire_d87_93),.data_out(wire_d87_94),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8808795(.data_in(wire_d87_94),.data_out(wire_d87_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8808796(.data_in(wire_d87_95),.data_out(wire_d87_96),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8808797(.data_in(wire_d87_96),.data_out(wire_d87_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8808798(.data_in(wire_d87_97),.data_out(wire_d87_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8808799(.data_in(wire_d87_98),.data_out(wire_d87_99),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance88087100(.data_in(wire_d87_99),.data_out(wire_d87_100),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance88087101(.data_in(wire_d87_100),.data_out(wire_d87_101),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance88087102(.data_in(wire_d87_101),.data_out(wire_d87_102),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance88087103(.data_in(wire_d87_102),.data_out(wire_d87_103),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance88087104(.data_in(wire_d87_103),.data_out(wire_d87_104),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance88087105(.data_in(wire_d87_104),.data_out(wire_d87_105),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance88087106(.data_in(wire_d87_105),.data_out(wire_d87_106),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance88087107(.data_in(wire_d87_106),.data_out(wire_d87_107),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance88087108(.data_in(wire_d87_107),.data_out(wire_d87_108),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance88087109(.data_in(wire_d87_108),.data_out(wire_d87_109),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance88087110(.data_in(wire_d87_109),.data_out(wire_d87_110),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance88087111(.data_in(wire_d87_110),.data_out(wire_d87_111),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance88087112(.data_in(wire_d87_111),.data_out(wire_d87_112),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance88087113(.data_in(wire_d87_112),.data_out(wire_d87_113),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance88087114(.data_in(wire_d87_113),.data_out(wire_d87_114),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance88087115(.data_in(wire_d87_114),.data_out(wire_d87_115),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance88087116(.data_in(wire_d87_115),.data_out(wire_d87_116),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance88087117(.data_in(wire_d87_116),.data_out(wire_d87_117),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance88087118(.data_in(wire_d87_117),.data_out(wire_d87_118),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance88087119(.data_in(wire_d87_118),.data_out(d_out87),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance890880(.data_in(d_in88),.data_out(wire_d88_0),.clk(clk),.rst(rst));            //channel 89
	decoder_top #(.WIDTH(WIDTH)) decoder_instance890881(.data_in(wire_d88_0),.data_out(wire_d88_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance890882(.data_in(wire_d88_1),.data_out(wire_d88_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance890883(.data_in(wire_d88_2),.data_out(wire_d88_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance890884(.data_in(wire_d88_3),.data_out(wire_d88_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance890885(.data_in(wire_d88_4),.data_out(wire_d88_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance890886(.data_in(wire_d88_5),.data_out(wire_d88_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance890887(.data_in(wire_d88_6),.data_out(wire_d88_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance890888(.data_in(wire_d88_7),.data_out(wire_d88_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance890889(.data_in(wire_d88_8),.data_out(wire_d88_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8908810(.data_in(wire_d88_9),.data_out(wire_d88_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8908811(.data_in(wire_d88_10),.data_out(wire_d88_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8908812(.data_in(wire_d88_11),.data_out(wire_d88_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8908813(.data_in(wire_d88_12),.data_out(wire_d88_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8908814(.data_in(wire_d88_13),.data_out(wire_d88_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8908815(.data_in(wire_d88_14),.data_out(wire_d88_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8908816(.data_in(wire_d88_15),.data_out(wire_d88_16),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8908817(.data_in(wire_d88_16),.data_out(wire_d88_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8908818(.data_in(wire_d88_17),.data_out(wire_d88_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8908819(.data_in(wire_d88_18),.data_out(wire_d88_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8908820(.data_in(wire_d88_19),.data_out(wire_d88_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8908821(.data_in(wire_d88_20),.data_out(wire_d88_21),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8908822(.data_in(wire_d88_21),.data_out(wire_d88_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8908823(.data_in(wire_d88_22),.data_out(wire_d88_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8908824(.data_in(wire_d88_23),.data_out(wire_d88_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8908825(.data_in(wire_d88_24),.data_out(wire_d88_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8908826(.data_in(wire_d88_25),.data_out(wire_d88_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8908827(.data_in(wire_d88_26),.data_out(wire_d88_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8908828(.data_in(wire_d88_27),.data_out(wire_d88_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8908829(.data_in(wire_d88_28),.data_out(wire_d88_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8908830(.data_in(wire_d88_29),.data_out(wire_d88_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8908831(.data_in(wire_d88_30),.data_out(wire_d88_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8908832(.data_in(wire_d88_31),.data_out(wire_d88_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8908833(.data_in(wire_d88_32),.data_out(wire_d88_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8908834(.data_in(wire_d88_33),.data_out(wire_d88_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8908835(.data_in(wire_d88_34),.data_out(wire_d88_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8908836(.data_in(wire_d88_35),.data_out(wire_d88_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8908837(.data_in(wire_d88_36),.data_out(wire_d88_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8908838(.data_in(wire_d88_37),.data_out(wire_d88_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8908839(.data_in(wire_d88_38),.data_out(wire_d88_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8908840(.data_in(wire_d88_39),.data_out(wire_d88_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8908841(.data_in(wire_d88_40),.data_out(wire_d88_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8908842(.data_in(wire_d88_41),.data_out(wire_d88_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8908843(.data_in(wire_d88_42),.data_out(wire_d88_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8908844(.data_in(wire_d88_43),.data_out(wire_d88_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8908845(.data_in(wire_d88_44),.data_out(wire_d88_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8908846(.data_in(wire_d88_45),.data_out(wire_d88_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8908847(.data_in(wire_d88_46),.data_out(wire_d88_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8908848(.data_in(wire_d88_47),.data_out(wire_d88_48),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8908849(.data_in(wire_d88_48),.data_out(wire_d88_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8908850(.data_in(wire_d88_49),.data_out(wire_d88_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8908851(.data_in(wire_d88_50),.data_out(wire_d88_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8908852(.data_in(wire_d88_51),.data_out(wire_d88_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8908853(.data_in(wire_d88_52),.data_out(wire_d88_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8908854(.data_in(wire_d88_53),.data_out(wire_d88_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8908855(.data_in(wire_d88_54),.data_out(wire_d88_55),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8908856(.data_in(wire_d88_55),.data_out(wire_d88_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8908857(.data_in(wire_d88_56),.data_out(wire_d88_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8908858(.data_in(wire_d88_57),.data_out(wire_d88_58),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8908859(.data_in(wire_d88_58),.data_out(wire_d88_59),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8908860(.data_in(wire_d88_59),.data_out(wire_d88_60),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8908861(.data_in(wire_d88_60),.data_out(wire_d88_61),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8908862(.data_in(wire_d88_61),.data_out(wire_d88_62),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8908863(.data_in(wire_d88_62),.data_out(wire_d88_63),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8908864(.data_in(wire_d88_63),.data_out(wire_d88_64),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8908865(.data_in(wire_d88_64),.data_out(wire_d88_65),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8908866(.data_in(wire_d88_65),.data_out(wire_d88_66),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8908867(.data_in(wire_d88_66),.data_out(wire_d88_67),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8908868(.data_in(wire_d88_67),.data_out(wire_d88_68),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8908869(.data_in(wire_d88_68),.data_out(wire_d88_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8908870(.data_in(wire_d88_69),.data_out(wire_d88_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8908871(.data_in(wire_d88_70),.data_out(wire_d88_71),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8908872(.data_in(wire_d88_71),.data_out(wire_d88_72),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8908873(.data_in(wire_d88_72),.data_out(wire_d88_73),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8908874(.data_in(wire_d88_73),.data_out(wire_d88_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8908875(.data_in(wire_d88_74),.data_out(wire_d88_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8908876(.data_in(wire_d88_75),.data_out(wire_d88_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8908877(.data_in(wire_d88_76),.data_out(wire_d88_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8908878(.data_in(wire_d88_77),.data_out(wire_d88_78),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8908879(.data_in(wire_d88_78),.data_out(wire_d88_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8908880(.data_in(wire_d88_79),.data_out(wire_d88_80),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8908881(.data_in(wire_d88_80),.data_out(wire_d88_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8908882(.data_in(wire_d88_81),.data_out(wire_d88_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8908883(.data_in(wire_d88_82),.data_out(wire_d88_83),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8908884(.data_in(wire_d88_83),.data_out(wire_d88_84),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8908885(.data_in(wire_d88_84),.data_out(wire_d88_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8908886(.data_in(wire_d88_85),.data_out(wire_d88_86),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8908887(.data_in(wire_d88_86),.data_out(wire_d88_87),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8908888(.data_in(wire_d88_87),.data_out(wire_d88_88),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8908889(.data_in(wire_d88_88),.data_out(wire_d88_89),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8908890(.data_in(wire_d88_89),.data_out(wire_d88_90),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8908891(.data_in(wire_d88_90),.data_out(wire_d88_91),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8908892(.data_in(wire_d88_91),.data_out(wire_d88_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8908893(.data_in(wire_d88_92),.data_out(wire_d88_93),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8908894(.data_in(wire_d88_93),.data_out(wire_d88_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8908895(.data_in(wire_d88_94),.data_out(wire_d88_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8908896(.data_in(wire_d88_95),.data_out(wire_d88_96),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8908897(.data_in(wire_d88_96),.data_out(wire_d88_97),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8908898(.data_in(wire_d88_97),.data_out(wire_d88_98),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8908899(.data_in(wire_d88_98),.data_out(wire_d88_99),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance89088100(.data_in(wire_d88_99),.data_out(wire_d88_100),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance89088101(.data_in(wire_d88_100),.data_out(wire_d88_101),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance89088102(.data_in(wire_d88_101),.data_out(wire_d88_102),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance89088103(.data_in(wire_d88_102),.data_out(wire_d88_103),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance89088104(.data_in(wire_d88_103),.data_out(wire_d88_104),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance89088105(.data_in(wire_d88_104),.data_out(wire_d88_105),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance89088106(.data_in(wire_d88_105),.data_out(wire_d88_106),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance89088107(.data_in(wire_d88_106),.data_out(wire_d88_107),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance89088108(.data_in(wire_d88_107),.data_out(wire_d88_108),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance89088109(.data_in(wire_d88_108),.data_out(wire_d88_109),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance89088110(.data_in(wire_d88_109),.data_out(wire_d88_110),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance89088111(.data_in(wire_d88_110),.data_out(wire_d88_111),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance89088112(.data_in(wire_d88_111),.data_out(wire_d88_112),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance89088113(.data_in(wire_d88_112),.data_out(wire_d88_113),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance89088114(.data_in(wire_d88_113),.data_out(wire_d88_114),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance89088115(.data_in(wire_d88_114),.data_out(wire_d88_115),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance89088116(.data_in(wire_d88_115),.data_out(wire_d88_116),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance89088117(.data_in(wire_d88_116),.data_out(wire_d88_117),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance89088118(.data_in(wire_d88_117),.data_out(wire_d88_118),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance89088119(.data_in(wire_d88_118),.data_out(d_out88),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance900890(.data_in(d_in89),.data_out(wire_d89_0),.clk(clk),.rst(rst));            //channel 90
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance900891(.data_in(wire_d89_0),.data_out(wire_d89_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance900892(.data_in(wire_d89_1),.data_out(wire_d89_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance900893(.data_in(wire_d89_2),.data_out(wire_d89_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance900894(.data_in(wire_d89_3),.data_out(wire_d89_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance900895(.data_in(wire_d89_4),.data_out(wire_d89_5),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance900896(.data_in(wire_d89_5),.data_out(wire_d89_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance900897(.data_in(wire_d89_6),.data_out(wire_d89_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance900898(.data_in(wire_d89_7),.data_out(wire_d89_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance900899(.data_in(wire_d89_8),.data_out(wire_d89_9),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9008910(.data_in(wire_d89_9),.data_out(wire_d89_10),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9008911(.data_in(wire_d89_10),.data_out(wire_d89_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9008912(.data_in(wire_d89_11),.data_out(wire_d89_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9008913(.data_in(wire_d89_12),.data_out(wire_d89_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9008914(.data_in(wire_d89_13),.data_out(wire_d89_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9008915(.data_in(wire_d89_14),.data_out(wire_d89_15),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9008916(.data_in(wire_d89_15),.data_out(wire_d89_16),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9008917(.data_in(wire_d89_16),.data_out(wire_d89_17),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9008918(.data_in(wire_d89_17),.data_out(wire_d89_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9008919(.data_in(wire_d89_18),.data_out(wire_d89_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9008920(.data_in(wire_d89_19),.data_out(wire_d89_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9008921(.data_in(wire_d89_20),.data_out(wire_d89_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9008922(.data_in(wire_d89_21),.data_out(wire_d89_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9008923(.data_in(wire_d89_22),.data_out(wire_d89_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9008924(.data_in(wire_d89_23),.data_out(wire_d89_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9008925(.data_in(wire_d89_24),.data_out(wire_d89_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9008926(.data_in(wire_d89_25),.data_out(wire_d89_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9008927(.data_in(wire_d89_26),.data_out(wire_d89_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9008928(.data_in(wire_d89_27),.data_out(wire_d89_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9008929(.data_in(wire_d89_28),.data_out(wire_d89_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9008930(.data_in(wire_d89_29),.data_out(wire_d89_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9008931(.data_in(wire_d89_30),.data_out(wire_d89_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9008932(.data_in(wire_d89_31),.data_out(wire_d89_32),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9008933(.data_in(wire_d89_32),.data_out(wire_d89_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9008934(.data_in(wire_d89_33),.data_out(wire_d89_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9008935(.data_in(wire_d89_34),.data_out(wire_d89_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9008936(.data_in(wire_d89_35),.data_out(wire_d89_36),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9008937(.data_in(wire_d89_36),.data_out(wire_d89_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9008938(.data_in(wire_d89_37),.data_out(wire_d89_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9008939(.data_in(wire_d89_38),.data_out(wire_d89_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9008940(.data_in(wire_d89_39),.data_out(wire_d89_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9008941(.data_in(wire_d89_40),.data_out(wire_d89_41),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9008942(.data_in(wire_d89_41),.data_out(wire_d89_42),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9008943(.data_in(wire_d89_42),.data_out(wire_d89_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9008944(.data_in(wire_d89_43),.data_out(wire_d89_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9008945(.data_in(wire_d89_44),.data_out(wire_d89_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9008946(.data_in(wire_d89_45),.data_out(wire_d89_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9008947(.data_in(wire_d89_46),.data_out(wire_d89_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9008948(.data_in(wire_d89_47),.data_out(wire_d89_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9008949(.data_in(wire_d89_48),.data_out(wire_d89_49),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9008950(.data_in(wire_d89_49),.data_out(wire_d89_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9008951(.data_in(wire_d89_50),.data_out(wire_d89_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9008952(.data_in(wire_d89_51),.data_out(wire_d89_52),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9008953(.data_in(wire_d89_52),.data_out(wire_d89_53),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9008954(.data_in(wire_d89_53),.data_out(wire_d89_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9008955(.data_in(wire_d89_54),.data_out(wire_d89_55),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9008956(.data_in(wire_d89_55),.data_out(wire_d89_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9008957(.data_in(wire_d89_56),.data_out(wire_d89_57),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9008958(.data_in(wire_d89_57),.data_out(wire_d89_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9008959(.data_in(wire_d89_58),.data_out(wire_d89_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9008960(.data_in(wire_d89_59),.data_out(wire_d89_60),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9008961(.data_in(wire_d89_60),.data_out(wire_d89_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9008962(.data_in(wire_d89_61),.data_out(wire_d89_62),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9008963(.data_in(wire_d89_62),.data_out(wire_d89_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9008964(.data_in(wire_d89_63),.data_out(wire_d89_64),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9008965(.data_in(wire_d89_64),.data_out(wire_d89_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9008966(.data_in(wire_d89_65),.data_out(wire_d89_66),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9008967(.data_in(wire_d89_66),.data_out(wire_d89_67),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9008968(.data_in(wire_d89_67),.data_out(wire_d89_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9008969(.data_in(wire_d89_68),.data_out(wire_d89_69),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9008970(.data_in(wire_d89_69),.data_out(wire_d89_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9008971(.data_in(wire_d89_70),.data_out(wire_d89_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9008972(.data_in(wire_d89_71),.data_out(wire_d89_72),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9008973(.data_in(wire_d89_72),.data_out(wire_d89_73),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9008974(.data_in(wire_d89_73),.data_out(wire_d89_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9008975(.data_in(wire_d89_74),.data_out(wire_d89_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9008976(.data_in(wire_d89_75),.data_out(wire_d89_76),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9008977(.data_in(wire_d89_76),.data_out(wire_d89_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9008978(.data_in(wire_d89_77),.data_out(wire_d89_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9008979(.data_in(wire_d89_78),.data_out(wire_d89_79),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9008980(.data_in(wire_d89_79),.data_out(wire_d89_80),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9008981(.data_in(wire_d89_80),.data_out(wire_d89_81),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9008982(.data_in(wire_d89_81),.data_out(wire_d89_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9008983(.data_in(wire_d89_82),.data_out(wire_d89_83),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9008984(.data_in(wire_d89_83),.data_out(wire_d89_84),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9008985(.data_in(wire_d89_84),.data_out(wire_d89_85),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9008986(.data_in(wire_d89_85),.data_out(wire_d89_86),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9008987(.data_in(wire_d89_86),.data_out(wire_d89_87),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9008988(.data_in(wire_d89_87),.data_out(wire_d89_88),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9008989(.data_in(wire_d89_88),.data_out(wire_d89_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9008990(.data_in(wire_d89_89),.data_out(wire_d89_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9008991(.data_in(wire_d89_90),.data_out(wire_d89_91),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9008992(.data_in(wire_d89_91),.data_out(wire_d89_92),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9008993(.data_in(wire_d89_92),.data_out(wire_d89_93),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9008994(.data_in(wire_d89_93),.data_out(wire_d89_94),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9008995(.data_in(wire_d89_94),.data_out(wire_d89_95),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9008996(.data_in(wire_d89_95),.data_out(wire_d89_96),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9008997(.data_in(wire_d89_96),.data_out(wire_d89_97),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9008998(.data_in(wire_d89_97),.data_out(wire_d89_98),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9008999(.data_in(wire_d89_98),.data_out(wire_d89_99),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance90089100(.data_in(wire_d89_99),.data_out(wire_d89_100),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance90089101(.data_in(wire_d89_100),.data_out(wire_d89_101),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance90089102(.data_in(wire_d89_101),.data_out(wire_d89_102),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance90089103(.data_in(wire_d89_102),.data_out(wire_d89_103),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance90089104(.data_in(wire_d89_103),.data_out(wire_d89_104),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance90089105(.data_in(wire_d89_104),.data_out(wire_d89_105),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance90089106(.data_in(wire_d89_105),.data_out(wire_d89_106),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance90089107(.data_in(wire_d89_106),.data_out(wire_d89_107),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance90089108(.data_in(wire_d89_107),.data_out(wire_d89_108),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance90089109(.data_in(wire_d89_108),.data_out(wire_d89_109),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance90089110(.data_in(wire_d89_109),.data_out(wire_d89_110),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance90089111(.data_in(wire_d89_110),.data_out(wire_d89_111),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance90089112(.data_in(wire_d89_111),.data_out(wire_d89_112),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance90089113(.data_in(wire_d89_112),.data_out(wire_d89_113),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance90089114(.data_in(wire_d89_113),.data_out(wire_d89_114),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance90089115(.data_in(wire_d89_114),.data_out(wire_d89_115),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance90089116(.data_in(wire_d89_115),.data_out(wire_d89_116),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance90089117(.data_in(wire_d89_116),.data_out(wire_d89_117),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance90089118(.data_in(wire_d89_117),.data_out(wire_d89_118),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance90089119(.data_in(wire_d89_118),.data_out(d_out89),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance910900(.data_in(d_in90),.data_out(wire_d90_0),.clk(clk),.rst(rst));            //channel 91
	register #(.WIDTH(WIDTH)) register_instance910901(.data_in(wire_d90_0),.data_out(wire_d90_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance910902(.data_in(wire_d90_1),.data_out(wire_d90_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance910903(.data_in(wire_d90_2),.data_out(wire_d90_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance910904(.data_in(wire_d90_3),.data_out(wire_d90_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance910905(.data_in(wire_d90_4),.data_out(wire_d90_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance910906(.data_in(wire_d90_5),.data_out(wire_d90_6),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance910907(.data_in(wire_d90_6),.data_out(wire_d90_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance910908(.data_in(wire_d90_7),.data_out(wire_d90_8),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance910909(.data_in(wire_d90_8),.data_out(wire_d90_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9109010(.data_in(wire_d90_9),.data_out(wire_d90_10),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9109011(.data_in(wire_d90_10),.data_out(wire_d90_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9109012(.data_in(wire_d90_11),.data_out(wire_d90_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9109013(.data_in(wire_d90_12),.data_out(wire_d90_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9109014(.data_in(wire_d90_13),.data_out(wire_d90_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9109015(.data_in(wire_d90_14),.data_out(wire_d90_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9109016(.data_in(wire_d90_15),.data_out(wire_d90_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9109017(.data_in(wire_d90_16),.data_out(wire_d90_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9109018(.data_in(wire_d90_17),.data_out(wire_d90_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9109019(.data_in(wire_d90_18),.data_out(wire_d90_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9109020(.data_in(wire_d90_19),.data_out(wire_d90_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9109021(.data_in(wire_d90_20),.data_out(wire_d90_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9109022(.data_in(wire_d90_21),.data_out(wire_d90_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9109023(.data_in(wire_d90_22),.data_out(wire_d90_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9109024(.data_in(wire_d90_23),.data_out(wire_d90_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9109025(.data_in(wire_d90_24),.data_out(wire_d90_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9109026(.data_in(wire_d90_25),.data_out(wire_d90_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9109027(.data_in(wire_d90_26),.data_out(wire_d90_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9109028(.data_in(wire_d90_27),.data_out(wire_d90_28),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9109029(.data_in(wire_d90_28),.data_out(wire_d90_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9109030(.data_in(wire_d90_29),.data_out(wire_d90_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9109031(.data_in(wire_d90_30),.data_out(wire_d90_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9109032(.data_in(wire_d90_31),.data_out(wire_d90_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9109033(.data_in(wire_d90_32),.data_out(wire_d90_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9109034(.data_in(wire_d90_33),.data_out(wire_d90_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9109035(.data_in(wire_d90_34),.data_out(wire_d90_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9109036(.data_in(wire_d90_35),.data_out(wire_d90_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9109037(.data_in(wire_d90_36),.data_out(wire_d90_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9109038(.data_in(wire_d90_37),.data_out(wire_d90_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9109039(.data_in(wire_d90_38),.data_out(wire_d90_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9109040(.data_in(wire_d90_39),.data_out(wire_d90_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9109041(.data_in(wire_d90_40),.data_out(wire_d90_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9109042(.data_in(wire_d90_41),.data_out(wire_d90_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9109043(.data_in(wire_d90_42),.data_out(wire_d90_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9109044(.data_in(wire_d90_43),.data_out(wire_d90_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9109045(.data_in(wire_d90_44),.data_out(wire_d90_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9109046(.data_in(wire_d90_45),.data_out(wire_d90_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9109047(.data_in(wire_d90_46),.data_out(wire_d90_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9109048(.data_in(wire_d90_47),.data_out(wire_d90_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9109049(.data_in(wire_d90_48),.data_out(wire_d90_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9109050(.data_in(wire_d90_49),.data_out(wire_d90_50),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9109051(.data_in(wire_d90_50),.data_out(wire_d90_51),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9109052(.data_in(wire_d90_51),.data_out(wire_d90_52),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9109053(.data_in(wire_d90_52),.data_out(wire_d90_53),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9109054(.data_in(wire_d90_53),.data_out(wire_d90_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9109055(.data_in(wire_d90_54),.data_out(wire_d90_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9109056(.data_in(wire_d90_55),.data_out(wire_d90_56),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9109057(.data_in(wire_d90_56),.data_out(wire_d90_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9109058(.data_in(wire_d90_57),.data_out(wire_d90_58),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9109059(.data_in(wire_d90_58),.data_out(wire_d90_59),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9109060(.data_in(wire_d90_59),.data_out(wire_d90_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9109061(.data_in(wire_d90_60),.data_out(wire_d90_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9109062(.data_in(wire_d90_61),.data_out(wire_d90_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9109063(.data_in(wire_d90_62),.data_out(wire_d90_63),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9109064(.data_in(wire_d90_63),.data_out(wire_d90_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9109065(.data_in(wire_d90_64),.data_out(wire_d90_65),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9109066(.data_in(wire_d90_65),.data_out(wire_d90_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9109067(.data_in(wire_d90_66),.data_out(wire_d90_67),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9109068(.data_in(wire_d90_67),.data_out(wire_d90_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9109069(.data_in(wire_d90_68),.data_out(wire_d90_69),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9109070(.data_in(wire_d90_69),.data_out(wire_d90_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9109071(.data_in(wire_d90_70),.data_out(wire_d90_71),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9109072(.data_in(wire_d90_71),.data_out(wire_d90_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9109073(.data_in(wire_d90_72),.data_out(wire_d90_73),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9109074(.data_in(wire_d90_73),.data_out(wire_d90_74),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9109075(.data_in(wire_d90_74),.data_out(wire_d90_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9109076(.data_in(wire_d90_75),.data_out(wire_d90_76),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9109077(.data_in(wire_d90_76),.data_out(wire_d90_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9109078(.data_in(wire_d90_77),.data_out(wire_d90_78),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9109079(.data_in(wire_d90_78),.data_out(wire_d90_79),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9109080(.data_in(wire_d90_79),.data_out(wire_d90_80),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9109081(.data_in(wire_d90_80),.data_out(wire_d90_81),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9109082(.data_in(wire_d90_81),.data_out(wire_d90_82),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9109083(.data_in(wire_d90_82),.data_out(wire_d90_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9109084(.data_in(wire_d90_83),.data_out(wire_d90_84),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9109085(.data_in(wire_d90_84),.data_out(wire_d90_85),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9109086(.data_in(wire_d90_85),.data_out(wire_d90_86),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9109087(.data_in(wire_d90_86),.data_out(wire_d90_87),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9109088(.data_in(wire_d90_87),.data_out(wire_d90_88),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9109089(.data_in(wire_d90_88),.data_out(wire_d90_89),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9109090(.data_in(wire_d90_89),.data_out(wire_d90_90),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9109091(.data_in(wire_d90_90),.data_out(wire_d90_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9109092(.data_in(wire_d90_91),.data_out(wire_d90_92),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9109093(.data_in(wire_d90_92),.data_out(wire_d90_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9109094(.data_in(wire_d90_93),.data_out(wire_d90_94),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9109095(.data_in(wire_d90_94),.data_out(wire_d90_95),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9109096(.data_in(wire_d90_95),.data_out(wire_d90_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9109097(.data_in(wire_d90_96),.data_out(wire_d90_97),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9109098(.data_in(wire_d90_97),.data_out(wire_d90_98),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9109099(.data_in(wire_d90_98),.data_out(wire_d90_99),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance91090100(.data_in(wire_d90_99),.data_out(wire_d90_100),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance91090101(.data_in(wire_d90_100),.data_out(wire_d90_101),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance91090102(.data_in(wire_d90_101),.data_out(wire_d90_102),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance91090103(.data_in(wire_d90_102),.data_out(wire_d90_103),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance91090104(.data_in(wire_d90_103),.data_out(wire_d90_104),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance91090105(.data_in(wire_d90_104),.data_out(wire_d90_105),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance91090106(.data_in(wire_d90_105),.data_out(wire_d90_106),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance91090107(.data_in(wire_d90_106),.data_out(wire_d90_107),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance91090108(.data_in(wire_d90_107),.data_out(wire_d90_108),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance91090109(.data_in(wire_d90_108),.data_out(wire_d90_109),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance91090110(.data_in(wire_d90_109),.data_out(wire_d90_110),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance91090111(.data_in(wire_d90_110),.data_out(wire_d90_111),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance91090112(.data_in(wire_d90_111),.data_out(wire_d90_112),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance91090113(.data_in(wire_d90_112),.data_out(wire_d90_113),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance91090114(.data_in(wire_d90_113),.data_out(wire_d90_114),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance91090115(.data_in(wire_d90_114),.data_out(wire_d90_115),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance91090116(.data_in(wire_d90_115),.data_out(wire_d90_116),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance91090117(.data_in(wire_d90_116),.data_out(wire_d90_117),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance91090118(.data_in(wire_d90_117),.data_out(wire_d90_118),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance91090119(.data_in(wire_d90_118),.data_out(d_out90),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance920910(.data_in(d_in91),.data_out(wire_d91_0),.clk(clk),.rst(rst));            //channel 92
	large_mux #(.WIDTH(WIDTH)) large_mux_instance920911(.data_in(wire_d91_0),.data_out(wire_d91_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance920912(.data_in(wire_d91_1),.data_out(wire_d91_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance920913(.data_in(wire_d91_2),.data_out(wire_d91_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance920914(.data_in(wire_d91_3),.data_out(wire_d91_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance920915(.data_in(wire_d91_4),.data_out(wire_d91_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance920916(.data_in(wire_d91_5),.data_out(wire_d91_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance920917(.data_in(wire_d91_6),.data_out(wire_d91_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance920918(.data_in(wire_d91_7),.data_out(wire_d91_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance920919(.data_in(wire_d91_8),.data_out(wire_d91_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9209110(.data_in(wire_d91_9),.data_out(wire_d91_10),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9209111(.data_in(wire_d91_10),.data_out(wire_d91_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9209112(.data_in(wire_d91_11),.data_out(wire_d91_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9209113(.data_in(wire_d91_12),.data_out(wire_d91_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9209114(.data_in(wire_d91_13),.data_out(wire_d91_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9209115(.data_in(wire_d91_14),.data_out(wire_d91_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9209116(.data_in(wire_d91_15),.data_out(wire_d91_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9209117(.data_in(wire_d91_16),.data_out(wire_d91_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9209118(.data_in(wire_d91_17),.data_out(wire_d91_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9209119(.data_in(wire_d91_18),.data_out(wire_d91_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9209120(.data_in(wire_d91_19),.data_out(wire_d91_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9209121(.data_in(wire_d91_20),.data_out(wire_d91_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9209122(.data_in(wire_d91_21),.data_out(wire_d91_22),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9209123(.data_in(wire_d91_22),.data_out(wire_d91_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9209124(.data_in(wire_d91_23),.data_out(wire_d91_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9209125(.data_in(wire_d91_24),.data_out(wire_d91_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9209126(.data_in(wire_d91_25),.data_out(wire_d91_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9209127(.data_in(wire_d91_26),.data_out(wire_d91_27),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9209128(.data_in(wire_d91_27),.data_out(wire_d91_28),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9209129(.data_in(wire_d91_28),.data_out(wire_d91_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9209130(.data_in(wire_d91_29),.data_out(wire_d91_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9209131(.data_in(wire_d91_30),.data_out(wire_d91_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9209132(.data_in(wire_d91_31),.data_out(wire_d91_32),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9209133(.data_in(wire_d91_32),.data_out(wire_d91_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9209134(.data_in(wire_d91_33),.data_out(wire_d91_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9209135(.data_in(wire_d91_34),.data_out(wire_d91_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9209136(.data_in(wire_d91_35),.data_out(wire_d91_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9209137(.data_in(wire_d91_36),.data_out(wire_d91_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9209138(.data_in(wire_d91_37),.data_out(wire_d91_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9209139(.data_in(wire_d91_38),.data_out(wire_d91_39),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9209140(.data_in(wire_d91_39),.data_out(wire_d91_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9209141(.data_in(wire_d91_40),.data_out(wire_d91_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9209142(.data_in(wire_d91_41),.data_out(wire_d91_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9209143(.data_in(wire_d91_42),.data_out(wire_d91_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9209144(.data_in(wire_d91_43),.data_out(wire_d91_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9209145(.data_in(wire_d91_44),.data_out(wire_d91_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9209146(.data_in(wire_d91_45),.data_out(wire_d91_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9209147(.data_in(wire_d91_46),.data_out(wire_d91_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9209148(.data_in(wire_d91_47),.data_out(wire_d91_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9209149(.data_in(wire_d91_48),.data_out(wire_d91_49),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9209150(.data_in(wire_d91_49),.data_out(wire_d91_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9209151(.data_in(wire_d91_50),.data_out(wire_d91_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9209152(.data_in(wire_d91_51),.data_out(wire_d91_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9209153(.data_in(wire_d91_52),.data_out(wire_d91_53),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9209154(.data_in(wire_d91_53),.data_out(wire_d91_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9209155(.data_in(wire_d91_54),.data_out(wire_d91_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9209156(.data_in(wire_d91_55),.data_out(wire_d91_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9209157(.data_in(wire_d91_56),.data_out(wire_d91_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9209158(.data_in(wire_d91_57),.data_out(wire_d91_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9209159(.data_in(wire_d91_58),.data_out(wire_d91_59),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9209160(.data_in(wire_d91_59),.data_out(wire_d91_60),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9209161(.data_in(wire_d91_60),.data_out(wire_d91_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9209162(.data_in(wire_d91_61),.data_out(wire_d91_62),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9209163(.data_in(wire_d91_62),.data_out(wire_d91_63),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9209164(.data_in(wire_d91_63),.data_out(wire_d91_64),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9209165(.data_in(wire_d91_64),.data_out(wire_d91_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9209166(.data_in(wire_d91_65),.data_out(wire_d91_66),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9209167(.data_in(wire_d91_66),.data_out(wire_d91_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9209168(.data_in(wire_d91_67),.data_out(wire_d91_68),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9209169(.data_in(wire_d91_68),.data_out(wire_d91_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9209170(.data_in(wire_d91_69),.data_out(wire_d91_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9209171(.data_in(wire_d91_70),.data_out(wire_d91_71),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9209172(.data_in(wire_d91_71),.data_out(wire_d91_72),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9209173(.data_in(wire_d91_72),.data_out(wire_d91_73),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9209174(.data_in(wire_d91_73),.data_out(wire_d91_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9209175(.data_in(wire_d91_74),.data_out(wire_d91_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9209176(.data_in(wire_d91_75),.data_out(wire_d91_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9209177(.data_in(wire_d91_76),.data_out(wire_d91_77),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9209178(.data_in(wire_d91_77),.data_out(wire_d91_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9209179(.data_in(wire_d91_78),.data_out(wire_d91_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9209180(.data_in(wire_d91_79),.data_out(wire_d91_80),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9209181(.data_in(wire_d91_80),.data_out(wire_d91_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9209182(.data_in(wire_d91_81),.data_out(wire_d91_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9209183(.data_in(wire_d91_82),.data_out(wire_d91_83),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9209184(.data_in(wire_d91_83),.data_out(wire_d91_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9209185(.data_in(wire_d91_84),.data_out(wire_d91_85),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9209186(.data_in(wire_d91_85),.data_out(wire_d91_86),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9209187(.data_in(wire_d91_86),.data_out(wire_d91_87),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9209188(.data_in(wire_d91_87),.data_out(wire_d91_88),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9209189(.data_in(wire_d91_88),.data_out(wire_d91_89),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9209190(.data_in(wire_d91_89),.data_out(wire_d91_90),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9209191(.data_in(wire_d91_90),.data_out(wire_d91_91),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9209192(.data_in(wire_d91_91),.data_out(wire_d91_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9209193(.data_in(wire_d91_92),.data_out(wire_d91_93),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9209194(.data_in(wire_d91_93),.data_out(wire_d91_94),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9209195(.data_in(wire_d91_94),.data_out(wire_d91_95),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9209196(.data_in(wire_d91_95),.data_out(wire_d91_96),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9209197(.data_in(wire_d91_96),.data_out(wire_d91_97),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9209198(.data_in(wire_d91_97),.data_out(wire_d91_98),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9209199(.data_in(wire_d91_98),.data_out(wire_d91_99),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance92091100(.data_in(wire_d91_99),.data_out(wire_d91_100),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance92091101(.data_in(wire_d91_100),.data_out(wire_d91_101),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance92091102(.data_in(wire_d91_101),.data_out(wire_d91_102),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance92091103(.data_in(wire_d91_102),.data_out(wire_d91_103),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance92091104(.data_in(wire_d91_103),.data_out(wire_d91_104),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance92091105(.data_in(wire_d91_104),.data_out(wire_d91_105),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance92091106(.data_in(wire_d91_105),.data_out(wire_d91_106),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance92091107(.data_in(wire_d91_106),.data_out(wire_d91_107),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance92091108(.data_in(wire_d91_107),.data_out(wire_d91_108),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance92091109(.data_in(wire_d91_108),.data_out(wire_d91_109),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance92091110(.data_in(wire_d91_109),.data_out(wire_d91_110),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance92091111(.data_in(wire_d91_110),.data_out(wire_d91_111),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance92091112(.data_in(wire_d91_111),.data_out(wire_d91_112),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance92091113(.data_in(wire_d91_112),.data_out(wire_d91_113),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance92091114(.data_in(wire_d91_113),.data_out(wire_d91_114),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance92091115(.data_in(wire_d91_114),.data_out(wire_d91_115),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance92091116(.data_in(wire_d91_115),.data_out(wire_d91_116),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance92091117(.data_in(wire_d91_116),.data_out(wire_d91_117),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance92091118(.data_in(wire_d91_117),.data_out(wire_d91_118),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance92091119(.data_in(wire_d91_118),.data_out(d_out91),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance930920(.data_in(d_in92),.data_out(wire_d92_0),.clk(clk),.rst(rst));            //channel 93
	encoder #(.WIDTH(WIDTH)) encoder_instance930921(.data_in(wire_d92_0),.data_out(wire_d92_1),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance930922(.data_in(wire_d92_1),.data_out(wire_d92_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance930923(.data_in(wire_d92_2),.data_out(wire_d92_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance930924(.data_in(wire_d92_3),.data_out(wire_d92_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance930925(.data_in(wire_d92_4),.data_out(wire_d92_5),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance930926(.data_in(wire_d92_5),.data_out(wire_d92_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance930927(.data_in(wire_d92_6),.data_out(wire_d92_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance930928(.data_in(wire_d92_7),.data_out(wire_d92_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance930929(.data_in(wire_d92_8),.data_out(wire_d92_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9309210(.data_in(wire_d92_9),.data_out(wire_d92_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9309211(.data_in(wire_d92_10),.data_out(wire_d92_11),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9309212(.data_in(wire_d92_11),.data_out(wire_d92_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9309213(.data_in(wire_d92_12),.data_out(wire_d92_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9309214(.data_in(wire_d92_13),.data_out(wire_d92_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9309215(.data_in(wire_d92_14),.data_out(wire_d92_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9309216(.data_in(wire_d92_15),.data_out(wire_d92_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9309217(.data_in(wire_d92_16),.data_out(wire_d92_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9309218(.data_in(wire_d92_17),.data_out(wire_d92_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9309219(.data_in(wire_d92_18),.data_out(wire_d92_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9309220(.data_in(wire_d92_19),.data_out(wire_d92_20),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9309221(.data_in(wire_d92_20),.data_out(wire_d92_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9309222(.data_in(wire_d92_21),.data_out(wire_d92_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9309223(.data_in(wire_d92_22),.data_out(wire_d92_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9309224(.data_in(wire_d92_23),.data_out(wire_d92_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9309225(.data_in(wire_d92_24),.data_out(wire_d92_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9309226(.data_in(wire_d92_25),.data_out(wire_d92_26),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9309227(.data_in(wire_d92_26),.data_out(wire_d92_27),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9309228(.data_in(wire_d92_27),.data_out(wire_d92_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9309229(.data_in(wire_d92_28),.data_out(wire_d92_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9309230(.data_in(wire_d92_29),.data_out(wire_d92_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9309231(.data_in(wire_d92_30),.data_out(wire_d92_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9309232(.data_in(wire_d92_31),.data_out(wire_d92_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9309233(.data_in(wire_d92_32),.data_out(wire_d92_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9309234(.data_in(wire_d92_33),.data_out(wire_d92_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9309235(.data_in(wire_d92_34),.data_out(wire_d92_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9309236(.data_in(wire_d92_35),.data_out(wire_d92_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9309237(.data_in(wire_d92_36),.data_out(wire_d92_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9309238(.data_in(wire_d92_37),.data_out(wire_d92_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9309239(.data_in(wire_d92_38),.data_out(wire_d92_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9309240(.data_in(wire_d92_39),.data_out(wire_d92_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9309241(.data_in(wire_d92_40),.data_out(wire_d92_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9309242(.data_in(wire_d92_41),.data_out(wire_d92_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9309243(.data_in(wire_d92_42),.data_out(wire_d92_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9309244(.data_in(wire_d92_43),.data_out(wire_d92_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9309245(.data_in(wire_d92_44),.data_out(wire_d92_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9309246(.data_in(wire_d92_45),.data_out(wire_d92_46),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9309247(.data_in(wire_d92_46),.data_out(wire_d92_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9309248(.data_in(wire_d92_47),.data_out(wire_d92_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9309249(.data_in(wire_d92_48),.data_out(wire_d92_49),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9309250(.data_in(wire_d92_49),.data_out(wire_d92_50),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9309251(.data_in(wire_d92_50),.data_out(wire_d92_51),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9309252(.data_in(wire_d92_51),.data_out(wire_d92_52),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9309253(.data_in(wire_d92_52),.data_out(wire_d92_53),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9309254(.data_in(wire_d92_53),.data_out(wire_d92_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9309255(.data_in(wire_d92_54),.data_out(wire_d92_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9309256(.data_in(wire_d92_55),.data_out(wire_d92_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9309257(.data_in(wire_d92_56),.data_out(wire_d92_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9309258(.data_in(wire_d92_57),.data_out(wire_d92_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9309259(.data_in(wire_d92_58),.data_out(wire_d92_59),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9309260(.data_in(wire_d92_59),.data_out(wire_d92_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9309261(.data_in(wire_d92_60),.data_out(wire_d92_61),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9309262(.data_in(wire_d92_61),.data_out(wire_d92_62),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9309263(.data_in(wire_d92_62),.data_out(wire_d92_63),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9309264(.data_in(wire_d92_63),.data_out(wire_d92_64),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9309265(.data_in(wire_d92_64),.data_out(wire_d92_65),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9309266(.data_in(wire_d92_65),.data_out(wire_d92_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9309267(.data_in(wire_d92_66),.data_out(wire_d92_67),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9309268(.data_in(wire_d92_67),.data_out(wire_d92_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9309269(.data_in(wire_d92_68),.data_out(wire_d92_69),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9309270(.data_in(wire_d92_69),.data_out(wire_d92_70),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9309271(.data_in(wire_d92_70),.data_out(wire_d92_71),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9309272(.data_in(wire_d92_71),.data_out(wire_d92_72),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9309273(.data_in(wire_d92_72),.data_out(wire_d92_73),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9309274(.data_in(wire_d92_73),.data_out(wire_d92_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9309275(.data_in(wire_d92_74),.data_out(wire_d92_75),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9309276(.data_in(wire_d92_75),.data_out(wire_d92_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9309277(.data_in(wire_d92_76),.data_out(wire_d92_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9309278(.data_in(wire_d92_77),.data_out(wire_d92_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9309279(.data_in(wire_d92_78),.data_out(wire_d92_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9309280(.data_in(wire_d92_79),.data_out(wire_d92_80),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9309281(.data_in(wire_d92_80),.data_out(wire_d92_81),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9309282(.data_in(wire_d92_81),.data_out(wire_d92_82),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9309283(.data_in(wire_d92_82),.data_out(wire_d92_83),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9309284(.data_in(wire_d92_83),.data_out(wire_d92_84),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9309285(.data_in(wire_d92_84),.data_out(wire_d92_85),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9309286(.data_in(wire_d92_85),.data_out(wire_d92_86),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9309287(.data_in(wire_d92_86),.data_out(wire_d92_87),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9309288(.data_in(wire_d92_87),.data_out(wire_d92_88),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9309289(.data_in(wire_d92_88),.data_out(wire_d92_89),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9309290(.data_in(wire_d92_89),.data_out(wire_d92_90),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9309291(.data_in(wire_d92_90),.data_out(wire_d92_91),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9309292(.data_in(wire_d92_91),.data_out(wire_d92_92),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9309293(.data_in(wire_d92_92),.data_out(wire_d92_93),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9309294(.data_in(wire_d92_93),.data_out(wire_d92_94),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9309295(.data_in(wire_d92_94),.data_out(wire_d92_95),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9309296(.data_in(wire_d92_95),.data_out(wire_d92_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9309297(.data_in(wire_d92_96),.data_out(wire_d92_97),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9309298(.data_in(wire_d92_97),.data_out(wire_d92_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9309299(.data_in(wire_d92_98),.data_out(wire_d92_99),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance93092100(.data_in(wire_d92_99),.data_out(wire_d92_100),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance93092101(.data_in(wire_d92_100),.data_out(wire_d92_101),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance93092102(.data_in(wire_d92_101),.data_out(wire_d92_102),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance93092103(.data_in(wire_d92_102),.data_out(wire_d92_103),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance93092104(.data_in(wire_d92_103),.data_out(wire_d92_104),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance93092105(.data_in(wire_d92_104),.data_out(wire_d92_105),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance93092106(.data_in(wire_d92_105),.data_out(wire_d92_106),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance93092107(.data_in(wire_d92_106),.data_out(wire_d92_107),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance93092108(.data_in(wire_d92_107),.data_out(wire_d92_108),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance93092109(.data_in(wire_d92_108),.data_out(wire_d92_109),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance93092110(.data_in(wire_d92_109),.data_out(wire_d92_110),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance93092111(.data_in(wire_d92_110),.data_out(wire_d92_111),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance93092112(.data_in(wire_d92_111),.data_out(wire_d92_112),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance93092113(.data_in(wire_d92_112),.data_out(wire_d92_113),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance93092114(.data_in(wire_d92_113),.data_out(wire_d92_114),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance93092115(.data_in(wire_d92_114),.data_out(wire_d92_115),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance93092116(.data_in(wire_d92_115),.data_out(wire_d92_116),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance93092117(.data_in(wire_d92_116),.data_out(wire_d92_117),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance93092118(.data_in(wire_d92_117),.data_out(wire_d92_118),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance93092119(.data_in(wire_d92_118),.data_out(d_out92),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance940930(.data_in(d_in93),.data_out(wire_d93_0),.clk(clk),.rst(rst));            //channel 94
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance940931(.data_in(wire_d93_0),.data_out(wire_d93_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance940932(.data_in(wire_d93_1),.data_out(wire_d93_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance940933(.data_in(wire_d93_2),.data_out(wire_d93_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance940934(.data_in(wire_d93_3),.data_out(wire_d93_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance940935(.data_in(wire_d93_4),.data_out(wire_d93_5),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance940936(.data_in(wire_d93_5),.data_out(wire_d93_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance940937(.data_in(wire_d93_6),.data_out(wire_d93_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance940938(.data_in(wire_d93_7),.data_out(wire_d93_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance940939(.data_in(wire_d93_8),.data_out(wire_d93_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9409310(.data_in(wire_d93_9),.data_out(wire_d93_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9409311(.data_in(wire_d93_10),.data_out(wire_d93_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9409312(.data_in(wire_d93_11),.data_out(wire_d93_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9409313(.data_in(wire_d93_12),.data_out(wire_d93_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9409314(.data_in(wire_d93_13),.data_out(wire_d93_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9409315(.data_in(wire_d93_14),.data_out(wire_d93_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9409316(.data_in(wire_d93_15),.data_out(wire_d93_16),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9409317(.data_in(wire_d93_16),.data_out(wire_d93_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9409318(.data_in(wire_d93_17),.data_out(wire_d93_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9409319(.data_in(wire_d93_18),.data_out(wire_d93_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9409320(.data_in(wire_d93_19),.data_out(wire_d93_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9409321(.data_in(wire_d93_20),.data_out(wire_d93_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9409322(.data_in(wire_d93_21),.data_out(wire_d93_22),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9409323(.data_in(wire_d93_22),.data_out(wire_d93_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9409324(.data_in(wire_d93_23),.data_out(wire_d93_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9409325(.data_in(wire_d93_24),.data_out(wire_d93_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9409326(.data_in(wire_d93_25),.data_out(wire_d93_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9409327(.data_in(wire_d93_26),.data_out(wire_d93_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9409328(.data_in(wire_d93_27),.data_out(wire_d93_28),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9409329(.data_in(wire_d93_28),.data_out(wire_d93_29),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9409330(.data_in(wire_d93_29),.data_out(wire_d93_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9409331(.data_in(wire_d93_30),.data_out(wire_d93_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9409332(.data_in(wire_d93_31),.data_out(wire_d93_32),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9409333(.data_in(wire_d93_32),.data_out(wire_d93_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9409334(.data_in(wire_d93_33),.data_out(wire_d93_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9409335(.data_in(wire_d93_34),.data_out(wire_d93_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9409336(.data_in(wire_d93_35),.data_out(wire_d93_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9409337(.data_in(wire_d93_36),.data_out(wire_d93_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9409338(.data_in(wire_d93_37),.data_out(wire_d93_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9409339(.data_in(wire_d93_38),.data_out(wire_d93_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9409340(.data_in(wire_d93_39),.data_out(wire_d93_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9409341(.data_in(wire_d93_40),.data_out(wire_d93_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9409342(.data_in(wire_d93_41),.data_out(wire_d93_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9409343(.data_in(wire_d93_42),.data_out(wire_d93_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9409344(.data_in(wire_d93_43),.data_out(wire_d93_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9409345(.data_in(wire_d93_44),.data_out(wire_d93_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9409346(.data_in(wire_d93_45),.data_out(wire_d93_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9409347(.data_in(wire_d93_46),.data_out(wire_d93_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9409348(.data_in(wire_d93_47),.data_out(wire_d93_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9409349(.data_in(wire_d93_48),.data_out(wire_d93_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9409350(.data_in(wire_d93_49),.data_out(wire_d93_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9409351(.data_in(wire_d93_50),.data_out(wire_d93_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9409352(.data_in(wire_d93_51),.data_out(wire_d93_52),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9409353(.data_in(wire_d93_52),.data_out(wire_d93_53),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9409354(.data_in(wire_d93_53),.data_out(wire_d93_54),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9409355(.data_in(wire_d93_54),.data_out(wire_d93_55),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9409356(.data_in(wire_d93_55),.data_out(wire_d93_56),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9409357(.data_in(wire_d93_56),.data_out(wire_d93_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9409358(.data_in(wire_d93_57),.data_out(wire_d93_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9409359(.data_in(wire_d93_58),.data_out(wire_d93_59),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9409360(.data_in(wire_d93_59),.data_out(wire_d93_60),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9409361(.data_in(wire_d93_60),.data_out(wire_d93_61),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9409362(.data_in(wire_d93_61),.data_out(wire_d93_62),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9409363(.data_in(wire_d93_62),.data_out(wire_d93_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9409364(.data_in(wire_d93_63),.data_out(wire_d93_64),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9409365(.data_in(wire_d93_64),.data_out(wire_d93_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9409366(.data_in(wire_d93_65),.data_out(wire_d93_66),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9409367(.data_in(wire_d93_66),.data_out(wire_d93_67),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9409368(.data_in(wire_d93_67),.data_out(wire_d93_68),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9409369(.data_in(wire_d93_68),.data_out(wire_d93_69),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9409370(.data_in(wire_d93_69),.data_out(wire_d93_70),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9409371(.data_in(wire_d93_70),.data_out(wire_d93_71),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9409372(.data_in(wire_d93_71),.data_out(wire_d93_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9409373(.data_in(wire_d93_72),.data_out(wire_d93_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9409374(.data_in(wire_d93_73),.data_out(wire_d93_74),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9409375(.data_in(wire_d93_74),.data_out(wire_d93_75),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9409376(.data_in(wire_d93_75),.data_out(wire_d93_76),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9409377(.data_in(wire_d93_76),.data_out(wire_d93_77),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9409378(.data_in(wire_d93_77),.data_out(wire_d93_78),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9409379(.data_in(wire_d93_78),.data_out(wire_d93_79),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9409380(.data_in(wire_d93_79),.data_out(wire_d93_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9409381(.data_in(wire_d93_80),.data_out(wire_d93_81),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9409382(.data_in(wire_d93_81),.data_out(wire_d93_82),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9409383(.data_in(wire_d93_82),.data_out(wire_d93_83),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9409384(.data_in(wire_d93_83),.data_out(wire_d93_84),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9409385(.data_in(wire_d93_84),.data_out(wire_d93_85),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9409386(.data_in(wire_d93_85),.data_out(wire_d93_86),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9409387(.data_in(wire_d93_86),.data_out(wire_d93_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9409388(.data_in(wire_d93_87),.data_out(wire_d93_88),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9409389(.data_in(wire_d93_88),.data_out(wire_d93_89),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9409390(.data_in(wire_d93_89),.data_out(wire_d93_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9409391(.data_in(wire_d93_90),.data_out(wire_d93_91),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9409392(.data_in(wire_d93_91),.data_out(wire_d93_92),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9409393(.data_in(wire_d93_92),.data_out(wire_d93_93),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9409394(.data_in(wire_d93_93),.data_out(wire_d93_94),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9409395(.data_in(wire_d93_94),.data_out(wire_d93_95),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9409396(.data_in(wire_d93_95),.data_out(wire_d93_96),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9409397(.data_in(wire_d93_96),.data_out(wire_d93_97),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9409398(.data_in(wire_d93_97),.data_out(wire_d93_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9409399(.data_in(wire_d93_98),.data_out(wire_d93_99),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance94093100(.data_in(wire_d93_99),.data_out(wire_d93_100),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance94093101(.data_in(wire_d93_100),.data_out(wire_d93_101),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance94093102(.data_in(wire_d93_101),.data_out(wire_d93_102),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance94093103(.data_in(wire_d93_102),.data_out(wire_d93_103),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance94093104(.data_in(wire_d93_103),.data_out(wire_d93_104),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance94093105(.data_in(wire_d93_104),.data_out(wire_d93_105),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance94093106(.data_in(wire_d93_105),.data_out(wire_d93_106),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance94093107(.data_in(wire_d93_106),.data_out(wire_d93_107),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance94093108(.data_in(wire_d93_107),.data_out(wire_d93_108),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance94093109(.data_in(wire_d93_108),.data_out(wire_d93_109),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance94093110(.data_in(wire_d93_109),.data_out(wire_d93_110),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance94093111(.data_in(wire_d93_110),.data_out(wire_d93_111),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance94093112(.data_in(wire_d93_111),.data_out(wire_d93_112),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance94093113(.data_in(wire_d93_112),.data_out(wire_d93_113),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance94093114(.data_in(wire_d93_113),.data_out(wire_d93_114),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance94093115(.data_in(wire_d93_114),.data_out(wire_d93_115),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance94093116(.data_in(wire_d93_115),.data_out(wire_d93_116),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance94093117(.data_in(wire_d93_116),.data_out(wire_d93_117),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance94093118(.data_in(wire_d93_117),.data_out(wire_d93_118),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance94093119(.data_in(wire_d93_118),.data_out(d_out93),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance950940(.data_in(d_in94),.data_out(wire_d94_0),.clk(clk),.rst(rst));            //channel 95
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance950941(.data_in(wire_d94_0),.data_out(wire_d94_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance950942(.data_in(wire_d94_1),.data_out(wire_d94_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance950943(.data_in(wire_d94_2),.data_out(wire_d94_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance950944(.data_in(wire_d94_3),.data_out(wire_d94_4),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance950945(.data_in(wire_d94_4),.data_out(wire_d94_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance950946(.data_in(wire_d94_5),.data_out(wire_d94_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance950947(.data_in(wire_d94_6),.data_out(wire_d94_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance950948(.data_in(wire_d94_7),.data_out(wire_d94_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance950949(.data_in(wire_d94_8),.data_out(wire_d94_9),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9509410(.data_in(wire_d94_9),.data_out(wire_d94_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9509411(.data_in(wire_d94_10),.data_out(wire_d94_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9509412(.data_in(wire_d94_11),.data_out(wire_d94_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9509413(.data_in(wire_d94_12),.data_out(wire_d94_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9509414(.data_in(wire_d94_13),.data_out(wire_d94_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9509415(.data_in(wire_d94_14),.data_out(wire_d94_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9509416(.data_in(wire_d94_15),.data_out(wire_d94_16),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9509417(.data_in(wire_d94_16),.data_out(wire_d94_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9509418(.data_in(wire_d94_17),.data_out(wire_d94_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9509419(.data_in(wire_d94_18),.data_out(wire_d94_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9509420(.data_in(wire_d94_19),.data_out(wire_d94_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9509421(.data_in(wire_d94_20),.data_out(wire_d94_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9509422(.data_in(wire_d94_21),.data_out(wire_d94_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9509423(.data_in(wire_d94_22),.data_out(wire_d94_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9509424(.data_in(wire_d94_23),.data_out(wire_d94_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9509425(.data_in(wire_d94_24),.data_out(wire_d94_25),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9509426(.data_in(wire_d94_25),.data_out(wire_d94_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9509427(.data_in(wire_d94_26),.data_out(wire_d94_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9509428(.data_in(wire_d94_27),.data_out(wire_d94_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9509429(.data_in(wire_d94_28),.data_out(wire_d94_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9509430(.data_in(wire_d94_29),.data_out(wire_d94_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9509431(.data_in(wire_d94_30),.data_out(wire_d94_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9509432(.data_in(wire_d94_31),.data_out(wire_d94_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9509433(.data_in(wire_d94_32),.data_out(wire_d94_33),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9509434(.data_in(wire_d94_33),.data_out(wire_d94_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9509435(.data_in(wire_d94_34),.data_out(wire_d94_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9509436(.data_in(wire_d94_35),.data_out(wire_d94_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9509437(.data_in(wire_d94_36),.data_out(wire_d94_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9509438(.data_in(wire_d94_37),.data_out(wire_d94_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9509439(.data_in(wire_d94_38),.data_out(wire_d94_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9509440(.data_in(wire_d94_39),.data_out(wire_d94_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9509441(.data_in(wire_d94_40),.data_out(wire_d94_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9509442(.data_in(wire_d94_41),.data_out(wire_d94_42),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9509443(.data_in(wire_d94_42),.data_out(wire_d94_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9509444(.data_in(wire_d94_43),.data_out(wire_d94_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9509445(.data_in(wire_d94_44),.data_out(wire_d94_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9509446(.data_in(wire_d94_45),.data_out(wire_d94_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9509447(.data_in(wire_d94_46),.data_out(wire_d94_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9509448(.data_in(wire_d94_47),.data_out(wire_d94_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9509449(.data_in(wire_d94_48),.data_out(wire_d94_49),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9509450(.data_in(wire_d94_49),.data_out(wire_d94_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9509451(.data_in(wire_d94_50),.data_out(wire_d94_51),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9509452(.data_in(wire_d94_51),.data_out(wire_d94_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9509453(.data_in(wire_d94_52),.data_out(wire_d94_53),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9509454(.data_in(wire_d94_53),.data_out(wire_d94_54),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9509455(.data_in(wire_d94_54),.data_out(wire_d94_55),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9509456(.data_in(wire_d94_55),.data_out(wire_d94_56),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9509457(.data_in(wire_d94_56),.data_out(wire_d94_57),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9509458(.data_in(wire_d94_57),.data_out(wire_d94_58),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9509459(.data_in(wire_d94_58),.data_out(wire_d94_59),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9509460(.data_in(wire_d94_59),.data_out(wire_d94_60),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9509461(.data_in(wire_d94_60),.data_out(wire_d94_61),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9509462(.data_in(wire_d94_61),.data_out(wire_d94_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9509463(.data_in(wire_d94_62),.data_out(wire_d94_63),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9509464(.data_in(wire_d94_63),.data_out(wire_d94_64),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9509465(.data_in(wire_d94_64),.data_out(wire_d94_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9509466(.data_in(wire_d94_65),.data_out(wire_d94_66),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9509467(.data_in(wire_d94_66),.data_out(wire_d94_67),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9509468(.data_in(wire_d94_67),.data_out(wire_d94_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9509469(.data_in(wire_d94_68),.data_out(wire_d94_69),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9509470(.data_in(wire_d94_69),.data_out(wire_d94_70),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9509471(.data_in(wire_d94_70),.data_out(wire_d94_71),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9509472(.data_in(wire_d94_71),.data_out(wire_d94_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9509473(.data_in(wire_d94_72),.data_out(wire_d94_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9509474(.data_in(wire_d94_73),.data_out(wire_d94_74),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9509475(.data_in(wire_d94_74),.data_out(wire_d94_75),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9509476(.data_in(wire_d94_75),.data_out(wire_d94_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9509477(.data_in(wire_d94_76),.data_out(wire_d94_77),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9509478(.data_in(wire_d94_77),.data_out(wire_d94_78),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9509479(.data_in(wire_d94_78),.data_out(wire_d94_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9509480(.data_in(wire_d94_79),.data_out(wire_d94_80),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9509481(.data_in(wire_d94_80),.data_out(wire_d94_81),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9509482(.data_in(wire_d94_81),.data_out(wire_d94_82),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9509483(.data_in(wire_d94_82),.data_out(wire_d94_83),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9509484(.data_in(wire_d94_83),.data_out(wire_d94_84),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9509485(.data_in(wire_d94_84),.data_out(wire_d94_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9509486(.data_in(wire_d94_85),.data_out(wire_d94_86),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9509487(.data_in(wire_d94_86),.data_out(wire_d94_87),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9509488(.data_in(wire_d94_87),.data_out(wire_d94_88),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9509489(.data_in(wire_d94_88),.data_out(wire_d94_89),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9509490(.data_in(wire_d94_89),.data_out(wire_d94_90),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9509491(.data_in(wire_d94_90),.data_out(wire_d94_91),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9509492(.data_in(wire_d94_91),.data_out(wire_d94_92),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9509493(.data_in(wire_d94_92),.data_out(wire_d94_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9509494(.data_in(wire_d94_93),.data_out(wire_d94_94),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9509495(.data_in(wire_d94_94),.data_out(wire_d94_95),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9509496(.data_in(wire_d94_95),.data_out(wire_d94_96),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9509497(.data_in(wire_d94_96),.data_out(wire_d94_97),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9509498(.data_in(wire_d94_97),.data_out(wire_d94_98),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9509499(.data_in(wire_d94_98),.data_out(wire_d94_99),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance95094100(.data_in(wire_d94_99),.data_out(wire_d94_100),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance95094101(.data_in(wire_d94_100),.data_out(wire_d94_101),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance95094102(.data_in(wire_d94_101),.data_out(wire_d94_102),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance95094103(.data_in(wire_d94_102),.data_out(wire_d94_103),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance95094104(.data_in(wire_d94_103),.data_out(wire_d94_104),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance95094105(.data_in(wire_d94_104),.data_out(wire_d94_105),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance95094106(.data_in(wire_d94_105),.data_out(wire_d94_106),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance95094107(.data_in(wire_d94_106),.data_out(wire_d94_107),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance95094108(.data_in(wire_d94_107),.data_out(wire_d94_108),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance95094109(.data_in(wire_d94_108),.data_out(wire_d94_109),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance95094110(.data_in(wire_d94_109),.data_out(wire_d94_110),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance95094111(.data_in(wire_d94_110),.data_out(wire_d94_111),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance95094112(.data_in(wire_d94_111),.data_out(wire_d94_112),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance95094113(.data_in(wire_d94_112),.data_out(wire_d94_113),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance95094114(.data_in(wire_d94_113),.data_out(wire_d94_114),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance95094115(.data_in(wire_d94_114),.data_out(wire_d94_115),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance95094116(.data_in(wire_d94_115),.data_out(wire_d94_116),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance95094117(.data_in(wire_d94_116),.data_out(wire_d94_117),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance95094118(.data_in(wire_d94_117),.data_out(wire_d94_118),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance95094119(.data_in(wire_d94_118),.data_out(d_out94),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance960950(.data_in(d_in95),.data_out(wire_d95_0),.clk(clk),.rst(rst));            //channel 96
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance960951(.data_in(wire_d95_0),.data_out(wire_d95_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance960952(.data_in(wire_d95_1),.data_out(wire_d95_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance960953(.data_in(wire_d95_2),.data_out(wire_d95_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance960954(.data_in(wire_d95_3),.data_out(wire_d95_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance960955(.data_in(wire_d95_4),.data_out(wire_d95_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance960956(.data_in(wire_d95_5),.data_out(wire_d95_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance960957(.data_in(wire_d95_6),.data_out(wire_d95_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance960958(.data_in(wire_d95_7),.data_out(wire_d95_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance960959(.data_in(wire_d95_8),.data_out(wire_d95_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9609510(.data_in(wire_d95_9),.data_out(wire_d95_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9609511(.data_in(wire_d95_10),.data_out(wire_d95_11),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9609512(.data_in(wire_d95_11),.data_out(wire_d95_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9609513(.data_in(wire_d95_12),.data_out(wire_d95_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9609514(.data_in(wire_d95_13),.data_out(wire_d95_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9609515(.data_in(wire_d95_14),.data_out(wire_d95_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9609516(.data_in(wire_d95_15),.data_out(wire_d95_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9609517(.data_in(wire_d95_16),.data_out(wire_d95_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9609518(.data_in(wire_d95_17),.data_out(wire_d95_18),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9609519(.data_in(wire_d95_18),.data_out(wire_d95_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9609520(.data_in(wire_d95_19),.data_out(wire_d95_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9609521(.data_in(wire_d95_20),.data_out(wire_d95_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9609522(.data_in(wire_d95_21),.data_out(wire_d95_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9609523(.data_in(wire_d95_22),.data_out(wire_d95_23),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9609524(.data_in(wire_d95_23),.data_out(wire_d95_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9609525(.data_in(wire_d95_24),.data_out(wire_d95_25),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9609526(.data_in(wire_d95_25),.data_out(wire_d95_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9609527(.data_in(wire_d95_26),.data_out(wire_d95_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9609528(.data_in(wire_d95_27),.data_out(wire_d95_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9609529(.data_in(wire_d95_28),.data_out(wire_d95_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9609530(.data_in(wire_d95_29),.data_out(wire_d95_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9609531(.data_in(wire_d95_30),.data_out(wire_d95_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9609532(.data_in(wire_d95_31),.data_out(wire_d95_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9609533(.data_in(wire_d95_32),.data_out(wire_d95_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9609534(.data_in(wire_d95_33),.data_out(wire_d95_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9609535(.data_in(wire_d95_34),.data_out(wire_d95_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9609536(.data_in(wire_d95_35),.data_out(wire_d95_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9609537(.data_in(wire_d95_36),.data_out(wire_d95_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9609538(.data_in(wire_d95_37),.data_out(wire_d95_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9609539(.data_in(wire_d95_38),.data_out(wire_d95_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9609540(.data_in(wire_d95_39),.data_out(wire_d95_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9609541(.data_in(wire_d95_40),.data_out(wire_d95_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9609542(.data_in(wire_d95_41),.data_out(wire_d95_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9609543(.data_in(wire_d95_42),.data_out(wire_d95_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9609544(.data_in(wire_d95_43),.data_out(wire_d95_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9609545(.data_in(wire_d95_44),.data_out(wire_d95_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9609546(.data_in(wire_d95_45),.data_out(wire_d95_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9609547(.data_in(wire_d95_46),.data_out(wire_d95_47),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9609548(.data_in(wire_d95_47),.data_out(wire_d95_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9609549(.data_in(wire_d95_48),.data_out(wire_d95_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9609550(.data_in(wire_d95_49),.data_out(wire_d95_50),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9609551(.data_in(wire_d95_50),.data_out(wire_d95_51),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9609552(.data_in(wire_d95_51),.data_out(wire_d95_52),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9609553(.data_in(wire_d95_52),.data_out(wire_d95_53),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9609554(.data_in(wire_d95_53),.data_out(wire_d95_54),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9609555(.data_in(wire_d95_54),.data_out(wire_d95_55),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9609556(.data_in(wire_d95_55),.data_out(wire_d95_56),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9609557(.data_in(wire_d95_56),.data_out(wire_d95_57),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9609558(.data_in(wire_d95_57),.data_out(wire_d95_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9609559(.data_in(wire_d95_58),.data_out(wire_d95_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9609560(.data_in(wire_d95_59),.data_out(wire_d95_60),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9609561(.data_in(wire_d95_60),.data_out(wire_d95_61),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9609562(.data_in(wire_d95_61),.data_out(wire_d95_62),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9609563(.data_in(wire_d95_62),.data_out(wire_d95_63),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9609564(.data_in(wire_d95_63),.data_out(wire_d95_64),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9609565(.data_in(wire_d95_64),.data_out(wire_d95_65),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9609566(.data_in(wire_d95_65),.data_out(wire_d95_66),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9609567(.data_in(wire_d95_66),.data_out(wire_d95_67),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9609568(.data_in(wire_d95_67),.data_out(wire_d95_68),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9609569(.data_in(wire_d95_68),.data_out(wire_d95_69),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9609570(.data_in(wire_d95_69),.data_out(wire_d95_70),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9609571(.data_in(wire_d95_70),.data_out(wire_d95_71),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9609572(.data_in(wire_d95_71),.data_out(wire_d95_72),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9609573(.data_in(wire_d95_72),.data_out(wire_d95_73),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9609574(.data_in(wire_d95_73),.data_out(wire_d95_74),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9609575(.data_in(wire_d95_74),.data_out(wire_d95_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9609576(.data_in(wire_d95_75),.data_out(wire_d95_76),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9609577(.data_in(wire_d95_76),.data_out(wire_d95_77),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9609578(.data_in(wire_d95_77),.data_out(wire_d95_78),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9609579(.data_in(wire_d95_78),.data_out(wire_d95_79),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9609580(.data_in(wire_d95_79),.data_out(wire_d95_80),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9609581(.data_in(wire_d95_80),.data_out(wire_d95_81),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9609582(.data_in(wire_d95_81),.data_out(wire_d95_82),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9609583(.data_in(wire_d95_82),.data_out(wire_d95_83),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9609584(.data_in(wire_d95_83),.data_out(wire_d95_84),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9609585(.data_in(wire_d95_84),.data_out(wire_d95_85),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9609586(.data_in(wire_d95_85),.data_out(wire_d95_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9609587(.data_in(wire_d95_86),.data_out(wire_d95_87),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9609588(.data_in(wire_d95_87),.data_out(wire_d95_88),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9609589(.data_in(wire_d95_88),.data_out(wire_d95_89),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9609590(.data_in(wire_d95_89),.data_out(wire_d95_90),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9609591(.data_in(wire_d95_90),.data_out(wire_d95_91),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9609592(.data_in(wire_d95_91),.data_out(wire_d95_92),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9609593(.data_in(wire_d95_92),.data_out(wire_d95_93),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9609594(.data_in(wire_d95_93),.data_out(wire_d95_94),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9609595(.data_in(wire_d95_94),.data_out(wire_d95_95),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9609596(.data_in(wire_d95_95),.data_out(wire_d95_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9609597(.data_in(wire_d95_96),.data_out(wire_d95_97),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9609598(.data_in(wire_d95_97),.data_out(wire_d95_98),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9609599(.data_in(wire_d95_98),.data_out(wire_d95_99),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance96095100(.data_in(wire_d95_99),.data_out(wire_d95_100),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance96095101(.data_in(wire_d95_100),.data_out(wire_d95_101),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance96095102(.data_in(wire_d95_101),.data_out(wire_d95_102),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance96095103(.data_in(wire_d95_102),.data_out(wire_d95_103),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance96095104(.data_in(wire_d95_103),.data_out(wire_d95_104),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance96095105(.data_in(wire_d95_104),.data_out(wire_d95_105),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance96095106(.data_in(wire_d95_105),.data_out(wire_d95_106),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance96095107(.data_in(wire_d95_106),.data_out(wire_d95_107),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance96095108(.data_in(wire_d95_107),.data_out(wire_d95_108),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance96095109(.data_in(wire_d95_108),.data_out(wire_d95_109),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance96095110(.data_in(wire_d95_109),.data_out(wire_d95_110),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance96095111(.data_in(wire_d95_110),.data_out(wire_d95_111),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance96095112(.data_in(wire_d95_111),.data_out(wire_d95_112),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance96095113(.data_in(wire_d95_112),.data_out(wire_d95_113),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance96095114(.data_in(wire_d95_113),.data_out(wire_d95_114),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance96095115(.data_in(wire_d95_114),.data_out(wire_d95_115),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance96095116(.data_in(wire_d95_115),.data_out(wire_d95_116),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance96095117(.data_in(wire_d95_116),.data_out(wire_d95_117),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance96095118(.data_in(wire_d95_117),.data_out(wire_d95_118),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance96095119(.data_in(wire_d95_118),.data_out(d_out95),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance970960(.data_in(d_in96),.data_out(wire_d96_0),.clk(clk),.rst(rst));            //channel 97
	invertion #(.WIDTH(WIDTH)) invertion_instance970961(.data_in(wire_d96_0),.data_out(wire_d96_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance970962(.data_in(wire_d96_1),.data_out(wire_d96_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance970963(.data_in(wire_d96_2),.data_out(wire_d96_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance970964(.data_in(wire_d96_3),.data_out(wire_d96_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance970965(.data_in(wire_d96_4),.data_out(wire_d96_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance970966(.data_in(wire_d96_5),.data_out(wire_d96_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance970967(.data_in(wire_d96_6),.data_out(wire_d96_7),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance970968(.data_in(wire_d96_7),.data_out(wire_d96_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance970969(.data_in(wire_d96_8),.data_out(wire_d96_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9709610(.data_in(wire_d96_9),.data_out(wire_d96_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9709611(.data_in(wire_d96_10),.data_out(wire_d96_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9709612(.data_in(wire_d96_11),.data_out(wire_d96_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9709613(.data_in(wire_d96_12),.data_out(wire_d96_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9709614(.data_in(wire_d96_13),.data_out(wire_d96_14),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9709615(.data_in(wire_d96_14),.data_out(wire_d96_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9709616(.data_in(wire_d96_15),.data_out(wire_d96_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9709617(.data_in(wire_d96_16),.data_out(wire_d96_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9709618(.data_in(wire_d96_17),.data_out(wire_d96_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9709619(.data_in(wire_d96_18),.data_out(wire_d96_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9709620(.data_in(wire_d96_19),.data_out(wire_d96_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9709621(.data_in(wire_d96_20),.data_out(wire_d96_21),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9709622(.data_in(wire_d96_21),.data_out(wire_d96_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9709623(.data_in(wire_d96_22),.data_out(wire_d96_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9709624(.data_in(wire_d96_23),.data_out(wire_d96_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9709625(.data_in(wire_d96_24),.data_out(wire_d96_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9709626(.data_in(wire_d96_25),.data_out(wire_d96_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9709627(.data_in(wire_d96_26),.data_out(wire_d96_27),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9709628(.data_in(wire_d96_27),.data_out(wire_d96_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9709629(.data_in(wire_d96_28),.data_out(wire_d96_29),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9709630(.data_in(wire_d96_29),.data_out(wire_d96_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9709631(.data_in(wire_d96_30),.data_out(wire_d96_31),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9709632(.data_in(wire_d96_31),.data_out(wire_d96_32),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9709633(.data_in(wire_d96_32),.data_out(wire_d96_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9709634(.data_in(wire_d96_33),.data_out(wire_d96_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9709635(.data_in(wire_d96_34),.data_out(wire_d96_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9709636(.data_in(wire_d96_35),.data_out(wire_d96_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9709637(.data_in(wire_d96_36),.data_out(wire_d96_37),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9709638(.data_in(wire_d96_37),.data_out(wire_d96_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9709639(.data_in(wire_d96_38),.data_out(wire_d96_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9709640(.data_in(wire_d96_39),.data_out(wire_d96_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9709641(.data_in(wire_d96_40),.data_out(wire_d96_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9709642(.data_in(wire_d96_41),.data_out(wire_d96_42),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9709643(.data_in(wire_d96_42),.data_out(wire_d96_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9709644(.data_in(wire_d96_43),.data_out(wire_d96_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9709645(.data_in(wire_d96_44),.data_out(wire_d96_45),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9709646(.data_in(wire_d96_45),.data_out(wire_d96_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9709647(.data_in(wire_d96_46),.data_out(wire_d96_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9709648(.data_in(wire_d96_47),.data_out(wire_d96_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9709649(.data_in(wire_d96_48),.data_out(wire_d96_49),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9709650(.data_in(wire_d96_49),.data_out(wire_d96_50),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9709651(.data_in(wire_d96_50),.data_out(wire_d96_51),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9709652(.data_in(wire_d96_51),.data_out(wire_d96_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9709653(.data_in(wire_d96_52),.data_out(wire_d96_53),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9709654(.data_in(wire_d96_53),.data_out(wire_d96_54),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9709655(.data_in(wire_d96_54),.data_out(wire_d96_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9709656(.data_in(wire_d96_55),.data_out(wire_d96_56),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9709657(.data_in(wire_d96_56),.data_out(wire_d96_57),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9709658(.data_in(wire_d96_57),.data_out(wire_d96_58),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9709659(.data_in(wire_d96_58),.data_out(wire_d96_59),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9709660(.data_in(wire_d96_59),.data_out(wire_d96_60),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9709661(.data_in(wire_d96_60),.data_out(wire_d96_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9709662(.data_in(wire_d96_61),.data_out(wire_d96_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9709663(.data_in(wire_d96_62),.data_out(wire_d96_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9709664(.data_in(wire_d96_63),.data_out(wire_d96_64),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9709665(.data_in(wire_d96_64),.data_out(wire_d96_65),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9709666(.data_in(wire_d96_65),.data_out(wire_d96_66),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9709667(.data_in(wire_d96_66),.data_out(wire_d96_67),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9709668(.data_in(wire_d96_67),.data_out(wire_d96_68),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9709669(.data_in(wire_d96_68),.data_out(wire_d96_69),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9709670(.data_in(wire_d96_69),.data_out(wire_d96_70),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9709671(.data_in(wire_d96_70),.data_out(wire_d96_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9709672(.data_in(wire_d96_71),.data_out(wire_d96_72),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9709673(.data_in(wire_d96_72),.data_out(wire_d96_73),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9709674(.data_in(wire_d96_73),.data_out(wire_d96_74),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9709675(.data_in(wire_d96_74),.data_out(wire_d96_75),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9709676(.data_in(wire_d96_75),.data_out(wire_d96_76),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9709677(.data_in(wire_d96_76),.data_out(wire_d96_77),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9709678(.data_in(wire_d96_77),.data_out(wire_d96_78),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9709679(.data_in(wire_d96_78),.data_out(wire_d96_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9709680(.data_in(wire_d96_79),.data_out(wire_d96_80),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9709681(.data_in(wire_d96_80),.data_out(wire_d96_81),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9709682(.data_in(wire_d96_81),.data_out(wire_d96_82),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9709683(.data_in(wire_d96_82),.data_out(wire_d96_83),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9709684(.data_in(wire_d96_83),.data_out(wire_d96_84),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9709685(.data_in(wire_d96_84),.data_out(wire_d96_85),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9709686(.data_in(wire_d96_85),.data_out(wire_d96_86),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9709687(.data_in(wire_d96_86),.data_out(wire_d96_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9709688(.data_in(wire_d96_87),.data_out(wire_d96_88),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9709689(.data_in(wire_d96_88),.data_out(wire_d96_89),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9709690(.data_in(wire_d96_89),.data_out(wire_d96_90),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9709691(.data_in(wire_d96_90),.data_out(wire_d96_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9709692(.data_in(wire_d96_91),.data_out(wire_d96_92),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9709693(.data_in(wire_d96_92),.data_out(wire_d96_93),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9709694(.data_in(wire_d96_93),.data_out(wire_d96_94),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9709695(.data_in(wire_d96_94),.data_out(wire_d96_95),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9709696(.data_in(wire_d96_95),.data_out(wire_d96_96),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9709697(.data_in(wire_d96_96),.data_out(wire_d96_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9709698(.data_in(wire_d96_97),.data_out(wire_d96_98),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9709699(.data_in(wire_d96_98),.data_out(wire_d96_99),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance97096100(.data_in(wire_d96_99),.data_out(wire_d96_100),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance97096101(.data_in(wire_d96_100),.data_out(wire_d96_101),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance97096102(.data_in(wire_d96_101),.data_out(wire_d96_102),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance97096103(.data_in(wire_d96_102),.data_out(wire_d96_103),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance97096104(.data_in(wire_d96_103),.data_out(wire_d96_104),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance97096105(.data_in(wire_d96_104),.data_out(wire_d96_105),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance97096106(.data_in(wire_d96_105),.data_out(wire_d96_106),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance97096107(.data_in(wire_d96_106),.data_out(wire_d96_107),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance97096108(.data_in(wire_d96_107),.data_out(wire_d96_108),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance97096109(.data_in(wire_d96_108),.data_out(wire_d96_109),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance97096110(.data_in(wire_d96_109),.data_out(wire_d96_110),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance97096111(.data_in(wire_d96_110),.data_out(wire_d96_111),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance97096112(.data_in(wire_d96_111),.data_out(wire_d96_112),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance97096113(.data_in(wire_d96_112),.data_out(wire_d96_113),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance97096114(.data_in(wire_d96_113),.data_out(wire_d96_114),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance97096115(.data_in(wire_d96_114),.data_out(wire_d96_115),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance97096116(.data_in(wire_d96_115),.data_out(wire_d96_116),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance97096117(.data_in(wire_d96_116),.data_out(wire_d96_117),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance97096118(.data_in(wire_d96_117),.data_out(wire_d96_118),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance97096119(.data_in(wire_d96_118),.data_out(d_out96),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance980970(.data_in(d_in97),.data_out(wire_d97_0),.clk(clk),.rst(rst));            //channel 98
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance980971(.data_in(wire_d97_0),.data_out(wire_d97_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance980972(.data_in(wire_d97_1),.data_out(wire_d97_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance980973(.data_in(wire_d97_2),.data_out(wire_d97_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance980974(.data_in(wire_d97_3),.data_out(wire_d97_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance980975(.data_in(wire_d97_4),.data_out(wire_d97_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance980976(.data_in(wire_d97_5),.data_out(wire_d97_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance980977(.data_in(wire_d97_6),.data_out(wire_d97_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance980978(.data_in(wire_d97_7),.data_out(wire_d97_8),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance980979(.data_in(wire_d97_8),.data_out(wire_d97_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9809710(.data_in(wire_d97_9),.data_out(wire_d97_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9809711(.data_in(wire_d97_10),.data_out(wire_d97_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9809712(.data_in(wire_d97_11),.data_out(wire_d97_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9809713(.data_in(wire_d97_12),.data_out(wire_d97_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9809714(.data_in(wire_d97_13),.data_out(wire_d97_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9809715(.data_in(wire_d97_14),.data_out(wire_d97_15),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9809716(.data_in(wire_d97_15),.data_out(wire_d97_16),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9809717(.data_in(wire_d97_16),.data_out(wire_d97_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9809718(.data_in(wire_d97_17),.data_out(wire_d97_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9809719(.data_in(wire_d97_18),.data_out(wire_d97_19),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9809720(.data_in(wire_d97_19),.data_out(wire_d97_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9809721(.data_in(wire_d97_20),.data_out(wire_d97_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9809722(.data_in(wire_d97_21),.data_out(wire_d97_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9809723(.data_in(wire_d97_22),.data_out(wire_d97_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9809724(.data_in(wire_d97_23),.data_out(wire_d97_24),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9809725(.data_in(wire_d97_24),.data_out(wire_d97_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9809726(.data_in(wire_d97_25),.data_out(wire_d97_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9809727(.data_in(wire_d97_26),.data_out(wire_d97_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9809728(.data_in(wire_d97_27),.data_out(wire_d97_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9809729(.data_in(wire_d97_28),.data_out(wire_d97_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9809730(.data_in(wire_d97_29),.data_out(wire_d97_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9809731(.data_in(wire_d97_30),.data_out(wire_d97_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9809732(.data_in(wire_d97_31),.data_out(wire_d97_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9809733(.data_in(wire_d97_32),.data_out(wire_d97_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9809734(.data_in(wire_d97_33),.data_out(wire_d97_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9809735(.data_in(wire_d97_34),.data_out(wire_d97_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9809736(.data_in(wire_d97_35),.data_out(wire_d97_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9809737(.data_in(wire_d97_36),.data_out(wire_d97_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9809738(.data_in(wire_d97_37),.data_out(wire_d97_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9809739(.data_in(wire_d97_38),.data_out(wire_d97_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9809740(.data_in(wire_d97_39),.data_out(wire_d97_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9809741(.data_in(wire_d97_40),.data_out(wire_d97_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9809742(.data_in(wire_d97_41),.data_out(wire_d97_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9809743(.data_in(wire_d97_42),.data_out(wire_d97_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9809744(.data_in(wire_d97_43),.data_out(wire_d97_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9809745(.data_in(wire_d97_44),.data_out(wire_d97_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9809746(.data_in(wire_d97_45),.data_out(wire_d97_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9809747(.data_in(wire_d97_46),.data_out(wire_d97_47),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9809748(.data_in(wire_d97_47),.data_out(wire_d97_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9809749(.data_in(wire_d97_48),.data_out(wire_d97_49),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9809750(.data_in(wire_d97_49),.data_out(wire_d97_50),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9809751(.data_in(wire_d97_50),.data_out(wire_d97_51),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9809752(.data_in(wire_d97_51),.data_out(wire_d97_52),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9809753(.data_in(wire_d97_52),.data_out(wire_d97_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9809754(.data_in(wire_d97_53),.data_out(wire_d97_54),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9809755(.data_in(wire_d97_54),.data_out(wire_d97_55),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9809756(.data_in(wire_d97_55),.data_out(wire_d97_56),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9809757(.data_in(wire_d97_56),.data_out(wire_d97_57),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9809758(.data_in(wire_d97_57),.data_out(wire_d97_58),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9809759(.data_in(wire_d97_58),.data_out(wire_d97_59),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9809760(.data_in(wire_d97_59),.data_out(wire_d97_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9809761(.data_in(wire_d97_60),.data_out(wire_d97_61),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9809762(.data_in(wire_d97_61),.data_out(wire_d97_62),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9809763(.data_in(wire_d97_62),.data_out(wire_d97_63),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9809764(.data_in(wire_d97_63),.data_out(wire_d97_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9809765(.data_in(wire_d97_64),.data_out(wire_d97_65),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9809766(.data_in(wire_d97_65),.data_out(wire_d97_66),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9809767(.data_in(wire_d97_66),.data_out(wire_d97_67),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9809768(.data_in(wire_d97_67),.data_out(wire_d97_68),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9809769(.data_in(wire_d97_68),.data_out(wire_d97_69),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9809770(.data_in(wire_d97_69),.data_out(wire_d97_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9809771(.data_in(wire_d97_70),.data_out(wire_d97_71),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9809772(.data_in(wire_d97_71),.data_out(wire_d97_72),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9809773(.data_in(wire_d97_72),.data_out(wire_d97_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9809774(.data_in(wire_d97_73),.data_out(wire_d97_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9809775(.data_in(wire_d97_74),.data_out(wire_d97_75),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9809776(.data_in(wire_d97_75),.data_out(wire_d97_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9809777(.data_in(wire_d97_76),.data_out(wire_d97_77),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9809778(.data_in(wire_d97_77),.data_out(wire_d97_78),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9809779(.data_in(wire_d97_78),.data_out(wire_d97_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9809780(.data_in(wire_d97_79),.data_out(wire_d97_80),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9809781(.data_in(wire_d97_80),.data_out(wire_d97_81),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9809782(.data_in(wire_d97_81),.data_out(wire_d97_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9809783(.data_in(wire_d97_82),.data_out(wire_d97_83),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9809784(.data_in(wire_d97_83),.data_out(wire_d97_84),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9809785(.data_in(wire_d97_84),.data_out(wire_d97_85),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9809786(.data_in(wire_d97_85),.data_out(wire_d97_86),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9809787(.data_in(wire_d97_86),.data_out(wire_d97_87),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9809788(.data_in(wire_d97_87),.data_out(wire_d97_88),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9809789(.data_in(wire_d97_88),.data_out(wire_d97_89),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9809790(.data_in(wire_d97_89),.data_out(wire_d97_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9809791(.data_in(wire_d97_90),.data_out(wire_d97_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9809792(.data_in(wire_d97_91),.data_out(wire_d97_92),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9809793(.data_in(wire_d97_92),.data_out(wire_d97_93),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9809794(.data_in(wire_d97_93),.data_out(wire_d97_94),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9809795(.data_in(wire_d97_94),.data_out(wire_d97_95),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9809796(.data_in(wire_d97_95),.data_out(wire_d97_96),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9809797(.data_in(wire_d97_96),.data_out(wire_d97_97),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9809798(.data_in(wire_d97_97),.data_out(wire_d97_98),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9809799(.data_in(wire_d97_98),.data_out(wire_d97_99),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance98097100(.data_in(wire_d97_99),.data_out(wire_d97_100),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance98097101(.data_in(wire_d97_100),.data_out(wire_d97_101),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance98097102(.data_in(wire_d97_101),.data_out(wire_d97_102),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance98097103(.data_in(wire_d97_102),.data_out(wire_d97_103),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance98097104(.data_in(wire_d97_103),.data_out(wire_d97_104),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance98097105(.data_in(wire_d97_104),.data_out(wire_d97_105),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance98097106(.data_in(wire_d97_105),.data_out(wire_d97_106),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance98097107(.data_in(wire_d97_106),.data_out(wire_d97_107),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance98097108(.data_in(wire_d97_107),.data_out(wire_d97_108),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance98097109(.data_in(wire_d97_108),.data_out(wire_d97_109),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance98097110(.data_in(wire_d97_109),.data_out(wire_d97_110),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance98097111(.data_in(wire_d97_110),.data_out(wire_d97_111),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance98097112(.data_in(wire_d97_111),.data_out(wire_d97_112),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance98097113(.data_in(wire_d97_112),.data_out(wire_d97_113),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance98097114(.data_in(wire_d97_113),.data_out(wire_d97_114),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance98097115(.data_in(wire_d97_114),.data_out(wire_d97_115),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance98097116(.data_in(wire_d97_115),.data_out(wire_d97_116),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance98097117(.data_in(wire_d97_116),.data_out(wire_d97_117),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance98097118(.data_in(wire_d97_117),.data_out(wire_d97_118),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance98097119(.data_in(wire_d97_118),.data_out(d_out97),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance990980(.data_in(d_in98),.data_out(wire_d98_0),.clk(clk),.rst(rst));            //channel 99
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance990981(.data_in(wire_d98_0),.data_out(wire_d98_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance990982(.data_in(wire_d98_1),.data_out(wire_d98_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance990983(.data_in(wire_d98_2),.data_out(wire_d98_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance990984(.data_in(wire_d98_3),.data_out(wire_d98_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance990985(.data_in(wire_d98_4),.data_out(wire_d98_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance990986(.data_in(wire_d98_5),.data_out(wire_d98_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance990987(.data_in(wire_d98_6),.data_out(wire_d98_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance990988(.data_in(wire_d98_7),.data_out(wire_d98_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance990989(.data_in(wire_d98_8),.data_out(wire_d98_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9909810(.data_in(wire_d98_9),.data_out(wire_d98_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9909811(.data_in(wire_d98_10),.data_out(wire_d98_11),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9909812(.data_in(wire_d98_11),.data_out(wire_d98_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9909813(.data_in(wire_d98_12),.data_out(wire_d98_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9909814(.data_in(wire_d98_13),.data_out(wire_d98_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9909815(.data_in(wire_d98_14),.data_out(wire_d98_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9909816(.data_in(wire_d98_15),.data_out(wire_d98_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9909817(.data_in(wire_d98_16),.data_out(wire_d98_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9909818(.data_in(wire_d98_17),.data_out(wire_d98_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9909819(.data_in(wire_d98_18),.data_out(wire_d98_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9909820(.data_in(wire_d98_19),.data_out(wire_d98_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9909821(.data_in(wire_d98_20),.data_out(wire_d98_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9909822(.data_in(wire_d98_21),.data_out(wire_d98_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9909823(.data_in(wire_d98_22),.data_out(wire_d98_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9909824(.data_in(wire_d98_23),.data_out(wire_d98_24),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9909825(.data_in(wire_d98_24),.data_out(wire_d98_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9909826(.data_in(wire_d98_25),.data_out(wire_d98_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9909827(.data_in(wire_d98_26),.data_out(wire_d98_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9909828(.data_in(wire_d98_27),.data_out(wire_d98_28),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9909829(.data_in(wire_d98_28),.data_out(wire_d98_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9909830(.data_in(wire_d98_29),.data_out(wire_d98_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9909831(.data_in(wire_d98_30),.data_out(wire_d98_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9909832(.data_in(wire_d98_31),.data_out(wire_d98_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9909833(.data_in(wire_d98_32),.data_out(wire_d98_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9909834(.data_in(wire_d98_33),.data_out(wire_d98_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9909835(.data_in(wire_d98_34),.data_out(wire_d98_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9909836(.data_in(wire_d98_35),.data_out(wire_d98_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9909837(.data_in(wire_d98_36),.data_out(wire_d98_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9909838(.data_in(wire_d98_37),.data_out(wire_d98_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9909839(.data_in(wire_d98_38),.data_out(wire_d98_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9909840(.data_in(wire_d98_39),.data_out(wire_d98_40),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9909841(.data_in(wire_d98_40),.data_out(wire_d98_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9909842(.data_in(wire_d98_41),.data_out(wire_d98_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9909843(.data_in(wire_d98_42),.data_out(wire_d98_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9909844(.data_in(wire_d98_43),.data_out(wire_d98_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9909845(.data_in(wire_d98_44),.data_out(wire_d98_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9909846(.data_in(wire_d98_45),.data_out(wire_d98_46),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9909847(.data_in(wire_d98_46),.data_out(wire_d98_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9909848(.data_in(wire_d98_47),.data_out(wire_d98_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9909849(.data_in(wire_d98_48),.data_out(wire_d98_49),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9909850(.data_in(wire_d98_49),.data_out(wire_d98_50),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9909851(.data_in(wire_d98_50),.data_out(wire_d98_51),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9909852(.data_in(wire_d98_51),.data_out(wire_d98_52),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9909853(.data_in(wire_d98_52),.data_out(wire_d98_53),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9909854(.data_in(wire_d98_53),.data_out(wire_d98_54),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9909855(.data_in(wire_d98_54),.data_out(wire_d98_55),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9909856(.data_in(wire_d98_55),.data_out(wire_d98_56),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9909857(.data_in(wire_d98_56),.data_out(wire_d98_57),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9909858(.data_in(wire_d98_57),.data_out(wire_d98_58),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9909859(.data_in(wire_d98_58),.data_out(wire_d98_59),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9909860(.data_in(wire_d98_59),.data_out(wire_d98_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9909861(.data_in(wire_d98_60),.data_out(wire_d98_61),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9909862(.data_in(wire_d98_61),.data_out(wire_d98_62),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9909863(.data_in(wire_d98_62),.data_out(wire_d98_63),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9909864(.data_in(wire_d98_63),.data_out(wire_d98_64),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9909865(.data_in(wire_d98_64),.data_out(wire_d98_65),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9909866(.data_in(wire_d98_65),.data_out(wire_d98_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9909867(.data_in(wire_d98_66),.data_out(wire_d98_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9909868(.data_in(wire_d98_67),.data_out(wire_d98_68),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9909869(.data_in(wire_d98_68),.data_out(wire_d98_69),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9909870(.data_in(wire_d98_69),.data_out(wire_d98_70),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9909871(.data_in(wire_d98_70),.data_out(wire_d98_71),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9909872(.data_in(wire_d98_71),.data_out(wire_d98_72),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9909873(.data_in(wire_d98_72),.data_out(wire_d98_73),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9909874(.data_in(wire_d98_73),.data_out(wire_d98_74),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9909875(.data_in(wire_d98_74),.data_out(wire_d98_75),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9909876(.data_in(wire_d98_75),.data_out(wire_d98_76),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9909877(.data_in(wire_d98_76),.data_out(wire_d98_77),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9909878(.data_in(wire_d98_77),.data_out(wire_d98_78),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9909879(.data_in(wire_d98_78),.data_out(wire_d98_79),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9909880(.data_in(wire_d98_79),.data_out(wire_d98_80),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9909881(.data_in(wire_d98_80),.data_out(wire_d98_81),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9909882(.data_in(wire_d98_81),.data_out(wire_d98_82),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9909883(.data_in(wire_d98_82),.data_out(wire_d98_83),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9909884(.data_in(wire_d98_83),.data_out(wire_d98_84),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9909885(.data_in(wire_d98_84),.data_out(wire_d98_85),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9909886(.data_in(wire_d98_85),.data_out(wire_d98_86),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9909887(.data_in(wire_d98_86),.data_out(wire_d98_87),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9909888(.data_in(wire_d98_87),.data_out(wire_d98_88),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9909889(.data_in(wire_d98_88),.data_out(wire_d98_89),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9909890(.data_in(wire_d98_89),.data_out(wire_d98_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9909891(.data_in(wire_d98_90),.data_out(wire_d98_91),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9909892(.data_in(wire_d98_91),.data_out(wire_d98_92),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9909893(.data_in(wire_d98_92),.data_out(wire_d98_93),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9909894(.data_in(wire_d98_93),.data_out(wire_d98_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9909895(.data_in(wire_d98_94),.data_out(wire_d98_95),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9909896(.data_in(wire_d98_95),.data_out(wire_d98_96),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9909897(.data_in(wire_d98_96),.data_out(wire_d98_97),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9909898(.data_in(wire_d98_97),.data_out(wire_d98_98),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9909899(.data_in(wire_d98_98),.data_out(wire_d98_99),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance99098100(.data_in(wire_d98_99),.data_out(wire_d98_100),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance99098101(.data_in(wire_d98_100),.data_out(wire_d98_101),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance99098102(.data_in(wire_d98_101),.data_out(wire_d98_102),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance99098103(.data_in(wire_d98_102),.data_out(wire_d98_103),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance99098104(.data_in(wire_d98_103),.data_out(wire_d98_104),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance99098105(.data_in(wire_d98_104),.data_out(wire_d98_105),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance99098106(.data_in(wire_d98_105),.data_out(wire_d98_106),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance99098107(.data_in(wire_d98_106),.data_out(wire_d98_107),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance99098108(.data_in(wire_d98_107),.data_out(wire_d98_108),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance99098109(.data_in(wire_d98_108),.data_out(wire_d98_109),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance99098110(.data_in(wire_d98_109),.data_out(wire_d98_110),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance99098111(.data_in(wire_d98_110),.data_out(wire_d98_111),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance99098112(.data_in(wire_d98_111),.data_out(wire_d98_112),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance99098113(.data_in(wire_d98_112),.data_out(wire_d98_113),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance99098114(.data_in(wire_d98_113),.data_out(wire_d98_114),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance99098115(.data_in(wire_d98_114),.data_out(wire_d98_115),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance99098116(.data_in(wire_d98_115),.data_out(wire_d98_116),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance99098117(.data_in(wire_d98_116),.data_out(wire_d98_117),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance99098118(.data_in(wire_d98_117),.data_out(wire_d98_118),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance99098119(.data_in(wire_d98_118),.data_out(d_out98),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance1000990(.data_in(d_in99),.data_out(wire_d99_0),.clk(clk),.rst(rst));            //channel 100
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1000991(.data_in(wire_d99_0),.data_out(wire_d99_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1000992(.data_in(wire_d99_1),.data_out(wire_d99_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1000993(.data_in(wire_d99_2),.data_out(wire_d99_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1000994(.data_in(wire_d99_3),.data_out(wire_d99_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1000995(.data_in(wire_d99_4),.data_out(wire_d99_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1000996(.data_in(wire_d99_5),.data_out(wire_d99_6),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1000997(.data_in(wire_d99_6),.data_out(wire_d99_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1000998(.data_in(wire_d99_7),.data_out(wire_d99_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1000999(.data_in(wire_d99_8),.data_out(wire_d99_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10009910(.data_in(wire_d99_9),.data_out(wire_d99_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10009911(.data_in(wire_d99_10),.data_out(wire_d99_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance10009912(.data_in(wire_d99_11),.data_out(wire_d99_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance10009913(.data_in(wire_d99_12),.data_out(wire_d99_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10009914(.data_in(wire_d99_13),.data_out(wire_d99_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance10009915(.data_in(wire_d99_14),.data_out(wire_d99_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10009916(.data_in(wire_d99_15),.data_out(wire_d99_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance10009917(.data_in(wire_d99_16),.data_out(wire_d99_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10009918(.data_in(wire_d99_17),.data_out(wire_d99_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance10009919(.data_in(wire_d99_18),.data_out(wire_d99_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance10009920(.data_in(wire_d99_19),.data_out(wire_d99_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10009921(.data_in(wire_d99_20),.data_out(wire_d99_21),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance10009922(.data_in(wire_d99_21),.data_out(wire_d99_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance10009923(.data_in(wire_d99_22),.data_out(wire_d99_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10009924(.data_in(wire_d99_23),.data_out(wire_d99_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance10009925(.data_in(wire_d99_24),.data_out(wire_d99_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10009926(.data_in(wire_d99_25),.data_out(wire_d99_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance10009927(.data_in(wire_d99_26),.data_out(wire_d99_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10009928(.data_in(wire_d99_27),.data_out(wire_d99_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance10009929(.data_in(wire_d99_28),.data_out(wire_d99_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10009930(.data_in(wire_d99_29),.data_out(wire_d99_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10009931(.data_in(wire_d99_30),.data_out(wire_d99_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10009932(.data_in(wire_d99_31),.data_out(wire_d99_32),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance10009933(.data_in(wire_d99_32),.data_out(wire_d99_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10009934(.data_in(wire_d99_33),.data_out(wire_d99_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10009935(.data_in(wire_d99_34),.data_out(wire_d99_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10009936(.data_in(wire_d99_35),.data_out(wire_d99_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10009937(.data_in(wire_d99_36),.data_out(wire_d99_37),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance10009938(.data_in(wire_d99_37),.data_out(wire_d99_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance10009939(.data_in(wire_d99_38),.data_out(wire_d99_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10009940(.data_in(wire_d99_39),.data_out(wire_d99_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance10009941(.data_in(wire_d99_40),.data_out(wire_d99_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance10009942(.data_in(wire_d99_41),.data_out(wire_d99_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10009943(.data_in(wire_d99_42),.data_out(wire_d99_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10009944(.data_in(wire_d99_43),.data_out(wire_d99_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10009945(.data_in(wire_d99_44),.data_out(wire_d99_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance10009946(.data_in(wire_d99_45),.data_out(wire_d99_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10009947(.data_in(wire_d99_46),.data_out(wire_d99_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance10009948(.data_in(wire_d99_47),.data_out(wire_d99_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance10009949(.data_in(wire_d99_48),.data_out(wire_d99_49),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance10009950(.data_in(wire_d99_49),.data_out(wire_d99_50),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10009951(.data_in(wire_d99_50),.data_out(wire_d99_51),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance10009952(.data_in(wire_d99_51),.data_out(wire_d99_52),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10009953(.data_in(wire_d99_52),.data_out(wire_d99_53),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10009954(.data_in(wire_d99_53),.data_out(wire_d99_54),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10009955(.data_in(wire_d99_54),.data_out(wire_d99_55),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance10009956(.data_in(wire_d99_55),.data_out(wire_d99_56),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance10009957(.data_in(wire_d99_56),.data_out(wire_d99_57),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10009958(.data_in(wire_d99_57),.data_out(wire_d99_58),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance10009959(.data_in(wire_d99_58),.data_out(wire_d99_59),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance10009960(.data_in(wire_d99_59),.data_out(wire_d99_60),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance10009961(.data_in(wire_d99_60),.data_out(wire_d99_61),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance10009962(.data_in(wire_d99_61),.data_out(wire_d99_62),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance10009963(.data_in(wire_d99_62),.data_out(wire_d99_63),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance10009964(.data_in(wire_d99_63),.data_out(wire_d99_64),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance10009965(.data_in(wire_d99_64),.data_out(wire_d99_65),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10009966(.data_in(wire_d99_65),.data_out(wire_d99_66),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance10009967(.data_in(wire_d99_66),.data_out(wire_d99_67),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance10009968(.data_in(wire_d99_67),.data_out(wire_d99_68),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10009969(.data_in(wire_d99_68),.data_out(wire_d99_69),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance10009970(.data_in(wire_d99_69),.data_out(wire_d99_70),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10009971(.data_in(wire_d99_70),.data_out(wire_d99_71),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance10009972(.data_in(wire_d99_71),.data_out(wire_d99_72),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10009973(.data_in(wire_d99_72),.data_out(wire_d99_73),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance10009974(.data_in(wire_d99_73),.data_out(wire_d99_74),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance10009975(.data_in(wire_d99_74),.data_out(wire_d99_75),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance10009976(.data_in(wire_d99_75),.data_out(wire_d99_76),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance10009977(.data_in(wire_d99_76),.data_out(wire_d99_77),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance10009978(.data_in(wire_d99_77),.data_out(wire_d99_78),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance10009979(.data_in(wire_d99_78),.data_out(wire_d99_79),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10009980(.data_in(wire_d99_79),.data_out(wire_d99_80),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance10009981(.data_in(wire_d99_80),.data_out(wire_d99_81),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10009982(.data_in(wire_d99_81),.data_out(wire_d99_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10009983(.data_in(wire_d99_82),.data_out(wire_d99_83),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance10009984(.data_in(wire_d99_83),.data_out(wire_d99_84),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10009985(.data_in(wire_d99_84),.data_out(wire_d99_85),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance10009986(.data_in(wire_d99_85),.data_out(wire_d99_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10009987(.data_in(wire_d99_86),.data_out(wire_d99_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10009988(.data_in(wire_d99_87),.data_out(wire_d99_88),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10009989(.data_in(wire_d99_88),.data_out(wire_d99_89),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10009990(.data_in(wire_d99_89),.data_out(wire_d99_90),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10009991(.data_in(wire_d99_90),.data_out(wire_d99_91),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10009992(.data_in(wire_d99_91),.data_out(wire_d99_92),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance10009993(.data_in(wire_d99_92),.data_out(wire_d99_93),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance10009994(.data_in(wire_d99_93),.data_out(wire_d99_94),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10009995(.data_in(wire_d99_94),.data_out(wire_d99_95),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance10009996(.data_in(wire_d99_95),.data_out(wire_d99_96),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance10009997(.data_in(wire_d99_96),.data_out(wire_d99_97),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10009998(.data_in(wire_d99_97),.data_out(wire_d99_98),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance10009999(.data_in(wire_d99_98),.data_out(wire_d99_99),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100099100(.data_in(wire_d99_99),.data_out(wire_d99_100),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100099101(.data_in(wire_d99_100),.data_out(wire_d99_101),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100099102(.data_in(wire_d99_101),.data_out(wire_d99_102),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100099103(.data_in(wire_d99_102),.data_out(wire_d99_103),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100099104(.data_in(wire_d99_103),.data_out(wire_d99_104),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100099105(.data_in(wire_d99_104),.data_out(wire_d99_105),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100099106(.data_in(wire_d99_105),.data_out(wire_d99_106),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100099107(.data_in(wire_d99_106),.data_out(wire_d99_107),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance100099108(.data_in(wire_d99_107),.data_out(wire_d99_108),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance100099109(.data_in(wire_d99_108),.data_out(wire_d99_109),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100099110(.data_in(wire_d99_109),.data_out(wire_d99_110),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100099111(.data_in(wire_d99_110),.data_out(wire_d99_111),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100099112(.data_in(wire_d99_111),.data_out(wire_d99_112),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100099113(.data_in(wire_d99_112),.data_out(wire_d99_113),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100099114(.data_in(wire_d99_113),.data_out(wire_d99_114),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100099115(.data_in(wire_d99_114),.data_out(wire_d99_115),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance100099116(.data_in(wire_d99_115),.data_out(wire_d99_116),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100099117(.data_in(wire_d99_116),.data_out(wire_d99_117),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100099118(.data_in(wire_d99_117),.data_out(wire_d99_118),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100099119(.data_in(wire_d99_118),.data_out(d_out99),.clk(clk),.rst(rst));


endmodule