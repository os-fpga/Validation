// `include "encoder.v"

module design48_10_100_top #(parameter WIDTH=32,CHANNEL=10) (clk, rst, in, out);

	localparam OUT_BUS=CHANNEL*WIDTH;
	input clk,rst;
	input [WIDTH-1:0] in;
	output [WIDTH-1:0] out;

	reg [WIDTH-1:0] d_in0;
	reg [WIDTH-1:0] d_in1;
	reg [WIDTH-1:0] d_in2;
	reg [WIDTH-1:0] d_in3;
	reg [WIDTH-1:0] d_in4;
	reg [WIDTH-1:0] d_in5;
	reg [WIDTH-1:0] d_in6;
	reg [WIDTH-1:0] d_in7;
	reg [WIDTH-1:0] d_in8;
	reg [WIDTH-1:0] d_in9;
	wire [WIDTH-1:0] d_out0;
	wire [WIDTH-1:0] d_out1;
	wire [WIDTH-1:0] d_out2;
	wire [WIDTH-1:0] d_out3;
	wire [WIDTH-1:0] d_out4;
	wire [WIDTH-1:0] d_out5;
	wire [WIDTH-1:0] d_out6;
	wire [WIDTH-1:0] d_out7;
	wire [WIDTH-1:0] d_out8;
	wire [WIDTH-1:0] d_out9;

	reg [OUT_BUS-1:0] tmp;

	always @ (posedge clk or posedge rst) begin
		if (rst)
			tmp <= 0;
		else
			tmp <= {tmp[OUT_BUS-(WIDTH-1):0],in};
	end

	always @ (posedge clk) begin
		d_in0 <= tmp[WIDTH-1:0];
		d_in1 <= tmp[(WIDTH*2)-1:WIDTH*1];
		d_in2 <= tmp[(WIDTH*3)-1:WIDTH*2];
		d_in3 <= tmp[(WIDTH*4)-1:WIDTH*3];
		d_in4 <= tmp[(WIDTH*5)-1:WIDTH*4];
		d_in5 <= tmp[(WIDTH*6)-1:WIDTH*5];
		d_in6 <= tmp[(WIDTH*7)-1:WIDTH*6];
		d_in7 <= tmp[(WIDTH*8)-1:WIDTH*7];
		d_in8 <= tmp[(WIDTH*9)-1:WIDTH*8];
		d_in9 <= tmp[(WIDTH*10)-1:WIDTH*9];
	end

	design48_10_100 #(.WIDTH(WIDTH)) design48_10_100_inst(.d_in0(d_in0),.d_in1(d_in1),.d_in2(d_in2),.d_in3(d_in3),.d_in4(d_in4),.d_in5(d_in5),.d_in6(d_in6),.d_in7(d_in7),.d_in8(d_in8),.d_in9(d_in9),.d_out0(d_out0),.d_out1(d_out1),.d_out2(d_out2),.d_out3(d_out3),.d_out4(d_out4),.d_out5(d_out5),.d_out6(d_out6),.d_out7(d_out7),.d_out8(d_out8),.d_out9(d_out9),.clk(clk),.rst(rst));

	assign out = d_out0^d_out1^d_out2^d_out3^d_out4^d_out5^d_out6^d_out7^d_out8^d_out9;

endmodule

module design48_10_100 #(parameter WIDTH=32) (d_in0, d_in1, d_in2, d_in3, d_in4, d_in5, d_in6, d_in7, d_in8, d_in9, d_out0, d_out1, d_out2, d_out3, d_out4, d_out5, d_out6, d_out7, d_out8, d_out9, clk, rst);
	input clk;
	input rst;
	input [WIDTH-1:0] d_in0; 
	input [WIDTH-1:0] d_in1; 
	input [WIDTH-1:0] d_in2; 
	input [WIDTH-1:0] d_in3; 
	input [WIDTH-1:0] d_in4; 
	input [WIDTH-1:0] d_in5; 
	input [WIDTH-1:0] d_in6; 
	input [WIDTH-1:0] d_in7; 
	input [WIDTH-1:0] d_in8; 
	input [WIDTH-1:0] d_in9; 
	output [WIDTH-1:0] d_out0; 
	output [WIDTH-1:0] d_out1; 
	output [WIDTH-1:0] d_out2; 
	output [WIDTH-1:0] d_out3; 
	output [WIDTH-1:0] d_out4; 
	output [WIDTH-1:0] d_out5; 
	output [WIDTH-1:0] d_out6; 
	output [WIDTH-1:0] d_out7; 
	output [WIDTH-1:0] d_out8; 
	output [WIDTH-1:0] d_out9; 

	wire [WIDTH-1:0] wire_d0_0;
	wire [WIDTH-1:0] wire_d0_1;
	wire [WIDTH-1:0] wire_d0_2;
	wire [WIDTH-1:0] wire_d0_3;
	wire [WIDTH-1:0] wire_d0_4;
	wire [WIDTH-1:0] wire_d0_5;
	wire [WIDTH-1:0] wire_d0_6;
	wire [WIDTH-1:0] wire_d0_7;
	wire [WIDTH-1:0] wire_d0_8;
	wire [WIDTH-1:0] wire_d0_9;
	wire [WIDTH-1:0] wire_d0_10;
	wire [WIDTH-1:0] wire_d0_11;
	wire [WIDTH-1:0] wire_d0_12;
	wire [WIDTH-1:0] wire_d0_13;
	wire [WIDTH-1:0] wire_d0_14;
	wire [WIDTH-1:0] wire_d0_15;
	wire [WIDTH-1:0] wire_d0_16;
	wire [WIDTH-1:0] wire_d0_17;
	wire [WIDTH-1:0] wire_d0_18;
	wire [WIDTH-1:0] wire_d0_19;
	wire [WIDTH-1:0] wire_d0_20;
	wire [WIDTH-1:0] wire_d0_21;
	wire [WIDTH-1:0] wire_d0_22;
	wire [WIDTH-1:0] wire_d0_23;
	wire [WIDTH-1:0] wire_d0_24;
	wire [WIDTH-1:0] wire_d0_25;
	wire [WIDTH-1:0] wire_d0_26;
	wire [WIDTH-1:0] wire_d0_27;
	wire [WIDTH-1:0] wire_d0_28;
	wire [WIDTH-1:0] wire_d0_29;
	wire [WIDTH-1:0] wire_d0_30;
	wire [WIDTH-1:0] wire_d0_31;
	wire [WIDTH-1:0] wire_d0_32;
	wire [WIDTH-1:0] wire_d0_33;
	wire [WIDTH-1:0] wire_d0_34;
	wire [WIDTH-1:0] wire_d0_35;
	wire [WIDTH-1:0] wire_d0_36;
	wire [WIDTH-1:0] wire_d0_37;
	wire [WIDTH-1:0] wire_d0_38;
	wire [WIDTH-1:0] wire_d0_39;
	wire [WIDTH-1:0] wire_d0_40;
	wire [WIDTH-1:0] wire_d0_41;
	wire [WIDTH-1:0] wire_d0_42;
	wire [WIDTH-1:0] wire_d0_43;
	wire [WIDTH-1:0] wire_d0_44;
	wire [WIDTH-1:0] wire_d0_45;
	wire [WIDTH-1:0] wire_d0_46;
	wire [WIDTH-1:0] wire_d0_47;
	wire [WIDTH-1:0] wire_d0_48;
	wire [WIDTH-1:0] wire_d0_49;
	wire [WIDTH-1:0] wire_d0_50;
	wire [WIDTH-1:0] wire_d0_51;
	wire [WIDTH-1:0] wire_d0_52;
	wire [WIDTH-1:0] wire_d0_53;
	wire [WIDTH-1:0] wire_d0_54;
	wire [WIDTH-1:0] wire_d0_55;
	wire [WIDTH-1:0] wire_d0_56;
	wire [WIDTH-1:0] wire_d0_57;
	wire [WIDTH-1:0] wire_d0_58;
	wire [WIDTH-1:0] wire_d0_59;
	wire [WIDTH-1:0] wire_d0_60;
	wire [WIDTH-1:0] wire_d0_61;
	wire [WIDTH-1:0] wire_d0_62;
	wire [WIDTH-1:0] wire_d0_63;
	wire [WIDTH-1:0] wire_d0_64;
	wire [WIDTH-1:0] wire_d0_65;
	wire [WIDTH-1:0] wire_d0_66;
	wire [WIDTH-1:0] wire_d0_67;
	wire [WIDTH-1:0] wire_d0_68;
	wire [WIDTH-1:0] wire_d0_69;
	wire [WIDTH-1:0] wire_d0_70;
	wire [WIDTH-1:0] wire_d0_71;
	wire [WIDTH-1:0] wire_d0_72;
	wire [WIDTH-1:0] wire_d0_73;
	wire [WIDTH-1:0] wire_d0_74;
	wire [WIDTH-1:0] wire_d0_75;
	wire [WIDTH-1:0] wire_d0_76;
	wire [WIDTH-1:0] wire_d0_77;
	wire [WIDTH-1:0] wire_d0_78;
	wire [WIDTH-1:0] wire_d0_79;
	wire [WIDTH-1:0] wire_d0_80;
	wire [WIDTH-1:0] wire_d0_81;
	wire [WIDTH-1:0] wire_d0_82;
	wire [WIDTH-1:0] wire_d0_83;
	wire [WIDTH-1:0] wire_d0_84;
	wire [WIDTH-1:0] wire_d0_85;
	wire [WIDTH-1:0] wire_d0_86;
	wire [WIDTH-1:0] wire_d0_87;
	wire [WIDTH-1:0] wire_d0_88;
	wire [WIDTH-1:0] wire_d0_89;
	wire [WIDTH-1:0] wire_d0_90;
	wire [WIDTH-1:0] wire_d0_91;
	wire [WIDTH-1:0] wire_d0_92;
	wire [WIDTH-1:0] wire_d0_93;
	wire [WIDTH-1:0] wire_d0_94;
	wire [WIDTH-1:0] wire_d0_95;
	wire [WIDTH-1:0] wire_d0_96;
	wire [WIDTH-1:0] wire_d0_97;
	wire [WIDTH-1:0] wire_d0_98;
	wire [WIDTH-1:0] wire_d1_0;
	wire [WIDTH-1:0] wire_d1_1;
	wire [WIDTH-1:0] wire_d1_2;
	wire [WIDTH-1:0] wire_d1_3;
	wire [WIDTH-1:0] wire_d1_4;
	wire [WIDTH-1:0] wire_d1_5;
	wire [WIDTH-1:0] wire_d1_6;
	wire [WIDTH-1:0] wire_d1_7;
	wire [WIDTH-1:0] wire_d1_8;
	wire [WIDTH-1:0] wire_d1_9;
	wire [WIDTH-1:0] wire_d1_10;
	wire [WIDTH-1:0] wire_d1_11;
	wire [WIDTH-1:0] wire_d1_12;
	wire [WIDTH-1:0] wire_d1_13;
	wire [WIDTH-1:0] wire_d1_14;
	wire [WIDTH-1:0] wire_d1_15;
	wire [WIDTH-1:0] wire_d1_16;
	wire [WIDTH-1:0] wire_d1_17;
	wire [WIDTH-1:0] wire_d1_18;
	wire [WIDTH-1:0] wire_d1_19;
	wire [WIDTH-1:0] wire_d1_20;
	wire [WIDTH-1:0] wire_d1_21;
	wire [WIDTH-1:0] wire_d1_22;
	wire [WIDTH-1:0] wire_d1_23;
	wire [WIDTH-1:0] wire_d1_24;
	wire [WIDTH-1:0] wire_d1_25;
	wire [WIDTH-1:0] wire_d1_26;
	wire [WIDTH-1:0] wire_d1_27;
	wire [WIDTH-1:0] wire_d1_28;
	wire [WIDTH-1:0] wire_d1_29;
	wire [WIDTH-1:0] wire_d1_30;
	wire [WIDTH-1:0] wire_d1_31;
	wire [WIDTH-1:0] wire_d1_32;
	wire [WIDTH-1:0] wire_d1_33;
	wire [WIDTH-1:0] wire_d1_34;
	wire [WIDTH-1:0] wire_d1_35;
	wire [WIDTH-1:0] wire_d1_36;
	wire [WIDTH-1:0] wire_d1_37;
	wire [WIDTH-1:0] wire_d1_38;
	wire [WIDTH-1:0] wire_d1_39;
	wire [WIDTH-1:0] wire_d1_40;
	wire [WIDTH-1:0] wire_d1_41;
	wire [WIDTH-1:0] wire_d1_42;
	wire [WIDTH-1:0] wire_d1_43;
	wire [WIDTH-1:0] wire_d1_44;
	wire [WIDTH-1:0] wire_d1_45;
	wire [WIDTH-1:0] wire_d1_46;
	wire [WIDTH-1:0] wire_d1_47;
	wire [WIDTH-1:0] wire_d1_48;
	wire [WIDTH-1:0] wire_d1_49;
	wire [WIDTH-1:0] wire_d1_50;
	wire [WIDTH-1:0] wire_d1_51;
	wire [WIDTH-1:0] wire_d1_52;
	wire [WIDTH-1:0] wire_d1_53;
	wire [WIDTH-1:0] wire_d1_54;
	wire [WIDTH-1:0] wire_d1_55;
	wire [WIDTH-1:0] wire_d1_56;
	wire [WIDTH-1:0] wire_d1_57;
	wire [WIDTH-1:0] wire_d1_58;
	wire [WIDTH-1:0] wire_d1_59;
	wire [WIDTH-1:0] wire_d1_60;
	wire [WIDTH-1:0] wire_d1_61;
	wire [WIDTH-1:0] wire_d1_62;
	wire [WIDTH-1:0] wire_d1_63;
	wire [WIDTH-1:0] wire_d1_64;
	wire [WIDTH-1:0] wire_d1_65;
	wire [WIDTH-1:0] wire_d1_66;
	wire [WIDTH-1:0] wire_d1_67;
	wire [WIDTH-1:0] wire_d1_68;
	wire [WIDTH-1:0] wire_d1_69;
	wire [WIDTH-1:0] wire_d1_70;
	wire [WIDTH-1:0] wire_d1_71;
	wire [WIDTH-1:0] wire_d1_72;
	wire [WIDTH-1:0] wire_d1_73;
	wire [WIDTH-1:0] wire_d1_74;
	wire [WIDTH-1:0] wire_d1_75;
	wire [WIDTH-1:0] wire_d1_76;
	wire [WIDTH-1:0] wire_d1_77;
	wire [WIDTH-1:0] wire_d1_78;
	wire [WIDTH-1:0] wire_d1_79;
	wire [WIDTH-1:0] wire_d1_80;
	wire [WIDTH-1:0] wire_d1_81;
	wire [WIDTH-1:0] wire_d1_82;
	wire [WIDTH-1:0] wire_d1_83;
	wire [WIDTH-1:0] wire_d1_84;
	wire [WIDTH-1:0] wire_d1_85;
	wire [WIDTH-1:0] wire_d1_86;
	wire [WIDTH-1:0] wire_d1_87;
	wire [WIDTH-1:0] wire_d1_88;
	wire [WIDTH-1:0] wire_d1_89;
	wire [WIDTH-1:0] wire_d1_90;
	wire [WIDTH-1:0] wire_d1_91;
	wire [WIDTH-1:0] wire_d1_92;
	wire [WIDTH-1:0] wire_d1_93;
	wire [WIDTH-1:0] wire_d1_94;
	wire [WIDTH-1:0] wire_d1_95;
	wire [WIDTH-1:0] wire_d1_96;
	wire [WIDTH-1:0] wire_d1_97;
	wire [WIDTH-1:0] wire_d1_98;
	wire [WIDTH-1:0] wire_d2_0;
	wire [WIDTH-1:0] wire_d2_1;
	wire [WIDTH-1:0] wire_d2_2;
	wire [WIDTH-1:0] wire_d2_3;
	wire [WIDTH-1:0] wire_d2_4;
	wire [WIDTH-1:0] wire_d2_5;
	wire [WIDTH-1:0] wire_d2_6;
	wire [WIDTH-1:0] wire_d2_7;
	wire [WIDTH-1:0] wire_d2_8;
	wire [WIDTH-1:0] wire_d2_9;
	wire [WIDTH-1:0] wire_d2_10;
	wire [WIDTH-1:0] wire_d2_11;
	wire [WIDTH-1:0] wire_d2_12;
	wire [WIDTH-1:0] wire_d2_13;
	wire [WIDTH-1:0] wire_d2_14;
	wire [WIDTH-1:0] wire_d2_15;
	wire [WIDTH-1:0] wire_d2_16;
	wire [WIDTH-1:0] wire_d2_17;
	wire [WIDTH-1:0] wire_d2_18;
	wire [WIDTH-1:0] wire_d2_19;
	wire [WIDTH-1:0] wire_d2_20;
	wire [WIDTH-1:0] wire_d2_21;
	wire [WIDTH-1:0] wire_d2_22;
	wire [WIDTH-1:0] wire_d2_23;
	wire [WIDTH-1:0] wire_d2_24;
	wire [WIDTH-1:0] wire_d2_25;
	wire [WIDTH-1:0] wire_d2_26;
	wire [WIDTH-1:0] wire_d2_27;
	wire [WIDTH-1:0] wire_d2_28;
	wire [WIDTH-1:0] wire_d2_29;
	wire [WIDTH-1:0] wire_d2_30;
	wire [WIDTH-1:0] wire_d2_31;
	wire [WIDTH-1:0] wire_d2_32;
	wire [WIDTH-1:0] wire_d2_33;
	wire [WIDTH-1:0] wire_d2_34;
	wire [WIDTH-1:0] wire_d2_35;
	wire [WIDTH-1:0] wire_d2_36;
	wire [WIDTH-1:0] wire_d2_37;
	wire [WIDTH-1:0] wire_d2_38;
	wire [WIDTH-1:0] wire_d2_39;
	wire [WIDTH-1:0] wire_d2_40;
	wire [WIDTH-1:0] wire_d2_41;
	wire [WIDTH-1:0] wire_d2_42;
	wire [WIDTH-1:0] wire_d2_43;
	wire [WIDTH-1:0] wire_d2_44;
	wire [WIDTH-1:0] wire_d2_45;
	wire [WIDTH-1:0] wire_d2_46;
	wire [WIDTH-1:0] wire_d2_47;
	wire [WIDTH-1:0] wire_d2_48;
	wire [WIDTH-1:0] wire_d2_49;
	wire [WIDTH-1:0] wire_d2_50;
	wire [WIDTH-1:0] wire_d2_51;
	wire [WIDTH-1:0] wire_d2_52;
	wire [WIDTH-1:0] wire_d2_53;
	wire [WIDTH-1:0] wire_d2_54;
	wire [WIDTH-1:0] wire_d2_55;
	wire [WIDTH-1:0] wire_d2_56;
	wire [WIDTH-1:0] wire_d2_57;
	wire [WIDTH-1:0] wire_d2_58;
	wire [WIDTH-1:0] wire_d2_59;
	wire [WIDTH-1:0] wire_d2_60;
	wire [WIDTH-1:0] wire_d2_61;
	wire [WIDTH-1:0] wire_d2_62;
	wire [WIDTH-1:0] wire_d2_63;
	wire [WIDTH-1:0] wire_d2_64;
	wire [WIDTH-1:0] wire_d2_65;
	wire [WIDTH-1:0] wire_d2_66;
	wire [WIDTH-1:0] wire_d2_67;
	wire [WIDTH-1:0] wire_d2_68;
	wire [WIDTH-1:0] wire_d2_69;
	wire [WIDTH-1:0] wire_d2_70;
	wire [WIDTH-1:0] wire_d2_71;
	wire [WIDTH-1:0] wire_d2_72;
	wire [WIDTH-1:0] wire_d2_73;
	wire [WIDTH-1:0] wire_d2_74;
	wire [WIDTH-1:0] wire_d2_75;
	wire [WIDTH-1:0] wire_d2_76;
	wire [WIDTH-1:0] wire_d2_77;
	wire [WIDTH-1:0] wire_d2_78;
	wire [WIDTH-1:0] wire_d2_79;
	wire [WIDTH-1:0] wire_d2_80;
	wire [WIDTH-1:0] wire_d2_81;
	wire [WIDTH-1:0] wire_d2_82;
	wire [WIDTH-1:0] wire_d2_83;
	wire [WIDTH-1:0] wire_d2_84;
	wire [WIDTH-1:0] wire_d2_85;
	wire [WIDTH-1:0] wire_d2_86;
	wire [WIDTH-1:0] wire_d2_87;
	wire [WIDTH-1:0] wire_d2_88;
	wire [WIDTH-1:0] wire_d2_89;
	wire [WIDTH-1:0] wire_d2_90;
	wire [WIDTH-1:0] wire_d2_91;
	wire [WIDTH-1:0] wire_d2_92;
	wire [WIDTH-1:0] wire_d2_93;
	wire [WIDTH-1:0] wire_d2_94;
	wire [WIDTH-1:0] wire_d2_95;
	wire [WIDTH-1:0] wire_d2_96;
	wire [WIDTH-1:0] wire_d2_97;
	wire [WIDTH-1:0] wire_d2_98;
	wire [WIDTH-1:0] wire_d3_0;
	wire [WIDTH-1:0] wire_d3_1;
	wire [WIDTH-1:0] wire_d3_2;
	wire [WIDTH-1:0] wire_d3_3;
	wire [WIDTH-1:0] wire_d3_4;
	wire [WIDTH-1:0] wire_d3_5;
	wire [WIDTH-1:0] wire_d3_6;
	wire [WIDTH-1:0] wire_d3_7;
	wire [WIDTH-1:0] wire_d3_8;
	wire [WIDTH-1:0] wire_d3_9;
	wire [WIDTH-1:0] wire_d3_10;
	wire [WIDTH-1:0] wire_d3_11;
	wire [WIDTH-1:0] wire_d3_12;
	wire [WIDTH-1:0] wire_d3_13;
	wire [WIDTH-1:0] wire_d3_14;
	wire [WIDTH-1:0] wire_d3_15;
	wire [WIDTH-1:0] wire_d3_16;
	wire [WIDTH-1:0] wire_d3_17;
	wire [WIDTH-1:0] wire_d3_18;
	wire [WIDTH-1:0] wire_d3_19;
	wire [WIDTH-1:0] wire_d3_20;
	wire [WIDTH-1:0] wire_d3_21;
	wire [WIDTH-1:0] wire_d3_22;
	wire [WIDTH-1:0] wire_d3_23;
	wire [WIDTH-1:0] wire_d3_24;
	wire [WIDTH-1:0] wire_d3_25;
	wire [WIDTH-1:0] wire_d3_26;
	wire [WIDTH-1:0] wire_d3_27;
	wire [WIDTH-1:0] wire_d3_28;
	wire [WIDTH-1:0] wire_d3_29;
	wire [WIDTH-1:0] wire_d3_30;
	wire [WIDTH-1:0] wire_d3_31;
	wire [WIDTH-1:0] wire_d3_32;
	wire [WIDTH-1:0] wire_d3_33;
	wire [WIDTH-1:0] wire_d3_34;
	wire [WIDTH-1:0] wire_d3_35;
	wire [WIDTH-1:0] wire_d3_36;
	wire [WIDTH-1:0] wire_d3_37;
	wire [WIDTH-1:0] wire_d3_38;
	wire [WIDTH-1:0] wire_d3_39;
	wire [WIDTH-1:0] wire_d3_40;
	wire [WIDTH-1:0] wire_d3_41;
	wire [WIDTH-1:0] wire_d3_42;
	wire [WIDTH-1:0] wire_d3_43;
	wire [WIDTH-1:0] wire_d3_44;
	wire [WIDTH-1:0] wire_d3_45;
	wire [WIDTH-1:0] wire_d3_46;
	wire [WIDTH-1:0] wire_d3_47;
	wire [WIDTH-1:0] wire_d3_48;
	wire [WIDTH-1:0] wire_d3_49;
	wire [WIDTH-1:0] wire_d3_50;
	wire [WIDTH-1:0] wire_d3_51;
	wire [WIDTH-1:0] wire_d3_52;
	wire [WIDTH-1:0] wire_d3_53;
	wire [WIDTH-1:0] wire_d3_54;
	wire [WIDTH-1:0] wire_d3_55;
	wire [WIDTH-1:0] wire_d3_56;
	wire [WIDTH-1:0] wire_d3_57;
	wire [WIDTH-1:0] wire_d3_58;
	wire [WIDTH-1:0] wire_d3_59;
	wire [WIDTH-1:0] wire_d3_60;
	wire [WIDTH-1:0] wire_d3_61;
	wire [WIDTH-1:0] wire_d3_62;
	wire [WIDTH-1:0] wire_d3_63;
	wire [WIDTH-1:0] wire_d3_64;
	wire [WIDTH-1:0] wire_d3_65;
	wire [WIDTH-1:0] wire_d3_66;
	wire [WIDTH-1:0] wire_d3_67;
	wire [WIDTH-1:0] wire_d3_68;
	wire [WIDTH-1:0] wire_d3_69;
	wire [WIDTH-1:0] wire_d3_70;
	wire [WIDTH-1:0] wire_d3_71;
	wire [WIDTH-1:0] wire_d3_72;
	wire [WIDTH-1:0] wire_d3_73;
	wire [WIDTH-1:0] wire_d3_74;
	wire [WIDTH-1:0] wire_d3_75;
	wire [WIDTH-1:0] wire_d3_76;
	wire [WIDTH-1:0] wire_d3_77;
	wire [WIDTH-1:0] wire_d3_78;
	wire [WIDTH-1:0] wire_d3_79;
	wire [WIDTH-1:0] wire_d3_80;
	wire [WIDTH-1:0] wire_d3_81;
	wire [WIDTH-1:0] wire_d3_82;
	wire [WIDTH-1:0] wire_d3_83;
	wire [WIDTH-1:0] wire_d3_84;
	wire [WIDTH-1:0] wire_d3_85;
	wire [WIDTH-1:0] wire_d3_86;
	wire [WIDTH-1:0] wire_d3_87;
	wire [WIDTH-1:0] wire_d3_88;
	wire [WIDTH-1:0] wire_d3_89;
	wire [WIDTH-1:0] wire_d3_90;
	wire [WIDTH-1:0] wire_d3_91;
	wire [WIDTH-1:0] wire_d3_92;
	wire [WIDTH-1:0] wire_d3_93;
	wire [WIDTH-1:0] wire_d3_94;
	wire [WIDTH-1:0] wire_d3_95;
	wire [WIDTH-1:0] wire_d3_96;
	wire [WIDTH-1:0] wire_d3_97;
	wire [WIDTH-1:0] wire_d3_98;
	wire [WIDTH-1:0] wire_d4_0;
	wire [WIDTH-1:0] wire_d4_1;
	wire [WIDTH-1:0] wire_d4_2;
	wire [WIDTH-1:0] wire_d4_3;
	wire [WIDTH-1:0] wire_d4_4;
	wire [WIDTH-1:0] wire_d4_5;
	wire [WIDTH-1:0] wire_d4_6;
	wire [WIDTH-1:0] wire_d4_7;
	wire [WIDTH-1:0] wire_d4_8;
	wire [WIDTH-1:0] wire_d4_9;
	wire [WIDTH-1:0] wire_d4_10;
	wire [WIDTH-1:0] wire_d4_11;
	wire [WIDTH-1:0] wire_d4_12;
	wire [WIDTH-1:0] wire_d4_13;
	wire [WIDTH-1:0] wire_d4_14;
	wire [WIDTH-1:0] wire_d4_15;
	wire [WIDTH-1:0] wire_d4_16;
	wire [WIDTH-1:0] wire_d4_17;
	wire [WIDTH-1:0] wire_d4_18;
	wire [WIDTH-1:0] wire_d4_19;
	wire [WIDTH-1:0] wire_d4_20;
	wire [WIDTH-1:0] wire_d4_21;
	wire [WIDTH-1:0] wire_d4_22;
	wire [WIDTH-1:0] wire_d4_23;
	wire [WIDTH-1:0] wire_d4_24;
	wire [WIDTH-1:0] wire_d4_25;
	wire [WIDTH-1:0] wire_d4_26;
	wire [WIDTH-1:0] wire_d4_27;
	wire [WIDTH-1:0] wire_d4_28;
	wire [WIDTH-1:0] wire_d4_29;
	wire [WIDTH-1:0] wire_d4_30;
	wire [WIDTH-1:0] wire_d4_31;
	wire [WIDTH-1:0] wire_d4_32;
	wire [WIDTH-1:0] wire_d4_33;
	wire [WIDTH-1:0] wire_d4_34;
	wire [WIDTH-1:0] wire_d4_35;
	wire [WIDTH-1:0] wire_d4_36;
	wire [WIDTH-1:0] wire_d4_37;
	wire [WIDTH-1:0] wire_d4_38;
	wire [WIDTH-1:0] wire_d4_39;
	wire [WIDTH-1:0] wire_d4_40;
	wire [WIDTH-1:0] wire_d4_41;
	wire [WIDTH-1:0] wire_d4_42;
	wire [WIDTH-1:0] wire_d4_43;
	wire [WIDTH-1:0] wire_d4_44;
	wire [WIDTH-1:0] wire_d4_45;
	wire [WIDTH-1:0] wire_d4_46;
	wire [WIDTH-1:0] wire_d4_47;
	wire [WIDTH-1:0] wire_d4_48;
	wire [WIDTH-1:0] wire_d4_49;
	wire [WIDTH-1:0] wire_d4_50;
	wire [WIDTH-1:0] wire_d4_51;
	wire [WIDTH-1:0] wire_d4_52;
	wire [WIDTH-1:0] wire_d4_53;
	wire [WIDTH-1:0] wire_d4_54;
	wire [WIDTH-1:0] wire_d4_55;
	wire [WIDTH-1:0] wire_d4_56;
	wire [WIDTH-1:0] wire_d4_57;
	wire [WIDTH-1:0] wire_d4_58;
	wire [WIDTH-1:0] wire_d4_59;
	wire [WIDTH-1:0] wire_d4_60;
	wire [WIDTH-1:0] wire_d4_61;
	wire [WIDTH-1:0] wire_d4_62;
	wire [WIDTH-1:0] wire_d4_63;
	wire [WIDTH-1:0] wire_d4_64;
	wire [WIDTH-1:0] wire_d4_65;
	wire [WIDTH-1:0] wire_d4_66;
	wire [WIDTH-1:0] wire_d4_67;
	wire [WIDTH-1:0] wire_d4_68;
	wire [WIDTH-1:0] wire_d4_69;
	wire [WIDTH-1:0] wire_d4_70;
	wire [WIDTH-1:0] wire_d4_71;
	wire [WIDTH-1:0] wire_d4_72;
	wire [WIDTH-1:0] wire_d4_73;
	wire [WIDTH-1:0] wire_d4_74;
	wire [WIDTH-1:0] wire_d4_75;
	wire [WIDTH-1:0] wire_d4_76;
	wire [WIDTH-1:0] wire_d4_77;
	wire [WIDTH-1:0] wire_d4_78;
	wire [WIDTH-1:0] wire_d4_79;
	wire [WIDTH-1:0] wire_d4_80;
	wire [WIDTH-1:0] wire_d4_81;
	wire [WIDTH-1:0] wire_d4_82;
	wire [WIDTH-1:0] wire_d4_83;
	wire [WIDTH-1:0] wire_d4_84;
	wire [WIDTH-1:0] wire_d4_85;
	wire [WIDTH-1:0] wire_d4_86;
	wire [WIDTH-1:0] wire_d4_87;
	wire [WIDTH-1:0] wire_d4_88;
	wire [WIDTH-1:0] wire_d4_89;
	wire [WIDTH-1:0] wire_d4_90;
	wire [WIDTH-1:0] wire_d4_91;
	wire [WIDTH-1:0] wire_d4_92;
	wire [WIDTH-1:0] wire_d4_93;
	wire [WIDTH-1:0] wire_d4_94;
	wire [WIDTH-1:0] wire_d4_95;
	wire [WIDTH-1:0] wire_d4_96;
	wire [WIDTH-1:0] wire_d4_97;
	wire [WIDTH-1:0] wire_d4_98;
	wire [WIDTH-1:0] wire_d5_0;
	wire [WIDTH-1:0] wire_d5_1;
	wire [WIDTH-1:0] wire_d5_2;
	wire [WIDTH-1:0] wire_d5_3;
	wire [WIDTH-1:0] wire_d5_4;
	wire [WIDTH-1:0] wire_d5_5;
	wire [WIDTH-1:0] wire_d5_6;
	wire [WIDTH-1:0] wire_d5_7;
	wire [WIDTH-1:0] wire_d5_8;
	wire [WIDTH-1:0] wire_d5_9;
	wire [WIDTH-1:0] wire_d5_10;
	wire [WIDTH-1:0] wire_d5_11;
	wire [WIDTH-1:0] wire_d5_12;
	wire [WIDTH-1:0] wire_d5_13;
	wire [WIDTH-1:0] wire_d5_14;
	wire [WIDTH-1:0] wire_d5_15;
	wire [WIDTH-1:0] wire_d5_16;
	wire [WIDTH-1:0] wire_d5_17;
	wire [WIDTH-1:0] wire_d5_18;
	wire [WIDTH-1:0] wire_d5_19;
	wire [WIDTH-1:0] wire_d5_20;
	wire [WIDTH-1:0] wire_d5_21;
	wire [WIDTH-1:0] wire_d5_22;
	wire [WIDTH-1:0] wire_d5_23;
	wire [WIDTH-1:0] wire_d5_24;
	wire [WIDTH-1:0] wire_d5_25;
	wire [WIDTH-1:0] wire_d5_26;
	wire [WIDTH-1:0] wire_d5_27;
	wire [WIDTH-1:0] wire_d5_28;
	wire [WIDTH-1:0] wire_d5_29;
	wire [WIDTH-1:0] wire_d5_30;
	wire [WIDTH-1:0] wire_d5_31;
	wire [WIDTH-1:0] wire_d5_32;
	wire [WIDTH-1:0] wire_d5_33;
	wire [WIDTH-1:0] wire_d5_34;
	wire [WIDTH-1:0] wire_d5_35;
	wire [WIDTH-1:0] wire_d5_36;
	wire [WIDTH-1:0] wire_d5_37;
	wire [WIDTH-1:0] wire_d5_38;
	wire [WIDTH-1:0] wire_d5_39;
	wire [WIDTH-1:0] wire_d5_40;
	wire [WIDTH-1:0] wire_d5_41;
	wire [WIDTH-1:0] wire_d5_42;
	wire [WIDTH-1:0] wire_d5_43;
	wire [WIDTH-1:0] wire_d5_44;
	wire [WIDTH-1:0] wire_d5_45;
	wire [WIDTH-1:0] wire_d5_46;
	wire [WIDTH-1:0] wire_d5_47;
	wire [WIDTH-1:0] wire_d5_48;
	wire [WIDTH-1:0] wire_d5_49;
	wire [WIDTH-1:0] wire_d5_50;
	wire [WIDTH-1:0] wire_d5_51;
	wire [WIDTH-1:0] wire_d5_52;
	wire [WIDTH-1:0] wire_d5_53;
	wire [WIDTH-1:0] wire_d5_54;
	wire [WIDTH-1:0] wire_d5_55;
	wire [WIDTH-1:0] wire_d5_56;
	wire [WIDTH-1:0] wire_d5_57;
	wire [WIDTH-1:0] wire_d5_58;
	wire [WIDTH-1:0] wire_d5_59;
	wire [WIDTH-1:0] wire_d5_60;
	wire [WIDTH-1:0] wire_d5_61;
	wire [WIDTH-1:0] wire_d5_62;
	wire [WIDTH-1:0] wire_d5_63;
	wire [WIDTH-1:0] wire_d5_64;
	wire [WIDTH-1:0] wire_d5_65;
	wire [WIDTH-1:0] wire_d5_66;
	wire [WIDTH-1:0] wire_d5_67;
	wire [WIDTH-1:0] wire_d5_68;
	wire [WIDTH-1:0] wire_d5_69;
	wire [WIDTH-1:0] wire_d5_70;
	wire [WIDTH-1:0] wire_d5_71;
	wire [WIDTH-1:0] wire_d5_72;
	wire [WIDTH-1:0] wire_d5_73;
	wire [WIDTH-1:0] wire_d5_74;
	wire [WIDTH-1:0] wire_d5_75;
	wire [WIDTH-1:0] wire_d5_76;
	wire [WIDTH-1:0] wire_d5_77;
	wire [WIDTH-1:0] wire_d5_78;
	wire [WIDTH-1:0] wire_d5_79;
	wire [WIDTH-1:0] wire_d5_80;
	wire [WIDTH-1:0] wire_d5_81;
	wire [WIDTH-1:0] wire_d5_82;
	wire [WIDTH-1:0] wire_d5_83;
	wire [WIDTH-1:0] wire_d5_84;
	wire [WIDTH-1:0] wire_d5_85;
	wire [WIDTH-1:0] wire_d5_86;
	wire [WIDTH-1:0] wire_d5_87;
	wire [WIDTH-1:0] wire_d5_88;
	wire [WIDTH-1:0] wire_d5_89;
	wire [WIDTH-1:0] wire_d5_90;
	wire [WIDTH-1:0] wire_d5_91;
	wire [WIDTH-1:0] wire_d5_92;
	wire [WIDTH-1:0] wire_d5_93;
	wire [WIDTH-1:0] wire_d5_94;
	wire [WIDTH-1:0] wire_d5_95;
	wire [WIDTH-1:0] wire_d5_96;
	wire [WIDTH-1:0] wire_d5_97;
	wire [WIDTH-1:0] wire_d5_98;
	wire [WIDTH-1:0] wire_d6_0;
	wire [WIDTH-1:0] wire_d6_1;
	wire [WIDTH-1:0] wire_d6_2;
	wire [WIDTH-1:0] wire_d6_3;
	wire [WIDTH-1:0] wire_d6_4;
	wire [WIDTH-1:0] wire_d6_5;
	wire [WIDTH-1:0] wire_d6_6;
	wire [WIDTH-1:0] wire_d6_7;
	wire [WIDTH-1:0] wire_d6_8;
	wire [WIDTH-1:0] wire_d6_9;
	wire [WIDTH-1:0] wire_d6_10;
	wire [WIDTH-1:0] wire_d6_11;
	wire [WIDTH-1:0] wire_d6_12;
	wire [WIDTH-1:0] wire_d6_13;
	wire [WIDTH-1:0] wire_d6_14;
	wire [WIDTH-1:0] wire_d6_15;
	wire [WIDTH-1:0] wire_d6_16;
	wire [WIDTH-1:0] wire_d6_17;
	wire [WIDTH-1:0] wire_d6_18;
	wire [WIDTH-1:0] wire_d6_19;
	wire [WIDTH-1:0] wire_d6_20;
	wire [WIDTH-1:0] wire_d6_21;
	wire [WIDTH-1:0] wire_d6_22;
	wire [WIDTH-1:0] wire_d6_23;
	wire [WIDTH-1:0] wire_d6_24;
	wire [WIDTH-1:0] wire_d6_25;
	wire [WIDTH-1:0] wire_d6_26;
	wire [WIDTH-1:0] wire_d6_27;
	wire [WIDTH-1:0] wire_d6_28;
	wire [WIDTH-1:0] wire_d6_29;
	wire [WIDTH-1:0] wire_d6_30;
	wire [WIDTH-1:0] wire_d6_31;
	wire [WIDTH-1:0] wire_d6_32;
	wire [WIDTH-1:0] wire_d6_33;
	wire [WIDTH-1:0] wire_d6_34;
	wire [WIDTH-1:0] wire_d6_35;
	wire [WIDTH-1:0] wire_d6_36;
	wire [WIDTH-1:0] wire_d6_37;
	wire [WIDTH-1:0] wire_d6_38;
	wire [WIDTH-1:0] wire_d6_39;
	wire [WIDTH-1:0] wire_d6_40;
	wire [WIDTH-1:0] wire_d6_41;
	wire [WIDTH-1:0] wire_d6_42;
	wire [WIDTH-1:0] wire_d6_43;
	wire [WIDTH-1:0] wire_d6_44;
	wire [WIDTH-1:0] wire_d6_45;
	wire [WIDTH-1:0] wire_d6_46;
	wire [WIDTH-1:0] wire_d6_47;
	wire [WIDTH-1:0] wire_d6_48;
	wire [WIDTH-1:0] wire_d6_49;
	wire [WIDTH-1:0] wire_d6_50;
	wire [WIDTH-1:0] wire_d6_51;
	wire [WIDTH-1:0] wire_d6_52;
	wire [WIDTH-1:0] wire_d6_53;
	wire [WIDTH-1:0] wire_d6_54;
	wire [WIDTH-1:0] wire_d6_55;
	wire [WIDTH-1:0] wire_d6_56;
	wire [WIDTH-1:0] wire_d6_57;
	wire [WIDTH-1:0] wire_d6_58;
	wire [WIDTH-1:0] wire_d6_59;
	wire [WIDTH-1:0] wire_d6_60;
	wire [WIDTH-1:0] wire_d6_61;
	wire [WIDTH-1:0] wire_d6_62;
	wire [WIDTH-1:0] wire_d6_63;
	wire [WIDTH-1:0] wire_d6_64;
	wire [WIDTH-1:0] wire_d6_65;
	wire [WIDTH-1:0] wire_d6_66;
	wire [WIDTH-1:0] wire_d6_67;
	wire [WIDTH-1:0] wire_d6_68;
	wire [WIDTH-1:0] wire_d6_69;
	wire [WIDTH-1:0] wire_d6_70;
	wire [WIDTH-1:0] wire_d6_71;
	wire [WIDTH-1:0] wire_d6_72;
	wire [WIDTH-1:0] wire_d6_73;
	wire [WIDTH-1:0] wire_d6_74;
	wire [WIDTH-1:0] wire_d6_75;
	wire [WIDTH-1:0] wire_d6_76;
	wire [WIDTH-1:0] wire_d6_77;
	wire [WIDTH-1:0] wire_d6_78;
	wire [WIDTH-1:0] wire_d6_79;
	wire [WIDTH-1:0] wire_d6_80;
	wire [WIDTH-1:0] wire_d6_81;
	wire [WIDTH-1:0] wire_d6_82;
	wire [WIDTH-1:0] wire_d6_83;
	wire [WIDTH-1:0] wire_d6_84;
	wire [WIDTH-1:0] wire_d6_85;
	wire [WIDTH-1:0] wire_d6_86;
	wire [WIDTH-1:0] wire_d6_87;
	wire [WIDTH-1:0] wire_d6_88;
	wire [WIDTH-1:0] wire_d6_89;
	wire [WIDTH-1:0] wire_d6_90;
	wire [WIDTH-1:0] wire_d6_91;
	wire [WIDTH-1:0] wire_d6_92;
	wire [WIDTH-1:0] wire_d6_93;
	wire [WIDTH-1:0] wire_d6_94;
	wire [WIDTH-1:0] wire_d6_95;
	wire [WIDTH-1:0] wire_d6_96;
	wire [WIDTH-1:0] wire_d6_97;
	wire [WIDTH-1:0] wire_d6_98;
	wire [WIDTH-1:0] wire_d7_0;
	wire [WIDTH-1:0] wire_d7_1;
	wire [WIDTH-1:0] wire_d7_2;
	wire [WIDTH-1:0] wire_d7_3;
	wire [WIDTH-1:0] wire_d7_4;
	wire [WIDTH-1:0] wire_d7_5;
	wire [WIDTH-1:0] wire_d7_6;
	wire [WIDTH-1:0] wire_d7_7;
	wire [WIDTH-1:0] wire_d7_8;
	wire [WIDTH-1:0] wire_d7_9;
	wire [WIDTH-1:0] wire_d7_10;
	wire [WIDTH-1:0] wire_d7_11;
	wire [WIDTH-1:0] wire_d7_12;
	wire [WIDTH-1:0] wire_d7_13;
	wire [WIDTH-1:0] wire_d7_14;
	wire [WIDTH-1:0] wire_d7_15;
	wire [WIDTH-1:0] wire_d7_16;
	wire [WIDTH-1:0] wire_d7_17;
	wire [WIDTH-1:0] wire_d7_18;
	wire [WIDTH-1:0] wire_d7_19;
	wire [WIDTH-1:0] wire_d7_20;
	wire [WIDTH-1:0] wire_d7_21;
	wire [WIDTH-1:0] wire_d7_22;
	wire [WIDTH-1:0] wire_d7_23;
	wire [WIDTH-1:0] wire_d7_24;
	wire [WIDTH-1:0] wire_d7_25;
	wire [WIDTH-1:0] wire_d7_26;
	wire [WIDTH-1:0] wire_d7_27;
	wire [WIDTH-1:0] wire_d7_28;
	wire [WIDTH-1:0] wire_d7_29;
	wire [WIDTH-1:0] wire_d7_30;
	wire [WIDTH-1:0] wire_d7_31;
	wire [WIDTH-1:0] wire_d7_32;
	wire [WIDTH-1:0] wire_d7_33;
	wire [WIDTH-1:0] wire_d7_34;
	wire [WIDTH-1:0] wire_d7_35;
	wire [WIDTH-1:0] wire_d7_36;
	wire [WIDTH-1:0] wire_d7_37;
	wire [WIDTH-1:0] wire_d7_38;
	wire [WIDTH-1:0] wire_d7_39;
	wire [WIDTH-1:0] wire_d7_40;
	wire [WIDTH-1:0] wire_d7_41;
	wire [WIDTH-1:0] wire_d7_42;
	wire [WIDTH-1:0] wire_d7_43;
	wire [WIDTH-1:0] wire_d7_44;
	wire [WIDTH-1:0] wire_d7_45;
	wire [WIDTH-1:0] wire_d7_46;
	wire [WIDTH-1:0] wire_d7_47;
	wire [WIDTH-1:0] wire_d7_48;
	wire [WIDTH-1:0] wire_d7_49;
	wire [WIDTH-1:0] wire_d7_50;
	wire [WIDTH-1:0] wire_d7_51;
	wire [WIDTH-1:0] wire_d7_52;
	wire [WIDTH-1:0] wire_d7_53;
	wire [WIDTH-1:0] wire_d7_54;
	wire [WIDTH-1:0] wire_d7_55;
	wire [WIDTH-1:0] wire_d7_56;
	wire [WIDTH-1:0] wire_d7_57;
	wire [WIDTH-1:0] wire_d7_58;
	wire [WIDTH-1:0] wire_d7_59;
	wire [WIDTH-1:0] wire_d7_60;
	wire [WIDTH-1:0] wire_d7_61;
	wire [WIDTH-1:0] wire_d7_62;
	wire [WIDTH-1:0] wire_d7_63;
	wire [WIDTH-1:0] wire_d7_64;
	wire [WIDTH-1:0] wire_d7_65;
	wire [WIDTH-1:0] wire_d7_66;
	wire [WIDTH-1:0] wire_d7_67;
	wire [WIDTH-1:0] wire_d7_68;
	wire [WIDTH-1:0] wire_d7_69;
	wire [WIDTH-1:0] wire_d7_70;
	wire [WIDTH-1:0] wire_d7_71;
	wire [WIDTH-1:0] wire_d7_72;
	wire [WIDTH-1:0] wire_d7_73;
	wire [WIDTH-1:0] wire_d7_74;
	wire [WIDTH-1:0] wire_d7_75;
	wire [WIDTH-1:0] wire_d7_76;
	wire [WIDTH-1:0] wire_d7_77;
	wire [WIDTH-1:0] wire_d7_78;
	wire [WIDTH-1:0] wire_d7_79;
	wire [WIDTH-1:0] wire_d7_80;
	wire [WIDTH-1:0] wire_d7_81;
	wire [WIDTH-1:0] wire_d7_82;
	wire [WIDTH-1:0] wire_d7_83;
	wire [WIDTH-1:0] wire_d7_84;
	wire [WIDTH-1:0] wire_d7_85;
	wire [WIDTH-1:0] wire_d7_86;
	wire [WIDTH-1:0] wire_d7_87;
	wire [WIDTH-1:0] wire_d7_88;
	wire [WIDTH-1:0] wire_d7_89;
	wire [WIDTH-1:0] wire_d7_90;
	wire [WIDTH-1:0] wire_d7_91;
	wire [WIDTH-1:0] wire_d7_92;
	wire [WIDTH-1:0] wire_d7_93;
	wire [WIDTH-1:0] wire_d7_94;
	wire [WIDTH-1:0] wire_d7_95;
	wire [WIDTH-1:0] wire_d7_96;
	wire [WIDTH-1:0] wire_d7_97;
	wire [WIDTH-1:0] wire_d7_98;
	wire [WIDTH-1:0] wire_d8_0;
	wire [WIDTH-1:0] wire_d8_1;
	wire [WIDTH-1:0] wire_d8_2;
	wire [WIDTH-1:0] wire_d8_3;
	wire [WIDTH-1:0] wire_d8_4;
	wire [WIDTH-1:0] wire_d8_5;
	wire [WIDTH-1:0] wire_d8_6;
	wire [WIDTH-1:0] wire_d8_7;
	wire [WIDTH-1:0] wire_d8_8;
	wire [WIDTH-1:0] wire_d8_9;
	wire [WIDTH-1:0] wire_d8_10;
	wire [WIDTH-1:0] wire_d8_11;
	wire [WIDTH-1:0] wire_d8_12;
	wire [WIDTH-1:0] wire_d8_13;
	wire [WIDTH-1:0] wire_d8_14;
	wire [WIDTH-1:0] wire_d8_15;
	wire [WIDTH-1:0] wire_d8_16;
	wire [WIDTH-1:0] wire_d8_17;
	wire [WIDTH-1:0] wire_d8_18;
	wire [WIDTH-1:0] wire_d8_19;
	wire [WIDTH-1:0] wire_d8_20;
	wire [WIDTH-1:0] wire_d8_21;
	wire [WIDTH-1:0] wire_d8_22;
	wire [WIDTH-1:0] wire_d8_23;
	wire [WIDTH-1:0] wire_d8_24;
	wire [WIDTH-1:0] wire_d8_25;
	wire [WIDTH-1:0] wire_d8_26;
	wire [WIDTH-1:0] wire_d8_27;
	wire [WIDTH-1:0] wire_d8_28;
	wire [WIDTH-1:0] wire_d8_29;
	wire [WIDTH-1:0] wire_d8_30;
	wire [WIDTH-1:0] wire_d8_31;
	wire [WIDTH-1:0] wire_d8_32;
	wire [WIDTH-1:0] wire_d8_33;
	wire [WIDTH-1:0] wire_d8_34;
	wire [WIDTH-1:0] wire_d8_35;
	wire [WIDTH-1:0] wire_d8_36;
	wire [WIDTH-1:0] wire_d8_37;
	wire [WIDTH-1:0] wire_d8_38;
	wire [WIDTH-1:0] wire_d8_39;
	wire [WIDTH-1:0] wire_d8_40;
	wire [WIDTH-1:0] wire_d8_41;
	wire [WIDTH-1:0] wire_d8_42;
	wire [WIDTH-1:0] wire_d8_43;
	wire [WIDTH-1:0] wire_d8_44;
	wire [WIDTH-1:0] wire_d8_45;
	wire [WIDTH-1:0] wire_d8_46;
	wire [WIDTH-1:0] wire_d8_47;
	wire [WIDTH-1:0] wire_d8_48;
	wire [WIDTH-1:0] wire_d8_49;
	wire [WIDTH-1:0] wire_d8_50;
	wire [WIDTH-1:0] wire_d8_51;
	wire [WIDTH-1:0] wire_d8_52;
	wire [WIDTH-1:0] wire_d8_53;
	wire [WIDTH-1:0] wire_d8_54;
	wire [WIDTH-1:0] wire_d8_55;
	wire [WIDTH-1:0] wire_d8_56;
	wire [WIDTH-1:0] wire_d8_57;
	wire [WIDTH-1:0] wire_d8_58;
	wire [WIDTH-1:0] wire_d8_59;
	wire [WIDTH-1:0] wire_d8_60;
	wire [WIDTH-1:0] wire_d8_61;
	wire [WIDTH-1:0] wire_d8_62;
	wire [WIDTH-1:0] wire_d8_63;
	wire [WIDTH-1:0] wire_d8_64;
	wire [WIDTH-1:0] wire_d8_65;
	wire [WIDTH-1:0] wire_d8_66;
	wire [WIDTH-1:0] wire_d8_67;
	wire [WIDTH-1:0] wire_d8_68;
	wire [WIDTH-1:0] wire_d8_69;
	wire [WIDTH-1:0] wire_d8_70;
	wire [WIDTH-1:0] wire_d8_71;
	wire [WIDTH-1:0] wire_d8_72;
	wire [WIDTH-1:0] wire_d8_73;
	wire [WIDTH-1:0] wire_d8_74;
	wire [WIDTH-1:0] wire_d8_75;
	wire [WIDTH-1:0] wire_d8_76;
	wire [WIDTH-1:0] wire_d8_77;
	wire [WIDTH-1:0] wire_d8_78;
	wire [WIDTH-1:0] wire_d8_79;
	wire [WIDTH-1:0] wire_d8_80;
	wire [WIDTH-1:0] wire_d8_81;
	wire [WIDTH-1:0] wire_d8_82;
	wire [WIDTH-1:0] wire_d8_83;
	wire [WIDTH-1:0] wire_d8_84;
	wire [WIDTH-1:0] wire_d8_85;
	wire [WIDTH-1:0] wire_d8_86;
	wire [WIDTH-1:0] wire_d8_87;
	wire [WIDTH-1:0] wire_d8_88;
	wire [WIDTH-1:0] wire_d8_89;
	wire [WIDTH-1:0] wire_d8_90;
	wire [WIDTH-1:0] wire_d8_91;
	wire [WIDTH-1:0] wire_d8_92;
	wire [WIDTH-1:0] wire_d8_93;
	wire [WIDTH-1:0] wire_d8_94;
	wire [WIDTH-1:0] wire_d8_95;
	wire [WIDTH-1:0] wire_d8_96;
	wire [WIDTH-1:0] wire_d8_97;
	wire [WIDTH-1:0] wire_d8_98;
	wire [WIDTH-1:0] wire_d9_0;
	wire [WIDTH-1:0] wire_d9_1;
	wire [WIDTH-1:0] wire_d9_2;
	wire [WIDTH-1:0] wire_d9_3;
	wire [WIDTH-1:0] wire_d9_4;
	wire [WIDTH-1:0] wire_d9_5;
	wire [WIDTH-1:0] wire_d9_6;
	wire [WIDTH-1:0] wire_d9_7;
	wire [WIDTH-1:0] wire_d9_8;
	wire [WIDTH-1:0] wire_d9_9;
	wire [WIDTH-1:0] wire_d9_10;
	wire [WIDTH-1:0] wire_d9_11;
	wire [WIDTH-1:0] wire_d9_12;
	wire [WIDTH-1:0] wire_d9_13;
	wire [WIDTH-1:0] wire_d9_14;
	wire [WIDTH-1:0] wire_d9_15;
	wire [WIDTH-1:0] wire_d9_16;
	wire [WIDTH-1:0] wire_d9_17;
	wire [WIDTH-1:0] wire_d9_18;
	wire [WIDTH-1:0] wire_d9_19;
	wire [WIDTH-1:0] wire_d9_20;
	wire [WIDTH-1:0] wire_d9_21;
	wire [WIDTH-1:0] wire_d9_22;
	wire [WIDTH-1:0] wire_d9_23;
	wire [WIDTH-1:0] wire_d9_24;
	wire [WIDTH-1:0] wire_d9_25;
	wire [WIDTH-1:0] wire_d9_26;
	wire [WIDTH-1:0] wire_d9_27;
	wire [WIDTH-1:0] wire_d9_28;
	wire [WIDTH-1:0] wire_d9_29;
	wire [WIDTH-1:0] wire_d9_30;
	wire [WIDTH-1:0] wire_d9_31;
	wire [WIDTH-1:0] wire_d9_32;
	wire [WIDTH-1:0] wire_d9_33;
	wire [WIDTH-1:0] wire_d9_34;
	wire [WIDTH-1:0] wire_d9_35;
	wire [WIDTH-1:0] wire_d9_36;
	wire [WIDTH-1:0] wire_d9_37;
	wire [WIDTH-1:0] wire_d9_38;
	wire [WIDTH-1:0] wire_d9_39;
	wire [WIDTH-1:0] wire_d9_40;
	wire [WIDTH-1:0] wire_d9_41;
	wire [WIDTH-1:0] wire_d9_42;
	wire [WIDTH-1:0] wire_d9_43;
	wire [WIDTH-1:0] wire_d9_44;
	wire [WIDTH-1:0] wire_d9_45;
	wire [WIDTH-1:0] wire_d9_46;
	wire [WIDTH-1:0] wire_d9_47;
	wire [WIDTH-1:0] wire_d9_48;
	wire [WIDTH-1:0] wire_d9_49;
	wire [WIDTH-1:0] wire_d9_50;
	wire [WIDTH-1:0] wire_d9_51;
	wire [WIDTH-1:0] wire_d9_52;
	wire [WIDTH-1:0] wire_d9_53;
	wire [WIDTH-1:0] wire_d9_54;
	wire [WIDTH-1:0] wire_d9_55;
	wire [WIDTH-1:0] wire_d9_56;
	wire [WIDTH-1:0] wire_d9_57;
	wire [WIDTH-1:0] wire_d9_58;
	wire [WIDTH-1:0] wire_d9_59;
	wire [WIDTH-1:0] wire_d9_60;
	wire [WIDTH-1:0] wire_d9_61;
	wire [WIDTH-1:0] wire_d9_62;
	wire [WIDTH-1:0] wire_d9_63;
	wire [WIDTH-1:0] wire_d9_64;
	wire [WIDTH-1:0] wire_d9_65;
	wire [WIDTH-1:0] wire_d9_66;
	wire [WIDTH-1:0] wire_d9_67;
	wire [WIDTH-1:0] wire_d9_68;
	wire [WIDTH-1:0] wire_d9_69;
	wire [WIDTH-1:0] wire_d9_70;
	wire [WIDTH-1:0] wire_d9_71;
	wire [WIDTH-1:0] wire_d9_72;
	wire [WIDTH-1:0] wire_d9_73;
	wire [WIDTH-1:0] wire_d9_74;
	wire [WIDTH-1:0] wire_d9_75;
	wire [WIDTH-1:0] wire_d9_76;
	wire [WIDTH-1:0] wire_d9_77;
	wire [WIDTH-1:0] wire_d9_78;
	wire [WIDTH-1:0] wire_d9_79;
	wire [WIDTH-1:0] wire_d9_80;
	wire [WIDTH-1:0] wire_d9_81;
	wire [WIDTH-1:0] wire_d9_82;
	wire [WIDTH-1:0] wire_d9_83;
	wire [WIDTH-1:0] wire_d9_84;
	wire [WIDTH-1:0] wire_d9_85;
	wire [WIDTH-1:0] wire_d9_86;
	wire [WIDTH-1:0] wire_d9_87;
	wire [WIDTH-1:0] wire_d9_88;
	wire [WIDTH-1:0] wire_d9_89;
	wire [WIDTH-1:0] wire_d9_90;
	wire [WIDTH-1:0] wire_d9_91;
	wire [WIDTH-1:0] wire_d9_92;
	wire [WIDTH-1:0] wire_d9_93;
	wire [WIDTH-1:0] wire_d9_94;
	wire [WIDTH-1:0] wire_d9_95;
	wire [WIDTH-1:0] wire_d9_96;
	wire [WIDTH-1:0] wire_d9_97;
	wire [WIDTH-1:0] wire_d9_98;

	encoder #(.WIDTH(WIDTH)) encoder_instance100(.data_in(d_in0),.data_out(wire_d0_0),.clk(clk),.rst(rst));            //channel 1
	encoder #(.WIDTH(WIDTH)) encoder_instance101(.data_in(wire_d0_0),.data_out(wire_d0_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance102(.data_in(wire_d0_1),.data_out(wire_d0_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance103(.data_in(wire_d0_2),.data_out(wire_d0_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance104(.data_in(wire_d0_3),.data_out(wire_d0_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance105(.data_in(wire_d0_4),.data_out(wire_d0_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance106(.data_in(wire_d0_5),.data_out(wire_d0_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance107(.data_in(wire_d0_6),.data_out(wire_d0_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance108(.data_in(wire_d0_7),.data_out(wire_d0_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance109(.data_in(wire_d0_8),.data_out(wire_d0_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1010(.data_in(wire_d0_9),.data_out(wire_d0_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1011(.data_in(wire_d0_10),.data_out(wire_d0_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1012(.data_in(wire_d0_11),.data_out(wire_d0_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1013(.data_in(wire_d0_12),.data_out(wire_d0_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1014(.data_in(wire_d0_13),.data_out(wire_d0_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1015(.data_in(wire_d0_14),.data_out(wire_d0_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1016(.data_in(wire_d0_15),.data_out(wire_d0_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1017(.data_in(wire_d0_16),.data_out(wire_d0_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1018(.data_in(wire_d0_17),.data_out(wire_d0_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1019(.data_in(wire_d0_18),.data_out(wire_d0_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1020(.data_in(wire_d0_19),.data_out(wire_d0_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1021(.data_in(wire_d0_20),.data_out(wire_d0_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1022(.data_in(wire_d0_21),.data_out(wire_d0_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1023(.data_in(wire_d0_22),.data_out(wire_d0_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1024(.data_in(wire_d0_23),.data_out(wire_d0_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1025(.data_in(wire_d0_24),.data_out(wire_d0_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1026(.data_in(wire_d0_25),.data_out(wire_d0_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1027(.data_in(wire_d0_26),.data_out(wire_d0_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1028(.data_in(wire_d0_27),.data_out(wire_d0_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1029(.data_in(wire_d0_28),.data_out(wire_d0_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1030(.data_in(wire_d0_29),.data_out(wire_d0_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1031(.data_in(wire_d0_30),.data_out(wire_d0_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1032(.data_in(wire_d0_31),.data_out(wire_d0_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1033(.data_in(wire_d0_32),.data_out(wire_d0_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1034(.data_in(wire_d0_33),.data_out(wire_d0_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1035(.data_in(wire_d0_34),.data_out(wire_d0_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1036(.data_in(wire_d0_35),.data_out(wire_d0_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1037(.data_in(wire_d0_36),.data_out(wire_d0_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1038(.data_in(wire_d0_37),.data_out(wire_d0_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1039(.data_in(wire_d0_38),.data_out(wire_d0_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1040(.data_in(wire_d0_39),.data_out(wire_d0_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1041(.data_in(wire_d0_40),.data_out(wire_d0_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1042(.data_in(wire_d0_41),.data_out(wire_d0_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1043(.data_in(wire_d0_42),.data_out(wire_d0_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1044(.data_in(wire_d0_43),.data_out(wire_d0_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1045(.data_in(wire_d0_44),.data_out(wire_d0_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1046(.data_in(wire_d0_45),.data_out(wire_d0_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1047(.data_in(wire_d0_46),.data_out(wire_d0_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1048(.data_in(wire_d0_47),.data_out(wire_d0_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1049(.data_in(wire_d0_48),.data_out(wire_d0_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1050(.data_in(wire_d0_49),.data_out(wire_d0_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1051(.data_in(wire_d0_50),.data_out(wire_d0_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1052(.data_in(wire_d0_51),.data_out(wire_d0_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1053(.data_in(wire_d0_52),.data_out(wire_d0_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1054(.data_in(wire_d0_53),.data_out(wire_d0_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1055(.data_in(wire_d0_54),.data_out(wire_d0_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1056(.data_in(wire_d0_55),.data_out(wire_d0_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1057(.data_in(wire_d0_56),.data_out(wire_d0_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1058(.data_in(wire_d0_57),.data_out(wire_d0_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1059(.data_in(wire_d0_58),.data_out(wire_d0_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1060(.data_in(wire_d0_59),.data_out(wire_d0_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1061(.data_in(wire_d0_60),.data_out(wire_d0_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1062(.data_in(wire_d0_61),.data_out(wire_d0_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1063(.data_in(wire_d0_62),.data_out(wire_d0_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1064(.data_in(wire_d0_63),.data_out(wire_d0_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1065(.data_in(wire_d0_64),.data_out(wire_d0_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1066(.data_in(wire_d0_65),.data_out(wire_d0_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1067(.data_in(wire_d0_66),.data_out(wire_d0_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1068(.data_in(wire_d0_67),.data_out(wire_d0_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1069(.data_in(wire_d0_68),.data_out(wire_d0_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1070(.data_in(wire_d0_69),.data_out(wire_d0_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1071(.data_in(wire_d0_70),.data_out(wire_d0_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1072(.data_in(wire_d0_71),.data_out(wire_d0_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1073(.data_in(wire_d0_72),.data_out(wire_d0_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1074(.data_in(wire_d0_73),.data_out(wire_d0_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1075(.data_in(wire_d0_74),.data_out(wire_d0_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1076(.data_in(wire_d0_75),.data_out(wire_d0_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1077(.data_in(wire_d0_76),.data_out(wire_d0_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1078(.data_in(wire_d0_77),.data_out(wire_d0_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1079(.data_in(wire_d0_78),.data_out(wire_d0_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1080(.data_in(wire_d0_79),.data_out(wire_d0_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1081(.data_in(wire_d0_80),.data_out(wire_d0_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1082(.data_in(wire_d0_81),.data_out(wire_d0_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1083(.data_in(wire_d0_82),.data_out(wire_d0_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1084(.data_in(wire_d0_83),.data_out(wire_d0_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1085(.data_in(wire_d0_84),.data_out(wire_d0_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1086(.data_in(wire_d0_85),.data_out(wire_d0_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1087(.data_in(wire_d0_86),.data_out(wire_d0_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1088(.data_in(wire_d0_87),.data_out(wire_d0_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1089(.data_in(wire_d0_88),.data_out(wire_d0_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1090(.data_in(wire_d0_89),.data_out(wire_d0_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1091(.data_in(wire_d0_90),.data_out(wire_d0_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1092(.data_in(wire_d0_91),.data_out(wire_d0_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1093(.data_in(wire_d0_92),.data_out(wire_d0_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1094(.data_in(wire_d0_93),.data_out(wire_d0_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1095(.data_in(wire_d0_94),.data_out(wire_d0_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1096(.data_in(wire_d0_95),.data_out(wire_d0_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1097(.data_in(wire_d0_96),.data_out(wire_d0_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1098(.data_in(wire_d0_97),.data_out(wire_d0_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1099(.data_in(wire_d0_98),.data_out(d_out0),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance210(.data_in(d_in1),.data_out(wire_d1_0),.clk(clk),.rst(rst));            //channel 2
	encoder #(.WIDTH(WIDTH)) encoder_instance211(.data_in(wire_d1_0),.data_out(wire_d1_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212(.data_in(wire_d1_1),.data_out(wire_d1_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance213(.data_in(wire_d1_2),.data_out(wire_d1_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance214(.data_in(wire_d1_3),.data_out(wire_d1_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance215(.data_in(wire_d1_4),.data_out(wire_d1_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance216(.data_in(wire_d1_5),.data_out(wire_d1_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance217(.data_in(wire_d1_6),.data_out(wire_d1_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance218(.data_in(wire_d1_7),.data_out(wire_d1_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance219(.data_in(wire_d1_8),.data_out(wire_d1_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2110(.data_in(wire_d1_9),.data_out(wire_d1_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2111(.data_in(wire_d1_10),.data_out(wire_d1_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2112(.data_in(wire_d1_11),.data_out(wire_d1_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2113(.data_in(wire_d1_12),.data_out(wire_d1_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2114(.data_in(wire_d1_13),.data_out(wire_d1_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2115(.data_in(wire_d1_14),.data_out(wire_d1_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2116(.data_in(wire_d1_15),.data_out(wire_d1_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2117(.data_in(wire_d1_16),.data_out(wire_d1_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2118(.data_in(wire_d1_17),.data_out(wire_d1_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2119(.data_in(wire_d1_18),.data_out(wire_d1_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2120(.data_in(wire_d1_19),.data_out(wire_d1_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2121(.data_in(wire_d1_20),.data_out(wire_d1_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2122(.data_in(wire_d1_21),.data_out(wire_d1_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2123(.data_in(wire_d1_22),.data_out(wire_d1_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2124(.data_in(wire_d1_23),.data_out(wire_d1_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2125(.data_in(wire_d1_24),.data_out(wire_d1_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2126(.data_in(wire_d1_25),.data_out(wire_d1_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2127(.data_in(wire_d1_26),.data_out(wire_d1_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2128(.data_in(wire_d1_27),.data_out(wire_d1_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2129(.data_in(wire_d1_28),.data_out(wire_d1_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2130(.data_in(wire_d1_29),.data_out(wire_d1_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2131(.data_in(wire_d1_30),.data_out(wire_d1_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2132(.data_in(wire_d1_31),.data_out(wire_d1_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2133(.data_in(wire_d1_32),.data_out(wire_d1_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2134(.data_in(wire_d1_33),.data_out(wire_d1_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2135(.data_in(wire_d1_34),.data_out(wire_d1_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2136(.data_in(wire_d1_35),.data_out(wire_d1_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2137(.data_in(wire_d1_36),.data_out(wire_d1_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2138(.data_in(wire_d1_37),.data_out(wire_d1_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2139(.data_in(wire_d1_38),.data_out(wire_d1_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2140(.data_in(wire_d1_39),.data_out(wire_d1_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2141(.data_in(wire_d1_40),.data_out(wire_d1_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2142(.data_in(wire_d1_41),.data_out(wire_d1_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2143(.data_in(wire_d1_42),.data_out(wire_d1_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2144(.data_in(wire_d1_43),.data_out(wire_d1_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2145(.data_in(wire_d1_44),.data_out(wire_d1_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2146(.data_in(wire_d1_45),.data_out(wire_d1_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2147(.data_in(wire_d1_46),.data_out(wire_d1_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2148(.data_in(wire_d1_47),.data_out(wire_d1_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2149(.data_in(wire_d1_48),.data_out(wire_d1_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2150(.data_in(wire_d1_49),.data_out(wire_d1_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2151(.data_in(wire_d1_50),.data_out(wire_d1_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2152(.data_in(wire_d1_51),.data_out(wire_d1_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2153(.data_in(wire_d1_52),.data_out(wire_d1_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2154(.data_in(wire_d1_53),.data_out(wire_d1_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2155(.data_in(wire_d1_54),.data_out(wire_d1_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2156(.data_in(wire_d1_55),.data_out(wire_d1_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2157(.data_in(wire_d1_56),.data_out(wire_d1_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2158(.data_in(wire_d1_57),.data_out(wire_d1_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2159(.data_in(wire_d1_58),.data_out(wire_d1_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2160(.data_in(wire_d1_59),.data_out(wire_d1_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2161(.data_in(wire_d1_60),.data_out(wire_d1_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2162(.data_in(wire_d1_61),.data_out(wire_d1_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2163(.data_in(wire_d1_62),.data_out(wire_d1_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2164(.data_in(wire_d1_63),.data_out(wire_d1_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2165(.data_in(wire_d1_64),.data_out(wire_d1_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2166(.data_in(wire_d1_65),.data_out(wire_d1_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2167(.data_in(wire_d1_66),.data_out(wire_d1_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2168(.data_in(wire_d1_67),.data_out(wire_d1_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2169(.data_in(wire_d1_68),.data_out(wire_d1_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2170(.data_in(wire_d1_69),.data_out(wire_d1_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2171(.data_in(wire_d1_70),.data_out(wire_d1_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2172(.data_in(wire_d1_71),.data_out(wire_d1_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2173(.data_in(wire_d1_72),.data_out(wire_d1_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2174(.data_in(wire_d1_73),.data_out(wire_d1_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2175(.data_in(wire_d1_74),.data_out(wire_d1_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2176(.data_in(wire_d1_75),.data_out(wire_d1_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2177(.data_in(wire_d1_76),.data_out(wire_d1_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2178(.data_in(wire_d1_77),.data_out(wire_d1_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2179(.data_in(wire_d1_78),.data_out(wire_d1_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2180(.data_in(wire_d1_79),.data_out(wire_d1_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2181(.data_in(wire_d1_80),.data_out(wire_d1_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2182(.data_in(wire_d1_81),.data_out(wire_d1_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2183(.data_in(wire_d1_82),.data_out(wire_d1_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2184(.data_in(wire_d1_83),.data_out(wire_d1_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2185(.data_in(wire_d1_84),.data_out(wire_d1_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2186(.data_in(wire_d1_85),.data_out(wire_d1_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2187(.data_in(wire_d1_86),.data_out(wire_d1_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2188(.data_in(wire_d1_87),.data_out(wire_d1_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2189(.data_in(wire_d1_88),.data_out(wire_d1_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2190(.data_in(wire_d1_89),.data_out(wire_d1_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2191(.data_in(wire_d1_90),.data_out(wire_d1_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2192(.data_in(wire_d1_91),.data_out(wire_d1_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2193(.data_in(wire_d1_92),.data_out(wire_d1_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2194(.data_in(wire_d1_93),.data_out(wire_d1_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2195(.data_in(wire_d1_94),.data_out(wire_d1_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2196(.data_in(wire_d1_95),.data_out(wire_d1_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2197(.data_in(wire_d1_96),.data_out(wire_d1_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2198(.data_in(wire_d1_97),.data_out(wire_d1_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2199(.data_in(wire_d1_98),.data_out(d_out1),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance320(.data_in(d_in2),.data_out(wire_d2_0),.clk(clk),.rst(rst));            //channel 3
	encoder #(.WIDTH(WIDTH)) encoder_instance321(.data_in(wire_d2_0),.data_out(wire_d2_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance322(.data_in(wire_d2_1),.data_out(wire_d2_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance323(.data_in(wire_d2_2),.data_out(wire_d2_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance324(.data_in(wire_d2_3),.data_out(wire_d2_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance325(.data_in(wire_d2_4),.data_out(wire_d2_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance326(.data_in(wire_d2_5),.data_out(wire_d2_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance327(.data_in(wire_d2_6),.data_out(wire_d2_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance328(.data_in(wire_d2_7),.data_out(wire_d2_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance329(.data_in(wire_d2_8),.data_out(wire_d2_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3210(.data_in(wire_d2_9),.data_out(wire_d2_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3211(.data_in(wire_d2_10),.data_out(wire_d2_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3212(.data_in(wire_d2_11),.data_out(wire_d2_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3213(.data_in(wire_d2_12),.data_out(wire_d2_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3214(.data_in(wire_d2_13),.data_out(wire_d2_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3215(.data_in(wire_d2_14),.data_out(wire_d2_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3216(.data_in(wire_d2_15),.data_out(wire_d2_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3217(.data_in(wire_d2_16),.data_out(wire_d2_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3218(.data_in(wire_d2_17),.data_out(wire_d2_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3219(.data_in(wire_d2_18),.data_out(wire_d2_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3220(.data_in(wire_d2_19),.data_out(wire_d2_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3221(.data_in(wire_d2_20),.data_out(wire_d2_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3222(.data_in(wire_d2_21),.data_out(wire_d2_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3223(.data_in(wire_d2_22),.data_out(wire_d2_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3224(.data_in(wire_d2_23),.data_out(wire_d2_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3225(.data_in(wire_d2_24),.data_out(wire_d2_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3226(.data_in(wire_d2_25),.data_out(wire_d2_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3227(.data_in(wire_d2_26),.data_out(wire_d2_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3228(.data_in(wire_d2_27),.data_out(wire_d2_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3229(.data_in(wire_d2_28),.data_out(wire_d2_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3230(.data_in(wire_d2_29),.data_out(wire_d2_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3231(.data_in(wire_d2_30),.data_out(wire_d2_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3232(.data_in(wire_d2_31),.data_out(wire_d2_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3233(.data_in(wire_d2_32),.data_out(wire_d2_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3234(.data_in(wire_d2_33),.data_out(wire_d2_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3235(.data_in(wire_d2_34),.data_out(wire_d2_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3236(.data_in(wire_d2_35),.data_out(wire_d2_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3237(.data_in(wire_d2_36),.data_out(wire_d2_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3238(.data_in(wire_d2_37),.data_out(wire_d2_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3239(.data_in(wire_d2_38),.data_out(wire_d2_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3240(.data_in(wire_d2_39),.data_out(wire_d2_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3241(.data_in(wire_d2_40),.data_out(wire_d2_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3242(.data_in(wire_d2_41),.data_out(wire_d2_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3243(.data_in(wire_d2_42),.data_out(wire_d2_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3244(.data_in(wire_d2_43),.data_out(wire_d2_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3245(.data_in(wire_d2_44),.data_out(wire_d2_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3246(.data_in(wire_d2_45),.data_out(wire_d2_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3247(.data_in(wire_d2_46),.data_out(wire_d2_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3248(.data_in(wire_d2_47),.data_out(wire_d2_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3249(.data_in(wire_d2_48),.data_out(wire_d2_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3250(.data_in(wire_d2_49),.data_out(wire_d2_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3251(.data_in(wire_d2_50),.data_out(wire_d2_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3252(.data_in(wire_d2_51),.data_out(wire_d2_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3253(.data_in(wire_d2_52),.data_out(wire_d2_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3254(.data_in(wire_d2_53),.data_out(wire_d2_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3255(.data_in(wire_d2_54),.data_out(wire_d2_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3256(.data_in(wire_d2_55),.data_out(wire_d2_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3257(.data_in(wire_d2_56),.data_out(wire_d2_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3258(.data_in(wire_d2_57),.data_out(wire_d2_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3259(.data_in(wire_d2_58),.data_out(wire_d2_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3260(.data_in(wire_d2_59),.data_out(wire_d2_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3261(.data_in(wire_d2_60),.data_out(wire_d2_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3262(.data_in(wire_d2_61),.data_out(wire_d2_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3263(.data_in(wire_d2_62),.data_out(wire_d2_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3264(.data_in(wire_d2_63),.data_out(wire_d2_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3265(.data_in(wire_d2_64),.data_out(wire_d2_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3266(.data_in(wire_d2_65),.data_out(wire_d2_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3267(.data_in(wire_d2_66),.data_out(wire_d2_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3268(.data_in(wire_d2_67),.data_out(wire_d2_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3269(.data_in(wire_d2_68),.data_out(wire_d2_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3270(.data_in(wire_d2_69),.data_out(wire_d2_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3271(.data_in(wire_d2_70),.data_out(wire_d2_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3272(.data_in(wire_d2_71),.data_out(wire_d2_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3273(.data_in(wire_d2_72),.data_out(wire_d2_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3274(.data_in(wire_d2_73),.data_out(wire_d2_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3275(.data_in(wire_d2_74),.data_out(wire_d2_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3276(.data_in(wire_d2_75),.data_out(wire_d2_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3277(.data_in(wire_d2_76),.data_out(wire_d2_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3278(.data_in(wire_d2_77),.data_out(wire_d2_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3279(.data_in(wire_d2_78),.data_out(wire_d2_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3280(.data_in(wire_d2_79),.data_out(wire_d2_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3281(.data_in(wire_d2_80),.data_out(wire_d2_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3282(.data_in(wire_d2_81),.data_out(wire_d2_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3283(.data_in(wire_d2_82),.data_out(wire_d2_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3284(.data_in(wire_d2_83),.data_out(wire_d2_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3285(.data_in(wire_d2_84),.data_out(wire_d2_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3286(.data_in(wire_d2_85),.data_out(wire_d2_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3287(.data_in(wire_d2_86),.data_out(wire_d2_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3288(.data_in(wire_d2_87),.data_out(wire_d2_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3289(.data_in(wire_d2_88),.data_out(wire_d2_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3290(.data_in(wire_d2_89),.data_out(wire_d2_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3291(.data_in(wire_d2_90),.data_out(wire_d2_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3292(.data_in(wire_d2_91),.data_out(wire_d2_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3293(.data_in(wire_d2_92),.data_out(wire_d2_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3294(.data_in(wire_d2_93),.data_out(wire_d2_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3295(.data_in(wire_d2_94),.data_out(wire_d2_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3296(.data_in(wire_d2_95),.data_out(wire_d2_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3297(.data_in(wire_d2_96),.data_out(wire_d2_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3298(.data_in(wire_d2_97),.data_out(wire_d2_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3299(.data_in(wire_d2_98),.data_out(d_out2),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance430(.data_in(d_in3),.data_out(wire_d3_0),.clk(clk),.rst(rst));            //channel 4
	encoder #(.WIDTH(WIDTH)) encoder_instance431(.data_in(wire_d3_0),.data_out(wire_d3_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance432(.data_in(wire_d3_1),.data_out(wire_d3_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance433(.data_in(wire_d3_2),.data_out(wire_d3_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance434(.data_in(wire_d3_3),.data_out(wire_d3_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance435(.data_in(wire_d3_4),.data_out(wire_d3_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance436(.data_in(wire_d3_5),.data_out(wire_d3_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance437(.data_in(wire_d3_6),.data_out(wire_d3_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance438(.data_in(wire_d3_7),.data_out(wire_d3_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance439(.data_in(wire_d3_8),.data_out(wire_d3_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4310(.data_in(wire_d3_9),.data_out(wire_d3_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4311(.data_in(wire_d3_10),.data_out(wire_d3_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4312(.data_in(wire_d3_11),.data_out(wire_d3_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4313(.data_in(wire_d3_12),.data_out(wire_d3_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4314(.data_in(wire_d3_13),.data_out(wire_d3_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4315(.data_in(wire_d3_14),.data_out(wire_d3_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4316(.data_in(wire_d3_15),.data_out(wire_d3_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4317(.data_in(wire_d3_16),.data_out(wire_d3_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4318(.data_in(wire_d3_17),.data_out(wire_d3_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4319(.data_in(wire_d3_18),.data_out(wire_d3_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4320(.data_in(wire_d3_19),.data_out(wire_d3_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4321(.data_in(wire_d3_20),.data_out(wire_d3_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4322(.data_in(wire_d3_21),.data_out(wire_d3_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4323(.data_in(wire_d3_22),.data_out(wire_d3_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4324(.data_in(wire_d3_23),.data_out(wire_d3_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4325(.data_in(wire_d3_24),.data_out(wire_d3_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4326(.data_in(wire_d3_25),.data_out(wire_d3_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4327(.data_in(wire_d3_26),.data_out(wire_d3_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4328(.data_in(wire_d3_27),.data_out(wire_d3_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4329(.data_in(wire_d3_28),.data_out(wire_d3_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4330(.data_in(wire_d3_29),.data_out(wire_d3_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4331(.data_in(wire_d3_30),.data_out(wire_d3_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4332(.data_in(wire_d3_31),.data_out(wire_d3_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4333(.data_in(wire_d3_32),.data_out(wire_d3_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4334(.data_in(wire_d3_33),.data_out(wire_d3_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4335(.data_in(wire_d3_34),.data_out(wire_d3_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4336(.data_in(wire_d3_35),.data_out(wire_d3_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4337(.data_in(wire_d3_36),.data_out(wire_d3_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4338(.data_in(wire_d3_37),.data_out(wire_d3_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4339(.data_in(wire_d3_38),.data_out(wire_d3_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4340(.data_in(wire_d3_39),.data_out(wire_d3_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4341(.data_in(wire_d3_40),.data_out(wire_d3_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4342(.data_in(wire_d3_41),.data_out(wire_d3_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4343(.data_in(wire_d3_42),.data_out(wire_d3_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4344(.data_in(wire_d3_43),.data_out(wire_d3_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4345(.data_in(wire_d3_44),.data_out(wire_d3_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4346(.data_in(wire_d3_45),.data_out(wire_d3_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4347(.data_in(wire_d3_46),.data_out(wire_d3_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4348(.data_in(wire_d3_47),.data_out(wire_d3_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4349(.data_in(wire_d3_48),.data_out(wire_d3_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4350(.data_in(wire_d3_49),.data_out(wire_d3_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4351(.data_in(wire_d3_50),.data_out(wire_d3_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4352(.data_in(wire_d3_51),.data_out(wire_d3_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4353(.data_in(wire_d3_52),.data_out(wire_d3_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4354(.data_in(wire_d3_53),.data_out(wire_d3_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4355(.data_in(wire_d3_54),.data_out(wire_d3_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4356(.data_in(wire_d3_55),.data_out(wire_d3_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4357(.data_in(wire_d3_56),.data_out(wire_d3_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4358(.data_in(wire_d3_57),.data_out(wire_d3_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4359(.data_in(wire_d3_58),.data_out(wire_d3_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4360(.data_in(wire_d3_59),.data_out(wire_d3_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4361(.data_in(wire_d3_60),.data_out(wire_d3_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4362(.data_in(wire_d3_61),.data_out(wire_d3_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4363(.data_in(wire_d3_62),.data_out(wire_d3_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4364(.data_in(wire_d3_63),.data_out(wire_d3_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4365(.data_in(wire_d3_64),.data_out(wire_d3_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4366(.data_in(wire_d3_65),.data_out(wire_d3_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4367(.data_in(wire_d3_66),.data_out(wire_d3_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4368(.data_in(wire_d3_67),.data_out(wire_d3_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4369(.data_in(wire_d3_68),.data_out(wire_d3_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4370(.data_in(wire_d3_69),.data_out(wire_d3_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4371(.data_in(wire_d3_70),.data_out(wire_d3_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4372(.data_in(wire_d3_71),.data_out(wire_d3_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4373(.data_in(wire_d3_72),.data_out(wire_d3_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4374(.data_in(wire_d3_73),.data_out(wire_d3_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4375(.data_in(wire_d3_74),.data_out(wire_d3_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4376(.data_in(wire_d3_75),.data_out(wire_d3_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4377(.data_in(wire_d3_76),.data_out(wire_d3_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4378(.data_in(wire_d3_77),.data_out(wire_d3_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4379(.data_in(wire_d3_78),.data_out(wire_d3_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4380(.data_in(wire_d3_79),.data_out(wire_d3_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4381(.data_in(wire_d3_80),.data_out(wire_d3_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4382(.data_in(wire_d3_81),.data_out(wire_d3_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4383(.data_in(wire_d3_82),.data_out(wire_d3_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4384(.data_in(wire_d3_83),.data_out(wire_d3_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4385(.data_in(wire_d3_84),.data_out(wire_d3_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4386(.data_in(wire_d3_85),.data_out(wire_d3_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4387(.data_in(wire_d3_86),.data_out(wire_d3_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4388(.data_in(wire_d3_87),.data_out(wire_d3_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4389(.data_in(wire_d3_88),.data_out(wire_d3_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4390(.data_in(wire_d3_89),.data_out(wire_d3_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4391(.data_in(wire_d3_90),.data_out(wire_d3_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4392(.data_in(wire_d3_91),.data_out(wire_d3_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4393(.data_in(wire_d3_92),.data_out(wire_d3_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4394(.data_in(wire_d3_93),.data_out(wire_d3_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4395(.data_in(wire_d3_94),.data_out(wire_d3_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4396(.data_in(wire_d3_95),.data_out(wire_d3_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4397(.data_in(wire_d3_96),.data_out(wire_d3_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4398(.data_in(wire_d3_97),.data_out(wire_d3_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4399(.data_in(wire_d3_98),.data_out(d_out3),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance540(.data_in(d_in4),.data_out(wire_d4_0),.clk(clk),.rst(rst));            //channel 5
	encoder #(.WIDTH(WIDTH)) encoder_instance541(.data_in(wire_d4_0),.data_out(wire_d4_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance542(.data_in(wire_d4_1),.data_out(wire_d4_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance543(.data_in(wire_d4_2),.data_out(wire_d4_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance544(.data_in(wire_d4_3),.data_out(wire_d4_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance545(.data_in(wire_d4_4),.data_out(wire_d4_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance546(.data_in(wire_d4_5),.data_out(wire_d4_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance547(.data_in(wire_d4_6),.data_out(wire_d4_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance548(.data_in(wire_d4_7),.data_out(wire_d4_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance549(.data_in(wire_d4_8),.data_out(wire_d4_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5410(.data_in(wire_d4_9),.data_out(wire_d4_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5411(.data_in(wire_d4_10),.data_out(wire_d4_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5412(.data_in(wire_d4_11),.data_out(wire_d4_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5413(.data_in(wire_d4_12),.data_out(wire_d4_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5414(.data_in(wire_d4_13),.data_out(wire_d4_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5415(.data_in(wire_d4_14),.data_out(wire_d4_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5416(.data_in(wire_d4_15),.data_out(wire_d4_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5417(.data_in(wire_d4_16),.data_out(wire_d4_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5418(.data_in(wire_d4_17),.data_out(wire_d4_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5419(.data_in(wire_d4_18),.data_out(wire_d4_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5420(.data_in(wire_d4_19),.data_out(wire_d4_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5421(.data_in(wire_d4_20),.data_out(wire_d4_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5422(.data_in(wire_d4_21),.data_out(wire_d4_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5423(.data_in(wire_d4_22),.data_out(wire_d4_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5424(.data_in(wire_d4_23),.data_out(wire_d4_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5425(.data_in(wire_d4_24),.data_out(wire_d4_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5426(.data_in(wire_d4_25),.data_out(wire_d4_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5427(.data_in(wire_d4_26),.data_out(wire_d4_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5428(.data_in(wire_d4_27),.data_out(wire_d4_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5429(.data_in(wire_d4_28),.data_out(wire_d4_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5430(.data_in(wire_d4_29),.data_out(wire_d4_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5431(.data_in(wire_d4_30),.data_out(wire_d4_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5432(.data_in(wire_d4_31),.data_out(wire_d4_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5433(.data_in(wire_d4_32),.data_out(wire_d4_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5434(.data_in(wire_d4_33),.data_out(wire_d4_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5435(.data_in(wire_d4_34),.data_out(wire_d4_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5436(.data_in(wire_d4_35),.data_out(wire_d4_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5437(.data_in(wire_d4_36),.data_out(wire_d4_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5438(.data_in(wire_d4_37),.data_out(wire_d4_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5439(.data_in(wire_d4_38),.data_out(wire_d4_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5440(.data_in(wire_d4_39),.data_out(wire_d4_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5441(.data_in(wire_d4_40),.data_out(wire_d4_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5442(.data_in(wire_d4_41),.data_out(wire_d4_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5443(.data_in(wire_d4_42),.data_out(wire_d4_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5444(.data_in(wire_d4_43),.data_out(wire_d4_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5445(.data_in(wire_d4_44),.data_out(wire_d4_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5446(.data_in(wire_d4_45),.data_out(wire_d4_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5447(.data_in(wire_d4_46),.data_out(wire_d4_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5448(.data_in(wire_d4_47),.data_out(wire_d4_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5449(.data_in(wire_d4_48),.data_out(wire_d4_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5450(.data_in(wire_d4_49),.data_out(wire_d4_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5451(.data_in(wire_d4_50),.data_out(wire_d4_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5452(.data_in(wire_d4_51),.data_out(wire_d4_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5453(.data_in(wire_d4_52),.data_out(wire_d4_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5454(.data_in(wire_d4_53),.data_out(wire_d4_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5455(.data_in(wire_d4_54),.data_out(wire_d4_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5456(.data_in(wire_d4_55),.data_out(wire_d4_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5457(.data_in(wire_d4_56),.data_out(wire_d4_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5458(.data_in(wire_d4_57),.data_out(wire_d4_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5459(.data_in(wire_d4_58),.data_out(wire_d4_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5460(.data_in(wire_d4_59),.data_out(wire_d4_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5461(.data_in(wire_d4_60),.data_out(wire_d4_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5462(.data_in(wire_d4_61),.data_out(wire_d4_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5463(.data_in(wire_d4_62),.data_out(wire_d4_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5464(.data_in(wire_d4_63),.data_out(wire_d4_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5465(.data_in(wire_d4_64),.data_out(wire_d4_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5466(.data_in(wire_d4_65),.data_out(wire_d4_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5467(.data_in(wire_d4_66),.data_out(wire_d4_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5468(.data_in(wire_d4_67),.data_out(wire_d4_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5469(.data_in(wire_d4_68),.data_out(wire_d4_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5470(.data_in(wire_d4_69),.data_out(wire_d4_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5471(.data_in(wire_d4_70),.data_out(wire_d4_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5472(.data_in(wire_d4_71),.data_out(wire_d4_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5473(.data_in(wire_d4_72),.data_out(wire_d4_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5474(.data_in(wire_d4_73),.data_out(wire_d4_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5475(.data_in(wire_d4_74),.data_out(wire_d4_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5476(.data_in(wire_d4_75),.data_out(wire_d4_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5477(.data_in(wire_d4_76),.data_out(wire_d4_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5478(.data_in(wire_d4_77),.data_out(wire_d4_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5479(.data_in(wire_d4_78),.data_out(wire_d4_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5480(.data_in(wire_d4_79),.data_out(wire_d4_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5481(.data_in(wire_d4_80),.data_out(wire_d4_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5482(.data_in(wire_d4_81),.data_out(wire_d4_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5483(.data_in(wire_d4_82),.data_out(wire_d4_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5484(.data_in(wire_d4_83),.data_out(wire_d4_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5485(.data_in(wire_d4_84),.data_out(wire_d4_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5486(.data_in(wire_d4_85),.data_out(wire_d4_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5487(.data_in(wire_d4_86),.data_out(wire_d4_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5488(.data_in(wire_d4_87),.data_out(wire_d4_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5489(.data_in(wire_d4_88),.data_out(wire_d4_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5490(.data_in(wire_d4_89),.data_out(wire_d4_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5491(.data_in(wire_d4_90),.data_out(wire_d4_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5492(.data_in(wire_d4_91),.data_out(wire_d4_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5493(.data_in(wire_d4_92),.data_out(wire_d4_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5494(.data_in(wire_d4_93),.data_out(wire_d4_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5495(.data_in(wire_d4_94),.data_out(wire_d4_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5496(.data_in(wire_d4_95),.data_out(wire_d4_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5497(.data_in(wire_d4_96),.data_out(wire_d4_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5498(.data_in(wire_d4_97),.data_out(wire_d4_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5499(.data_in(wire_d4_98),.data_out(d_out4),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance650(.data_in(d_in5),.data_out(wire_d5_0),.clk(clk),.rst(rst));            //channel 6
	encoder #(.WIDTH(WIDTH)) encoder_instance651(.data_in(wire_d5_0),.data_out(wire_d5_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance652(.data_in(wire_d5_1),.data_out(wire_d5_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance653(.data_in(wire_d5_2),.data_out(wire_d5_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance654(.data_in(wire_d5_3),.data_out(wire_d5_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance655(.data_in(wire_d5_4),.data_out(wire_d5_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance656(.data_in(wire_d5_5),.data_out(wire_d5_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance657(.data_in(wire_d5_6),.data_out(wire_d5_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance658(.data_in(wire_d5_7),.data_out(wire_d5_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance659(.data_in(wire_d5_8),.data_out(wire_d5_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6510(.data_in(wire_d5_9),.data_out(wire_d5_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6511(.data_in(wire_d5_10),.data_out(wire_d5_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6512(.data_in(wire_d5_11),.data_out(wire_d5_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6513(.data_in(wire_d5_12),.data_out(wire_d5_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6514(.data_in(wire_d5_13),.data_out(wire_d5_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6515(.data_in(wire_d5_14),.data_out(wire_d5_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6516(.data_in(wire_d5_15),.data_out(wire_d5_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6517(.data_in(wire_d5_16),.data_out(wire_d5_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6518(.data_in(wire_d5_17),.data_out(wire_d5_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6519(.data_in(wire_d5_18),.data_out(wire_d5_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6520(.data_in(wire_d5_19),.data_out(wire_d5_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6521(.data_in(wire_d5_20),.data_out(wire_d5_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6522(.data_in(wire_d5_21),.data_out(wire_d5_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6523(.data_in(wire_d5_22),.data_out(wire_d5_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6524(.data_in(wire_d5_23),.data_out(wire_d5_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6525(.data_in(wire_d5_24),.data_out(wire_d5_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6526(.data_in(wire_d5_25),.data_out(wire_d5_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6527(.data_in(wire_d5_26),.data_out(wire_d5_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6528(.data_in(wire_d5_27),.data_out(wire_d5_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6529(.data_in(wire_d5_28),.data_out(wire_d5_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6530(.data_in(wire_d5_29),.data_out(wire_d5_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6531(.data_in(wire_d5_30),.data_out(wire_d5_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6532(.data_in(wire_d5_31),.data_out(wire_d5_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6533(.data_in(wire_d5_32),.data_out(wire_d5_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6534(.data_in(wire_d5_33),.data_out(wire_d5_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6535(.data_in(wire_d5_34),.data_out(wire_d5_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6536(.data_in(wire_d5_35),.data_out(wire_d5_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6537(.data_in(wire_d5_36),.data_out(wire_d5_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6538(.data_in(wire_d5_37),.data_out(wire_d5_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6539(.data_in(wire_d5_38),.data_out(wire_d5_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6540(.data_in(wire_d5_39),.data_out(wire_d5_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6541(.data_in(wire_d5_40),.data_out(wire_d5_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6542(.data_in(wire_d5_41),.data_out(wire_d5_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6543(.data_in(wire_d5_42),.data_out(wire_d5_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6544(.data_in(wire_d5_43),.data_out(wire_d5_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6545(.data_in(wire_d5_44),.data_out(wire_d5_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6546(.data_in(wire_d5_45),.data_out(wire_d5_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6547(.data_in(wire_d5_46),.data_out(wire_d5_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6548(.data_in(wire_d5_47),.data_out(wire_d5_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6549(.data_in(wire_d5_48),.data_out(wire_d5_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6550(.data_in(wire_d5_49),.data_out(wire_d5_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6551(.data_in(wire_d5_50),.data_out(wire_d5_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6552(.data_in(wire_d5_51),.data_out(wire_d5_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6553(.data_in(wire_d5_52),.data_out(wire_d5_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6554(.data_in(wire_d5_53),.data_out(wire_d5_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6555(.data_in(wire_d5_54),.data_out(wire_d5_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6556(.data_in(wire_d5_55),.data_out(wire_d5_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6557(.data_in(wire_d5_56),.data_out(wire_d5_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6558(.data_in(wire_d5_57),.data_out(wire_d5_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6559(.data_in(wire_d5_58),.data_out(wire_d5_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6560(.data_in(wire_d5_59),.data_out(wire_d5_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6561(.data_in(wire_d5_60),.data_out(wire_d5_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6562(.data_in(wire_d5_61),.data_out(wire_d5_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6563(.data_in(wire_d5_62),.data_out(wire_d5_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6564(.data_in(wire_d5_63),.data_out(wire_d5_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6565(.data_in(wire_d5_64),.data_out(wire_d5_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6566(.data_in(wire_d5_65),.data_out(wire_d5_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6567(.data_in(wire_d5_66),.data_out(wire_d5_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6568(.data_in(wire_d5_67),.data_out(wire_d5_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6569(.data_in(wire_d5_68),.data_out(wire_d5_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6570(.data_in(wire_d5_69),.data_out(wire_d5_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6571(.data_in(wire_d5_70),.data_out(wire_d5_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6572(.data_in(wire_d5_71),.data_out(wire_d5_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6573(.data_in(wire_d5_72),.data_out(wire_d5_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6574(.data_in(wire_d5_73),.data_out(wire_d5_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6575(.data_in(wire_d5_74),.data_out(wire_d5_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6576(.data_in(wire_d5_75),.data_out(wire_d5_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6577(.data_in(wire_d5_76),.data_out(wire_d5_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6578(.data_in(wire_d5_77),.data_out(wire_d5_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6579(.data_in(wire_d5_78),.data_out(wire_d5_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6580(.data_in(wire_d5_79),.data_out(wire_d5_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6581(.data_in(wire_d5_80),.data_out(wire_d5_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6582(.data_in(wire_d5_81),.data_out(wire_d5_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6583(.data_in(wire_d5_82),.data_out(wire_d5_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6584(.data_in(wire_d5_83),.data_out(wire_d5_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6585(.data_in(wire_d5_84),.data_out(wire_d5_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6586(.data_in(wire_d5_85),.data_out(wire_d5_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6587(.data_in(wire_d5_86),.data_out(wire_d5_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6588(.data_in(wire_d5_87),.data_out(wire_d5_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6589(.data_in(wire_d5_88),.data_out(wire_d5_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6590(.data_in(wire_d5_89),.data_out(wire_d5_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6591(.data_in(wire_d5_90),.data_out(wire_d5_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6592(.data_in(wire_d5_91),.data_out(wire_d5_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6593(.data_in(wire_d5_92),.data_out(wire_d5_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6594(.data_in(wire_d5_93),.data_out(wire_d5_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6595(.data_in(wire_d5_94),.data_out(wire_d5_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6596(.data_in(wire_d5_95),.data_out(wire_d5_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6597(.data_in(wire_d5_96),.data_out(wire_d5_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6598(.data_in(wire_d5_97),.data_out(wire_d5_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6599(.data_in(wire_d5_98),.data_out(d_out5),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance760(.data_in(d_in6),.data_out(wire_d6_0),.clk(clk),.rst(rst));            //channel 7
	encoder #(.WIDTH(WIDTH)) encoder_instance761(.data_in(wire_d6_0),.data_out(wire_d6_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance762(.data_in(wire_d6_1),.data_out(wire_d6_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance763(.data_in(wire_d6_2),.data_out(wire_d6_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance764(.data_in(wire_d6_3),.data_out(wire_d6_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance765(.data_in(wire_d6_4),.data_out(wire_d6_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance766(.data_in(wire_d6_5),.data_out(wire_d6_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance767(.data_in(wire_d6_6),.data_out(wire_d6_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance768(.data_in(wire_d6_7),.data_out(wire_d6_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance769(.data_in(wire_d6_8),.data_out(wire_d6_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7610(.data_in(wire_d6_9),.data_out(wire_d6_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7611(.data_in(wire_d6_10),.data_out(wire_d6_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7612(.data_in(wire_d6_11),.data_out(wire_d6_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7613(.data_in(wire_d6_12),.data_out(wire_d6_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7614(.data_in(wire_d6_13),.data_out(wire_d6_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7615(.data_in(wire_d6_14),.data_out(wire_d6_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7616(.data_in(wire_d6_15),.data_out(wire_d6_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7617(.data_in(wire_d6_16),.data_out(wire_d6_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7618(.data_in(wire_d6_17),.data_out(wire_d6_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7619(.data_in(wire_d6_18),.data_out(wire_d6_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7620(.data_in(wire_d6_19),.data_out(wire_d6_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7621(.data_in(wire_d6_20),.data_out(wire_d6_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7622(.data_in(wire_d6_21),.data_out(wire_d6_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7623(.data_in(wire_d6_22),.data_out(wire_d6_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7624(.data_in(wire_d6_23),.data_out(wire_d6_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7625(.data_in(wire_d6_24),.data_out(wire_d6_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7626(.data_in(wire_d6_25),.data_out(wire_d6_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7627(.data_in(wire_d6_26),.data_out(wire_d6_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7628(.data_in(wire_d6_27),.data_out(wire_d6_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7629(.data_in(wire_d6_28),.data_out(wire_d6_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7630(.data_in(wire_d6_29),.data_out(wire_d6_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7631(.data_in(wire_d6_30),.data_out(wire_d6_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7632(.data_in(wire_d6_31),.data_out(wire_d6_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7633(.data_in(wire_d6_32),.data_out(wire_d6_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7634(.data_in(wire_d6_33),.data_out(wire_d6_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7635(.data_in(wire_d6_34),.data_out(wire_d6_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7636(.data_in(wire_d6_35),.data_out(wire_d6_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7637(.data_in(wire_d6_36),.data_out(wire_d6_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7638(.data_in(wire_d6_37),.data_out(wire_d6_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7639(.data_in(wire_d6_38),.data_out(wire_d6_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7640(.data_in(wire_d6_39),.data_out(wire_d6_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7641(.data_in(wire_d6_40),.data_out(wire_d6_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7642(.data_in(wire_d6_41),.data_out(wire_d6_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7643(.data_in(wire_d6_42),.data_out(wire_d6_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7644(.data_in(wire_d6_43),.data_out(wire_d6_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7645(.data_in(wire_d6_44),.data_out(wire_d6_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7646(.data_in(wire_d6_45),.data_out(wire_d6_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7647(.data_in(wire_d6_46),.data_out(wire_d6_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7648(.data_in(wire_d6_47),.data_out(wire_d6_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7649(.data_in(wire_d6_48),.data_out(wire_d6_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7650(.data_in(wire_d6_49),.data_out(wire_d6_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7651(.data_in(wire_d6_50),.data_out(wire_d6_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7652(.data_in(wire_d6_51),.data_out(wire_d6_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7653(.data_in(wire_d6_52),.data_out(wire_d6_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7654(.data_in(wire_d6_53),.data_out(wire_d6_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7655(.data_in(wire_d6_54),.data_out(wire_d6_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7656(.data_in(wire_d6_55),.data_out(wire_d6_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7657(.data_in(wire_d6_56),.data_out(wire_d6_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7658(.data_in(wire_d6_57),.data_out(wire_d6_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7659(.data_in(wire_d6_58),.data_out(wire_d6_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7660(.data_in(wire_d6_59),.data_out(wire_d6_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7661(.data_in(wire_d6_60),.data_out(wire_d6_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7662(.data_in(wire_d6_61),.data_out(wire_d6_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7663(.data_in(wire_d6_62),.data_out(wire_d6_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7664(.data_in(wire_d6_63),.data_out(wire_d6_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7665(.data_in(wire_d6_64),.data_out(wire_d6_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7666(.data_in(wire_d6_65),.data_out(wire_d6_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7667(.data_in(wire_d6_66),.data_out(wire_d6_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7668(.data_in(wire_d6_67),.data_out(wire_d6_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7669(.data_in(wire_d6_68),.data_out(wire_d6_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7670(.data_in(wire_d6_69),.data_out(wire_d6_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7671(.data_in(wire_d6_70),.data_out(wire_d6_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7672(.data_in(wire_d6_71),.data_out(wire_d6_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7673(.data_in(wire_d6_72),.data_out(wire_d6_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7674(.data_in(wire_d6_73),.data_out(wire_d6_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7675(.data_in(wire_d6_74),.data_out(wire_d6_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7676(.data_in(wire_d6_75),.data_out(wire_d6_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7677(.data_in(wire_d6_76),.data_out(wire_d6_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7678(.data_in(wire_d6_77),.data_out(wire_d6_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7679(.data_in(wire_d6_78),.data_out(wire_d6_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7680(.data_in(wire_d6_79),.data_out(wire_d6_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7681(.data_in(wire_d6_80),.data_out(wire_d6_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7682(.data_in(wire_d6_81),.data_out(wire_d6_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7683(.data_in(wire_d6_82),.data_out(wire_d6_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7684(.data_in(wire_d6_83),.data_out(wire_d6_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7685(.data_in(wire_d6_84),.data_out(wire_d6_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7686(.data_in(wire_d6_85),.data_out(wire_d6_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7687(.data_in(wire_d6_86),.data_out(wire_d6_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7688(.data_in(wire_d6_87),.data_out(wire_d6_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7689(.data_in(wire_d6_88),.data_out(wire_d6_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7690(.data_in(wire_d6_89),.data_out(wire_d6_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7691(.data_in(wire_d6_90),.data_out(wire_d6_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7692(.data_in(wire_d6_91),.data_out(wire_d6_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7693(.data_in(wire_d6_92),.data_out(wire_d6_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7694(.data_in(wire_d6_93),.data_out(wire_d6_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7695(.data_in(wire_d6_94),.data_out(wire_d6_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7696(.data_in(wire_d6_95),.data_out(wire_d6_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7697(.data_in(wire_d6_96),.data_out(wire_d6_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7698(.data_in(wire_d6_97),.data_out(wire_d6_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7699(.data_in(wire_d6_98),.data_out(d_out6),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance870(.data_in(d_in7),.data_out(wire_d7_0),.clk(clk),.rst(rst));            //channel 8
	encoder #(.WIDTH(WIDTH)) encoder_instance871(.data_in(wire_d7_0),.data_out(wire_d7_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance872(.data_in(wire_d7_1),.data_out(wire_d7_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance873(.data_in(wire_d7_2),.data_out(wire_d7_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance874(.data_in(wire_d7_3),.data_out(wire_d7_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance875(.data_in(wire_d7_4),.data_out(wire_d7_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance876(.data_in(wire_d7_5),.data_out(wire_d7_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance877(.data_in(wire_d7_6),.data_out(wire_d7_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance878(.data_in(wire_d7_7),.data_out(wire_d7_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance879(.data_in(wire_d7_8),.data_out(wire_d7_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8710(.data_in(wire_d7_9),.data_out(wire_d7_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8711(.data_in(wire_d7_10),.data_out(wire_d7_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8712(.data_in(wire_d7_11),.data_out(wire_d7_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8713(.data_in(wire_d7_12),.data_out(wire_d7_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8714(.data_in(wire_d7_13),.data_out(wire_d7_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8715(.data_in(wire_d7_14),.data_out(wire_d7_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8716(.data_in(wire_d7_15),.data_out(wire_d7_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8717(.data_in(wire_d7_16),.data_out(wire_d7_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8718(.data_in(wire_d7_17),.data_out(wire_d7_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8719(.data_in(wire_d7_18),.data_out(wire_d7_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8720(.data_in(wire_d7_19),.data_out(wire_d7_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8721(.data_in(wire_d7_20),.data_out(wire_d7_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8722(.data_in(wire_d7_21),.data_out(wire_d7_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8723(.data_in(wire_d7_22),.data_out(wire_d7_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8724(.data_in(wire_d7_23),.data_out(wire_d7_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8725(.data_in(wire_d7_24),.data_out(wire_d7_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8726(.data_in(wire_d7_25),.data_out(wire_d7_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8727(.data_in(wire_d7_26),.data_out(wire_d7_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8728(.data_in(wire_d7_27),.data_out(wire_d7_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8729(.data_in(wire_d7_28),.data_out(wire_d7_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8730(.data_in(wire_d7_29),.data_out(wire_d7_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8731(.data_in(wire_d7_30),.data_out(wire_d7_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8732(.data_in(wire_d7_31),.data_out(wire_d7_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8733(.data_in(wire_d7_32),.data_out(wire_d7_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8734(.data_in(wire_d7_33),.data_out(wire_d7_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8735(.data_in(wire_d7_34),.data_out(wire_d7_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8736(.data_in(wire_d7_35),.data_out(wire_d7_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8737(.data_in(wire_d7_36),.data_out(wire_d7_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8738(.data_in(wire_d7_37),.data_out(wire_d7_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8739(.data_in(wire_d7_38),.data_out(wire_d7_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8740(.data_in(wire_d7_39),.data_out(wire_d7_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8741(.data_in(wire_d7_40),.data_out(wire_d7_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8742(.data_in(wire_d7_41),.data_out(wire_d7_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8743(.data_in(wire_d7_42),.data_out(wire_d7_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8744(.data_in(wire_d7_43),.data_out(wire_d7_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8745(.data_in(wire_d7_44),.data_out(wire_d7_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8746(.data_in(wire_d7_45),.data_out(wire_d7_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8747(.data_in(wire_d7_46),.data_out(wire_d7_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8748(.data_in(wire_d7_47),.data_out(wire_d7_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8749(.data_in(wire_d7_48),.data_out(wire_d7_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8750(.data_in(wire_d7_49),.data_out(wire_d7_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8751(.data_in(wire_d7_50),.data_out(wire_d7_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8752(.data_in(wire_d7_51),.data_out(wire_d7_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8753(.data_in(wire_d7_52),.data_out(wire_d7_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8754(.data_in(wire_d7_53),.data_out(wire_d7_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8755(.data_in(wire_d7_54),.data_out(wire_d7_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8756(.data_in(wire_d7_55),.data_out(wire_d7_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8757(.data_in(wire_d7_56),.data_out(wire_d7_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8758(.data_in(wire_d7_57),.data_out(wire_d7_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8759(.data_in(wire_d7_58),.data_out(wire_d7_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8760(.data_in(wire_d7_59),.data_out(wire_d7_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8761(.data_in(wire_d7_60),.data_out(wire_d7_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8762(.data_in(wire_d7_61),.data_out(wire_d7_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8763(.data_in(wire_d7_62),.data_out(wire_d7_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8764(.data_in(wire_d7_63),.data_out(wire_d7_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8765(.data_in(wire_d7_64),.data_out(wire_d7_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8766(.data_in(wire_d7_65),.data_out(wire_d7_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8767(.data_in(wire_d7_66),.data_out(wire_d7_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8768(.data_in(wire_d7_67),.data_out(wire_d7_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8769(.data_in(wire_d7_68),.data_out(wire_d7_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8770(.data_in(wire_d7_69),.data_out(wire_d7_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8771(.data_in(wire_d7_70),.data_out(wire_d7_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8772(.data_in(wire_d7_71),.data_out(wire_d7_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8773(.data_in(wire_d7_72),.data_out(wire_d7_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8774(.data_in(wire_d7_73),.data_out(wire_d7_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8775(.data_in(wire_d7_74),.data_out(wire_d7_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8776(.data_in(wire_d7_75),.data_out(wire_d7_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8777(.data_in(wire_d7_76),.data_out(wire_d7_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8778(.data_in(wire_d7_77),.data_out(wire_d7_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8779(.data_in(wire_d7_78),.data_out(wire_d7_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8780(.data_in(wire_d7_79),.data_out(wire_d7_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8781(.data_in(wire_d7_80),.data_out(wire_d7_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8782(.data_in(wire_d7_81),.data_out(wire_d7_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8783(.data_in(wire_d7_82),.data_out(wire_d7_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8784(.data_in(wire_d7_83),.data_out(wire_d7_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8785(.data_in(wire_d7_84),.data_out(wire_d7_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8786(.data_in(wire_d7_85),.data_out(wire_d7_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8787(.data_in(wire_d7_86),.data_out(wire_d7_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8788(.data_in(wire_d7_87),.data_out(wire_d7_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8789(.data_in(wire_d7_88),.data_out(wire_d7_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8790(.data_in(wire_d7_89),.data_out(wire_d7_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8791(.data_in(wire_d7_90),.data_out(wire_d7_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8792(.data_in(wire_d7_91),.data_out(wire_d7_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8793(.data_in(wire_d7_92),.data_out(wire_d7_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8794(.data_in(wire_d7_93),.data_out(wire_d7_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8795(.data_in(wire_d7_94),.data_out(wire_d7_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8796(.data_in(wire_d7_95),.data_out(wire_d7_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8797(.data_in(wire_d7_96),.data_out(wire_d7_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8798(.data_in(wire_d7_97),.data_out(wire_d7_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8799(.data_in(wire_d7_98),.data_out(d_out7),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance980(.data_in(d_in8),.data_out(wire_d8_0),.clk(clk),.rst(rst));            //channel 9
	encoder #(.WIDTH(WIDTH)) encoder_instance981(.data_in(wire_d8_0),.data_out(wire_d8_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance982(.data_in(wire_d8_1),.data_out(wire_d8_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance983(.data_in(wire_d8_2),.data_out(wire_d8_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance984(.data_in(wire_d8_3),.data_out(wire_d8_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance985(.data_in(wire_d8_4),.data_out(wire_d8_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance986(.data_in(wire_d8_5),.data_out(wire_d8_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance987(.data_in(wire_d8_6),.data_out(wire_d8_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance988(.data_in(wire_d8_7),.data_out(wire_d8_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance989(.data_in(wire_d8_8),.data_out(wire_d8_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9810(.data_in(wire_d8_9),.data_out(wire_d8_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9811(.data_in(wire_d8_10),.data_out(wire_d8_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9812(.data_in(wire_d8_11),.data_out(wire_d8_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9813(.data_in(wire_d8_12),.data_out(wire_d8_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9814(.data_in(wire_d8_13),.data_out(wire_d8_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9815(.data_in(wire_d8_14),.data_out(wire_d8_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9816(.data_in(wire_d8_15),.data_out(wire_d8_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9817(.data_in(wire_d8_16),.data_out(wire_d8_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9818(.data_in(wire_d8_17),.data_out(wire_d8_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9819(.data_in(wire_d8_18),.data_out(wire_d8_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9820(.data_in(wire_d8_19),.data_out(wire_d8_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9821(.data_in(wire_d8_20),.data_out(wire_d8_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9822(.data_in(wire_d8_21),.data_out(wire_d8_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9823(.data_in(wire_d8_22),.data_out(wire_d8_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9824(.data_in(wire_d8_23),.data_out(wire_d8_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9825(.data_in(wire_d8_24),.data_out(wire_d8_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9826(.data_in(wire_d8_25),.data_out(wire_d8_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9827(.data_in(wire_d8_26),.data_out(wire_d8_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9828(.data_in(wire_d8_27),.data_out(wire_d8_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9829(.data_in(wire_d8_28),.data_out(wire_d8_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9830(.data_in(wire_d8_29),.data_out(wire_d8_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9831(.data_in(wire_d8_30),.data_out(wire_d8_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9832(.data_in(wire_d8_31),.data_out(wire_d8_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9833(.data_in(wire_d8_32),.data_out(wire_d8_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9834(.data_in(wire_d8_33),.data_out(wire_d8_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9835(.data_in(wire_d8_34),.data_out(wire_d8_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9836(.data_in(wire_d8_35),.data_out(wire_d8_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9837(.data_in(wire_d8_36),.data_out(wire_d8_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9838(.data_in(wire_d8_37),.data_out(wire_d8_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9839(.data_in(wire_d8_38),.data_out(wire_d8_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9840(.data_in(wire_d8_39),.data_out(wire_d8_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9841(.data_in(wire_d8_40),.data_out(wire_d8_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9842(.data_in(wire_d8_41),.data_out(wire_d8_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9843(.data_in(wire_d8_42),.data_out(wire_d8_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9844(.data_in(wire_d8_43),.data_out(wire_d8_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9845(.data_in(wire_d8_44),.data_out(wire_d8_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9846(.data_in(wire_d8_45),.data_out(wire_d8_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9847(.data_in(wire_d8_46),.data_out(wire_d8_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9848(.data_in(wire_d8_47),.data_out(wire_d8_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9849(.data_in(wire_d8_48),.data_out(wire_d8_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9850(.data_in(wire_d8_49),.data_out(wire_d8_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9851(.data_in(wire_d8_50),.data_out(wire_d8_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9852(.data_in(wire_d8_51),.data_out(wire_d8_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9853(.data_in(wire_d8_52),.data_out(wire_d8_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9854(.data_in(wire_d8_53),.data_out(wire_d8_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9855(.data_in(wire_d8_54),.data_out(wire_d8_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9856(.data_in(wire_d8_55),.data_out(wire_d8_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9857(.data_in(wire_d8_56),.data_out(wire_d8_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9858(.data_in(wire_d8_57),.data_out(wire_d8_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9859(.data_in(wire_d8_58),.data_out(wire_d8_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9860(.data_in(wire_d8_59),.data_out(wire_d8_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9861(.data_in(wire_d8_60),.data_out(wire_d8_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9862(.data_in(wire_d8_61),.data_out(wire_d8_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9863(.data_in(wire_d8_62),.data_out(wire_d8_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9864(.data_in(wire_d8_63),.data_out(wire_d8_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9865(.data_in(wire_d8_64),.data_out(wire_d8_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9866(.data_in(wire_d8_65),.data_out(wire_d8_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9867(.data_in(wire_d8_66),.data_out(wire_d8_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9868(.data_in(wire_d8_67),.data_out(wire_d8_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9869(.data_in(wire_d8_68),.data_out(wire_d8_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9870(.data_in(wire_d8_69),.data_out(wire_d8_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9871(.data_in(wire_d8_70),.data_out(wire_d8_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9872(.data_in(wire_d8_71),.data_out(wire_d8_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9873(.data_in(wire_d8_72),.data_out(wire_d8_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9874(.data_in(wire_d8_73),.data_out(wire_d8_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9875(.data_in(wire_d8_74),.data_out(wire_d8_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9876(.data_in(wire_d8_75),.data_out(wire_d8_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9877(.data_in(wire_d8_76),.data_out(wire_d8_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9878(.data_in(wire_d8_77),.data_out(wire_d8_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9879(.data_in(wire_d8_78),.data_out(wire_d8_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9880(.data_in(wire_d8_79),.data_out(wire_d8_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9881(.data_in(wire_d8_80),.data_out(wire_d8_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9882(.data_in(wire_d8_81),.data_out(wire_d8_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9883(.data_in(wire_d8_82),.data_out(wire_d8_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9884(.data_in(wire_d8_83),.data_out(wire_d8_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9885(.data_in(wire_d8_84),.data_out(wire_d8_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9886(.data_in(wire_d8_85),.data_out(wire_d8_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9887(.data_in(wire_d8_86),.data_out(wire_d8_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9888(.data_in(wire_d8_87),.data_out(wire_d8_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9889(.data_in(wire_d8_88),.data_out(wire_d8_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9890(.data_in(wire_d8_89),.data_out(wire_d8_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9891(.data_in(wire_d8_90),.data_out(wire_d8_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9892(.data_in(wire_d8_91),.data_out(wire_d8_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9893(.data_in(wire_d8_92),.data_out(wire_d8_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9894(.data_in(wire_d8_93),.data_out(wire_d8_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9895(.data_in(wire_d8_94),.data_out(wire_d8_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9896(.data_in(wire_d8_95),.data_out(wire_d8_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9897(.data_in(wire_d8_96),.data_out(wire_d8_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9898(.data_in(wire_d8_97),.data_out(wire_d8_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9899(.data_in(wire_d8_98),.data_out(d_out8),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance10090(.data_in(d_in9),.data_out(wire_d9_0),.clk(clk),.rst(rst));            //channel 10
	encoder #(.WIDTH(WIDTH)) encoder_instance10091(.data_in(wire_d9_0),.data_out(wire_d9_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10092(.data_in(wire_d9_1),.data_out(wire_d9_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10093(.data_in(wire_d9_2),.data_out(wire_d9_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10094(.data_in(wire_d9_3),.data_out(wire_d9_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10095(.data_in(wire_d9_4),.data_out(wire_d9_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10096(.data_in(wire_d9_5),.data_out(wire_d9_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10097(.data_in(wire_d9_6),.data_out(wire_d9_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10098(.data_in(wire_d9_7),.data_out(wire_d9_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10099(.data_in(wire_d9_8),.data_out(wire_d9_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100910(.data_in(wire_d9_9),.data_out(wire_d9_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100911(.data_in(wire_d9_10),.data_out(wire_d9_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100912(.data_in(wire_d9_11),.data_out(wire_d9_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100913(.data_in(wire_d9_12),.data_out(wire_d9_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100914(.data_in(wire_d9_13),.data_out(wire_d9_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100915(.data_in(wire_d9_14),.data_out(wire_d9_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100916(.data_in(wire_d9_15),.data_out(wire_d9_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100917(.data_in(wire_d9_16),.data_out(wire_d9_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100918(.data_in(wire_d9_17),.data_out(wire_d9_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100919(.data_in(wire_d9_18),.data_out(wire_d9_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100920(.data_in(wire_d9_19),.data_out(wire_d9_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100921(.data_in(wire_d9_20),.data_out(wire_d9_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100922(.data_in(wire_d9_21),.data_out(wire_d9_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100923(.data_in(wire_d9_22),.data_out(wire_d9_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100924(.data_in(wire_d9_23),.data_out(wire_d9_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100925(.data_in(wire_d9_24),.data_out(wire_d9_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100926(.data_in(wire_d9_25),.data_out(wire_d9_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100927(.data_in(wire_d9_26),.data_out(wire_d9_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100928(.data_in(wire_d9_27),.data_out(wire_d9_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100929(.data_in(wire_d9_28),.data_out(wire_d9_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100930(.data_in(wire_d9_29),.data_out(wire_d9_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100931(.data_in(wire_d9_30),.data_out(wire_d9_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100932(.data_in(wire_d9_31),.data_out(wire_d9_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100933(.data_in(wire_d9_32),.data_out(wire_d9_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100934(.data_in(wire_d9_33),.data_out(wire_d9_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100935(.data_in(wire_d9_34),.data_out(wire_d9_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100936(.data_in(wire_d9_35),.data_out(wire_d9_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100937(.data_in(wire_d9_36),.data_out(wire_d9_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100938(.data_in(wire_d9_37),.data_out(wire_d9_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100939(.data_in(wire_d9_38),.data_out(wire_d9_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100940(.data_in(wire_d9_39),.data_out(wire_d9_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100941(.data_in(wire_d9_40),.data_out(wire_d9_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100942(.data_in(wire_d9_41),.data_out(wire_d9_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100943(.data_in(wire_d9_42),.data_out(wire_d9_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100944(.data_in(wire_d9_43),.data_out(wire_d9_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100945(.data_in(wire_d9_44),.data_out(wire_d9_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100946(.data_in(wire_d9_45),.data_out(wire_d9_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100947(.data_in(wire_d9_46),.data_out(wire_d9_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100948(.data_in(wire_d9_47),.data_out(wire_d9_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100949(.data_in(wire_d9_48),.data_out(wire_d9_49),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100950(.data_in(wire_d9_49),.data_out(wire_d9_50),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100951(.data_in(wire_d9_50),.data_out(wire_d9_51),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100952(.data_in(wire_d9_51),.data_out(wire_d9_52),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100953(.data_in(wire_d9_52),.data_out(wire_d9_53),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100954(.data_in(wire_d9_53),.data_out(wire_d9_54),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100955(.data_in(wire_d9_54),.data_out(wire_d9_55),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100956(.data_in(wire_d9_55),.data_out(wire_d9_56),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100957(.data_in(wire_d9_56),.data_out(wire_d9_57),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100958(.data_in(wire_d9_57),.data_out(wire_d9_58),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100959(.data_in(wire_d9_58),.data_out(wire_d9_59),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100960(.data_in(wire_d9_59),.data_out(wire_d9_60),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100961(.data_in(wire_d9_60),.data_out(wire_d9_61),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100962(.data_in(wire_d9_61),.data_out(wire_d9_62),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100963(.data_in(wire_d9_62),.data_out(wire_d9_63),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100964(.data_in(wire_d9_63),.data_out(wire_d9_64),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100965(.data_in(wire_d9_64),.data_out(wire_d9_65),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100966(.data_in(wire_d9_65),.data_out(wire_d9_66),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100967(.data_in(wire_d9_66),.data_out(wire_d9_67),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100968(.data_in(wire_d9_67),.data_out(wire_d9_68),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100969(.data_in(wire_d9_68),.data_out(wire_d9_69),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100970(.data_in(wire_d9_69),.data_out(wire_d9_70),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100971(.data_in(wire_d9_70),.data_out(wire_d9_71),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100972(.data_in(wire_d9_71),.data_out(wire_d9_72),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100973(.data_in(wire_d9_72),.data_out(wire_d9_73),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100974(.data_in(wire_d9_73),.data_out(wire_d9_74),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100975(.data_in(wire_d9_74),.data_out(wire_d9_75),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100976(.data_in(wire_d9_75),.data_out(wire_d9_76),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100977(.data_in(wire_d9_76),.data_out(wire_d9_77),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100978(.data_in(wire_d9_77),.data_out(wire_d9_78),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100979(.data_in(wire_d9_78),.data_out(wire_d9_79),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100980(.data_in(wire_d9_79),.data_out(wire_d9_80),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100981(.data_in(wire_d9_80),.data_out(wire_d9_81),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100982(.data_in(wire_d9_81),.data_out(wire_d9_82),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100983(.data_in(wire_d9_82),.data_out(wire_d9_83),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100984(.data_in(wire_d9_83),.data_out(wire_d9_84),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100985(.data_in(wire_d9_84),.data_out(wire_d9_85),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100986(.data_in(wire_d9_85),.data_out(wire_d9_86),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100987(.data_in(wire_d9_86),.data_out(wire_d9_87),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100988(.data_in(wire_d9_87),.data_out(wire_d9_88),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100989(.data_in(wire_d9_88),.data_out(wire_d9_89),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100990(.data_in(wire_d9_89),.data_out(wire_d9_90),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100991(.data_in(wire_d9_90),.data_out(wire_d9_91),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100992(.data_in(wire_d9_91),.data_out(wire_d9_92),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100993(.data_in(wire_d9_92),.data_out(wire_d9_93),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100994(.data_in(wire_d9_93),.data_out(wire_d9_94),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100995(.data_in(wire_d9_94),.data_out(wire_d9_95),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100996(.data_in(wire_d9_95),.data_out(wire_d9_96),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100997(.data_in(wire_d9_96),.data_out(wire_d9_97),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100998(.data_in(wire_d9_97),.data_out(wire_d9_98),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100999(.data_in(wire_d9_98),.data_out(d_out9),.clk(clk),.rst(rst));


endmodule