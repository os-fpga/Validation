
module co_sim_shift_register_512bit;

  parameter CLK_PERIOD = 2;
  parameter WIDTH = 512;

  reg clk;
  reg reset;
  reg shift_in;

  wire [WIDTH-1:0] out_reg,out_reg_netlist;

  integer mismatch=0;

  shift_register_512bit golden (.clk(clk),.reset(reset),.shift_in(shift_in),.out_reg(out_reg));
  `ifdef PNR
    shift_register_512bit_post_route netlist (
clk ,
reset ,
shift_in ,
out_reg_netlist[0] ,
out_reg_netlist[1] ,
out_reg_netlist[2] ,
out_reg_netlist[3] ,
out_reg_netlist[4] ,
out_reg_netlist[5] ,
out_reg_netlist[6] ,
out_reg_netlist[7] ,
out_reg_netlist[8] ,
out_reg_netlist[9] ,
out_reg_netlist[10] ,
out_reg_netlist[11] ,
out_reg_netlist[12] ,
out_reg_netlist[13] ,
out_reg_netlist[14] ,
out_reg_netlist[15] ,
out_reg_netlist[16] ,
out_reg_netlist[17] ,
out_reg_netlist[18] ,
out_reg_netlist[19] ,
out_reg_netlist[20] ,
out_reg_netlist[21] ,
out_reg_netlist[22] ,
out_reg_netlist[23] ,
out_reg_netlist[24] ,
out_reg_netlist[25] ,
out_reg_netlist[26] ,
out_reg_netlist[27] ,
out_reg_netlist[28] ,
out_reg_netlist[29] ,
out_reg_netlist[30] ,
out_reg_netlist[31] ,
out_reg_netlist[32] ,
out_reg_netlist[33] ,
out_reg_netlist[34] ,
out_reg_netlist[35] ,
out_reg_netlist[36] ,
out_reg_netlist[37] ,
out_reg_netlist[38] ,
out_reg_netlist[39] ,
out_reg_netlist[40] ,
out_reg_netlist[41] ,
out_reg_netlist[42] ,
out_reg_netlist[43] ,
out_reg_netlist[44] ,
out_reg_netlist[45] ,
out_reg_netlist[46] ,
out_reg_netlist[47] ,
out_reg_netlist[48] ,
out_reg_netlist[49] ,
out_reg_netlist[50] ,
out_reg_netlist[51] ,
out_reg_netlist[52] ,
out_reg_netlist[53] ,
out_reg_netlist[54] ,
out_reg_netlist[55] ,
out_reg_netlist[56] ,
out_reg_netlist[57] ,
out_reg_netlist[58] ,
out_reg_netlist[59] ,
out_reg_netlist[60] ,
out_reg_netlist[61] ,
out_reg_netlist[62] ,
out_reg_netlist[63] ,
out_reg_netlist[64] ,
out_reg_netlist[65] ,
out_reg_netlist[66] ,
out_reg_netlist[67] ,
out_reg_netlist[68] ,
out_reg_netlist[69] ,
out_reg_netlist[70] ,
out_reg_netlist[71] ,
out_reg_netlist[72] ,
out_reg_netlist[73] ,
out_reg_netlist[74] ,
out_reg_netlist[75] ,
out_reg_netlist[76] ,
out_reg_netlist[77] ,
out_reg_netlist[78] ,
out_reg_netlist[79] ,
out_reg_netlist[80] ,
out_reg_netlist[81] ,
out_reg_netlist[82] ,
out_reg_netlist[83] ,
out_reg_netlist[84] ,
out_reg_netlist[85] ,
out_reg_netlist[86] ,
out_reg_netlist[87] ,
out_reg_netlist[88] ,
out_reg_netlist[89] ,
out_reg_netlist[90] ,
out_reg_netlist[91] ,
out_reg_netlist[92] ,
out_reg_netlist[93] ,
out_reg_netlist[94] ,
out_reg_netlist[95] ,
out_reg_netlist[96] ,
out_reg_netlist[97] ,
out_reg_netlist[98] ,
out_reg_netlist[99] ,
out_reg_netlist[100] ,
out_reg_netlist[101] ,
out_reg_netlist[102] ,
out_reg_netlist[103] ,
out_reg_netlist[104] ,
out_reg_netlist[105] ,
out_reg_netlist[106] ,
out_reg_netlist[107] ,
out_reg_netlist[108] ,
out_reg_netlist[109] ,
out_reg_netlist[110] ,
out_reg_netlist[111] ,
out_reg_netlist[112] ,
out_reg_netlist[113] ,
out_reg_netlist[114] ,
out_reg_netlist[115] ,
out_reg_netlist[116] ,
out_reg_netlist[117] ,
out_reg_netlist[118] ,
out_reg_netlist[119] ,
out_reg_netlist[120] ,
out_reg_netlist[121] ,
out_reg_netlist[122] ,
out_reg_netlist[123] ,
out_reg_netlist[124] ,
out_reg_netlist[125] ,
out_reg_netlist[126] ,
out_reg_netlist[127] ,
out_reg_netlist[128] ,
out_reg_netlist[129] ,
out_reg_netlist[130] ,
out_reg_netlist[131] ,
out_reg_netlist[132] ,
out_reg_netlist[133] ,
out_reg_netlist[134] ,
out_reg_netlist[135] ,
out_reg_netlist[136] ,
out_reg_netlist[137] ,
out_reg_netlist[138] ,
out_reg_netlist[139] ,
out_reg_netlist[140] ,
out_reg_netlist[141] ,
out_reg_netlist[142] ,
out_reg_netlist[143] ,
out_reg_netlist[144] ,
out_reg_netlist[145] ,
out_reg_netlist[146] ,
out_reg_netlist[147] ,
out_reg_netlist[148] ,
out_reg_netlist[149] ,
out_reg_netlist[150] ,
out_reg_netlist[151] ,
out_reg_netlist[152] ,
out_reg_netlist[153] ,
out_reg_netlist[154] ,
out_reg_netlist[155] ,
out_reg_netlist[156] ,
out_reg_netlist[157] ,
out_reg_netlist[158] ,
out_reg_netlist[159] ,
out_reg_netlist[160] ,
out_reg_netlist[161] ,
out_reg_netlist[162] ,
out_reg_netlist[163] ,
out_reg_netlist[164] ,
out_reg_netlist[165] ,
out_reg_netlist[166] ,
out_reg_netlist[167] ,
out_reg_netlist[168] ,
out_reg_netlist[169] ,
out_reg_netlist[170] ,
out_reg_netlist[171] ,
out_reg_netlist[172] ,
out_reg_netlist[173] ,
out_reg_netlist[174] ,
out_reg_netlist[175] ,
out_reg_netlist[176] ,
out_reg_netlist[177] ,
out_reg_netlist[178] ,
out_reg_netlist[179] ,
out_reg_netlist[180] ,
out_reg_netlist[181] ,
out_reg_netlist[182] ,
out_reg_netlist[183] ,
out_reg_netlist[184] ,
out_reg_netlist[185] ,
out_reg_netlist[186] ,
out_reg_netlist[187] ,
out_reg_netlist[188] ,
out_reg_netlist[189] ,
out_reg_netlist[190] ,
out_reg_netlist[191] ,
out_reg_netlist[192] ,
out_reg_netlist[193] ,
out_reg_netlist[194] ,
out_reg_netlist[195] ,
out_reg_netlist[196] ,
out_reg_netlist[197] ,
out_reg_netlist[198] ,
out_reg_netlist[199] ,
out_reg_netlist[200] ,
out_reg_netlist[201] ,
out_reg_netlist[202] ,
out_reg_netlist[203] ,
out_reg_netlist[204] ,
out_reg_netlist[205] ,
out_reg_netlist[206] ,
out_reg_netlist[207] ,
out_reg_netlist[208] ,
out_reg_netlist[209] ,
out_reg_netlist[210] ,
out_reg_netlist[211] ,
out_reg_netlist[212] ,
out_reg_netlist[213] ,
out_reg_netlist[214] ,
out_reg_netlist[215] ,
out_reg_netlist[216] ,
out_reg_netlist[217] ,
out_reg_netlist[218] ,
out_reg_netlist[219] ,
out_reg_netlist[220] ,
out_reg_netlist[221] ,
out_reg_netlist[222] ,
out_reg_netlist[223] ,
out_reg_netlist[224] ,
out_reg_netlist[225] ,
out_reg_netlist[226] ,
out_reg_netlist[227] ,
out_reg_netlist[228] ,
out_reg_netlist[229] ,
out_reg_netlist[230] ,
out_reg_netlist[231] ,
out_reg_netlist[232] ,
out_reg_netlist[233] ,
out_reg_netlist[234] ,
out_reg_netlist[235] ,
out_reg_netlist[236] ,
out_reg_netlist[237] ,
out_reg_netlist[238] ,
out_reg_netlist[239] ,
out_reg_netlist[240] ,
out_reg_netlist[241] ,
out_reg_netlist[242] ,
out_reg_netlist[243] ,
out_reg_netlist[244] ,
out_reg_netlist[245] ,
out_reg_netlist[246] ,
out_reg_netlist[247] ,
out_reg_netlist[248] ,
out_reg_netlist[249] ,
out_reg_netlist[250] ,
out_reg_netlist[251] ,
out_reg_netlist[252] ,
out_reg_netlist[253] ,
out_reg_netlist[254] ,
out_reg_netlist[255] ,
out_reg_netlist[256] ,
out_reg_netlist[257] ,
out_reg_netlist[258] ,
out_reg_netlist[259] ,
out_reg_netlist[260] ,
out_reg_netlist[261] ,
out_reg_netlist[262] ,
out_reg_netlist[263] ,
out_reg_netlist[264] ,
out_reg_netlist[265] ,
out_reg_netlist[266] ,
out_reg_netlist[267] ,
out_reg_netlist[268] ,
out_reg_netlist[269] ,
out_reg_netlist[270] ,
out_reg_netlist[271] ,
out_reg_netlist[272] ,
out_reg_netlist[273] ,
out_reg_netlist[274] ,
out_reg_netlist[275] ,
out_reg_netlist[276] ,
out_reg_netlist[277] ,
out_reg_netlist[278] ,
out_reg_netlist[279] ,
out_reg_netlist[280] ,
out_reg_netlist[281] ,
out_reg_netlist[282] ,
out_reg_netlist[283] ,
out_reg_netlist[284] ,
out_reg_netlist[285] ,
out_reg_netlist[286] ,
out_reg_netlist[287] ,
out_reg_netlist[288] ,
out_reg_netlist[289] ,
out_reg_netlist[290] ,
out_reg_netlist[291] ,
out_reg_netlist[292] ,
out_reg_netlist[293] ,
out_reg_netlist[294] ,
out_reg_netlist[295] ,
out_reg_netlist[296] ,
out_reg_netlist[297] ,
out_reg_netlist[298] ,
out_reg_netlist[299] ,
out_reg_netlist[300] ,
out_reg_netlist[301] ,
out_reg_netlist[302] ,
out_reg_netlist[303] ,
out_reg_netlist[304] ,
out_reg_netlist[305] ,
out_reg_netlist[306] ,
out_reg_netlist[307] ,
out_reg_netlist[308] ,
out_reg_netlist[309] ,
out_reg_netlist[310] ,
out_reg_netlist[311] ,
out_reg_netlist[312] ,
out_reg_netlist[313] ,
out_reg_netlist[314] ,
out_reg_netlist[315] ,
out_reg_netlist[316] ,
out_reg_netlist[317] ,
out_reg_netlist[318] ,
out_reg_netlist[319] ,
out_reg_netlist[320] ,
out_reg_netlist[321] ,
out_reg_netlist[322] ,
out_reg_netlist[323] ,
out_reg_netlist[324] ,
out_reg_netlist[325] ,
out_reg_netlist[326] ,
out_reg_netlist[327] ,
out_reg_netlist[328] ,
out_reg_netlist[329] ,
out_reg_netlist[330] ,
out_reg_netlist[331] ,
out_reg_netlist[332] ,
out_reg_netlist[333] ,
out_reg_netlist[334] ,
out_reg_netlist[335] ,
out_reg_netlist[336] ,
out_reg_netlist[337] ,
out_reg_netlist[338] ,
out_reg_netlist[339] ,
out_reg_netlist[340] ,
out_reg_netlist[341] ,
out_reg_netlist[342] ,
out_reg_netlist[343] ,
out_reg_netlist[344] ,
out_reg_netlist[345] ,
out_reg_netlist[346] ,
out_reg_netlist[347] ,
out_reg_netlist[348] ,
out_reg_netlist[349] ,
out_reg_netlist[350] ,
out_reg_netlist[351] ,
out_reg_netlist[352] ,
out_reg_netlist[353] ,
out_reg_netlist[354] ,
out_reg_netlist[355] ,
out_reg_netlist[356] ,
out_reg_netlist[357] ,
out_reg_netlist[358] ,
out_reg_netlist[359] ,
out_reg_netlist[360] ,
out_reg_netlist[361] ,
out_reg_netlist[362] ,
out_reg_netlist[363] ,
out_reg_netlist[364] ,
out_reg_netlist[365] ,
out_reg_netlist[366] ,
out_reg_netlist[367] ,
out_reg_netlist[368] ,
out_reg_netlist[369] ,
out_reg_netlist[370] ,
out_reg_netlist[371] ,
out_reg_netlist[372] ,
out_reg_netlist[373] ,
out_reg_netlist[374] ,
out_reg_netlist[375] ,
out_reg_netlist[376] ,
out_reg_netlist[377] ,
out_reg_netlist[378] ,
out_reg_netlist[379] ,
out_reg_netlist[380] ,
out_reg_netlist[381] ,
out_reg_netlist[382] ,
out_reg_netlist[383] ,
out_reg_netlist[384] ,
out_reg_netlist[385] ,
out_reg_netlist[386] ,
out_reg_netlist[387] ,
out_reg_netlist[388] ,
out_reg_netlist[389] ,
out_reg_netlist[390] ,
out_reg_netlist[391] ,
out_reg_netlist[392] ,
out_reg_netlist[393] ,
out_reg_netlist[394] ,
out_reg_netlist[395] ,
out_reg_netlist[396] ,
out_reg_netlist[397] ,
out_reg_netlist[398] ,
out_reg_netlist[399] ,
out_reg_netlist[400] ,
out_reg_netlist[401] ,
out_reg_netlist[402] ,
out_reg_netlist[403] ,
out_reg_netlist[404] ,
out_reg_netlist[405] ,
out_reg_netlist[406] ,
out_reg_netlist[407] ,
out_reg_netlist[408] ,
out_reg_netlist[409] ,
out_reg_netlist[410] ,
out_reg_netlist[411] ,
out_reg_netlist[412] ,
out_reg_netlist[413] ,
out_reg_netlist[414] ,
out_reg_netlist[415] ,
out_reg_netlist[416] ,
out_reg_netlist[417] ,
out_reg_netlist[418] ,
out_reg_netlist[419] ,
out_reg_netlist[420] ,
out_reg_netlist[421] ,
out_reg_netlist[422] ,
out_reg_netlist[423] ,
out_reg_netlist[424] ,
out_reg_netlist[425] ,
out_reg_netlist[426] ,
out_reg_netlist[427] ,
out_reg_netlist[428] ,
out_reg_netlist[429] ,
out_reg_netlist[430] ,
out_reg_netlist[431] ,
out_reg_netlist[432] ,
out_reg_netlist[433] ,
out_reg_netlist[434] ,
out_reg_netlist[435] ,
out_reg_netlist[436] ,
out_reg_netlist[437] ,
out_reg_netlist[438] ,
out_reg_netlist[439] ,
out_reg_netlist[440] ,
out_reg_netlist[441] ,
out_reg_netlist[442] ,
out_reg_netlist[443] ,
out_reg_netlist[444] ,
out_reg_netlist[445] ,
out_reg_netlist[446] ,
out_reg_netlist[447] ,
out_reg_netlist[448] ,
out_reg_netlist[449] ,
out_reg_netlist[450] ,
out_reg_netlist[451] ,
out_reg_netlist[452] ,
out_reg_netlist[453] ,
out_reg_netlist[454] ,
out_reg_netlist[455] ,
out_reg_netlist[456] ,
out_reg_netlist[457] ,
out_reg_netlist[458] ,
out_reg_netlist[459] ,
out_reg_netlist[460] ,
out_reg_netlist[461] ,
out_reg_netlist[462] ,
out_reg_netlist[463] ,
out_reg_netlist[464] ,
out_reg_netlist[465] ,
out_reg_netlist[466] ,
out_reg_netlist[467] ,
out_reg_netlist[468] ,
out_reg_netlist[469] ,
out_reg_netlist[470] ,
out_reg_netlist[471] ,
out_reg_netlist[472] ,
out_reg_netlist[473] ,
out_reg_netlist[474] ,
out_reg_netlist[475] ,
out_reg_netlist[476] ,
out_reg_netlist[477] ,
out_reg_netlist[478] ,
out_reg_netlist[479] ,
out_reg_netlist[480] ,
out_reg_netlist[481] ,
out_reg_netlist[482] ,
out_reg_netlist[483] ,
out_reg_netlist[484] ,
out_reg_netlist[485] ,
out_reg_netlist[486] ,
out_reg_netlist[487] ,
out_reg_netlist[488] ,
out_reg_netlist[489] ,
out_reg_netlist[490] ,
out_reg_netlist[491] ,
out_reg_netlist[492] ,
out_reg_netlist[493] ,
out_reg_netlist[494] ,
out_reg_netlist[495] ,
out_reg_netlist[496] ,
out_reg_netlist[497] ,
out_reg_netlist[498] ,
out_reg_netlist[499] ,
out_reg_netlist[500] ,
out_reg_netlist[501] ,
out_reg_netlist[502] ,
out_reg_netlist[503] ,
out_reg_netlist[504] ,
out_reg_netlist[505] ,
out_reg_netlist[506] ,
out_reg_netlist[507] ,
out_reg_netlist[508] ,
out_reg_netlist[509] ,
out_reg_netlist[510] ,
out_reg_netlist[511]
  );
  `else
    shift_register_512bit_post_synth netlist (.clk(clk),.reset(reset),.shift_in(shift_in),.out_reg(out_reg_netlist));
  `endif 

  always #((CLK_PERIOD/2)) clk = ~clk;

  initial begin
    clk = 0;
    reset = 1;
    shift_in = 0;

    #20 reset = 0;
    display_stimulus();

    repeat(1500)@(negedge clk) begin
        shift_in = $random;
        @(negedge clk);
        display_stimulus();
        @(negedge clk);
        compare();
    end

    repeat(10)@(negedge clk);

    if(mismatch == 0)
      $display("\n**** All Comparison Matched ***\nSimulation Passed");
    else
      $display("%0d comparison(s) mismatched\nError: Simulation Failed", mismatch);

    $finish;
  end

  task compare();
  	if(out_reg !== out_reg_netlist) begin
    	$display("Data Mismatch. Golden: %0d, Netlist: %0d, Time: %0t", out_reg, out_reg_netlist, $time);
    	mismatch = mismatch+1;
 	end
  	else
  		$display("Data Matched. Golden: %0d, Netlist: %0d, Time: %0t", out_reg, out_reg_netlist, $time);
  endtask

  task display_stimulus();
  	$display ($time,," Test stimulus is: inpt=%0d", out_reg);
  endtask

  initial begin
    $dumpfile("tb.vcd");
    $dumpvars;
  end
endmodule 
