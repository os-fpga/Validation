// system.v

// Generated using ACDS version 12.0 178 at 2012.07.10.20:23:16

`timescale 1 ps / 1 ps
module system (
		output wire [29:0]  ddr_address,         //      ddr.address
		output wire [31:0]  ddr_byteenable,      //         .byteenable
		output wire [5:0]   ddr_burstcount,      //         .burstcount
		output wire         ddr_write,           //         .write
		output wire [255:0] ddr_writedata,       //         .writedata
		output wire         ddr_read,            //         .read
		input  wire [255:0] ddr_readdata,        //         .readdata
		input  wire         ddr_readdatavalid,   //         .readdatavalid
		input  wire         ddr_waitrequest,     //         .waitrequest
		output wire         ddr_burstbegin,      //         .burstbegin
		input  wire         reset_reset,         //    reset.reset
		input  wire [31:0]  usb_address,         //      usb.address
		input  wire         usb_address_ready,   //         .address_ready
		input  wire [31:0]  usb_writedata,       //         .writedata
		input  wire         usb_writedata_ready, //         .writedata_ready
		output wire [31:0]  usb_readdata,        //         .readdata
		output wire         usb_readdata_ready,  //         .readdata_ready
		output wire         usb_address_want,    //         .address_want
		output wire         usb_writedata_want,  //         .writedata_want
		input  wire         usb_readdata_want,   //         .readdata_want
		input  wire         comp_clk_clk,        // comp_clk.clk
		input  wire         ddr_clk_clk          //  ddr_clk.clk
	);

	wire          lu_ddr_waitrequest;                                                              // lu_ddr_translator:av_waitrequest -> lu:ddr_waitrequest
	wire    [5:0] lu_ddr_burstcount;                                                               // lu:ddr_size -> lu_ddr_translator:av_burstcount
	wire   [29:0] lu_ddr_address;                                                                  // lu:ddr_address -> lu_ddr_translator:av_address
	wire  [255:0] lu_ddr_writedata;                                                                // lu:ddr_writedata -> lu_ddr_translator:av_writedata
	wire          lu_ddr_write;                                                                    // lu:ddr_write -> lu_ddr_translator:av_write
	wire          lu_ddr_read;                                                                     // lu:ddr_read -> lu_ddr_translator:av_read
	wire  [255:0] lu_ddr_readdata;                                                                 // lu_ddr_translator:av_readdata -> lu:ddr_rdata
	wire          lu_ddr_readdatavalid;                                                            // lu_ddr_translator:av_readdatavalid -> lu:ddr_rdatavalid
	wire   [31:0] lu_ddr_byteenable;                                                               // lu:ddr_byteenable -> lu_ddr_translator:av_byteenable
	wire          ports2avalon_master_waitrequest;                                                 // ports2avalon_master_translator:av_waitrequest -> ports2avalon:waitrequest
	wire   [31:0] ports2avalon_master_writedata;                                                   // ports2avalon:writedata -> ports2avalon_master_translator:av_writedata
	wire   [31:0] ports2avalon_master_address;                                                     // ports2avalon:address -> ports2avalon_master_translator:av_address
	wire          ports2avalon_master_write;                                                       // ports2avalon:write -> ports2avalon_master_translator:av_write
	wire          ports2avalon_master_read;                                                        // ports2avalon:read -> ports2avalon_master_translator:av_read
	wire   [31:0] ports2avalon_master_readdata;                                                    // ports2avalon_master_translator:av_readdata -> ports2avalon:readdata
	wire          export_s_translator_avalon_anti_slave_0_waitrequest;                             // export:s_waitrequest -> export_s_translator:av_waitrequest
	wire    [5:0] export_s_translator_avalon_anti_slave_0_burstcount;                              // export_s_translator:av_burstcount -> export:s_burstcount
	wire  [255:0] export_s_translator_avalon_anti_slave_0_writedata;                               // export_s_translator:av_writedata -> export:s_writedata
	wire   [24:0] export_s_translator_avalon_anti_slave_0_address;                                 // export_s_translator:av_address -> export:s_address
	wire          export_s_translator_avalon_anti_slave_0_write;                                   // export_s_translator:av_write -> export:s_write
	wire          export_s_translator_avalon_anti_slave_0_beginbursttransfer;                      // export_s_translator:av_beginbursttransfer -> export:s_burstbegin
	wire          export_s_translator_avalon_anti_slave_0_read;                                    // export_s_translator:av_read -> export:s_read
	wire  [255:0] export_s_translator_avalon_anti_slave_0_readdata;                                // export:s_readdata -> export_s_translator:av_readdata
	wire          export_s_translator_avalon_anti_slave_0_readdatavalid;                           // export:s_readdatavalid -> export_s_translator:av_readdatavalid
	wire   [31:0] export_s_translator_avalon_anti_slave_0_byteenable;                              // export_s_translator:av_byteenable -> export:s_byteenable
	wire          lu_s_translator_avalon_anti_slave_0_waitrequest;                                 // lu:s_waitrequest -> lu_s_translator:av_waitrequest
	wire   [31:0] lu_s_translator_avalon_anti_slave_0_writedata;                                   // lu_s_translator:av_writedata -> lu:s_writedata
	wire    [1:0] lu_s_translator_avalon_anti_slave_0_address;                                     // lu_s_translator:av_address -> lu:s_address
	wire          lu_s_translator_avalon_anti_slave_0_write;                                       // lu_s_translator:av_write -> lu:s_write
	wire          lu_s_translator_avalon_anti_slave_0_read;                                        // lu_s_translator:av_read -> lu:s_read
	wire   [31:0] lu_s_translator_avalon_anti_slave_0_readdata;                                    // lu:s_readdata -> lu_s_translator:av_readdata
	wire          lu_ddr_translator_avalon_universal_master_0_waitrequest;                         // lu_ddr_translator_avalon_universal_master_0_agent:av_waitrequest -> lu_ddr_translator:uav_waitrequest
	wire   [10:0] lu_ddr_translator_avalon_universal_master_0_burstcount;                          // lu_ddr_translator:uav_burstcount -> lu_ddr_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [255:0] lu_ddr_translator_avalon_universal_master_0_writedata;                           // lu_ddr_translator:uav_writedata -> lu_ddr_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] lu_ddr_translator_avalon_universal_master_0_address;                             // lu_ddr_translator:uav_address -> lu_ddr_translator_avalon_universal_master_0_agent:av_address
	wire          lu_ddr_translator_avalon_universal_master_0_lock;                                // lu_ddr_translator:uav_lock -> lu_ddr_translator_avalon_universal_master_0_agent:av_lock
	wire          lu_ddr_translator_avalon_universal_master_0_write;                               // lu_ddr_translator:uav_write -> lu_ddr_translator_avalon_universal_master_0_agent:av_write
	wire          lu_ddr_translator_avalon_universal_master_0_read;                                // lu_ddr_translator:uav_read -> lu_ddr_translator_avalon_universal_master_0_agent:av_read
	wire  [255:0] lu_ddr_translator_avalon_universal_master_0_readdata;                            // lu_ddr_translator_avalon_universal_master_0_agent:av_readdata -> lu_ddr_translator:uav_readdata
	wire          lu_ddr_translator_avalon_universal_master_0_debugaccess;                         // lu_ddr_translator:uav_debugaccess -> lu_ddr_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [31:0] lu_ddr_translator_avalon_universal_master_0_byteenable;                          // lu_ddr_translator:uav_byteenable -> lu_ddr_translator_avalon_universal_master_0_agent:av_byteenable
	wire          lu_ddr_translator_avalon_universal_master_0_readdatavalid;                       // lu_ddr_translator_avalon_universal_master_0_agent:av_readdatavalid -> lu_ddr_translator:uav_readdatavalid
	wire          ports2avalon_master_translator_avalon_universal_master_0_waitrequest;            // ports2avalon_master_translator_avalon_universal_master_0_agent:av_waitrequest -> ports2avalon_master_translator:uav_waitrequest
	wire    [2:0] ports2avalon_master_translator_avalon_universal_master_0_burstcount;             // ports2avalon_master_translator:uav_burstcount -> ports2avalon_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] ports2avalon_master_translator_avalon_universal_master_0_writedata;              // ports2avalon_master_translator:uav_writedata -> ports2avalon_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] ports2avalon_master_translator_avalon_universal_master_0_address;                // ports2avalon_master_translator:uav_address -> ports2avalon_master_translator_avalon_universal_master_0_agent:av_address
	wire          ports2avalon_master_translator_avalon_universal_master_0_lock;                   // ports2avalon_master_translator:uav_lock -> ports2avalon_master_translator_avalon_universal_master_0_agent:av_lock
	wire          ports2avalon_master_translator_avalon_universal_master_0_write;                  // ports2avalon_master_translator:uav_write -> ports2avalon_master_translator_avalon_universal_master_0_agent:av_write
	wire          ports2avalon_master_translator_avalon_universal_master_0_read;                   // ports2avalon_master_translator:uav_read -> ports2avalon_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] ports2avalon_master_translator_avalon_universal_master_0_readdata;               // ports2avalon_master_translator_avalon_universal_master_0_agent:av_readdata -> ports2avalon_master_translator:uav_readdata
	wire          ports2avalon_master_translator_avalon_universal_master_0_debugaccess;            // ports2avalon_master_translator:uav_debugaccess -> ports2avalon_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] ports2avalon_master_translator_avalon_universal_master_0_byteenable;             // ports2avalon_master_translator:uav_byteenable -> ports2avalon_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          ports2avalon_master_translator_avalon_universal_master_0_readdatavalid;          // ports2avalon_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> ports2avalon_master_translator:uav_readdatavalid
	wire          export_s_translator_avalon_universal_slave_0_agent_m0_waitrequest;               // export_s_translator:uav_waitrequest -> export_s_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [10:0] export_s_translator_avalon_universal_slave_0_agent_m0_burstcount;                // export_s_translator_avalon_universal_slave_0_agent:m0_burstcount -> export_s_translator:uav_burstcount
	wire  [255:0] export_s_translator_avalon_universal_slave_0_agent_m0_writedata;                 // export_s_translator_avalon_universal_slave_0_agent:m0_writedata -> export_s_translator:uav_writedata
	wire   [31:0] export_s_translator_avalon_universal_slave_0_agent_m0_address;                   // export_s_translator_avalon_universal_slave_0_agent:m0_address -> export_s_translator:uav_address
	wire          export_s_translator_avalon_universal_slave_0_agent_m0_write;                     // export_s_translator_avalon_universal_slave_0_agent:m0_write -> export_s_translator:uav_write
	wire          export_s_translator_avalon_universal_slave_0_agent_m0_lock;                      // export_s_translator_avalon_universal_slave_0_agent:m0_lock -> export_s_translator:uav_lock
	wire          export_s_translator_avalon_universal_slave_0_agent_m0_read;                      // export_s_translator_avalon_universal_slave_0_agent:m0_read -> export_s_translator:uav_read
	wire  [255:0] export_s_translator_avalon_universal_slave_0_agent_m0_readdata;                  // export_s_translator:uav_readdata -> export_s_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          export_s_translator_avalon_universal_slave_0_agent_m0_readdatavalid;             // export_s_translator:uav_readdatavalid -> export_s_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          export_s_translator_avalon_universal_slave_0_agent_m0_debugaccess;               // export_s_translator_avalon_universal_slave_0_agent:m0_debugaccess -> export_s_translator:uav_debugaccess
	wire   [31:0] export_s_translator_avalon_universal_slave_0_agent_m0_byteenable;                // export_s_translator_avalon_universal_slave_0_agent:m0_byteenable -> export_s_translator:uav_byteenable
	wire          export_s_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;        // export_s_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> export_s_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          export_s_translator_avalon_universal_slave_0_agent_rf_source_valid;              // export_s_translator_avalon_universal_slave_0_agent:rf_source_valid -> export_s_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          export_s_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;      // export_s_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> export_s_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [367:0] export_s_translator_avalon_universal_slave_0_agent_rf_source_data;               // export_s_translator_avalon_universal_slave_0_agent:rf_source_data -> export_s_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          export_s_translator_avalon_universal_slave_0_agent_rf_source_ready;              // export_s_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> export_s_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          export_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;     // export_s_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> export_s_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          export_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;           // export_s_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> export_s_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          export_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;   // export_s_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> export_s_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [367:0] export_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;            // export_s_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> export_s_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          export_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;           // export_s_translator_avalon_universal_slave_0_agent:rf_sink_ready -> export_s_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          export_s_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;         // export_s_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> export_s_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [255:0] export_s_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;          // export_s_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> export_s_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          export_s_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;         // export_s_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> export_s_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          lu_s_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // lu_s_translator:uav_waitrequest -> lu_s_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] lu_s_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // lu_s_translator_avalon_universal_slave_0_agent:m0_burstcount -> lu_s_translator:uav_burstcount
	wire   [31:0] lu_s_translator_avalon_universal_slave_0_agent_m0_writedata;                     // lu_s_translator_avalon_universal_slave_0_agent:m0_writedata -> lu_s_translator:uav_writedata
	wire   [31:0] lu_s_translator_avalon_universal_slave_0_agent_m0_address;                       // lu_s_translator_avalon_universal_slave_0_agent:m0_address -> lu_s_translator:uav_address
	wire          lu_s_translator_avalon_universal_slave_0_agent_m0_write;                         // lu_s_translator_avalon_universal_slave_0_agent:m0_write -> lu_s_translator:uav_write
	wire          lu_s_translator_avalon_universal_slave_0_agent_m0_lock;                          // lu_s_translator_avalon_universal_slave_0_agent:m0_lock -> lu_s_translator:uav_lock
	wire          lu_s_translator_avalon_universal_slave_0_agent_m0_read;                          // lu_s_translator_avalon_universal_slave_0_agent:m0_read -> lu_s_translator:uav_read
	wire   [31:0] lu_s_translator_avalon_universal_slave_0_agent_m0_readdata;                      // lu_s_translator:uav_readdata -> lu_s_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          lu_s_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // lu_s_translator:uav_readdatavalid -> lu_s_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          lu_s_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // lu_s_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lu_s_translator:uav_debugaccess
	wire    [3:0] lu_s_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // lu_s_translator_avalon_universal_slave_0_agent:m0_byteenable -> lu_s_translator:uav_byteenable
	wire          lu_s_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // lu_s_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          lu_s_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // lu_s_translator_avalon_universal_slave_0_agent:rf_source_valid -> lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          lu_s_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // lu_s_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [115:0] lu_s_translator_avalon_universal_slave_0_agent_rf_source_data;                   // lu_s_translator_avalon_universal_slave_0_agent:rf_source_data -> lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          lu_s_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lu_s_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lu_s_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lu_s_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lu_s_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [115:0] lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lu_s_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // lu_s_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          lu_s_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // lu_s_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lu_s_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] lu_s_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // lu_s_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lu_s_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          lu_s_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // lu_s_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lu_s_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          lu_ddr_translator_avalon_universal_master_0_agent_cp_endofpacket;                // lu_ddr_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          lu_ddr_translator_avalon_universal_master_0_agent_cp_valid;                      // lu_ddr_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          lu_ddr_translator_avalon_universal_master_0_agent_cp_startofpacket;              // lu_ddr_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [366:0] lu_ddr_translator_avalon_universal_master_0_agent_cp_data;                       // lu_ddr_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          lu_ddr_translator_avalon_universal_master_0_agent_cp_ready;                      // addr_router:sink_ready -> lu_ddr_translator_avalon_universal_master_0_agent:cp_ready
	wire          ports2avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket;   // ports2avalon_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          ports2avalon_master_translator_avalon_universal_master_0_agent_cp_valid;         // ports2avalon_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          ports2avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket; // ports2avalon_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [114:0] ports2avalon_master_translator_avalon_universal_master_0_agent_cp_data;          // ports2avalon_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          ports2avalon_master_translator_avalon_universal_master_0_agent_cp_ready;         // addr_router_001:sink_ready -> ports2avalon_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          addr_router_src_endofpacket;                                                     // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          addr_router_src_valid;                                                           // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire          addr_router_src_startofpacket;                                                   // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [366:0] addr_router_src_data;                                                            // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire    [1:0] addr_router_src_channel;                                                         // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire          addr_router_src_ready;                                                           // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire          mux_pipeline_003_source0_ready;                                                  // lu_ddr_translator_avalon_universal_master_0_agent:rp_ready -> mux_pipeline_003:out_ready
	wire          addr_router_001_src_endofpacket;                                                 // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                       // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                               // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [114:0] addr_router_001_src_data;                                                        // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire    [1:0] addr_router_001_src_channel;                                                     // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                       // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                // rsp_xbar_mux_001:src_endofpacket -> ports2avalon_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                      // rsp_xbar_mux_001:src_valid -> ports2avalon_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                              // rsp_xbar_mux_001:src_startofpacket -> ports2avalon_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [114:0] rsp_xbar_mux_001_src_data;                                                       // rsp_xbar_mux_001:src_data -> ports2avalon_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [1:0] rsp_xbar_mux_001_src_channel;                                                    // rsp_xbar_mux_001:src_channel -> ports2avalon_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_001_src_ready;                                                      // ports2avalon_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire          id_router_src_endofpacket;                                                       // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                             // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                     // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [366:0] id_router_src_data;                                                              // id_router:src_data -> rsp_xbar_demux:sink_data
	wire    [1:0] id_router_src_channel;                                                           // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                             // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          id_router_001_src_endofpacket;                                                   // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                         // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                 // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [114:0] id_router_001_src_data;                                                          // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire    [1:0] id_router_001_src_channel;                                                       // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                         // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                             // cmd_xbar_demux_001:src0_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                   // cmd_xbar_demux_001:src0_valid -> width_adapter:in_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                           // cmd_xbar_demux_001:src0_startofpacket -> width_adapter:in_startofpacket
	wire  [114:0] cmd_xbar_demux_001_src0_data;                                                    // cmd_xbar_demux_001:src0_data -> width_adapter:in_data
	wire    [1:0] cmd_xbar_demux_001_src0_channel;                                                 // cmd_xbar_demux_001:src0_channel -> width_adapter:in_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                   // width_adapter:in_ready -> cmd_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                 // rsp_xbar_demux:src1_endofpacket -> width_adapter_001:in_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                       // rsp_xbar_demux:src1_valid -> width_adapter_001:in_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                               // rsp_xbar_demux:src1_startofpacket -> width_adapter_001:in_startofpacket
	wire  [366:0] rsp_xbar_demux_src1_data;                                                        // rsp_xbar_demux:src1_data -> width_adapter_001:in_data
	wire    [1:0] rsp_xbar_demux_src1_channel;                                                     // rsp_xbar_demux:src1_channel -> width_adapter_001:in_channel
	wire          rsp_xbar_demux_src1_ready;                                                       // width_adapter_001:in_ready -> rsp_xbar_demux:src1_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                    // cmd_xbar_mux:src_endofpacket -> agent_pipeline:in_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                          // cmd_xbar_mux:src_valid -> agent_pipeline:in_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                  // cmd_xbar_mux:src_startofpacket -> agent_pipeline:in_startofpacket
	wire  [366:0] cmd_xbar_mux_src_data;                                                           // cmd_xbar_mux:src_data -> agent_pipeline:in_data
	wire    [1:0] cmd_xbar_mux_src_channel;                                                        // cmd_xbar_mux:src_channel -> agent_pipeline:in_channel
	wire          cmd_xbar_mux_src_ready;                                                          // agent_pipeline:in_ready -> cmd_xbar_mux:src_ready
	wire          agent_pipeline_source0_endofpacket;                                              // agent_pipeline:out_endofpacket -> export_s_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_source0_valid;                                                    // agent_pipeline:out_valid -> export_s_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_source0_startofpacket;                                            // agent_pipeline:out_startofpacket -> export_s_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [366:0] agent_pipeline_source0_data;                                                     // agent_pipeline:out_data -> export_s_translator_avalon_universal_slave_0_agent:cp_data
	wire    [1:0] agent_pipeline_source0_channel;                                                  // agent_pipeline:out_channel -> export_s_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_source0_ready;                                                    // export_s_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline:out_ready
	wire          agent_pipeline_001_source0_endofpacket;                                          // agent_pipeline_001:out_endofpacket -> id_router:sink_endofpacket
	wire          agent_pipeline_001_source0_valid;                                                // agent_pipeline_001:out_valid -> id_router:sink_valid
	wire          agent_pipeline_001_source0_startofpacket;                                        // agent_pipeline_001:out_startofpacket -> id_router:sink_startofpacket
	wire  [366:0] agent_pipeline_001_source0_data;                                                 // agent_pipeline_001:out_data -> id_router:sink_data
	wire          agent_pipeline_001_source0_ready;                                                // id_router:sink_ready -> agent_pipeline_001:out_ready
	wire          export_s_translator_avalon_universal_slave_0_agent_rp_endofpacket;               // export_s_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_001:in_endofpacket
	wire          export_s_translator_avalon_universal_slave_0_agent_rp_valid;                     // export_s_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_001:in_valid
	wire          export_s_translator_avalon_universal_slave_0_agent_rp_startofpacket;             // export_s_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_001:in_startofpacket
	wire  [366:0] export_s_translator_avalon_universal_slave_0_agent_rp_data;                      // export_s_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_001:in_data
	wire          export_s_translator_avalon_universal_slave_0_agent_rp_ready;                     // agent_pipeline_001:in_ready -> export_s_translator_avalon_universal_slave_0_agent:rp_ready
	wire          mux_pipeline_002_source0_ready;                                                  // agent_pipeline_002:in_ready -> mux_pipeline_002:out_ready
	wire          agent_pipeline_002_source0_endofpacket;                                          // agent_pipeline_002:out_endofpacket -> lu_s_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_002_source0_valid;                                                // agent_pipeline_002:out_valid -> lu_s_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_002_source0_startofpacket;                                        // agent_pipeline_002:out_startofpacket -> lu_s_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [114:0] agent_pipeline_002_source0_data;                                                 // agent_pipeline_002:out_data -> lu_s_translator_avalon_universal_slave_0_agent:cp_data
	wire    [1:0] agent_pipeline_002_source0_channel;                                              // agent_pipeline_002:out_channel -> lu_s_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_002_source0_ready;                                                // lu_s_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_002:out_ready
	wire          agent_pipeline_003_source0_endofpacket;                                          // agent_pipeline_003:out_endofpacket -> id_router_001:sink_endofpacket
	wire          agent_pipeline_003_source0_valid;                                                // agent_pipeline_003:out_valid -> id_router_001:sink_valid
	wire          agent_pipeline_003_source0_startofpacket;                                        // agent_pipeline_003:out_startofpacket -> id_router_001:sink_startofpacket
	wire  [114:0] agent_pipeline_003_source0_data;                                                 // agent_pipeline_003:out_data -> id_router_001:sink_data
	wire          agent_pipeline_003_source0_ready;                                                // id_router_001:sink_ready -> agent_pipeline_003:out_ready
	wire          lu_s_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // lu_s_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_003:in_endofpacket
	wire          lu_s_translator_avalon_universal_slave_0_agent_rp_valid;                         // lu_s_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_003:in_valid
	wire          lu_s_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // lu_s_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_003:in_startofpacket
	wire  [114:0] lu_s_translator_avalon_universal_slave_0_agent_rp_data;                          // lu_s_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_003:in_data
	wire          lu_s_translator_avalon_universal_slave_0_agent_rp_ready;                         // agent_pipeline_003:in_ready -> lu_s_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_demux_src0_endofpacket;                                                 // cmd_xbar_demux:src0_endofpacket -> mux_pipeline:in_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                       // cmd_xbar_demux:src0_valid -> mux_pipeline:in_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                               // cmd_xbar_demux:src0_startofpacket -> mux_pipeline:in_startofpacket
	wire  [366:0] cmd_xbar_demux_src0_data;                                                        // cmd_xbar_demux:src0_data -> mux_pipeline:in_data
	wire    [1:0] cmd_xbar_demux_src0_channel;                                                     // cmd_xbar_demux:src0_channel -> mux_pipeline:in_channel
	wire          cmd_xbar_demux_src0_ready;                                                       // mux_pipeline:in_ready -> cmd_xbar_demux:src0_ready
	wire          mux_pipeline_source0_endofpacket;                                                // mux_pipeline:out_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          mux_pipeline_source0_valid;                                                      // mux_pipeline:out_valid -> cmd_xbar_mux:sink0_valid
	wire          mux_pipeline_source0_startofpacket;                                              // mux_pipeline:out_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [366:0] mux_pipeline_source0_data;                                                       // mux_pipeline:out_data -> cmd_xbar_mux:sink0_data
	wire    [1:0] mux_pipeline_source0_channel;                                                    // mux_pipeline:out_channel -> cmd_xbar_mux:sink0_channel
	wire          mux_pipeline_source0_ready;                                                      // cmd_xbar_mux:sink0_ready -> mux_pipeline:out_ready
	wire          width_adapter_src_endofpacket;                                                   // width_adapter:out_endofpacket -> mux_pipeline_001:in_endofpacket
	wire          width_adapter_src_valid;                                                         // width_adapter:out_valid -> mux_pipeline_001:in_valid
	wire          width_adapter_src_startofpacket;                                                 // width_adapter:out_startofpacket -> mux_pipeline_001:in_startofpacket
	wire  [366:0] width_adapter_src_data;                                                          // width_adapter:out_data -> mux_pipeline_001:in_data
	wire          width_adapter_src_ready;                                                         // mux_pipeline_001:in_ready -> width_adapter:out_ready
	wire    [1:0] width_adapter_src_channel;                                                       // width_adapter:out_channel -> mux_pipeline_001:in_channel
	wire          mux_pipeline_001_source0_endofpacket;                                            // mux_pipeline_001:out_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          mux_pipeline_001_source0_valid;                                                  // mux_pipeline_001:out_valid -> cmd_xbar_mux:sink1_valid
	wire          mux_pipeline_001_source0_startofpacket;                                          // mux_pipeline_001:out_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [366:0] mux_pipeline_001_source0_data;                                                   // mux_pipeline_001:out_data -> cmd_xbar_mux:sink1_data
	wire    [1:0] mux_pipeline_001_source0_channel;                                                // mux_pipeline_001:out_channel -> cmd_xbar_mux:sink1_channel
	wire          mux_pipeline_001_source0_ready;                                                  // cmd_xbar_mux:sink1_ready -> mux_pipeline_001:out_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                             // cmd_xbar_demux_001:src1_endofpacket -> mux_pipeline_002:in_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                   // cmd_xbar_demux_001:src1_valid -> mux_pipeline_002:in_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                           // cmd_xbar_demux_001:src1_startofpacket -> mux_pipeline_002:in_startofpacket
	wire  [114:0] cmd_xbar_demux_001_src1_data;                                                    // cmd_xbar_demux_001:src1_data -> mux_pipeline_002:in_data
	wire    [1:0] cmd_xbar_demux_001_src1_channel;                                                 // cmd_xbar_demux_001:src1_channel -> mux_pipeline_002:in_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                   // mux_pipeline_002:in_ready -> cmd_xbar_demux_001:src1_ready
	wire          mux_pipeline_002_source0_endofpacket;                                            // mux_pipeline_002:out_endofpacket -> agent_pipeline_002:in_endofpacket
	wire          mux_pipeline_002_source0_valid;                                                  // mux_pipeline_002:out_valid -> agent_pipeline_002:in_valid
	wire          mux_pipeline_002_source0_startofpacket;                                          // mux_pipeline_002:out_startofpacket -> agent_pipeline_002:in_startofpacket
	wire  [114:0] mux_pipeline_002_source0_data;                                                   // mux_pipeline_002:out_data -> agent_pipeline_002:in_data
	wire    [1:0] mux_pipeline_002_source0_channel;                                                // mux_pipeline_002:out_channel -> agent_pipeline_002:in_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                 // rsp_xbar_demux:src0_endofpacket -> mux_pipeline_003:in_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                       // rsp_xbar_demux:src0_valid -> mux_pipeline_003:in_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                               // rsp_xbar_demux:src0_startofpacket -> mux_pipeline_003:in_startofpacket
	wire  [366:0] rsp_xbar_demux_src0_data;                                                        // rsp_xbar_demux:src0_data -> mux_pipeline_003:in_data
	wire    [1:0] rsp_xbar_demux_src0_channel;                                                     // rsp_xbar_demux:src0_channel -> mux_pipeline_003:in_channel
	wire          rsp_xbar_demux_src0_ready;                                                       // mux_pipeline_003:in_ready -> rsp_xbar_demux:src0_ready
	wire          mux_pipeline_003_source0_endofpacket;                                            // mux_pipeline_003:out_endofpacket -> lu_ddr_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          mux_pipeline_003_source0_valid;                                                  // mux_pipeline_003:out_valid -> lu_ddr_translator_avalon_universal_master_0_agent:rp_valid
	wire          mux_pipeline_003_source0_startofpacket;                                          // mux_pipeline_003:out_startofpacket -> lu_ddr_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [366:0] mux_pipeline_003_source0_data;                                                   // mux_pipeline_003:out_data -> lu_ddr_translator_avalon_universal_master_0_agent:rp_data
	wire    [1:0] mux_pipeline_003_source0_channel;                                                // mux_pipeline_003:out_channel -> lu_ddr_translator_avalon_universal_master_0_agent:rp_channel
	wire          width_adapter_001_src_endofpacket;                                               // width_adapter_001:out_endofpacket -> mux_pipeline_004:in_endofpacket
	wire          width_adapter_001_src_valid;                                                     // width_adapter_001:out_valid -> mux_pipeline_004:in_valid
	wire          width_adapter_001_src_startofpacket;                                             // width_adapter_001:out_startofpacket -> mux_pipeline_004:in_startofpacket
	wire  [114:0] width_adapter_001_src_data;                                                      // width_adapter_001:out_data -> mux_pipeline_004:in_data
	wire          width_adapter_001_src_ready;                                                     // mux_pipeline_004:in_ready -> width_adapter_001:out_ready
	wire    [1:0] width_adapter_001_src_channel;                                                   // width_adapter_001:out_channel -> mux_pipeline_004:in_channel
	wire          mux_pipeline_004_source0_endofpacket;                                            // mux_pipeline_004:out_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          mux_pipeline_004_source0_valid;                                                  // mux_pipeline_004:out_valid -> rsp_xbar_mux_001:sink0_valid
	wire          mux_pipeline_004_source0_startofpacket;                                          // mux_pipeline_004:out_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [114:0] mux_pipeline_004_source0_data;                                                   // mux_pipeline_004:out_data -> rsp_xbar_mux_001:sink0_data
	wire    [1:0] mux_pipeline_004_source0_channel;                                                // mux_pipeline_004:out_channel -> rsp_xbar_mux_001:sink0_channel
	wire          mux_pipeline_004_source0_ready;                                                  // rsp_xbar_mux_001:sink0_ready -> mux_pipeline_004:out_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                             // rsp_xbar_demux_001:src0_endofpacket -> mux_pipeline_005:in_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                   // rsp_xbar_demux_001:src0_valid -> mux_pipeline_005:in_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                           // rsp_xbar_demux_001:src0_startofpacket -> mux_pipeline_005:in_startofpacket
	wire  [114:0] rsp_xbar_demux_001_src0_data;                                                    // rsp_xbar_demux_001:src0_data -> mux_pipeline_005:in_data
	wire    [1:0] rsp_xbar_demux_001_src0_channel;                                                 // rsp_xbar_demux_001:src0_channel -> mux_pipeline_005:in_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                   // mux_pipeline_005:in_ready -> rsp_xbar_demux_001:src0_ready
	wire          mux_pipeline_005_source0_endofpacket;                                            // mux_pipeline_005:out_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          mux_pipeline_005_source0_valid;                                                  // mux_pipeline_005:out_valid -> rsp_xbar_mux_001:sink1_valid
	wire          mux_pipeline_005_source0_startofpacket;                                          // mux_pipeline_005:out_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [114:0] mux_pipeline_005_source0_data;                                                   // mux_pipeline_005:out_data -> rsp_xbar_mux_001:sink1_data
	wire    [1:0] mux_pipeline_005_source0_channel;                                                // mux_pipeline_005:out_channel -> rsp_xbar_mux_001:sink1_channel
	wire          mux_pipeline_005_source0_ready;                                                  // rsp_xbar_mux_001:sink1_ready -> mux_pipeline_005:out_ready

	ports2avalon #(
		.ADDRESS_WIDTH (32)
	) ports2avalon (
		.clk                 (ddr_clk_clk),                     //  clock.clk
		.reset_n             (~reset_reset),                    //  reset.reset_n
		.address             (ports2avalon_master_address),     // master.address
		.read                (ports2avalon_master_read),        //       .read
		.readdata            (ports2avalon_master_readdata),    //       .readdata
		.write               (ports2avalon_master_write),       //       .write
		.writedata           (ports2avalon_master_writedata),   //       .writedata
		.waitrequest         (ports2avalon_master_waitrequest), //       .waitrequest
		.usb_address         (usb_address),                     //    usb.export
		.usb_address_ready   (usb_address_ready),               //       .export
		.usb_writedata       (usb_writedata),                   //       .export
		.usb_writedata_ready (usb_writedata_ready),             //       .export
		.usb_readdata        (usb_readdata),                    //       .export
		.usb_readdata_ready  (usb_readdata_ready),              //       .export
		.usb_address_want    (usb_address_want),                //       .export
		.usb_writedata_want  (usb_writedata_want),              //       .export
		.usb_readdata_want   (usb_readdata_want)                //       .export
	);

	lu_qsys_wrapper #(
		.BURSTLEN      (6),
		.ADDRESS_WIDTH (30)
	) lu (
		.ddr_byteenable  (lu_ddr_byteenable),                               //      ddr.byteenable
		.ddr_read        (lu_ddr_read),                                     //         .read
		.ddr_size        (lu_ddr_burstcount),                               //         .burstcount
		.ddr_writedata   (lu_ddr_writedata),                                //         .writedata
		.ddr_write       (lu_ddr_write),                                    //         .write
		.ddr_rdata       (lu_ddr_readdata),                                 //         .readdata
		.ddr_rdatavalid  (lu_ddr_readdatavalid),                            //         .readdatavalid
		.ddr_waitrequest (lu_ddr_waitrequest),                              //         .waitrequest
		.ddr_address     (lu_ddr_address),                                  //         .address
		.s_address       (lu_s_translator_avalon_anti_slave_0_address),     //        s.address
		.s_writedata     (lu_s_translator_avalon_anti_slave_0_writedata),   //         .writedata
		.s_readdata      (lu_s_translator_avalon_anti_slave_0_readdata),    //         .readdata
		.s_read          (lu_s_translator_avalon_anti_slave_0_read),        //         .read
		.s_write         (lu_s_translator_avalon_anti_slave_0_write),       //         .write
		.s_waitrequest   (lu_s_translator_avalon_anti_slave_0_waitrequest), //         .waitrequest
		.ddr_clk         (ddr_clk_clk),                                     //  ddr_clk.clk
		.comp_clk        (comp_clk_clk),                                    // comp_clk.clk
		.reset           (reset_reset)                                      //    reset.reset
	);

	export_master #(
		.DWIDTH     (256),
		.AWIDTH_S   (25),
		.AWIDTH_M   (30),
		.BYTEWIDTH  (32),
		.BURSTWIDTH (6)
	) export_inst (
		.clk             (ddr_clk_clk),                                                //    clock.clk
		.reset           (reset_reset),                                                //    reset.reset
		.s_address       (export_s_translator_avalon_anti_slave_0_address),            //        s.address
		.s_byteenable    (export_s_translator_avalon_anti_slave_0_byteenable),         //         .byteenable
		.s_burstcount    (export_s_translator_avalon_anti_slave_0_burstcount),         //         .burstcount
		.s_write         (export_s_translator_avalon_anti_slave_0_write),              //         .write
		.s_writedata     (export_s_translator_avalon_anti_slave_0_writedata),          //         .writedata
		.s_read          (export_s_translator_avalon_anti_slave_0_read),               //         .read
		.s_readdata      (export_s_translator_avalon_anti_slave_0_readdata),           //         .readdata
		.s_readdatavalid (export_s_translator_avalon_anti_slave_0_readdatavalid),      //         .readdatavalid
		.s_waitrequest   (export_s_translator_avalon_anti_slave_0_waitrequest),        //         .waitrequest
		.s_burstbegin    (export_s_translator_avalon_anti_slave_0_beginbursttransfer), //         .beginbursttransfer
		.m_address       (ddr_address),                                                // m_export.export
		.m_byteenable    (ddr_byteenable),                                             //         .export
		.m_burstcount    (ddr_burstcount),                                             //         .export
		.m_write         (ddr_write),                                                  //         .export
		.m_writedata     (ddr_writedata),                                              //         .export
		.m_read          (ddr_read),                                                   //         .export
		.m_readdata      (ddr_readdata),                                               //         .export
		.m_readdatavalid (ddr_readdatavalid),                                          //         .export
		.m_waitrequest   (ddr_waitrequest),                                            //         .export
		.m_burstbegin    (ddr_burstbegin)                                              //         .export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (30),
		.AV_DATA_W                   (256),
		.AV_BURSTCOUNT_W             (6),
		.AV_BYTEENABLE_W             (32),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (11),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (32),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) lu_ddr_translator (
		.clk                   (ddr_clk_clk),                                               //                       clk.clk
		.reset                 (reset_reset),                                               //                     reset.reset
		.uav_address           (lu_ddr_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (lu_ddr_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (lu_ddr_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (lu_ddr_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (lu_ddr_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (lu_ddr_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (lu_ddr_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (lu_ddr_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (lu_ddr_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (lu_ddr_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (lu_ddr_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (lu_ddr_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (lu_ddr_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (lu_ddr_burstcount),                                         //                          .burstcount
		.av_byteenable         (lu_ddr_byteenable),                                         //                          .byteenable
		.av_read               (lu_ddr_read),                                               //                          .read
		.av_readdata           (lu_ddr_readdata),                                           //                          .readdata
		.av_readdatavalid      (lu_ddr_readdatavalid),                                      //                          .readdatavalid
		.av_write              (lu_ddr_write),                                              //                          .write
		.av_writedata          (lu_ddr_writedata),                                          //                          .writedata
		.av_beginbursttransfer (1'b0),                                                      //               (terminated)
		.av_begintransfer      (1'b0),                                                      //               (terminated)
		.av_chipselect         (1'b0),                                                      //               (terminated)
		.av_lock               (1'b0),                                                      //               (terminated)
		.av_debugaccess        (1'b0),                                                      //               (terminated)
		.uav_clken             (),                                                          //               (terminated)
		.av_clken              (1'b1)                                                       //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) ports2avalon_master_translator (
		.clk                   (ddr_clk_clk),                                                            //                       clk.clk
		.reset                 (reset_reset),                                                            //                     reset.reset
		.uav_address           (ports2avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (ports2avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (ports2avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (ports2avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (ports2avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (ports2avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (ports2avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (ports2avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (ports2avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (ports2avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (ports2avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (ports2avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (ports2avalon_master_waitrequest),                                        //                          .waitrequest
		.av_read               (ports2avalon_master_read),                                               //                          .read
		.av_readdata           (ports2avalon_master_readdata),                                           //                          .readdata
		.av_write              (ports2avalon_master_write),                                              //                          .write
		.av_writedata          (ports2avalon_master_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                   //               (terminated)
		.av_byteenable         (4'b1111),                                                                //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                   //               (terminated)
		.av_begintransfer      (1'b0),                                                                   //               (terminated)
		.av_chipselect         (1'b0),                                                                   //               (terminated)
		.av_readdatavalid      (),                                                                       //               (terminated)
		.av_lock               (1'b0),                                                                   //               (terminated)
		.av_debugaccess        (1'b0),                                                                   //               (terminated)
		.uav_clken             (),                                                                       //               (terminated)
		.av_clken              (1'b1)                                                                    //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (25),
		.AV_DATA_W                      (256),
		.UAV_DATA_W                     (256),
		.AV_BURSTCOUNT_W                (6),
		.AV_BYTEENABLE_W                (32),
		.UAV_BYTEENABLE_W               (32),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (11),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (32),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) export_s_translator (
		.clk                   (ddr_clk_clk),                                                         //                      clk.clk
		.reset                 (reset_reset),                                                         //                    reset.reset
		.uav_address           (export_s_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (export_s_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (export_s_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (export_s_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (export_s_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (export_s_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (export_s_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (export_s_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (export_s_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (export_s_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (export_s_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (export_s_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (export_s_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (export_s_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (export_s_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (export_s_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_beginbursttransfer (export_s_translator_avalon_anti_slave_0_beginbursttransfer),          //                         .beginbursttransfer
		.av_burstcount         (export_s_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (export_s_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (export_s_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (export_s_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                    //              (terminated)
		.av_lock               (),                                                                    //              (terminated)
		.av_chipselect         (),                                                                    //              (terminated)
		.av_clken              (),                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                //              (terminated)
		.av_debugaccess        (),                                                                    //              (terminated)
		.av_outputenable       ()                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lu_s_translator (
		.clk                   (ddr_clk_clk),                                                     //                      clk.clk
		.reset                 (reset_reset),                                                     //                    reset.reset
		.uav_address           (lu_s_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (lu_s_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (lu_s_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (lu_s_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (lu_s_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (lu_s_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (lu_s_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (lu_s_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (lu_s_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (lu_s_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (lu_s_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (lu_s_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (lu_s_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (lu_s_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (lu_s_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (lu_s_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (lu_s_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                //              (terminated)
		.av_burstcount         (),                                                                //              (terminated)
		.av_byteenable         (),                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                            //              (terminated)
		.av_writebyteenable    (),                                                                //              (terminated)
		.av_lock               (),                                                                //              (terminated)
		.av_chipselect         (),                                                                //              (terminated)
		.av_clken              (),                                                                //              (terminated)
		.uav_clken             (1'b0),                                                            //              (terminated)
		.av_debugaccess        (),                                                                //              (terminated)
		.av_outputenable       ()                                                                 //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (360),
		.PKT_PROTECTION_L          (358),
		.PKT_BEGIN_BURST           (354),
		.PKT_BURSTWRAP_H           (347),
		.PKT_BURSTWRAP_L           (337),
		.PKT_BURST_SIZE_H          (350),
		.PKT_BURST_SIZE_L          (348),
		.PKT_BURST_TYPE_H          (352),
		.PKT_BURST_TYPE_L          (351),
		.PKT_BYTE_CNT_H            (336),
		.PKT_BYTE_CNT_L            (326),
		.PKT_ADDR_H                (319),
		.PKT_ADDR_L                (288),
		.PKT_TRANS_COMPRESSED_READ (320),
		.PKT_TRANS_POSTED          (321),
		.PKT_TRANS_WRITE           (322),
		.PKT_TRANS_READ            (323),
		.PKT_TRANS_LOCK            (324),
		.PKT_TRANS_EXCLUSIVE       (325),
		.PKT_DATA_H                (255),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (287),
		.PKT_BYTEEN_L              (256),
		.PKT_SRC_ID_H              (355),
		.PKT_SRC_ID_L              (355),
		.PKT_DEST_ID_H             (356),
		.PKT_DEST_ID_L             (356),
		.PKT_THREAD_ID_H           (357),
		.PKT_THREAD_ID_L           (357),
		.PKT_CACHE_H               (364),
		.PKT_CACHE_L               (361),
		.PKT_ADDR_SIDEBAND_H       (353),
		.PKT_ADDR_SIDEBAND_L       (353),
		.ST_DATA_W                 (367),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (11),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (2047),
		.CACHE_VALUE               (4'b0000)
	) lu_ddr_translator_avalon_universal_master_0_agent (
		.clk              (ddr_clk_clk),                                                        //       clk.clk
		.reset            (reset_reset),                                                        // clk_reset.reset
		.av_address       (lu_ddr_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (lu_ddr_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (lu_ddr_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (lu_ddr_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (lu_ddr_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (lu_ddr_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (lu_ddr_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (lu_ddr_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (lu_ddr_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (lu_ddr_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (lu_ddr_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (lu_ddr_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (lu_ddr_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (lu_ddr_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (lu_ddr_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (lu_ddr_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (mux_pipeline_003_source0_valid),                                     //        rp.valid
		.rp_data          (mux_pipeline_003_source0_data),                                      //          .data
		.rp_channel       (mux_pipeline_003_source0_channel),                                   //          .channel
		.rp_startofpacket (mux_pipeline_003_source0_startofpacket),                             //          .startofpacket
		.rp_endofpacket   (mux_pipeline_003_source0_endofpacket),                               //          .endofpacket
		.rp_ready         (mux_pipeline_003_source0_ready)                                      //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (108),
		.PKT_PROTECTION_L          (106),
		.PKT_BEGIN_BURST           (102),
		.PKT_BURSTWRAP_H           (95),
		.PKT_BURSTWRAP_L           (85),
		.PKT_BURST_SIZE_H          (98),
		.PKT_BURST_SIZE_L          (96),
		.PKT_BURST_TYPE_H          (100),
		.PKT_BURST_TYPE_L          (99),
		.PKT_BYTE_CNT_H            (84),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (103),
		.PKT_SRC_ID_L              (103),
		.PKT_DEST_ID_H             (104),
		.PKT_DEST_ID_L             (104),
		.PKT_THREAD_ID_H           (105),
		.PKT_THREAD_ID_L           (105),
		.PKT_CACHE_H               (112),
		.PKT_CACHE_L               (109),
		.PKT_ADDR_SIDEBAND_H       (101),
		.PKT_ADDR_SIDEBAND_L       (101),
		.ST_DATA_W                 (115),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (1),
		.BURSTWRAP_VALUE           (2047),
		.CACHE_VALUE               (4'b0000)
	) ports2avalon_master_translator_avalon_universal_master_0_agent (
		.clk              (ddr_clk_clk),                                                                     //       clk.clk
		.reset            (reset_reset),                                                                     // clk_reset.reset
		.av_address       (ports2avalon_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (ports2avalon_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (ports2avalon_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (ports2avalon_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (ports2avalon_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (ports2avalon_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (ports2avalon_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (ports2avalon_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (ports2avalon_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (ports2avalon_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (ports2avalon_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (ports2avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (ports2avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (ports2avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (ports2avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (ports2avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_001_src_valid),                                                      //        rp.valid
		.rp_data          (rsp_xbar_mux_001_src_data),                                                       //          .data
		.rp_channel       (rsp_xbar_mux_001_src_channel),                                                    //          .channel
		.rp_startofpacket (rsp_xbar_mux_001_src_startofpacket),                                              //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_001_src_endofpacket),                                                //          .endofpacket
		.rp_ready         (rsp_xbar_mux_001_src_ready)                                                       //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (255),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (354),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (287),
		.PKT_BYTEEN_L              (256),
		.PKT_ADDR_H                (319),
		.PKT_ADDR_L                (288),
		.PKT_TRANS_COMPRESSED_READ (320),
		.PKT_TRANS_POSTED          (321),
		.PKT_TRANS_WRITE           (322),
		.PKT_TRANS_READ            (323),
		.PKT_TRANS_LOCK            (324),
		.PKT_SRC_ID_H              (355),
		.PKT_SRC_ID_L              (355),
		.PKT_DEST_ID_H             (356),
		.PKT_DEST_ID_L             (356),
		.PKT_BURSTWRAP_H           (347),
		.PKT_BURSTWRAP_L           (337),
		.PKT_BYTE_CNT_H            (336),
		.PKT_BYTE_CNT_L            (326),
		.PKT_PROTECTION_H          (360),
		.PKT_PROTECTION_L          (358),
		.PKT_RESPONSE_STATUS_H     (366),
		.PKT_RESPONSE_STATUS_L     (365),
		.PKT_BURST_SIZE_H          (350),
		.PKT_BURST_SIZE_L          (348),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (367),
		.AVS_BURSTCOUNT_W          (11),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) export_s_translator_avalon_universal_slave_0_agent (
		.clk                     (ddr_clk_clk),                                                                   //             clk.clk
		.reset                   (reset_reset),                                                                   //       clk_reset.reset
		.m0_address              (export_s_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (export_s_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (export_s_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (export_s_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (export_s_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (export_s_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (export_s_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (export_s_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (export_s_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (export_s_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (export_s_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (export_s_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (export_s_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (export_s_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (export_s_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (export_s_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_source0_ready),                                                  //              cp.ready
		.cp_valid                (agent_pipeline_source0_valid),                                                  //                .valid
		.cp_data                 (agent_pipeline_source0_data),                                                   //                .data
		.cp_startofpacket        (agent_pipeline_source0_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (agent_pipeline_source0_endofpacket),                                            //                .endofpacket
		.cp_channel              (agent_pipeline_source0_channel),                                                //                .channel
		.rf_sink_ready           (export_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (export_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (export_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (export_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (export_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (export_s_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (export_s_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (export_s_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (export_s_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (export_s_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (export_s_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (export_s_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (export_s_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (export_s_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (export_s_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (export_s_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (368),
		.FIFO_DEPTH          (65),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) export_s_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (ddr_clk_clk),                                                                   //       clk.clk
		.reset             (reset_reset),                                                                   // clk_reset.reset
		.in_data           (export_s_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (export_s_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (export_s_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (export_s_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (export_s_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (export_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (export_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (export_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (export_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (export_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (102),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (103),
		.PKT_SRC_ID_L              (103),
		.PKT_DEST_ID_H             (104),
		.PKT_DEST_ID_L             (104),
		.PKT_BURSTWRAP_H           (95),
		.PKT_BURSTWRAP_L           (85),
		.PKT_BYTE_CNT_H            (84),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (108),
		.PKT_PROTECTION_L          (106),
		.PKT_RESPONSE_STATUS_H     (114),
		.PKT_RESPONSE_STATUS_L     (113),
		.PKT_BURST_SIZE_H          (98),
		.PKT_BURST_SIZE_L          (96),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (115),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) lu_s_translator_avalon_universal_slave_0_agent (
		.clk                     (ddr_clk_clk),                                                               //             clk.clk
		.reset                   (reset_reset),                                                               //       clk_reset.reset
		.m0_address              (lu_s_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lu_s_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lu_s_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lu_s_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lu_s_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lu_s_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lu_s_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lu_s_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lu_s_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lu_s_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lu_s_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lu_s_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lu_s_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lu_s_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lu_s_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lu_s_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_002_source0_ready),                                          //              cp.ready
		.cp_valid                (agent_pipeline_002_source0_valid),                                          //                .valid
		.cp_data                 (agent_pipeline_002_source0_data),                                           //                .data
		.cp_startofpacket        (agent_pipeline_002_source0_startofpacket),                                  //                .startofpacket
		.cp_endofpacket          (agent_pipeline_002_source0_endofpacket),                                    //                .endofpacket
		.cp_channel              (agent_pipeline_002_source0_channel),                                        //                .channel
		.rf_sink_ready           (lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lu_s_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lu_s_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lu_s_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lu_s_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lu_s_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lu_s_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lu_s_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lu_s_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lu_s_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lu_s_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lu_s_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (116),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (ddr_clk_clk),                                                               //       clk.clk
		.reset             (reset_reset),                                                               // clk_reset.reset
		.in_data           (lu_s_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lu_s_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lu_s_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lu_s_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lu_s_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lu_s_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                     // (terminated)
		.csr_read          (1'b0),                                                                      // (terminated)
		.csr_write         (1'b0),                                                                      // (terminated)
		.csr_readdata      (),                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                      // (terminated)
		.almost_full_data  (),                                                                          // (terminated)
		.almost_empty_data (),                                                                          // (terminated)
		.in_empty          (1'b0),                                                                      // (terminated)
		.out_empty         (),                                                                          // (terminated)
		.in_error          (1'b0),                                                                      // (terminated)
		.out_error         (),                                                                          // (terminated)
		.in_channel        (1'b0),                                                                      // (terminated)
		.out_channel       ()                                                                           // (terminated)
	);

	system_addr_router addr_router (
		.sink_ready         (lu_ddr_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (lu_ddr_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (lu_ddr_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (lu_ddr_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lu_ddr_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (ddr_clk_clk),                                                        //       clk.clk
		.reset              (reset_reset),                                                        // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                              //       src.ready
		.src_valid          (addr_router_src_valid),                                              //          .valid
		.src_data           (addr_router_src_data),                                               //          .data
		.src_channel        (addr_router_src_channel),                                            //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                         //          .endofpacket
	);

	system_addr_router_001 addr_router_001 (
		.sink_ready         (ports2avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (ports2avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (ports2avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (ports2avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ports2avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (ddr_clk_clk),                                                                     //       clk.clk
		.reset              (reset_reset),                                                                     // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                       //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                       //          .valid
		.src_data           (addr_router_001_src_data),                                                        //          .data
		.src_channel        (addr_router_001_src_channel),                                                     //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                  //          .endofpacket
	);

	system_id_router id_router (
		.sink_ready         (agent_pipeline_001_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_001_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_001_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_001_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_001_source0_endofpacket),   //          .endofpacket
		.clk                (ddr_clk_clk),                              //       clk.clk
		.reset              (reset_reset),                              // clk_reset.reset
		.src_ready          (id_router_src_ready),                      //       src.ready
		.src_valid          (id_router_src_valid),                      //          .valid
		.src_data           (id_router_src_data),                       //          .data
		.src_channel        (id_router_src_channel),                    //          .channel
		.src_startofpacket  (id_router_src_startofpacket),              //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                 //          .endofpacket
	);

	system_id_router_001 id_router_001 (
		.sink_ready         (agent_pipeline_003_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_003_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_003_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_003_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_003_source0_endofpacket),   //          .endofpacket
		.clk                (ddr_clk_clk),                              //       clk.clk
		.reset              (reset_reset),                              // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                  //       src.ready
		.src_valid          (id_router_001_src_valid),                  //          .valid
		.src_data           (id_router_001_src_data),                   //          .data
		.src_channel        (id_router_001_src_channel),                //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)             //          .endofpacket
	);

	system_cmd_xbar_demux cmd_xbar_demux (
		.clk                (ddr_clk_clk),                       //       clk.clk
		.reset              (reset_reset),                       // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket)    //          .endofpacket
	);

	system_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (ddr_clk_clk),                           //       clk.clk
		.reset              (reset_reset),                           // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	system_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (ddr_clk_clk),                            //       clk.clk
		.reset               (reset_reset),                            // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                 //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                 //          .valid
		.src_data            (cmd_xbar_mux_src_data),                  //          .data
		.src_channel         (cmd_xbar_mux_src_channel),               //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),         //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),           //          .endofpacket
		.sink0_ready         (mux_pipeline_source0_ready),             //     sink0.ready
		.sink0_valid         (mux_pipeline_source0_valid),             //          .valid
		.sink0_channel       (mux_pipeline_source0_channel),           //          .channel
		.sink0_data          (mux_pipeline_source0_data),              //          .data
		.sink0_startofpacket (mux_pipeline_source0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (mux_pipeline_source0_endofpacket),       //          .endofpacket
		.sink1_ready         (mux_pipeline_001_source0_ready),         //     sink1.ready
		.sink1_valid         (mux_pipeline_001_source0_valid),         //          .valid
		.sink1_channel       (mux_pipeline_001_source0_channel),       //          .channel
		.sink1_data          (mux_pipeline_001_source0_data),          //          .data
		.sink1_startofpacket (mux_pipeline_001_source0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (mux_pipeline_001_source0_endofpacket)    //          .endofpacket
	);

	system_rsp_xbar_demux rsp_xbar_demux (
		.clk                (ddr_clk_clk),                       //       clk.clk
		.reset              (reset_reset),                       // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	system_rsp_xbar_demux_001 rsp_xbar_demux_001 (
		.clk                (ddr_clk_clk),                           //       clk.clk
		.reset              (reset_reset),                           // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	system_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (ddr_clk_clk),                            //       clk.clk
		.reset               (reset_reset),                            // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),             //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),             //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),              //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),           //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),       //          .endofpacket
		.sink0_ready         (mux_pipeline_004_source0_ready),         //     sink0.ready
		.sink0_valid         (mux_pipeline_004_source0_valid),         //          .valid
		.sink0_channel       (mux_pipeline_004_source0_channel),       //          .channel
		.sink0_data          (mux_pipeline_004_source0_data),          //          .data
		.sink0_startofpacket (mux_pipeline_004_source0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (mux_pipeline_004_source0_endofpacket),   //          .endofpacket
		.sink1_ready         (mux_pipeline_005_source0_ready),         //     sink1.ready
		.sink1_valid         (mux_pipeline_005_source0_valid),         //          .valid
		.sink1_channel       (mux_pipeline_005_source0_channel),       //          .channel
		.sink1_data          (mux_pipeline_005_source0_data),          //          .data
		.sink1_startofpacket (mux_pipeline_005_source0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (mux_pipeline_005_source0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (84),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (95),
		.IN_PKT_BURSTWRAP_L            (85),
		.IN_PKT_BURST_SIZE_H           (98),
		.IN_PKT_BURST_SIZE_L           (96),
		.IN_PKT_RESPONSE_STATUS_H      (114),
		.IN_PKT_RESPONSE_STATUS_L      (113),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (100),
		.IN_PKT_BURST_TYPE_L           (99),
		.IN_ST_DATA_W                  (115),
		.OUT_PKT_ADDR_H                (319),
		.OUT_PKT_ADDR_L                (288),
		.OUT_PKT_DATA_H                (255),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (287),
		.OUT_PKT_BYTEEN_L              (256),
		.OUT_PKT_BYTE_CNT_H            (336),
		.OUT_PKT_BYTE_CNT_L            (326),
		.OUT_PKT_TRANS_COMPRESSED_READ (320),
		.OUT_PKT_BURST_SIZE_H          (350),
		.OUT_PKT_BURST_SIZE_L          (348),
		.OUT_PKT_RESPONSE_STATUS_H     (366),
		.OUT_PKT_RESPONSE_STATUS_L     (365),
		.OUT_PKT_TRANS_EXCLUSIVE       (325),
		.OUT_PKT_BURST_TYPE_H          (352),
		.OUT_PKT_BURST_TYPE_L          (351),
		.OUT_ST_DATA_W                 (367),
		.ST_CHANNEL_W                  (2),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk                  (ddr_clk_clk),                           //       clk.clk
		.reset                (reset_reset),                           // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src0_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src0_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src0_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src0_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),         //       src.endofpacket
		.out_data             (width_adapter_src_data),                //          .data
		.out_channel          (width_adapter_src_channel),             //          .channel
		.out_valid            (width_adapter_src_valid),               //          .valid
		.out_ready            (width_adapter_src_ready),               //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),       //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (319),
		.IN_PKT_ADDR_L                 (288),
		.IN_PKT_DATA_H                 (255),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (287),
		.IN_PKT_BYTEEN_L               (256),
		.IN_PKT_BYTE_CNT_H             (336),
		.IN_PKT_BYTE_CNT_L             (326),
		.IN_PKT_TRANS_COMPRESSED_READ  (320),
		.IN_PKT_BURSTWRAP_H            (347),
		.IN_PKT_BURSTWRAP_L            (337),
		.IN_PKT_BURST_SIZE_H           (350),
		.IN_PKT_BURST_SIZE_L           (348),
		.IN_PKT_RESPONSE_STATUS_H      (366),
		.IN_PKT_RESPONSE_STATUS_L      (365),
		.IN_PKT_TRANS_EXCLUSIVE        (325),
		.IN_PKT_BURST_TYPE_H           (352),
		.IN_PKT_BURST_TYPE_L           (351),
		.IN_ST_DATA_W                  (367),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (84),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (98),
		.OUT_PKT_BURST_SIZE_L          (96),
		.OUT_PKT_RESPONSE_STATUS_H     (114),
		.OUT_PKT_RESPONSE_STATUS_L     (113),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (100),
		.OUT_PKT_BURST_TYPE_L          (99),
		.OUT_ST_DATA_W                 (115),
		.ST_CHANNEL_W                  (2),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_001 (
		.clk                  (ddr_clk_clk),                         //       clk.clk
		.reset                (reset_reset),                         // clk_reset.reset
		.in_valid             (rsp_xbar_demux_src1_valid),           //      sink.valid
		.in_channel           (rsp_xbar_demux_src1_channel),         //          .channel
		.in_startofpacket     (rsp_xbar_demux_src1_startofpacket),   //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_src1_endofpacket),     //          .endofpacket
		.in_ready             (rsp_xbar_demux_src1_ready),           //          .ready
		.in_data              (rsp_xbar_demux_src1_data),            //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (367),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (2),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline (
		.clk               (ddr_clk_clk),                          //       cr0.clk
		.reset             (reset_reset),                          // cr0_reset.reset
		.in_ready          (cmd_xbar_mux_src_ready),               //     sink0.ready
		.in_valid          (cmd_xbar_mux_src_valid),               //          .valid
		.in_startofpacket  (cmd_xbar_mux_src_startofpacket),       //          .startofpacket
		.in_endofpacket    (cmd_xbar_mux_src_endofpacket),         //          .endofpacket
		.in_data           (cmd_xbar_mux_src_data),                //          .data
		.in_channel        (cmd_xbar_mux_src_channel),             //          .channel
		.out_ready         (agent_pipeline_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_source0_data),          //          .data
		.out_channel       (agent_pipeline_source0_channel),       //          .channel
		.in_empty          (1'b0),                                 // (terminated)
		.out_empty         (),                                     // (terminated)
		.out_error         (),                                     // (terminated)
		.in_error          (1'b0)                                  // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (367),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_001 (
		.clk               (ddr_clk_clk),                                                         //       cr0.clk
		.reset             (reset_reset),                                                         // cr0_reset.reset
		.in_ready          (export_s_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (export_s_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (export_s_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (export_s_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (export_s_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_001_source0_ready),                                    //   source0.ready
		.out_valid         (agent_pipeline_001_source0_valid),                                    //          .valid
		.out_startofpacket (agent_pipeline_001_source0_startofpacket),                            //          .startofpacket
		.out_endofpacket   (agent_pipeline_001_source0_endofpacket),                              //          .endofpacket
		.out_data          (agent_pipeline_001_source0_data),                                     //          .data
		.in_empty          (1'b0),                                                                // (terminated)
		.out_empty         (),                                                                    // (terminated)
		.out_error         (),                                                                    // (terminated)
		.in_error          (1'b0),                                                                // (terminated)
		.out_channel       (),                                                                    // (terminated)
		.in_channel        (1'b0)                                                                 // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (115),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (2),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_002 (
		.clk               (ddr_clk_clk),                              //       cr0.clk
		.reset             (reset_reset),                              // cr0_reset.reset
		.in_ready          (mux_pipeline_002_source0_ready),           //     sink0.ready
		.in_valid          (mux_pipeline_002_source0_valid),           //          .valid
		.in_startofpacket  (mux_pipeline_002_source0_startofpacket),   //          .startofpacket
		.in_endofpacket    (mux_pipeline_002_source0_endofpacket),     //          .endofpacket
		.in_data           (mux_pipeline_002_source0_data),            //          .data
		.in_channel        (mux_pipeline_002_source0_channel),         //          .channel
		.out_ready         (agent_pipeline_002_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_002_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_002_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_002_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_002_source0_data),          //          .data
		.out_channel       (agent_pipeline_002_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (115),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_003 (
		.clk               (ddr_clk_clk),                                                     //       cr0.clk
		.reset             (reset_reset),                                                     // cr0_reset.reset
		.in_ready          (lu_s_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (lu_s_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (lu_s_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (lu_s_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (lu_s_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_003_source0_ready),                                //   source0.ready
		.out_valid         (agent_pipeline_003_source0_valid),                                //          .valid
		.out_startofpacket (agent_pipeline_003_source0_startofpacket),                        //          .startofpacket
		.out_endofpacket   (agent_pipeline_003_source0_endofpacket),                          //          .endofpacket
		.out_data          (agent_pipeline_003_source0_data),                                 //          .data
		.in_empty          (1'b0),                                                            // (terminated)
		.out_empty         (),                                                                // (terminated)
		.out_error         (),                                                                // (terminated)
		.in_error          (1'b0),                                                            // (terminated)
		.out_channel       (),                                                                // (terminated)
		.in_channel        (1'b0)                                                             // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (367),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (2),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline (
		.clk               (ddr_clk_clk),                        //       cr0.clk
		.reset             (reset_reset),                        // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src0_ready),          //     sink0.ready
		.in_valid          (cmd_xbar_demux_src0_valid),          //          .valid
		.in_startofpacket  (cmd_xbar_demux_src0_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src0_endofpacket),    //          .endofpacket
		.in_data           (cmd_xbar_demux_src0_data),           //          .data
		.in_channel        (cmd_xbar_demux_src0_channel),        //          .channel
		.out_ready         (mux_pipeline_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_source0_data),          //          .data
		.out_channel       (mux_pipeline_source0_channel),       //          .channel
		.in_empty          (1'b0),                               // (terminated)
		.out_empty         (),                                   // (terminated)
		.out_error         (),                                   // (terminated)
		.in_error          (1'b0)                                // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (367),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (2),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_001 (
		.clk               (ddr_clk_clk),                            //       cr0.clk
		.reset             (reset_reset),                            // cr0_reset.reset
		.in_ready          (width_adapter_src_ready),                //     sink0.ready
		.in_valid          (width_adapter_src_valid),                //          .valid
		.in_startofpacket  (width_adapter_src_startofpacket),        //          .startofpacket
		.in_endofpacket    (width_adapter_src_endofpacket),          //          .endofpacket
		.in_data           (width_adapter_src_data),                 //          .data
		.in_channel        (width_adapter_src_channel),              //          .channel
		.out_ready         (mux_pipeline_001_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_001_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_001_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_001_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_001_source0_data),          //          .data
		.out_channel       (mux_pipeline_001_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (115),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (2),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_002 (
		.clk               (ddr_clk_clk),                            //       cr0.clk
		.reset             (reset_reset),                            // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_001_src1_ready),          //     sink0.ready
		.in_valid          (cmd_xbar_demux_001_src1_valid),          //          .valid
		.in_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //          .endofpacket
		.in_data           (cmd_xbar_demux_001_src1_data),           //          .data
		.in_channel        (cmd_xbar_demux_001_src1_channel),        //          .channel
		.out_ready         (mux_pipeline_002_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_002_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_002_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_002_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_002_source0_data),          //          .data
		.out_channel       (mux_pipeline_002_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (367),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (2),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_003 (
		.clk               (ddr_clk_clk),                            //       cr0.clk
		.reset             (reset_reset),                            // cr0_reset.reset
		.in_ready          (rsp_xbar_demux_src0_ready),              //     sink0.ready
		.in_valid          (rsp_xbar_demux_src0_valid),              //          .valid
		.in_startofpacket  (rsp_xbar_demux_src0_startofpacket),      //          .startofpacket
		.in_endofpacket    (rsp_xbar_demux_src0_endofpacket),        //          .endofpacket
		.in_data           (rsp_xbar_demux_src0_data),               //          .data
		.in_channel        (rsp_xbar_demux_src0_channel),            //          .channel
		.out_ready         (mux_pipeline_003_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_003_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_003_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_003_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_003_source0_data),          //          .data
		.out_channel       (mux_pipeline_003_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (115),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (2),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_004 (
		.clk               (ddr_clk_clk),                            //       cr0.clk
		.reset             (reset_reset),                            // cr0_reset.reset
		.in_ready          (width_adapter_001_src_ready),            //     sink0.ready
		.in_valid          (width_adapter_001_src_valid),            //          .valid
		.in_startofpacket  (width_adapter_001_src_startofpacket),    //          .startofpacket
		.in_endofpacket    (width_adapter_001_src_endofpacket),      //          .endofpacket
		.in_data           (width_adapter_001_src_data),             //          .data
		.in_channel        (width_adapter_001_src_channel),          //          .channel
		.out_ready         (mux_pipeline_004_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_004_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_004_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_004_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_004_source0_data),          //          .data
		.out_channel       (mux_pipeline_004_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (115),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (2),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) mux_pipeline_005 (
		.clk               (ddr_clk_clk),                            //       cr0.clk
		.reset             (reset_reset),                            // cr0_reset.reset
		.in_ready          (rsp_xbar_demux_001_src0_ready),          //     sink0.ready
		.in_valid          (rsp_xbar_demux_001_src0_valid),          //          .valid
		.in_startofpacket  (rsp_xbar_demux_001_src0_startofpacket),  //          .startofpacket
		.in_endofpacket    (rsp_xbar_demux_001_src0_endofpacket),    //          .endofpacket
		.in_data           (rsp_xbar_demux_001_src0_data),           //          .data
		.in_channel        (rsp_xbar_demux_001_src0_channel),        //          .channel
		.out_ready         (mux_pipeline_005_source0_ready),         //   source0.ready
		.out_valid         (mux_pipeline_005_source0_valid),         //          .valid
		.out_startofpacket (mux_pipeline_005_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (mux_pipeline_005_source0_endofpacket),   //          .endofpacket
		.out_data          (mux_pipeline_005_source0_data),          //          .data
		.out_channel       (mux_pipeline_005_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

endmodule
