// hh_system.v

// Generated using ACDS version 12.0 178 at 2012.07.10.17:46:07

`timescale 1 ps / 1 ps
module hh_system (
		input  wire        reset_reset_n,                      //              reset.reset_n
		input  wire        clk_clk,                            //                clk.clk
		input  wire [31:0] ports2avalon_0_usb_address,         // ports2avalon_0_usb.address
		input  wire        ports2avalon_0_usb_address_ready,   //                   .address_ready
		input  wire [31:0] ports2avalon_0_usb_writedata,       //                   .writedata
		input  wire        ports2avalon_0_usb_writedata_ready, //                   .writedata_ready
		output wire [31:0] ports2avalon_0_usb_readdata,        //                   .readdata
		output wire        ports2avalon_0_usb_readdata_ready,  //                   .readdata_ready
		output wire        ports2avalon_0_usb_address_want,    //                   .address_want
		output wire        ports2avalon_0_usb_writedata_want,  //                   .writedata_want
		input  wire        ports2avalon_0_usb_readdata_want    //                   .readdata_want
	);

	wire          hh_core_0_outputdata_source_valid;                                                        // hh_core_0:o_valid -> timing_adapter:in_valid
	wire   [31:0] hh_core_0_outputdata_source_data;                                                         // hh_core_0:o_data -> timing_adapter:in_data
	wire          hh_core_0_outputdata_source_ready;                                                        // timing_adapter:in_ready -> hh_core_0:i_ready
	wire          timing_adapter_out_valid;                                                                 // timing_adapter:out_valid -> output_data:avalonst_sink_valid
	wire   [31:0] timing_adapter_out_data;                                                                  // timing_adapter:out_data -> output_data:avalonst_sink_data
	wire          timing_adapter_out_ready;                                                                 // output_data:avalonst_sink_ready -> timing_adapter:out_ready
	wire          input_data_out_valid;                                                                     // input_data:avalonst_source_valid -> timing_adapter_1:in_valid
	wire   [31:0] input_data_out_data;                                                                      // input_data:avalonst_source_data -> timing_adapter_1:in_data
	wire          input_data_out_ready;                                                                     // timing_adapter_1:in_ready -> input_data:avalonst_source_ready
	wire          timing_adapter_1_out_valid;                                                               // timing_adapter_1:out_valid -> hh_core_0:i_valid
	wire   [31:0] timing_adapter_1_out_data;                                                                // timing_adapter_1:out_data -> hh_core_0:i_data
	wire          timing_adapter_1_out_ready;                                                               // hh_core_0:o_ready -> timing_adapter_1:out_ready
	wire          ports2avalon_0_master_waitrequest;                                                        // ports2avalon_0_master_translator:av_waitrequest -> ports2avalon_0:waitrequest
	wire   [31:0] ports2avalon_0_master_writedata;                                                          // ports2avalon_0:writedata -> ports2avalon_0_master_translator:av_writedata
	wire   [31:0] ports2avalon_0_master_address;                                                            // ports2avalon_0:address -> ports2avalon_0_master_translator:av_address
	wire          ports2avalon_0_master_write;                                                              // ports2avalon_0:write -> ports2avalon_0_master_translator:av_write
	wire          ports2avalon_0_master_read;                                                               // ports2avalon_0:read -> ports2avalon_0_master_translator:av_read
	wire   [31:0] ports2avalon_0_master_readdata;                                                           // ports2avalon_0_master_translator:av_readdata -> ports2avalon_0:readdata
	wire          output_data_out_translator_avalon_anti_slave_0_waitrequest;                               // output_data:avalonmm_read_slave_waitrequest -> output_data_out_translator:av_waitrequest
	wire          output_data_out_translator_avalon_anti_slave_0_address;                                   // output_data_out_translator:av_address -> output_data:avalonmm_read_slave_address
	wire          output_data_out_translator_avalon_anti_slave_0_read;                                      // output_data_out_translator:av_read -> output_data:avalonmm_read_slave_read
	wire   [31:0] output_data_out_translator_avalon_anti_slave_0_readdata;                                  // output_data:avalonmm_read_slave_readdata -> output_data_out_translator:av_readdata
	wire          input_data_in_translator_avalon_anti_slave_0_waitrequest;                                 // input_data:avalonmm_write_slave_waitrequest -> input_data_in_translator:av_waitrequest
	wire   [31:0] input_data_in_translator_avalon_anti_slave_0_writedata;                                   // input_data_in_translator:av_writedata -> input_data:avalonmm_write_slave_writedata
	wire          input_data_in_translator_avalon_anti_slave_0_address;                                     // input_data_in_translator:av_address -> input_data:avalonmm_write_slave_address
	wire          input_data_in_translator_avalon_anti_slave_0_write;                                       // input_data_in_translator:av_write -> input_data:avalonmm_write_slave_write
	wire          hh_core_0_ctrl_port_translator_avalon_anti_slave_0_waitrequest;                           // hh_core_0:o_waitrequest -> hh_core_0_ctrl_port_translator:av_waitrequest
	wire   [31:0] hh_core_0_ctrl_port_translator_avalon_anti_slave_0_writedata;                             // hh_core_0_ctrl_port_translator:av_writedata -> hh_core_0:i_writedata
	wire    [1:0] hh_core_0_ctrl_port_translator_avalon_anti_slave_0_address;                               // hh_core_0_ctrl_port_translator:av_address -> hh_core_0:i_address
	wire          hh_core_0_ctrl_port_translator_avalon_anti_slave_0_write;                                 // hh_core_0_ctrl_port_translator:av_write -> hh_core_0:i_write
	wire          hh_core_0_ctrl_port_translator_avalon_anti_slave_0_read;                                  // hh_core_0_ctrl_port_translator:av_read -> hh_core_0:i_read
	wire   [31:0] hh_core_0_ctrl_port_translator_avalon_anti_slave_0_readdata;                              // hh_core_0:o_readdata -> hh_core_0_ctrl_port_translator:av_readdata
	wire   [31:0] input_data_in_csr_translator_avalon_anti_slave_0_writedata;                               // input_data_in_csr_translator:av_writedata -> input_data:wrclk_control_slave_writedata
	wire    [2:0] input_data_in_csr_translator_avalon_anti_slave_0_address;                                 // input_data_in_csr_translator:av_address -> input_data:wrclk_control_slave_address
	wire          input_data_in_csr_translator_avalon_anti_slave_0_write;                                   // input_data_in_csr_translator:av_write -> input_data:wrclk_control_slave_write
	wire          input_data_in_csr_translator_avalon_anti_slave_0_read;                                    // input_data_in_csr_translator:av_read -> input_data:wrclk_control_slave_read
	wire   [31:0] input_data_in_csr_translator_avalon_anti_slave_0_readdata;                                // input_data:wrclk_control_slave_readdata -> input_data_in_csr_translator:av_readdata
	wire   [31:0] output_data_in_csr_translator_avalon_anti_slave_0_writedata;                              // output_data_in_csr_translator:av_writedata -> output_data:wrclk_control_slave_writedata
	wire    [2:0] output_data_in_csr_translator_avalon_anti_slave_0_address;                                // output_data_in_csr_translator:av_address -> output_data:wrclk_control_slave_address
	wire          output_data_in_csr_translator_avalon_anti_slave_0_write;                                  // output_data_in_csr_translator:av_write -> output_data:wrclk_control_slave_write
	wire          output_data_in_csr_translator_avalon_anti_slave_0_read;                                   // output_data_in_csr_translator:av_read -> output_data:wrclk_control_slave_read
	wire   [31:0] output_data_in_csr_translator_avalon_anti_slave_0_readdata;                               // output_data:wrclk_control_slave_readdata -> output_data_in_csr_translator:av_readdata
	wire          ports2avalon_0_master_translator_avalon_universal_master_0_waitrequest;                   // ports2avalon_0_master_translator_avalon_universal_master_0_agent:av_waitrequest -> ports2avalon_0_master_translator:uav_waitrequest
	wire    [2:0] ports2avalon_0_master_translator_avalon_universal_master_0_burstcount;                    // ports2avalon_0_master_translator:uav_burstcount -> ports2avalon_0_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] ports2avalon_0_master_translator_avalon_universal_master_0_writedata;                     // ports2avalon_0_master_translator:uav_writedata -> ports2avalon_0_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] ports2avalon_0_master_translator_avalon_universal_master_0_address;                       // ports2avalon_0_master_translator:uav_address -> ports2avalon_0_master_translator_avalon_universal_master_0_agent:av_address
	wire          ports2avalon_0_master_translator_avalon_universal_master_0_lock;                          // ports2avalon_0_master_translator:uav_lock -> ports2avalon_0_master_translator_avalon_universal_master_0_agent:av_lock
	wire          ports2avalon_0_master_translator_avalon_universal_master_0_write;                         // ports2avalon_0_master_translator:uav_write -> ports2avalon_0_master_translator_avalon_universal_master_0_agent:av_write
	wire          ports2avalon_0_master_translator_avalon_universal_master_0_read;                          // ports2avalon_0_master_translator:uav_read -> ports2avalon_0_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] ports2avalon_0_master_translator_avalon_universal_master_0_readdata;                      // ports2avalon_0_master_translator_avalon_universal_master_0_agent:av_readdata -> ports2avalon_0_master_translator:uav_readdata
	wire          ports2avalon_0_master_translator_avalon_universal_master_0_debugaccess;                   // ports2avalon_0_master_translator:uav_debugaccess -> ports2avalon_0_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] ports2avalon_0_master_translator_avalon_universal_master_0_byteenable;                    // ports2avalon_0_master_translator:uav_byteenable -> ports2avalon_0_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          ports2avalon_0_master_translator_avalon_universal_master_0_readdatavalid;                 // ports2avalon_0_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> ports2avalon_0_master_translator:uav_readdatavalid
	wire          output_data_out_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // output_data_out_translator:uav_waitrequest -> output_data_out_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] output_data_out_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // output_data_out_translator_avalon_universal_slave_0_agent:m0_burstcount -> output_data_out_translator:uav_burstcount
	wire   [31:0] output_data_out_translator_avalon_universal_slave_0_agent_m0_writedata;                   // output_data_out_translator_avalon_universal_slave_0_agent:m0_writedata -> output_data_out_translator:uav_writedata
	wire   [31:0] output_data_out_translator_avalon_universal_slave_0_agent_m0_address;                     // output_data_out_translator_avalon_universal_slave_0_agent:m0_address -> output_data_out_translator:uav_address
	wire          output_data_out_translator_avalon_universal_slave_0_agent_m0_write;                       // output_data_out_translator_avalon_universal_slave_0_agent:m0_write -> output_data_out_translator:uav_write
	wire          output_data_out_translator_avalon_universal_slave_0_agent_m0_lock;                        // output_data_out_translator_avalon_universal_slave_0_agent:m0_lock -> output_data_out_translator:uav_lock
	wire          output_data_out_translator_avalon_universal_slave_0_agent_m0_read;                        // output_data_out_translator_avalon_universal_slave_0_agent:m0_read -> output_data_out_translator:uav_read
	wire   [31:0] output_data_out_translator_avalon_universal_slave_0_agent_m0_readdata;                    // output_data_out_translator:uav_readdata -> output_data_out_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          output_data_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // output_data_out_translator:uav_readdatavalid -> output_data_out_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          output_data_out_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // output_data_out_translator_avalon_universal_slave_0_agent:m0_debugaccess -> output_data_out_translator:uav_debugaccess
	wire    [3:0] output_data_out_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // output_data_out_translator_avalon_universal_slave_0_agent:m0_byteenable -> output_data_out_translator:uav_byteenable
	wire          output_data_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // output_data_out_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          output_data_out_translator_avalon_universal_slave_0_agent_rf_source_valid;                // output_data_out_translator_avalon_universal_slave_0_agent:rf_source_valid -> output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          output_data_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // output_data_out_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] output_data_out_translator_avalon_universal_slave_0_agent_rf_source_data;                 // output_data_out_translator_avalon_universal_slave_0_agent:rf_source_data -> output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          output_data_out_translator_avalon_universal_slave_0_agent_rf_source_ready;                // output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> output_data_out_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> output_data_out_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> output_data_out_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> output_data_out_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> output_data_out_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // output_data_out_translator_avalon_universal_slave_0_agent:rf_sink_ready -> output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          output_data_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // output_data_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> output_data_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] output_data_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // output_data_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> output_data_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          output_data_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // output_data_out_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> output_data_out_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          input_data_in_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // input_data_in_translator:uav_waitrequest -> input_data_in_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] input_data_in_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // input_data_in_translator_avalon_universal_slave_0_agent:m0_burstcount -> input_data_in_translator:uav_burstcount
	wire   [31:0] input_data_in_translator_avalon_universal_slave_0_agent_m0_writedata;                     // input_data_in_translator_avalon_universal_slave_0_agent:m0_writedata -> input_data_in_translator:uav_writedata
	wire   [31:0] input_data_in_translator_avalon_universal_slave_0_agent_m0_address;                       // input_data_in_translator_avalon_universal_slave_0_agent:m0_address -> input_data_in_translator:uav_address
	wire          input_data_in_translator_avalon_universal_slave_0_agent_m0_write;                         // input_data_in_translator_avalon_universal_slave_0_agent:m0_write -> input_data_in_translator:uav_write
	wire          input_data_in_translator_avalon_universal_slave_0_agent_m0_lock;                          // input_data_in_translator_avalon_universal_slave_0_agent:m0_lock -> input_data_in_translator:uav_lock
	wire          input_data_in_translator_avalon_universal_slave_0_agent_m0_read;                          // input_data_in_translator_avalon_universal_slave_0_agent:m0_read -> input_data_in_translator:uav_read
	wire   [31:0] input_data_in_translator_avalon_universal_slave_0_agent_m0_readdata;                      // input_data_in_translator:uav_readdata -> input_data_in_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          input_data_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // input_data_in_translator:uav_readdatavalid -> input_data_in_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          input_data_in_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // input_data_in_translator_avalon_universal_slave_0_agent:m0_debugaccess -> input_data_in_translator:uav_debugaccess
	wire    [3:0] input_data_in_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // input_data_in_translator_avalon_universal_slave_0_agent:m0_byteenable -> input_data_in_translator:uav_byteenable
	wire          input_data_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // input_data_in_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          input_data_in_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // input_data_in_translator_avalon_universal_slave_0_agent:rf_source_valid -> input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          input_data_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // input_data_in_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] input_data_in_translator_avalon_universal_slave_0_agent_rf_source_data;                   // input_data_in_translator_avalon_universal_slave_0_agent:rf_source_data -> input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          input_data_in_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> input_data_in_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> input_data_in_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> input_data_in_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> input_data_in_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> input_data_in_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // input_data_in_translator_avalon_universal_slave_0_agent:rf_sink_ready -> input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          input_data_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // input_data_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> input_data_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] input_data_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // input_data_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> input_data_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          input_data_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // input_data_in_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> input_data_in_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // hh_core_0_ctrl_port_translator:uav_waitrequest -> hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_burstcount;              // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> hh_core_0_ctrl_port_translator:uav_burstcount
	wire   [31:0] hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_writedata;               // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:m0_writedata -> hh_core_0_ctrl_port_translator:uav_writedata
	wire   [31:0] hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_address;                 // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:m0_address -> hh_core_0_ctrl_port_translator:uav_address
	wire          hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_write;                   // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:m0_write -> hh_core_0_ctrl_port_translator:uav_write
	wire          hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_lock;                    // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:m0_lock -> hh_core_0_ctrl_port_translator:uav_lock
	wire          hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_read;                    // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:m0_read -> hh_core_0_ctrl_port_translator:uav_read
	wire   [31:0] hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_readdata;                // hh_core_0_ctrl_port_translator:uav_readdata -> hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // hh_core_0_ctrl_port_translator:uav_readdatavalid -> hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hh_core_0_ctrl_port_translator:uav_debugaccess
	wire    [3:0] hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_byteenable;              // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> hh_core_0_ctrl_port_translator:uav_byteenable
	wire          hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rf_source_valid;            // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rf_source_data;             // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:rf_source_data -> hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rf_source_ready;            // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;               // input_data_in_csr_translator:uav_waitrequest -> input_data_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                // input_data_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> input_data_in_csr_translator:uav_burstcount
	wire   [31:0] input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                 // input_data_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> input_data_in_csr_translator:uav_writedata
	wire   [31:0] input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                   // input_data_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> input_data_in_csr_translator:uav_address
	wire          input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                     // input_data_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> input_data_in_csr_translator:uav_write
	wire          input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                      // input_data_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> input_data_in_csr_translator:uav_lock
	wire          input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                      // input_data_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> input_data_in_csr_translator:uav_read
	wire   [31:0] input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                  // input_data_in_csr_translator:uav_readdata -> input_data_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;             // input_data_in_csr_translator:uav_readdatavalid -> input_data_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;               // input_data_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> input_data_in_csr_translator:uav_debugaccess
	wire    [3:0] input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                // input_data_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> input_data_in_csr_translator:uav_byteenable
	wire          input_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;        // input_data_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          input_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;              // input_data_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          input_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;      // input_data_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] input_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;               // input_data_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          input_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;              // input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> input_data_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;     // input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> input_data_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;           // input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> input_data_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;   // input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> input_data_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;            // input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> input_data_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;           // input_data_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          input_data_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;         // input_data_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> input_data_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] input_data_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;          // input_data_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> input_data_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          input_data_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;         // input_data_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> input_data_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // output_data_in_csr_translator:uav_waitrequest -> output_data_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;               // output_data_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> output_data_in_csr_translator:uav_burstcount
	wire   [31:0] output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                // output_data_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> output_data_in_csr_translator:uav_writedata
	wire   [31:0] output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                  // output_data_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> output_data_in_csr_translator:uav_address
	wire          output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                    // output_data_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> output_data_in_csr_translator:uav_write
	wire          output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                     // output_data_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> output_data_in_csr_translator:uav_lock
	wire          output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                     // output_data_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> output_data_in_csr_translator:uav_read
	wire   [31:0] output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                 // output_data_in_csr_translator:uav_readdata -> output_data_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // output_data_in_csr_translator:uav_readdatavalid -> output_data_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // output_data_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> output_data_in_csr_translator:uav_debugaccess
	wire    [3:0] output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;               // output_data_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> output_data_in_csr_translator:uav_byteenable
	wire          output_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // output_data_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          output_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;             // output_data_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          output_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // output_data_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] output_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;              // output_data_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          output_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;             // output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> output_data_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> output_data_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> output_data_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> output_data_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> output_data_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // output_data_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          output_data_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // output_data_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> output_data_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] output_data_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // output_data_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> output_data_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          output_data_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // output_data_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> output_data_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ports2avalon_0_master_translator_avalon_universal_master_0_agent_cp_endofpacket;          // ports2avalon_0_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          ports2avalon_0_master_translator_avalon_universal_master_0_agent_cp_valid;                // ports2avalon_0_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          ports2avalon_0_master_translator_avalon_universal_master_0_agent_cp_startofpacket;        // ports2avalon_0_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [102:0] ports2avalon_0_master_translator_avalon_universal_master_0_agent_cp_data;                 // ports2avalon_0_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          ports2avalon_0_master_translator_avalon_universal_master_0_agent_cp_ready;                // addr_router:sink_ready -> ports2avalon_0_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          output_data_out_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // output_data_out_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          output_data_out_translator_avalon_universal_slave_0_agent_rp_valid;                       // output_data_out_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          output_data_out_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // output_data_out_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [102:0] output_data_out_translator_avalon_universal_slave_0_agent_rp_data;                        // output_data_out_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          output_data_out_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router:sink_ready -> output_data_out_translator_avalon_universal_slave_0_agent:rp_ready
	wire          input_data_in_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // input_data_in_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          input_data_in_translator_avalon_universal_slave_0_agent_rp_valid;                         // input_data_in_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          input_data_in_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // input_data_in_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [102:0] input_data_in_translator_avalon_universal_slave_0_agent_rp_data;                          // input_data_in_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          input_data_in_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_001:sink_ready -> input_data_in_translator_avalon_universal_slave_0_agent:rp_ready
	wire          hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rp_valid;                   // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [102:0] hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rp_data;                    // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_002:sink_ready -> hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:rp_ready
	wire          input_data_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;               // input_data_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          input_data_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                     // input_data_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          input_data_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;             // input_data_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [102:0] input_data_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                      // input_data_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          input_data_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                     // id_router_003:sink_ready -> input_data_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          output_data_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // output_data_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          output_data_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                    // output_data_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          output_data_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // output_data_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [102:0] output_data_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                     // output_data_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          output_data_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_004:sink_ready -> output_data_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          rst_controller_reset_out_reset;                                                           // rst_controller:reset_out -> [addr_router:reset, cmd_xbar_demux:reset, hh_core_0:reset, hh_core_0_ctrl_port_translator:reset, hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:reset, hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, input_data:reset_n, input_data_in_csr_translator:reset, input_data_in_csr_translator_avalon_universal_slave_0_agent:reset, input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, input_data_in_translator:reset, input_data_in_translator_avalon_universal_slave_0_agent:reset, input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, output_data:reset_n, output_data_in_csr_translator:reset, output_data_in_csr_translator_avalon_universal_slave_0_agent:reset, output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, output_data_out_translator:reset, output_data_out_translator_avalon_universal_slave_0_agent:reset, output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ports2avalon_0_master_translator:reset, ports2avalon_0_master_translator_avalon_universal_master_0_agent:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_mux:reset, timing_adapter:reset_n, timing_adapter_1:reset_n]
	wire          cmd_xbar_demux_src0_endofpacket;                                                          // cmd_xbar_demux:src0_endofpacket -> output_data_out_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                // cmd_xbar_demux:src0_valid -> output_data_out_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                        // cmd_xbar_demux:src0_startofpacket -> output_data_out_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_src0_data;                                                                 // cmd_xbar_demux:src0_data -> output_data_out_translator_avalon_universal_slave_0_agent:cp_data
	wire    [4:0] cmd_xbar_demux_src0_channel;                                                              // cmd_xbar_demux:src0_channel -> output_data_out_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_src1_endofpacket;                                                          // cmd_xbar_demux:src1_endofpacket -> input_data_in_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                // cmd_xbar_demux:src1_valid -> input_data_in_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                        // cmd_xbar_demux:src1_startofpacket -> input_data_in_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_src1_data;                                                                 // cmd_xbar_demux:src1_data -> input_data_in_translator_avalon_universal_slave_0_agent:cp_data
	wire    [4:0] cmd_xbar_demux_src1_channel;                                                              // cmd_xbar_demux:src1_channel -> input_data_in_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_src2_endofpacket;                                                          // cmd_xbar_demux:src2_endofpacket -> hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                // cmd_xbar_demux:src2_valid -> hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                        // cmd_xbar_demux:src2_startofpacket -> hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_src2_data;                                                                 // cmd_xbar_demux:src2_data -> hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:cp_data
	wire    [4:0] cmd_xbar_demux_src2_channel;                                                              // cmd_xbar_demux:src2_channel -> hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_src3_endofpacket;                                                          // cmd_xbar_demux:src3_endofpacket -> input_data_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src3_valid;                                                                // cmd_xbar_demux:src3_valid -> input_data_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src3_startofpacket;                                                        // cmd_xbar_demux:src3_startofpacket -> input_data_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_src3_data;                                                                 // cmd_xbar_demux:src3_data -> input_data_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire    [4:0] cmd_xbar_demux_src3_channel;                                                              // cmd_xbar_demux:src3_channel -> input_data_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_src4_endofpacket;                                                          // cmd_xbar_demux:src4_endofpacket -> output_data_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src4_valid;                                                                // cmd_xbar_demux:src4_valid -> output_data_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src4_startofpacket;                                                        // cmd_xbar_demux:src4_startofpacket -> output_data_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_src4_data;                                                                 // cmd_xbar_demux:src4_data -> output_data_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire    [4:0] cmd_xbar_demux_src4_channel;                                                              // cmd_xbar_demux:src4_channel -> output_data_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                          // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                        // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [102:0] rsp_xbar_demux_src0_data;                                                                 // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire    [4:0] rsp_xbar_demux_src0_channel;                                                              // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                      // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                            // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                    // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [102:0] rsp_xbar_demux_001_src0_data;                                                             // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire    [4:0] rsp_xbar_demux_001_src0_channel;                                                          // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                            // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                      // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                            // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                    // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [102:0] rsp_xbar_demux_002_src0_data;                                                             // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire    [4:0] rsp_xbar_demux_002_src0_channel;                                                          // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                            // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                      // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                            // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                    // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [102:0] rsp_xbar_demux_003_src0_data;                                                             // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire    [4:0] rsp_xbar_demux_003_src0_channel;                                                          // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                            // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                      // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                            // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                    // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [102:0] rsp_xbar_demux_004_src0_data;                                                             // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire    [4:0] rsp_xbar_demux_004_src0_channel;                                                          // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                            // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          addr_router_src_endofpacket;                                                              // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          addr_router_src_valid;                                                                    // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire          addr_router_src_startofpacket;                                                            // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [102:0] addr_router_src_data;                                                                     // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire    [4:0] addr_router_src_channel;                                                                  // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire          addr_router_src_ready;                                                                    // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                             // rsp_xbar_mux:src_endofpacket -> ports2avalon_0_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                   // rsp_xbar_mux:src_valid -> ports2avalon_0_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                           // rsp_xbar_mux:src_startofpacket -> ports2avalon_0_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [102:0] rsp_xbar_mux_src_data;                                                                    // rsp_xbar_mux:src_data -> ports2avalon_0_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [4:0] rsp_xbar_mux_src_channel;                                                                 // rsp_xbar_mux:src_channel -> ports2avalon_0_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_src_ready;                                                                   // ports2avalon_0_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire          cmd_xbar_demux_src0_ready;                                                                // output_data_out_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src0_ready
	wire          id_router_src_endofpacket;                                                                // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                      // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                              // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [102:0] id_router_src_data;                                                                       // id_router:src_data -> rsp_xbar_demux:sink_data
	wire    [4:0] id_router_src_channel;                                                                    // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                      // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_demux_src1_ready;                                                                // input_data_in_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src1_ready
	wire          id_router_001_src_endofpacket;                                                            // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                  // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                          // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [102:0] id_router_001_src_data;                                                                   // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire    [4:0] id_router_001_src_channel;                                                                // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                  // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_demux_src2_ready;                                                                // hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src2_ready
	wire          id_router_002_src_endofpacket;                                                            // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                  // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                          // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [102:0] id_router_002_src_data;                                                                   // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire    [4:0] id_router_002_src_channel;                                                                // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                  // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_demux_src3_ready;                                                                // input_data_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src3_ready
	wire          id_router_003_src_endofpacket;                                                            // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                  // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                          // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [102:0] id_router_003_src_data;                                                                   // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire    [4:0] id_router_003_src_channel;                                                                // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                  // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_src4_ready;                                                                // output_data_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src4_ready
	wire          id_router_004_src_endofpacket;                                                            // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                  // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                          // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [102:0] id_router_004_src_data;                                                                   // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire    [4:0] id_router_004_src_channel;                                                                // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                  // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready

	hh_core hh_core_0 (
		.clk           (clk_clk),                                                        //             clock.clk
		.reset         (rst_controller_reset_out_reset),                                 //             reset.reset
		.i_writedata   (hh_core_0_ctrl_port_translator_avalon_anti_slave_0_writedata),   //         ctrl_port.writedata
		.i_address     (hh_core_0_ctrl_port_translator_avalon_anti_slave_0_address),     //                  .address
		.o_readdata    (hh_core_0_ctrl_port_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.i_read        (hh_core_0_ctrl_port_translator_avalon_anti_slave_0_read),        //                  .read
		.i_write       (hh_core_0_ctrl_port_translator_avalon_anti_slave_0_write),       //                  .write
		.o_waitrequest (hh_core_0_ctrl_port_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.i_data        (timing_adapter_1_out_data),                                      //    inputdata_sink.data
		.o_ready       (timing_adapter_1_out_ready),                                     //                  .ready
		.i_valid       (timing_adapter_1_out_valid),                                     //                  .valid
		.o_data        (hh_core_0_outputdata_source_data),                               // outputdata_source.data
		.i_ready       (hh_core_0_outputdata_source_ready),                              //                  .ready
		.o_valid       (hh_core_0_outputdata_source_valid)                               //                  .valid
	);

	ports2avalon #(
		.ADDRESS_WIDTH (32)
	) ports2avalon_0 (
		.clk                 (clk_clk),                            //  clock.clk
		.reset_n             (reset_reset_n),                      //  reset.reset_n
		.address             (ports2avalon_0_master_address),      // master.address
		.read                (ports2avalon_0_master_read),         //       .read
		.readdata            (ports2avalon_0_master_readdata),     //       .readdata
		.write               (ports2avalon_0_master_write),        //       .write
		.writedata           (ports2avalon_0_master_writedata),    //       .writedata
		.waitrequest         (ports2avalon_0_master_waitrequest),  //       .waitrequest
		.usb_address         (ports2avalon_0_usb_address),         //    usb.export
		.usb_address_ready   (ports2avalon_0_usb_address_ready),   //       .export
		.usb_writedata       (ports2avalon_0_usb_writedata),       //       .export
		.usb_writedata_ready (ports2avalon_0_usb_writedata_ready), //       .export
		.usb_readdata        (ports2avalon_0_usb_readdata),        //       .export
		.usb_readdata_ready  (ports2avalon_0_usb_readdata_ready),  //       .export
		.usb_address_want    (ports2avalon_0_usb_address_want),    //       .export
		.usb_writedata_want  (ports2avalon_0_usb_writedata_want),  //       .export
		.usb_readdata_want   (ports2avalon_0_usb_readdata_want)    //       .export
	);

	hh_system_input_data input_data (
		.wrclock                          (clk_clk),                                                    //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),                            // reset_in.reset_n
		.avalonmm_write_slave_writedata   (input_data_in_translator_avalon_anti_slave_0_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (input_data_in_translator_avalon_anti_slave_0_write),         //         .write
		.avalonmm_write_slave_address     (input_data_in_translator_avalon_anti_slave_0_address),       //         .address
		.avalonmm_write_slave_waitrequest (input_data_in_translator_avalon_anti_slave_0_waitrequest),   //         .waitrequest
		.wrclk_control_slave_address      (input_data_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read         (input_data_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata    (input_data_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write        (input_data_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata     (input_data_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.avalonst_source_valid            (input_data_out_valid),                                       //      out.valid
		.avalonst_source_data             (input_data_out_data),                                        //         .data
		.avalonst_source_ready            (input_data_out_ready)                                        //         .ready
	);

	hh_system_output_data output_data (
		.wrclock                         (clk_clk),                                                     //   clk_in.clk
		.reset_n                         (~rst_controller_reset_out_reset),                             // reset_in.reset_n
		.avalonst_sink_valid             (timing_adapter_out_valid),                                    //       in.valid
		.avalonst_sink_data              (timing_adapter_out_data),                                     //         .data
		.avalonst_sink_ready             (timing_adapter_out_ready),                                    //         .ready
		.wrclk_control_slave_address     (output_data_in_csr_translator_avalon_anti_slave_0_address),   //   in_csr.address
		.wrclk_control_slave_read        (output_data_in_csr_translator_avalon_anti_slave_0_read),      //         .read
		.wrclk_control_slave_writedata   (output_data_in_csr_translator_avalon_anti_slave_0_writedata), //         .writedata
		.wrclk_control_slave_write       (output_data_in_csr_translator_avalon_anti_slave_0_write),     //         .write
		.wrclk_control_slave_readdata    (output_data_in_csr_translator_avalon_anti_slave_0_readdata),  //         .readdata
		.wrclk_control_slave_irq         (),                                                            //   in_irq.irq
		.avalonmm_read_slave_readdata    (output_data_out_translator_avalon_anti_slave_0_readdata),     //      out.readdata
		.avalonmm_read_slave_read        (output_data_out_translator_avalon_anti_slave_0_read),         //         .read
		.avalonmm_read_slave_address     (output_data_out_translator_avalon_anti_slave_0_address),      //         .address
		.avalonmm_read_slave_waitrequest (output_data_out_translator_avalon_anti_slave_0_waitrequest)   //         .waitrequest
	);

	hh_system_timing_adapter timing_adapter (
		.clk       (clk_clk),                           //   clk.clk
		.reset_n   (~rst_controller_reset_out_reset),   // reset.reset_n
		.in_ready  (hh_core_0_outputdata_source_ready), //    in.ready
		.in_valid  (hh_core_0_outputdata_source_valid), //      .valid
		.in_data   (hh_core_0_outputdata_source_data),  //      .data
		.out_ready (timing_adapter_out_ready),          //   out.ready
		.out_valid (timing_adapter_out_valid),          //      .valid
		.out_data  (timing_adapter_out_data)            //      .data
	);

	hh_system_timing_adapter_1 timing_adapter_1 (
		.clk       (clk_clk),                         //   clk.clk
		.reset_n   (~rst_controller_reset_out_reset), // reset.reset_n
		.in_ready  (input_data_out_ready),            //    in.ready
		.in_valid  (input_data_out_valid),            //      .valid
		.in_data   (input_data_out_data),             //      .data
		.out_ready (timing_adapter_1_out_ready),      //   out.ready
		.out_valid (timing_adapter_1_out_valid),      //      .valid
		.out_data  (timing_adapter_1_out_data)        //      .data
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) ports2avalon_0_master_translator (
		.clk                   (clk_clk),                                                                  //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                           //                     reset.reset
		.uav_address           (ports2avalon_0_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (ports2avalon_0_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (ports2avalon_0_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (ports2avalon_0_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (ports2avalon_0_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (ports2avalon_0_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (ports2avalon_0_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (ports2avalon_0_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (ports2avalon_0_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (ports2avalon_0_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (ports2avalon_0_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (ports2avalon_0_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (ports2avalon_0_master_waitrequest),                                        //                          .waitrequest
		.av_read               (ports2avalon_0_master_read),                                               //                          .read
		.av_readdata           (ports2avalon_0_master_readdata),                                           //                          .readdata
		.av_write              (ports2avalon_0_master_write),                                              //                          .write
		.av_writedata          (ports2avalon_0_master_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                     //               (terminated)
		.av_byteenable         (4'b1111),                                                                  //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                     //               (terminated)
		.av_begintransfer      (1'b0),                                                                     //               (terminated)
		.av_chipselect         (1'b0),                                                                     //               (terminated)
		.av_readdatavalid      (),                                                                         //               (terminated)
		.av_lock               (1'b0),                                                                     //               (terminated)
		.av_debugaccess        (1'b0),                                                                     //               (terminated)
		.uav_clken             (),                                                                         //               (terminated)
		.av_clken              (1'b1)                                                                      //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) output_data_out_translator (
		.clk                   (clk_clk),                                                                    //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                             //                    reset.reset
		.uav_address           (output_data_out_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (output_data_out_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (output_data_out_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (output_data_out_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (output_data_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (output_data_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (output_data_out_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (output_data_out_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (output_data_out_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (output_data_out_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (output_data_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (output_data_out_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_read               (output_data_out_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (output_data_out_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (output_data_out_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_write              (),                                                                           //              (terminated)
		.av_writedata          (),                                                                           //              (terminated)
		.av_begintransfer      (),                                                                           //              (terminated)
		.av_beginbursttransfer (),                                                                           //              (terminated)
		.av_burstcount         (),                                                                           //              (terminated)
		.av_byteenable         (),                                                                           //              (terminated)
		.av_readdatavalid      (1'b0),                                                                       //              (terminated)
		.av_writebyteenable    (),                                                                           //              (terminated)
		.av_lock               (),                                                                           //              (terminated)
		.av_chipselect         (),                                                                           //              (terminated)
		.av_clken              (),                                                                           //              (terminated)
		.uav_clken             (1'b0),                                                                       //              (terminated)
		.av_debugaccess        (),                                                                           //              (terminated)
		.av_outputenable       ()                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) input_data_in_translator (
		.clk                   (clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address           (input_data_in_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (input_data_in_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (input_data_in_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (input_data_in_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (input_data_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (input_data_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (input_data_in_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (input_data_in_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (input_data_in_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (input_data_in_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (input_data_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (input_data_in_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (input_data_in_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_writedata          (input_data_in_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (input_data_in_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_read               (),                                                                         //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                     //              (terminated)
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hh_core_0_ctrl_port_translator (
		.clk                   (clk_clk),                                                                        //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (hh_core_0_ctrl_port_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (hh_core_0_ctrl_port_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (hh_core_0_ctrl_port_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (hh_core_0_ctrl_port_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (hh_core_0_ctrl_port_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (hh_core_0_ctrl_port_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_byteenable         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.av_chipselect         (),                                                                               //              (terminated)
		.av_clken              (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) input_data_in_csr_translator (
		.clk                   (clk_clk),                                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                               //                    reset.reset
		.uav_address           (input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (input_data_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (input_data_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (input_data_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (input_data_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (input_data_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) output_data_in_csr_translator (
		.clk                   (clk_clk),                                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                //                    reset.reset
		.uav_address           (output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (output_data_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (output_data_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (output_data_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (output_data_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (output_data_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_waitrequest        (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_BEGIN_BURST           (86),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (90),
		.PKT_THREAD_ID_H           (93),
		.PKT_THREAD_ID_L           (93),
		.PKT_CACHE_H               (100),
		.PKT_CACHE_L               (97),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.ST_DATA_W                 (103),
		.ST_CHANNEL_W              (5),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) ports2avalon_0_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                           //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.av_address       (ports2avalon_0_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (ports2avalon_0_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (ports2avalon_0_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (ports2avalon_0_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (ports2avalon_0_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (ports2avalon_0_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (ports2avalon_0_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (ports2avalon_0_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (ports2avalon_0_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (ports2avalon_0_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (ports2avalon_0_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (ports2avalon_0_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (ports2avalon_0_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (ports2avalon_0_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (ports2avalon_0_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (ports2avalon_0_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_src_valid),                                                            //        rp.valid
		.rp_data          (rsp_xbar_mux_src_data),                                                             //          .data
		.rp_channel       (rsp_xbar_mux_src_channel),                                                          //          .channel
		.rp_startofpacket (rsp_xbar_mux_src_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_src_endofpacket),                                                      //          .endofpacket
		.rp_ready         (rsp_xbar_mux_src_ready)                                                             //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (90),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) output_data_out_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (output_data_out_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (output_data_out_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (output_data_out_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (output_data_out_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (output_data_out_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (output_data_out_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (output_data_out_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (output_data_out_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (output_data_out_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (output_data_out_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (output_data_out_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (output_data_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (output_data_out_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (output_data_out_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (output_data_out_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (output_data_out_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src0_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_src0_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_src0_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_src0_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src0_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src0_channel),                                                          //                .channel
		.rf_sink_ready           (output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (output_data_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (output_data_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (output_data_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (output_data_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (output_data_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (output_data_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (output_data_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (output_data_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (output_data_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (output_data_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (output_data_out_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (output_data_out_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (output_data_out_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (output_data_out_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (output_data_out_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (output_data_out_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (output_data_out_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (90),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) input_data_in_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (input_data_in_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (input_data_in_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (input_data_in_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (input_data_in_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (input_data_in_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (input_data_in_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (input_data_in_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (input_data_in_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (input_data_in_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (input_data_in_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (input_data_in_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (input_data_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (input_data_in_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (input_data_in_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (input_data_in_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (input_data_in_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src1_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_src1_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_src1_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_src1_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src1_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src1_channel),                                                        //                .channel
		.rf_sink_ready           (input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (input_data_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (input_data_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (input_data_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (input_data_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (input_data_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (input_data_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (input_data_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (input_data_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (input_data_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (input_data_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (input_data_in_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (input_data_in_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (input_data_in_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (input_data_in_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (input_data_in_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (input_data_in_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (input_data_in_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (90),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src2_ready),                                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_src2_valid),                                                                //                .valid
		.cp_data                 (cmd_xbar_demux_src2_data),                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_src2_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src2_endofpacket),                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src2_channel),                                                              //                .channel
		.rf_sink_ready           (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (90),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) input_data_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (input_data_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (input_data_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (input_data_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (input_data_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (input_data_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (input_data_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src3_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_src3_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_src3_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_src3_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src3_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src3_channel),                                                            //                .channel
		.rf_sink_ready           (input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (input_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (input_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (input_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (input_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (input_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (input_data_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (input_data_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (input_data_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (input_data_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (input_data_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (input_data_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (input_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (input_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (input_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (input_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (input_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (input_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (86),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (89),
		.PKT_SRC_ID_L              (87),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (90),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) output_data_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (output_data_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (output_data_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (output_data_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (output_data_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (output_data_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (output_data_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src4_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_src4_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_demux_src4_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_src4_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src4_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src4_channel),                                                             //                .channel
		.rf_sink_ready           (output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (output_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (output_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (output_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (output_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (output_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (output_data_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (output_data_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (output_data_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (output_data_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (output_data_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (output_data_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (output_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (output_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (output_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (output_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (output_data_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (output_data_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	hh_system_addr_router addr_router (
		.sink_ready         (ports2avalon_0_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (ports2avalon_0_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (ports2avalon_0_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (ports2avalon_0_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ports2avalon_0_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_src_valid),                                                             //          .valid
		.src_data           (addr_router_src_data),                                                              //          .data
		.src_channel        (addr_router_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                        //          .endofpacket
	);

	hh_system_id_router id_router (
		.sink_ready         (output_data_out_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (output_data_out_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (output_data_out_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (output_data_out_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (output_data_out_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                        //       src.ready
		.src_valid          (id_router_src_valid),                                                        //          .valid
		.src_data           (id_router_src_data),                                                         //          .data
		.src_channel        (id_router_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                   //          .endofpacket
	);

	hh_system_id_router id_router_001 (
		.sink_ready         (input_data_in_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (input_data_in_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (input_data_in_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (input_data_in_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (input_data_in_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                  //       src.ready
		.src_valid          (id_router_001_src_valid),                                                  //          .valid
		.src_data           (id_router_001_src_data),                                                   //          .data
		.src_channel        (id_router_001_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                             //          .endofpacket
	);

	hh_system_id_router id_router_002 (
		.sink_ready         (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hh_core_0_ctrl_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                        //       src.ready
		.src_valid          (id_router_002_src_valid),                                                        //          .valid
		.src_data           (id_router_002_src_data),                                                         //          .data
		.src_channel        (id_router_002_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                   //          .endofpacket
	);

	hh_system_id_router id_router_003 (
		.sink_ready         (input_data_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (input_data_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (input_data_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (input_data_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (input_data_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                      //       src.ready
		.src_valid          (id_router_003_src_valid),                                                      //          .valid
		.src_data           (id_router_003_src_data),                                                       //          .data
		.src_channel        (id_router_003_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                 //          .endofpacket
	);

	hh_system_id_router id_router_004 (
		.sink_ready         (output_data_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (output_data_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (output_data_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (output_data_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (output_data_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                       //       src.ready
		.src_valid          (id_router_004_src_valid),                                                       //          .valid
		.src_data           (id_router_004_src_data),                                                        //          .data
		.src_channel        (id_router_004_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                  //          .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	hh_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket),   //          .endofpacket
		.src4_ready         (cmd_xbar_demux_src4_ready),         //      src4.ready
		.src4_valid         (cmd_xbar_demux_src4_valid),         //          .valid
		.src4_data          (cmd_xbar_demux_src4_data),          //          .data
		.src4_channel       (cmd_xbar_demux_src4_channel),       //          .channel
		.src4_startofpacket (cmd_xbar_demux_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_src4_endofpacket)    //          .endofpacket
	);

	hh_system_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)    //          .endofpacket
	);

	hh_system_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	hh_system_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	hh_system_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	hh_system_rsp_xbar_demux rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	hh_system_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

endmodule
