//`timescale 1 ps/ 1 ps 
///////////////////////////////////////////////////////////////// 
// Company: 
// Engineer: 
// Create Date: 2022-06-22 14:14:28
// Design Name: 
// Module Name: i2c_master_defines
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision: 
// Additional Comments:
// 
///////////////////////////////////////////////////////////////// 

`define I2C_CMD_NOP   4'b0000
`define I2C_CMD_START 4'b0001
`define I2C_CMD_STOP  4'b0010
`define I2C_CMD_WRITE 4'b0100
`define I2C_CMD_READ  4'b1000


