
module co_sim_tdp_256x16;

    reg clkA, clkB, weA, weB;
    reg [3:0] addrA, addrB;
    reg [255:0] dinA, dinB;
    wire [255:0] doutA, doutB, doutA_net, doutB_net;

    integer mismatch=0;
    reg [6:0]cycle, i;

    tdp_256x16 golden(.*);
    `ifdef PNR
        tdp_256x16_post_route netlist( clkA ,
    clkB ,
    weA ,
    weB ,
    addrA[0] ,
    addrA[1] ,
    addrA[2] ,
    addrA[3] ,
    addrB[0] ,
    addrB[1] ,
    addrB[2] ,
    addrB[3] ,
    dinA[0] ,
    dinA[1] ,
    dinA[2] ,
    dinA[3] ,
    dinA[4] ,
    dinA[5] ,
    dinA[6] ,
    dinA[7] ,
    dinA[8] ,
    dinA[9] ,
    dinA[10] ,
    dinA[11] ,
    dinA[12] ,
    dinA[13] ,
    dinA[14] ,
    dinA[15] ,
    dinA[16] ,
    dinA[17] ,
    dinA[18] ,
    dinA[19] ,
    dinA[20] ,
    dinA[21] ,
    dinA[22] ,
    dinA[23] ,
    dinA[24] ,
    dinA[25] ,
    dinA[26] ,
    dinA[27] ,
    dinA[28] ,
    dinA[29] ,
    dinA[30] ,
    dinA[31] ,
    dinA[32] ,
    dinA[33] ,
    dinA[34] ,
    dinA[35] ,
    dinA[36] ,
    dinA[37] ,
    dinA[38] ,
    dinA[39] ,
    dinA[40] ,
    dinA[41] ,
    dinA[42] ,
    dinA[43] ,
    dinA[44] ,
    dinA[45] ,
    dinA[46] ,
    dinA[47] ,
    dinA[48] ,
    dinA[49] ,
    dinA[50] ,
    dinA[51] ,
    dinA[52] ,
    dinA[53] ,
    dinA[54] ,
    dinA[55] ,
    dinA[56] ,
    dinA[57] ,
    dinA[58] ,
    dinA[59] ,
    dinA[60] ,
    dinA[61] ,
    dinA[62] ,
    dinA[63] ,
    dinA[64] ,
    dinA[65] ,
    dinA[66] ,
    dinA[67] ,
    dinA[68] ,
    dinA[69] ,
    dinA[70] ,
    dinA[71] ,
    dinA[72] ,
    dinA[73] ,
    dinA[74] ,
    dinA[75] ,
    dinA[76] ,
    dinA[77] ,
    dinA[78] ,
    dinA[79] ,
    dinA[80] ,
    dinA[81] ,
    dinA[82] ,
    dinA[83] ,
    dinA[84] ,
    dinA[85] ,
    dinA[86] ,
    dinA[87] ,
    dinA[88] ,
    dinA[89] ,
    dinA[90] ,
    dinA[91] ,
    dinA[92] ,
    dinA[93] ,
    dinA[94] ,
    dinA[95] ,
    dinA[96] ,
    dinA[97] ,
    dinA[98] ,
    dinA[99] ,
    dinA[100] ,
    dinA[101] ,
    dinA[102] ,
    dinA[103] ,
    dinA[104] ,
    dinA[105] ,
    dinA[106] ,
    dinA[107] ,
    dinA[108] ,
    dinA[109] ,
    dinA[110] ,
    dinA[111] ,
    dinA[112] ,
    dinA[113] ,
    dinA[114] ,
    dinA[115] ,
    dinA[116] ,
    dinA[117] ,
    dinA[118] ,
    dinA[119] ,
    dinA[120] ,
    dinA[121] ,
    dinA[122] ,
    dinA[123] ,
    dinA[124] ,
    dinA[125] ,
    dinA[126] ,
    dinA[127] ,
    dinA[128] ,
    dinA[129] ,
    dinA[130] ,
    dinA[131] ,
    dinA[132] ,
    dinA[133] ,
    dinA[134] ,
    dinA[135] ,
    dinA[136] ,
    dinA[137] ,
    dinA[138] ,
    dinA[139] ,
    dinA[140] ,
    dinA[141] ,
    dinA[142] ,
    dinA[143] ,
    dinA[144] ,
    dinA[145] ,
    dinA[146] ,
    dinA[147] ,
    dinA[148] ,
    dinA[149] ,
    dinA[150] ,
    dinA[151] ,
    dinA[152] ,
    dinA[153] ,
    dinA[154] ,
    dinA[155] ,
    dinA[156] ,
    dinA[157] ,
    dinA[158] ,
    dinA[159] ,
    dinA[160] ,
    dinA[161] ,
    dinA[162] ,
    dinA[163] ,
    dinA[164] ,
    dinA[165] ,
    dinA[166] ,
    dinA[167] ,
    dinA[168] ,
    dinA[169] ,
    dinA[170] ,
    dinA[171] ,
    dinA[172] ,
    dinA[173] ,
    dinA[174] ,
    dinA[175] ,
    dinA[176] ,
    dinA[177] ,
    dinA[178] ,
    dinA[179] ,
    dinA[180] ,
    dinA[181] ,
    dinA[182] ,
    dinA[183] ,
    dinA[184] ,
    dinA[185] ,
    dinA[186] ,
    dinA[187] ,
    dinA[188] ,
    dinA[189] ,
    dinA[190] ,
    dinA[191] ,
    dinA[192] ,
    dinA[193] ,
    dinA[194] ,
    dinA[195] ,
    dinA[196] ,
    dinA[197] ,
    dinA[198] ,
    dinA[199] ,
    dinA[200] ,
    dinA[201] ,
    dinA[202] ,
    dinA[203] ,
    dinA[204] ,
    dinA[205] ,
    dinA[206] ,
    dinA[207] ,
    dinA[208] ,
    dinA[209] ,
    dinA[210] ,
    dinA[211] ,
    dinA[212] ,
    dinA[213] ,
    dinA[214] ,
    dinA[215] ,
    dinA[216] ,
    dinA[217] ,
    dinA[218] ,
    dinA[219] ,
    dinA[220] ,
    dinA[221] ,
    dinA[222] ,
    dinA[223] ,
    dinA[224] ,
    dinA[225] ,
    dinA[226] ,
    dinA[227] ,
    dinA[228] ,
    dinA[229] ,
    dinA[230] ,
    dinA[231] ,
    dinA[232] ,
    dinA[233] ,
    dinA[234] ,
    dinA[235] ,
    dinA[236] ,
    dinA[237] ,
    dinA[238] ,
    dinA[239] ,
    dinA[240] ,
    dinA[241] ,
    dinA[242] ,
    dinA[243] ,
    dinA[244] ,
    dinA[245] ,
    dinA[246] ,
    dinA[247] ,
    dinA[248] ,
    dinA[249] ,
    dinA[250] ,
    dinA[251] ,
    dinA[252] ,
    dinA[253] ,
    dinA[254] ,
    dinA[255] ,
    dinB[0] ,
    dinB[1] ,
    dinB[2] ,
    dinB[3] ,
    dinB[4] ,
    dinB[5] ,
    dinB[6] ,
    dinB[7] ,
    dinB[8] ,
    dinB[9] ,
    dinB[10] ,
    dinB[11] ,
    dinB[12] ,
    dinB[13] ,
    dinB[14] ,
    dinB[15] ,
    dinB[16] ,
    dinB[17] ,
    dinB[18] ,
    dinB[19] ,
    dinB[20] ,
    dinB[21] ,
    dinB[22] ,
    dinB[23] ,
    dinB[24] ,
    dinB[25] ,
    dinB[26] ,
    dinB[27] ,
    dinB[28] ,
    dinB[29] ,
    dinB[30] ,
    dinB[31] ,
    dinB[32] ,
    dinB[33] ,
    dinB[34] ,
    dinB[35] ,
    dinB[36] ,
    dinB[37] ,
    dinB[38] ,
    dinB[39] ,
    dinB[40] ,
    dinB[41] ,
    dinB[42] ,
    dinB[43] ,
    dinB[44] ,
    dinB[45] ,
    dinB[46] ,
    dinB[47] ,
    dinB[48] ,
    dinB[49] ,
    dinB[50] ,
    dinB[51] ,
    dinB[52] ,
    dinB[53] ,
    dinB[54] ,
    dinB[55] ,
    dinB[56] ,
    dinB[57] ,
    dinB[58] ,
    dinB[59] ,
    dinB[60] ,
    dinB[61] ,
    dinB[62] ,
    dinB[63] ,
    dinB[64] ,
    dinB[65] ,
    dinB[66] ,
    dinB[67] ,
    dinB[68] ,
    dinB[69] ,
    dinB[70] ,
    dinB[71] ,
    dinB[72] ,
    dinB[73] ,
    dinB[74] ,
    dinB[75] ,
    dinB[76] ,
    dinB[77] ,
    dinB[78] ,
    dinB[79] ,
    dinB[80] ,
    dinB[81] ,
    dinB[82] ,
    dinB[83] ,
    dinB[84] ,
    dinB[85] ,
    dinB[86] ,
    dinB[87] ,
    dinB[88] ,
    dinB[89] ,
    dinB[90] ,
    dinB[91] ,
    dinB[92] ,
    dinB[93] ,
    dinB[94] ,
    dinB[95] ,
    dinB[96] ,
    dinB[97] ,
    dinB[98] ,
    dinB[99] ,
    dinB[100] ,
    dinB[101] ,
    dinB[102] ,
    dinB[103] ,
    dinB[104] ,
    dinB[105] ,
    dinB[106] ,
    dinB[107] ,
    dinB[108] ,
    dinB[109] ,
    dinB[110] ,
    dinB[111] ,
    dinB[112] ,
    dinB[113] ,
    dinB[114] ,
    dinB[115] ,
    dinB[116] ,
    dinB[117] ,
    dinB[118] ,
    dinB[119] ,
    dinB[120] ,
    dinB[121] ,
    dinB[122] ,
    dinB[123] ,
    dinB[124] ,
    dinB[125] ,
    dinB[126] ,
    dinB[127] ,
    dinB[128] ,
    dinB[129] ,
    dinB[130] ,
    dinB[131] ,
    dinB[132] ,
    dinB[133] ,
    dinB[134] ,
    dinB[135] ,
    dinB[136] ,
    dinB[137] ,
    dinB[138] ,
    dinB[139] ,
    dinB[140] ,
    dinB[141] ,
    dinB[142] ,
    dinB[143] ,
    dinB[144] ,
    dinB[145] ,
    dinB[146] ,
    dinB[147] ,
    dinB[148] ,
    dinB[149] ,
    dinB[150] ,
    dinB[151] ,
    dinB[152] ,
    dinB[153] ,
    dinB[154] ,
    dinB[155] ,
    dinB[156] ,
    dinB[157] ,
    dinB[158] ,
    dinB[159] ,
    dinB[160] ,
    dinB[161] ,
    dinB[162] ,
    dinB[163] ,
    dinB[164] ,
    dinB[165] ,
    dinB[166] ,
    dinB[167] ,
    dinB[168] ,
    dinB[169] ,
    dinB[170] ,
    dinB[171] ,
    dinB[172] ,
    dinB[173] ,
    dinB[174] ,
    dinB[175] ,
    dinB[176] ,
    dinB[177] ,
    dinB[178] ,
    dinB[179] ,
    dinB[180] ,
    dinB[181] ,
    dinB[182] ,
    dinB[183] ,
    dinB[184] ,
    dinB[185] ,
    dinB[186] ,
    dinB[187] ,
    dinB[188] ,
    dinB[189] ,
    dinB[190] ,
    dinB[191] ,
    dinB[192] ,
    dinB[193] ,
    dinB[194] ,
    dinB[195] ,
    dinB[196] ,
    dinB[197] ,
    dinB[198] ,
    dinB[199] ,
    dinB[200] ,
    dinB[201] ,
    dinB[202] ,
    dinB[203] ,
    dinB[204] ,
    dinB[205] ,
    dinB[206] ,
    dinB[207] ,
    dinB[208] ,
    dinB[209] ,
    dinB[210] ,
    dinB[211] ,
    dinB[212] ,
    dinB[213] ,
    dinB[214] ,
    dinB[215] ,
    dinB[216] ,
    dinB[217] ,
    dinB[218] ,
    dinB[219] ,
    dinB[220] ,
    dinB[221] ,
    dinB[222] ,
    dinB[223] ,
    dinB[224] ,
    dinB[225] ,
    dinB[226] ,
    dinB[227] ,
    dinB[228] ,
    dinB[229] ,
    dinB[230] ,
    dinB[231] ,
    dinB[232] ,
    dinB[233] ,
    dinB[234] ,
    dinB[235] ,
    dinB[236] ,
    dinB[237] ,
    dinB[238] ,
    dinB[239] ,
    dinB[240] ,
    dinB[241] ,
    dinB[242] ,
    dinB[243] ,
    dinB[244] ,
    dinB[245] ,
    dinB[246] ,
    dinB[247] ,
    dinB[248] ,
    dinB[249] ,
    dinB[250] ,
    dinB[251] ,
    dinB[252] ,
    dinB[253] ,
    dinB[254] ,
    dinB[255] ,
    doutA_net[0] ,
    doutB_net[255] ,
    doutA_net[1] ,
    doutA_net[2] ,
    doutA_net[3] ,
    doutA_net[4] ,
    doutA_net[5] ,
    doutA_net[6] ,
    doutA_net[7] ,
    doutA_net[8] ,
    doutA_net[9] ,
    doutA_net[10] ,
    doutA_net[11] ,
    doutA_net[12] ,
    doutA_net[13] ,
    doutA_net[14] ,
    doutA_net[15] ,
    doutA_net[16] ,
    doutA_net[17] ,
    doutA_net[36] ,
    doutA_net[37] ,
    doutA_net[38] ,
    doutA_net[39] ,
    doutA_net[40] ,
    doutA_net[41] ,
    doutA_net[42] ,
    doutA_net[43] ,
    doutA_net[44] ,
    doutA_net[45] ,
    doutA_net[46] ,
    doutA_net[47] ,
    doutA_net[48] ,
    doutA_net[49] ,
    doutA_net[50] ,
    doutA_net[51] ,
    doutA_net[52] ,
    doutA_net[53] ,
    doutA_net[72] ,
    doutA_net[73] ,
    doutA_net[74] ,
    doutA_net[75] ,
    doutA_net[76] ,
    doutA_net[77] ,
    doutA_net[78] ,
    doutA_net[79] ,
    doutA_net[80] ,
    doutA_net[81] ,
    doutA_net[82] ,
    doutA_net[83] ,
    doutA_net[84] ,
    doutA_net[85] ,
    doutA_net[86] ,
    doutA_net[87] ,
    doutA_net[88] ,
    doutA_net[89] ,
    doutA_net[108] ,
    doutA_net[109] ,
    doutA_net[110] ,
    doutA_net[111] ,
    doutA_net[112] ,
    doutA_net[113] ,
    doutA_net[114] ,
    doutA_net[115] ,
    doutA_net[116] ,
    doutA_net[117] ,
    doutA_net[118] ,
    doutA_net[119] ,
    doutA_net[120] ,
    doutA_net[121] ,
    doutA_net[122] ,
    doutA_net[123] ,
    doutA_net[124] ,
    doutA_net[125] ,
    doutA_net[144] ,
    doutA_net[145] ,
    doutA_net[146] ,
    doutA_net[147] ,
    doutA_net[148] ,
    doutA_net[149] ,
    doutA_net[150] ,
    doutA_net[151] ,
    doutA_net[152] ,
    doutA_net[153] ,
    doutA_net[154] ,
    doutA_net[155] ,
    doutA_net[156] ,
    doutA_net[157] ,
    doutA_net[158] ,
    doutA_net[159] ,
    doutA_net[160] ,
    doutA_net[161] ,
    doutA_net[180] ,
    doutA_net[181] ,
    doutA_net[182] ,
    doutA_net[183] ,
    doutA_net[184] ,
    doutA_net[185] ,
    doutA_net[186] ,
    doutA_net[187] ,
    doutA_net[188] ,
    doutA_net[189] ,
    doutA_net[190] ,
    doutA_net[191] ,
    doutA_net[192] ,
    doutA_net[193] ,
    doutA_net[194] ,
    doutA_net[195] ,
    doutA_net[196] ,
    doutA_net[197] ,
    doutA_net[216] ,
    doutA_net[217] ,
    doutA_net[218] ,
    doutA_net[219] ,
    doutA_net[220] ,
    doutA_net[221] ,
    doutA_net[222] ,
    doutA_net[223] ,
    doutA_net[224] ,
    doutA_net[225] ,
    doutA_net[226] ,
    doutA_net[227] ,
    doutA_net[228] ,
    doutA_net[229] ,
    doutA_net[230] ,
    doutA_net[231] ,
    doutA_net[232] ,
    doutA_net[233] ,
    doutA_net[252] ,
    doutA_net[253] ,
    doutA_net[254] ,
    doutA_net[255] ,
    doutB_net[0] ,
    doutB_net[1] ,
    doutB_net[2] ,
    doutB_net[3] ,
    doutB_net[4] ,
    doutB_net[5] ,
    doutB_net[6] ,
    doutB_net[7] ,
    doutB_net[8] ,
    doutB_net[9] ,
    doutB_net[10] ,
    doutB_net[11] ,
    doutB_net[12] ,
    doutB_net[13] ,
    doutB_net[14] ,
    doutB_net[15] ,
    doutB_net[16] ,
    doutB_net[17] ,
    doutB_net[36] ,
    doutB_net[37] ,
    doutB_net[38] ,
    doutB_net[39] ,
    doutB_net[40] ,
    doutB_net[41] ,
    doutB_net[42] ,
    doutB_net[43] ,
    doutB_net[44] ,
    doutB_net[45] ,
    doutB_net[46] ,
    doutB_net[47] ,
    doutB_net[48] ,
    doutB_net[49] ,
    doutB_net[50] ,
    doutB_net[51] ,
    doutB_net[52] ,
    doutB_net[53] ,
    doutB_net[72] ,
    doutB_net[73] ,
    doutB_net[74] ,
    doutB_net[75] ,
    doutB_net[76] ,
    doutB_net[77] ,
    doutB_net[78] ,
    doutB_net[79] ,
    doutB_net[80] ,
    doutB_net[81] ,
    doutB_net[82] ,
    doutB_net[83] ,
    doutB_net[84] ,
    doutB_net[85] ,
    doutB_net[86] ,
    doutB_net[87] ,
    doutB_net[88] ,
    doutB_net[89] ,
    doutB_net[108] ,
    doutB_net[109] ,
    doutB_net[110] ,
    doutB_net[111] ,
    doutB_net[112] ,
    doutB_net[113] ,
    doutB_net[114] ,
    doutB_net[115] ,
    doutB_net[116] ,
    doutB_net[117] ,
    doutB_net[118] ,
    doutB_net[119] ,
    doutB_net[120] ,
    doutB_net[121] ,
    doutB_net[122] ,
    doutB_net[123] ,
    doutB_net[124] ,
    doutB_net[125] ,
    doutB_net[144] ,
    doutB_net[145] ,
    doutB_net[146] ,
    doutB_net[147] ,
    doutB_net[148] ,
    doutB_net[149] ,
    doutB_net[150] ,
    doutB_net[151] ,
    doutB_net[152] ,
    doutB_net[153] ,
    doutB_net[154] ,
    doutB_net[155] ,
    doutB_net[156] ,
    doutB_net[157] ,
    doutB_net[158] ,
    doutB_net[159] ,
    doutB_net[160] ,
    doutB_net[161] ,
    doutB_net[180] ,
    doutB_net[181] ,
    doutB_net[182] ,
    doutB_net[183] ,
    doutB_net[184] ,
    doutB_net[185] ,
    doutB_net[186] ,
    doutB_net[187] ,
    doutB_net[188] ,
    doutB_net[189] ,
    doutB_net[190] ,
    doutB_net[191] ,
    doutB_net[192] ,
    doutB_net[193] ,
    doutB_net[194] ,
    doutB_net[195] ,
    doutB_net[196] ,
    doutB_net[197] ,
    doutB_net[216] ,
    doutB_net[217] ,
    doutB_net[218] ,
    doutB_net[219] ,
    doutB_net[220] ,
    doutB_net[221] ,
    doutB_net[222] ,
    doutB_net[223] ,
    doutB_net[224] ,
    doutB_net[225] ,
    doutB_net[226] ,
    doutB_net[227] ,
    doutB_net[228] ,
    doutB_net[229] ,
    doutB_net[230] ,
    doutB_net[231] ,
    doutB_net[232] ,
    doutB_net[233] ,
    doutB_net[252] ,
    doutB_net[253] ,
    doutB_net[254] ,
    doutA_net[18] ,
    doutA_net[19] ,
    doutA_net[20] ,
    doutA_net[21] ,
    doutA_net[22] ,
    doutA_net[23] ,
    doutA_net[24] ,
    doutA_net[25] ,
    doutA_net[26] ,
    doutA_net[27] ,
    doutA_net[28] ,
    doutA_net[29] ,
    doutA_net[30] ,
    doutA_net[31] ,
    doutA_net[32] ,
    doutA_net[33] ,
    doutA_net[34] ,
    doutA_net[35] ,
    doutA_net[54] ,
    doutA_net[55] ,
    doutA_net[56] ,
    doutA_net[57] ,
    doutA_net[58] ,
    doutA_net[59] ,
    doutA_net[60] ,
    doutA_net[61] ,
    doutA_net[62] ,
    doutA_net[63] ,
    doutA_net[64] ,
    doutA_net[65] ,
    doutA_net[66] ,
    doutA_net[67] ,
    doutA_net[68] ,
    doutA_net[69] ,
    doutA_net[70] ,
    doutA_net[71] ,
    doutA_net[90] ,
    doutA_net[91] ,
    doutA_net[92] ,
    doutA_net[93] ,
    doutA_net[94] ,
    doutA_net[95] ,
    doutA_net[96] ,
    doutA_net[97] ,
    doutA_net[98] ,
    doutA_net[99] ,
    doutA_net[100] ,
    doutA_net[101] ,
    doutA_net[102] ,
    doutA_net[103] ,
    doutA_net[104] ,
    doutA_net[105] ,
    doutA_net[106] ,
    doutA_net[107] ,
    doutA_net[126] ,
    doutA_net[127] ,
    doutA_net[128] ,
    doutA_net[129] ,
    doutA_net[130] ,
    doutA_net[131] ,
    doutA_net[132] ,
    doutA_net[133] ,
    doutA_net[134] ,
    doutA_net[135] ,
    doutA_net[136] ,
    doutA_net[137] ,
    doutA_net[138] ,
    doutA_net[139] ,
    doutA_net[140] ,
    doutA_net[141] ,
    doutA_net[142] ,
    doutA_net[143] ,
    doutA_net[162] ,
    doutA_net[163] ,
    doutA_net[164] ,
    doutA_net[165] ,
    doutA_net[166] ,
    doutA_net[167] ,
    doutA_net[168] ,
    doutA_net[169] ,
    doutA_net[170] ,
    doutA_net[171] ,
    doutA_net[172] ,
    doutA_net[173] ,
    doutA_net[174] ,
    doutA_net[175] ,
    doutA_net[176] ,
    doutA_net[177] ,
    doutA_net[178] ,
    doutA_net[179] ,
    doutA_net[198] ,
    doutA_net[199] ,
    doutA_net[200] ,
    doutA_net[201] ,
    doutA_net[202] ,
    doutA_net[203] ,
    doutA_net[204] ,
    doutA_net[205] ,
    doutA_net[206] ,
    doutA_net[207] ,
    doutA_net[208] ,
    doutA_net[209] ,
    doutA_net[210] ,
    doutA_net[211] ,
    doutA_net[212] ,
    doutA_net[213] ,
    doutA_net[214] ,
    doutA_net[215] ,
    doutA_net[234] ,
    doutA_net[235] ,
    doutA_net[236] ,
    doutA_net[237] ,
    doutA_net[238] ,
    doutA_net[239] ,
    doutA_net[240] ,
    doutA_net[241] ,
    doutA_net[242] ,
    doutA_net[243] ,
    doutA_net[244] ,
    doutA_net[245] ,
    doutA_net[246] ,
    doutA_net[247] ,
    doutA_net[248] ,
    doutA_net[249] ,
    doutA_net[250] ,
    doutA_net[251] ,
    doutB_net[18] ,
    doutB_net[19] ,
    doutB_net[20] ,
    doutB_net[21] ,
    doutB_net[22] ,
    doutB_net[23] ,
    doutB_net[24] ,
    doutB_net[25] ,
    doutB_net[26] ,
    doutB_net[27] ,
    doutB_net[28] ,
    doutB_net[29] ,
    doutB_net[30] ,
    doutB_net[31] ,
    doutB_net[32] ,
    doutB_net[33] ,
    doutB_net[34] ,
    doutB_net[35] ,
    doutB_net[54] ,
    doutB_net[55] ,
    doutB_net[56] ,
    doutB_net[57] ,
    doutB_net[58] ,
    doutB_net[59] ,
    doutB_net[60] ,
    doutB_net[61] ,
    doutB_net[62] ,
    doutB_net[63] ,
    doutB_net[64] ,
    doutB_net[65] ,
    doutB_net[66] ,
    doutB_net[67] ,
    doutB_net[68] ,
    doutB_net[69] ,
    doutB_net[70] ,
    doutB_net[71] ,
    doutB_net[90] ,
    doutB_net[91] ,
    doutB_net[92] ,
    doutB_net[93] ,
    doutB_net[94] ,
    doutB_net[95] ,
    doutB_net[96] ,
    doutB_net[97] ,
    doutB_net[98] ,
    doutB_net[99] ,
    doutB_net[100] ,
    doutB_net[101] ,
    doutB_net[102] ,
    doutB_net[103] ,
    doutB_net[104] ,
    doutB_net[105] ,
    doutB_net[106] ,
    doutB_net[107] ,
    doutB_net[126] ,
    doutB_net[127] ,
    doutB_net[128] ,
    doutB_net[129] ,
    doutB_net[130] ,
    doutB_net[131] ,
    doutB_net[132] ,
    doutB_net[133] ,
    doutB_net[134] ,
    doutB_net[135] ,
    doutB_net[136] ,
    doutB_net[137] ,
    doutB_net[138] ,
    doutB_net[139] ,
    doutB_net[140] ,
    doutB_net[141] ,
    doutB_net[142] ,
    doutB_net[143] ,
    doutB_net[162] ,
    doutB_net[163] ,
    doutB_net[164] ,
    doutB_net[165] ,
    doutB_net[166] ,
    doutB_net[167] ,
    doutB_net[168] ,
    doutB_net[169] ,
    doutB_net[170] ,
    doutB_net[171] ,
    doutB_net[172] ,
    doutB_net[173] ,
    doutB_net[174] ,
    doutB_net[175] ,
    doutB_net[176] ,
    doutB_net[177] ,
    doutB_net[178] ,
    doutB_net[179] ,
    doutB_net[198] ,
    doutB_net[199] ,
    doutB_net[200] ,
    doutB_net[201] ,
    doutB_net[202] ,
    doutB_net[203] ,
    doutB_net[204] ,
    doutB_net[205] ,
    doutB_net[206] ,
    doutB_net[207] ,
    doutB_net[208] ,
    doutB_net[209] ,
    doutB_net[210] ,
    doutB_net[211] ,
    doutB_net[212] ,
    doutB_net[213] ,
    doutB_net[214] ,
    doutB_net[215] ,
    doutB_net[234] ,
    doutB_net[235] ,
    doutB_net[236] ,
    doutB_net[237] ,
    doutB_net[238] ,
    doutB_net[239] ,
    doutB_net[240] ,
    doutB_net[241] ,
    doutB_net[242] ,
    doutB_net[243] ,
    doutB_net[244] ,
    doutB_net[245] ,
    doutB_net[246] ,
    doutB_net[247] ,
    doutB_net[248] ,
    doutB_net[249] ,
    doutB_net[250] ,
    doutB_net[251] );
    `else
        tdp_256x16_post_synth netlist(.*, .doutA(doutA_net), .doutB(doutB_net));
    `endif


    
    //clock//
    initial begin
        clkA = 1'b0;
        forever #10 clkA = ~clkA;
    end
    initial begin
        clkB = 1'b0;
        forever #5 clkB = ~clkB;
    end
    initial begin
        for(integer i = 0; i<16; i=i+1) begin 
            golden.ram[i] ='b0;
        end 
    end

    initial begin

    {weA,weB, addrA,addrB, dinA, dinB, cycle, i} = 0;
 
 
    repeat (1) @ (negedge clkA);
    addrA <= 'd1; addrB <= 'd2; weA <=1'b1; weB <=1'b1; dinA<= {$random}; dinB<= {$random};
    compare(cycle);
    repeat (1) @ (negedge clkA);
    addrA <= 'd1; addrB <= 'd2; weA <=1'b0; weB <=1'b0; dinA<= {$random}; dinB<= {$random};
    compare(cycle);

    for (integer i=0; i<512; i=i+1)begin
        repeat (1) @ (negedge clkA)

        addrA <= $urandom_range(0,7); addrB <= $urandom_range(8,15); weA <=1'b1; weB <=1'b1; dinA<= {$random}; dinB<= {$random};
        cycle = cycle +1;
     
        compare(cycle);

    end

    for (integer i=0; i<512; i=i+1)begin
        repeat (1) @ (negedge clkB)

        addrA <= $urandom_range(0,7); addrB <= $urandom_range(8,15); weA <=1'b0; weB <=1'b0; dinA<= {$random}; dinB<= {$random};
        cycle = cycle +1;
     
        compare(cycle);

    end

    for (integer i=0; i<512; i=i+1)begin
        repeat (1) @ (negedge clkA)

        addrA <= $urandom_range(0,7); addrB <= $urandom_range(8,15); weA <=1'b0; weB <=1'b1; dinA<= {$random}; dinB<= {$random};
        cycle = cycle +1;
     
        compare(cycle);

    end

    for (integer i=0; i<512; i=i+1)begin
        repeat (1) @ (negedge clkB)

        addrA <= $urandom_range(0,7); addrB <= $urandom_range(8,15); weA <=1'b1; weB <=1'b0; dinA<= {$random}; dinB<= {$random};
        cycle = cycle +1;
     
        compare(cycle);

    end
    
    //random
    for (integer i=0; i<512; i=i+1)begin
        repeat (1) @ (negedge clkA)
        addrA <=$urandom_range(8,15); addrB <= $urandom_range(0,7); weA <={$random}; weB <={$random}; dinA<= {$random}; dinB<= {$random};
        cycle = cycle +1;
       
        compare(cycle);
    end
    if(mismatch == 0)
        $display("\n**** All Comparison Matched ***\nSimulation Passed");
    else
        $display("%0d comparison(s) mismatched\nERROR: SIM: Simulation Failed", mismatch);
    

    repeat (10) @(negedge clkA); $finish;
    end

    task compare(input integer cycle);
    //$display("\n Comparison at cycle %0d", cycle);
    if(doutA !== doutA_net) begin
        $display("doutA mismatch. Golden: %0h, Netlist: %0h, Time: %0t", doutA, doutA_net,$time);
        mismatch = mismatch+1;
    end

     if(doutB !== doutB_net) begin
        $display("doutB mismatch. Golden: %0h, Netlist: %0h, Time: %0t", doutB, doutB_net,$time);
        mismatch = mismatch+1;
    end
    
    
    endtask


initial begin
    $dumpfile("tb.vcd");
    $dumpvars;
end
endmodule