
module co_sim_tdp_512x10;

    reg clkA, clkB, weA, weB;
    reg [3:0] addrA, addrB;
    reg [511:0] dinA, dinB;
    wire [511:0] doutA, doutB, doutA_net, doutB_net;

    integer mismatch=0;
    reg [6:0]cycle, i;

    tdp_512x10 golden(.*);
     `ifdef PNR
        tdp_512x10_post_route netlist( 
      input \clkA ,
    input \clkB ,
    input \weA ,
    input \weB ,
    input \addrA[0] ,
    input \addrA[1] ,
    input \addrA[2] ,
    input \addrA[3] ,
    input \addrB[0] ,
    input \addrB[1] ,
    input \addrB[2] ,
    input \addrB[3] ,
    input \dinA[0] ,
    input \dinA[1] ,
    input \dinA[2] ,
    input \dinA[3] ,
    input \dinA[4] ,
    input \dinA[5] ,
    input \dinA[6] ,
    input \dinA[7] ,
    input \dinA[8] ,
    input \dinA[9] ,
    input \dinA[10] ,
    input \dinA[11] ,
    input \dinA[12] ,
    input \dinA[13] ,
    input \dinA[14] ,
    input \dinA[15] ,
    input \dinA[16] ,
    input \dinA[17] ,
    input \dinA[18] ,
    input \dinA[19] ,
    input \dinA[20] ,
    input \dinA[21] ,
    input \dinA[22] ,
    input \dinA[23] ,
    input \dinA[24] ,
    input \dinA[25] ,
    input \dinA[26] ,
    input \dinA[27] ,
    input \dinA[28] ,
    input \dinA[29] ,
    input \dinA[30] ,
    input \dinA[31] ,
    input \dinA[32] ,
    input \dinA[33] ,
    input \dinA[34] ,
    input \dinA[35] ,
    input \dinA[36] ,
    input \dinA[37] ,
    input \dinA[38] ,
    input \dinA[39] ,
    input \dinA[40] ,
    input \dinA[41] ,
    input \dinA[42] ,
    input \dinA[43] ,
    input \dinA[44] ,
    input \dinA[45] ,
    input \dinA[46] ,
    input \dinA[47] ,
    input \dinA[48] ,
    input \dinA[49] ,
    input \dinA[50] ,
    input \dinA[51] ,
    input \dinA[52] ,
    input \dinA[53] ,
    input \dinA[54] ,
    input \dinA[55] ,
    input \dinA[56] ,
    input \dinA[57] ,
    input \dinA[58] ,
    input \dinA[59] ,
    input \dinA[60] ,
    input \dinA[61] ,
    input \dinA[62] ,
    input \dinA[63] ,
    input \dinA[64] ,
    input \dinA[65] ,
    input \dinA[66] ,
    input \dinA[67] ,
    input \dinA[68] ,
    input \dinA[69] ,
    input \dinA[70] ,
    input \dinA[71] ,
    input \dinA[72] ,
    input \dinA[73] ,
    input \dinA[74] ,
    input \dinA[75] ,
    input \dinA[76] ,
    input \dinA[77] ,
    input \dinA[78] ,
    input \dinA[79] ,
    input \dinA[80] ,
    input \dinA[81] ,
    input \dinA[82] ,
    input \dinA[83] ,
    input \dinA[84] ,
    input \dinA[85] ,
    input \dinA[86] ,
    input \dinA[87] ,
    input \dinA[88] ,
    input \dinA[89] ,
    input \dinA[90] ,
    input \dinA[91] ,
    input \dinA[92] ,
    input \dinA[93] ,
    input \dinA[94] ,
    input \dinA[95] ,
    input \dinA[96] ,
    input \dinA[97] ,
    input \dinA[98] ,
    input \dinA[99] ,
    input \dinA[100] ,
    input \dinA[101] ,
    input \dinA[102] ,
    input \dinA[103] ,
    input \dinA[104] ,
    input \dinA[105] ,
    input \dinA[106] ,
    input \dinA[107] ,
    input \dinA[108] ,
    input \dinA[109] ,
    input \dinA[110] ,
    input \dinA[111] ,
    input \dinA[112] ,
    input \dinA[113] ,
    input \dinA[114] ,
    input \dinA[115] ,
    input \dinA[116] ,
    input \dinA[117] ,
    input \dinA[118] ,
    input \dinA[119] ,
    input \dinA[120] ,
    input \dinA[121] ,
    input \dinA[122] ,
    input \dinA[123] ,
    input \dinA[124] ,
    input \dinA[125] ,
    input \dinA[126] ,
    input \dinA[127] ,
    input \dinA[128] ,
    input \dinA[129] ,
    input \dinA[130] ,
    input \dinA[131] ,
    input \dinA[132] ,
    input \dinA[133] ,
    input \dinA[134] ,
    input \dinA[135] ,
    input \dinA[136] ,
    input \dinA[137] ,
    input \dinA[138] ,
    input \dinA[139] ,
    input \dinA[140] ,
    input \dinA[141] ,
    input \dinA[142] ,
    input \dinA[143] ,
    input \dinA[144] ,
    input \dinA[145] ,
    input \dinA[146] ,
    input \dinA[147] ,
    input \dinA[148] ,
    input \dinA[149] ,
    input \dinA[150] ,
    input \dinA[151] ,
    input \dinA[152] ,
    input \dinA[153] ,
    input \dinA[154] ,
    input \dinA[155] ,
    input \dinA[156] ,
    input \dinA[157] ,
    input \dinA[158] ,
    input \dinA[159] ,
    input \dinA[160] ,
    input \dinA[161] ,
    input \dinA[162] ,
    input \dinA[163] ,
    input \dinA[164] ,
    input \dinA[165] ,
    input \dinA[166] ,
    input \dinA[167] ,
    input \dinA[168] ,
    input \dinA[169] ,
    input \dinA[170] ,
    input \dinA[171] ,
    input \dinA[172] ,
    input \dinA[173] ,
    input \dinA[174] ,
    input \dinA[175] ,
    input \dinA[176] ,
    input \dinA[177] ,
    input \dinA[178] ,
    input \dinA[179] ,
    input \dinA[180] ,
    input \dinA[181] ,
    input \dinA[182] ,
    input \dinA[183] ,
    input \dinA[184] ,
    input \dinA[185] ,
    input \dinA[186] ,
    input \dinA[187] ,
    input \dinA[188] ,
    input \dinA[189] ,
    input \dinA[190] ,
    input \dinA[191] ,
    input \dinA[192] ,
    input \dinA[193] ,
    input \dinA[194] ,
    input \dinA[195] ,
    input \dinA[196] ,
    input \dinA[197] ,
    input \dinA[198] ,
    input \dinA[199] ,
    input \dinA[200] ,
    input \dinA[201] ,
    input \dinA[202] ,
    input \dinA[203] ,
    input \dinA[204] ,
    input \dinA[205] ,
    input \dinA[206] ,
    input \dinA[207] ,
    input \dinA[208] ,
    input \dinA[209] ,
    input \dinA[210] ,
    input \dinA[211] ,
    input \dinA[212] ,
    input \dinA[213] ,
    input \dinA[214] ,
    input \dinA[215] ,
    input \dinA[216] ,
    input \dinA[217] ,
    input \dinA[218] ,
    input \dinA[219] ,
    input \dinA[220] ,
    input \dinA[221] ,
    input \dinA[222] ,
    input \dinA[223] ,
    input \dinA[224] ,
    input \dinA[225] ,
    input \dinA[226] ,
    input \dinA[227] ,
    input \dinA[228] ,
    input \dinA[229] ,
    input \dinA[230] ,
    input \dinA[231] ,
    input \dinA[232] ,
    input \dinA[233] ,
    input \dinA[234] ,
    input \dinA[235] ,
    input \dinA[236] ,
    input \dinA[237] ,
    input \dinA[238] ,
    input \dinA[239] ,
    input \dinA[240] ,
    input \dinA[241] ,
    input \dinA[242] ,
    input \dinA[243] ,
    input \dinA[244] ,
    input \dinA[245] ,
    input \dinA[246] ,
    input \dinA[247] ,
    input \dinA[248] ,
    input \dinA[249] ,
    input \dinA[250] ,
    input \dinA[251] ,
    input \dinA[252] ,
    input \dinA[253] ,
    input \dinA[254] ,
    input \dinA[255] ,
    input \dinA[256] ,
    input \dinA[257] ,
    input \dinA[258] ,
    input \dinA[259] ,
    input \dinA[260] ,
    input \dinA[261] ,
    input \dinA[262] ,
    input \dinA[263] ,
    input \dinA[264] ,
    input \dinA[265] ,
    input \dinA[266] ,
    input \dinA[267] ,
    input \dinA[268] ,
    input \dinA[269] ,
    input \dinA[270] ,
    input \dinA[271] ,
    input \dinA[272] ,
    input \dinA[273] ,
    input \dinA[274] ,
    input \dinA[275] ,
    input \dinA[276] ,
    input \dinA[277] ,
    input \dinA[278] ,
    input \dinA[279] ,
    input \dinA[280] ,
    input \dinA[281] ,
    input \dinA[282] ,
    input \dinA[283] ,
    input \dinA[284] ,
    input \dinA[285] ,
    input \dinA[286] ,
    input \dinA[287] ,
    input \dinA[288] ,
    input \dinA[289] ,
    input \dinA[290] ,
    input \dinA[291] ,
    input \dinA[292] ,
    input \dinA[293] ,
    input \dinA[294] ,
    input \dinA[295] ,
    input \dinA[296] ,
    input \dinA[297] ,
    input \dinA[298] ,
    input \dinA[299] ,
    input \dinA[300] ,
    input \dinA[301] ,
    input \dinA[302] ,
    input \dinA[303] ,
    input \dinA[304] ,
    input \dinA[305] ,
    input \dinA[306] ,
    input \dinA[307] ,
    input \dinA[308] ,
    input \dinA[309] ,
    input \dinA[310] ,
    input \dinA[311] ,
    input \dinA[312] ,
    input \dinA[313] ,
    input \dinA[314] ,
    input \dinA[315] ,
    input \dinA[316] ,
    input \dinA[317] ,
    input \dinA[318] ,
    input \dinA[319] ,
    input \dinA[320] ,
    input \dinA[321] ,
    input \dinA[322] ,
    input \dinA[323] ,
    input \dinA[324] ,
    input \dinA[325] ,
    input \dinA[326] ,
    input \dinA[327] ,
    input \dinA[328] ,
    input \dinA[329] ,
    input \dinA[330] ,
    input \dinA[331] ,
    input \dinA[332] ,
    input \dinA[333] ,
    input \dinA[334] ,
    input \dinA[335] ,
    input \dinA[336] ,
    input \dinA[337] ,
    input \dinA[338] ,
    input \dinA[339] ,
    input \dinA[340] ,
    input \dinA[341] ,
    input \dinA[342] ,
    input \dinA[343] ,
    input \dinA[344] ,
    input \dinA[345] ,
    input \dinA[346] ,
    input \dinA[347] ,
    input \dinA[348] ,
    input \dinA[349] ,
    input \dinA[350] ,
    input \dinA[351] ,
    input \dinA[352] ,
    input \dinA[353] ,
    input \dinA[354] ,
    input \dinA[355] ,
    input \dinA[356] ,
    input \dinA[357] ,
    input \dinA[358] ,
    input \dinA[359] ,
    input \dinA[360] ,
    input \dinA[361] ,
    input \dinA[362] ,
    input \dinA[363] ,
    input \dinA[364] ,
    input \dinA[365] ,
    input \dinA[366] ,
    input \dinA[367] ,
    input \dinA[368] ,
    input \dinA[369] ,
    input \dinA[370] ,
    input \dinA[371] ,
    input \dinA[372] ,
    input \dinA[373] ,
    input \dinA[374] ,
    input \dinA[375] ,
    input \dinA[376] ,
    input \dinA[377] ,
    input \dinA[378] ,
    input \dinA[379] ,
    input \dinA[380] ,
    input \dinA[381] ,
    input \dinA[382] ,
    input \dinA[383] ,
    input \dinA[384] ,
    input \dinA[385] ,
    input \dinA[386] ,
    input \dinA[387] ,
    input \dinA[388] ,
    input \dinA[389] ,
    input \dinA[390] ,
    input \dinA[391] ,
    input \dinA[392] ,
    input \dinA[393] ,
    input \dinA[394] ,
    input \dinA[395] ,
    input \dinA[396] ,
    input \dinA[397] ,
    input \dinA[398] ,
    input \dinA[399] ,
    input \dinA[400] ,
    input \dinA[401] ,
    input \dinA[402] ,
    input \dinA[403] ,
    input \dinA[404] ,
    input \dinA[405] ,
    input \dinA[406] ,
    input \dinA[407] ,
    input \dinA[408] ,
    input \dinA[409] ,
    input \dinA[410] ,
    input \dinA[411] ,
    input \dinA[412] ,
    input \dinA[413] ,
    input \dinA[414] ,
    input \dinA[415] ,
    input \dinA[416] ,
    input \dinA[417] ,
    input \dinA[418] ,
    input \dinA[419] ,
    input \dinA[420] ,
    input \dinA[421] ,
    input \dinA[422] ,
    input \dinA[423] ,
    input \dinA[424] ,
    input \dinA[425] ,
    input \dinA[426] ,
    input \dinA[427] ,
    input \dinA[428] ,
    input \dinA[429] ,
    input \dinA[430] ,
    input \dinA[431] ,
    input \dinA[432] ,
    input \dinA[433] ,
    input \dinA[434] ,
    input \dinA[435] ,
    input \dinA[436] ,
    input \dinA[437] ,
    input \dinA[438] ,
    input \dinA[439] ,
    input \dinA[440] ,
    input \dinA[441] ,
    input \dinA[442] ,
    input \dinA[443] ,
    input \dinA[444] ,
    input \dinA[445] ,
    input \dinA[446] ,
    input \dinA[447] ,
    input \dinA[448] ,
    input \dinA[449] ,
    input \dinA[450] ,
    input \dinA[451] ,
    input \dinA[452] ,
    input \dinA[453] ,
    input \dinA[454] ,
    input \dinA[455] ,
    input \dinA[456] ,
    input \dinA[457] ,
    input \dinA[458] ,
    input \dinA[459] ,
    input \dinA[460] ,
    input \dinA[461] ,
    input \dinA[462] ,
    input \dinA[463] ,
    input \dinA[464] ,
    input \dinA[465] ,
    input \dinA[466] ,
    input \dinA[467] ,
    input \dinA[468] ,
    input \dinA[469] ,
    input \dinA[470] ,
    input \dinA[471] ,
    input \dinA[472] ,
    input \dinA[473] ,
    input \dinA[474] ,
    input \dinA[475] ,
    input \dinA[476] ,
    input \dinA[477] ,
    input \dinA[478] ,
    input \dinA[479] ,
    input \dinA[480] ,
    input \dinA[481] ,
    input \dinA[482] ,
    input \dinA[483] ,
    input \dinA[484] ,
    input \dinA[485] ,
    input \dinA[486] ,
    input \dinA[487] ,
    input \dinA[488] ,
    input \dinA[489] ,
    input \dinA[490] ,
    input \dinA[491] ,
    input \dinA[492] ,
    input \dinA[493] ,
    input \dinA[494] ,
    input \dinA[495] ,
    input \dinA[496] ,
    input \dinA[497] ,
    input \dinA[498] ,
    input \dinA[499] ,
    input \dinA[500] ,
    input \dinA[501] ,
    input \dinA[502] ,
    input \dinA[503] ,
    input \dinA[504] ,
    input \dinA[505] ,
    input \dinA[506] ,
    input \dinA[507] ,
    input \dinA[508] ,
    input \dinA[509] ,
    input \dinA[510] ,
    input \dinA[511] ,
    input \dinB[0] ,
    input \dinB[1] ,
    input \dinB[2] ,
    input \dinB[3] ,
    input \dinB[4] ,
    input \dinB[5] ,
    input \dinB[6] ,
    input \dinB[7] ,
    input \dinB[8] ,
    input \dinB[9] ,
    input \dinB[10] ,
    input \dinB[11] ,
    input \dinB[12] ,
    input \dinB[13] ,
    input \dinB[14] ,
    input \dinB[15] ,
    input \dinB[16] ,
    input \dinB[17] ,
    input \dinB[18] ,
    input \dinB[19] ,
    input \dinB[20] ,
    input \dinB[21] ,
    input \dinB[22] ,
    input \dinB[23] ,
    input \dinB[24] ,
    input \dinB[25] ,
    input \dinB[26] ,
    input \dinB[27] ,
    input \dinB[28] ,
    input \dinB[29] ,
    input \dinB[30] ,
    input \dinB[31] ,
    input \dinB[32] ,
    input \dinB[33] ,
    input \dinB[34] ,
    input \dinB[35] ,
    input \dinB[36] ,
    input \dinB[37] ,
    input \dinB[38] ,
    input \dinB[39] ,
    input \dinB[40] ,
    input \dinB[41] ,
    input \dinB[42] ,
    input \dinB[43] ,
    input \dinB[44] ,
    input \dinB[45] ,
    input \dinB[46] ,
    input \dinB[47] ,
    input \dinB[48] ,
    input \dinB[49] ,
    input \dinB[50] ,
    input \dinB[51] ,
    input \dinB[52] ,
    input \dinB[53] ,
    input \dinB[54] ,
    input \dinB[55] ,
    input \dinB[56] ,
    input \dinB[57] ,
    input \dinB[58] ,
    input \dinB[59] ,
    input \dinB[60] ,
    input \dinB[61] ,
    input \dinB[62] ,
    input \dinB[63] ,
    input \dinB[64] ,
    input \dinB[65] ,
    input \dinB[66] ,
    input \dinB[67] ,
    input \dinB[68] ,
    input \dinB[69] ,
    input \dinB[70] ,
    input \dinB[71] ,
    input \dinB[72] ,
    input \dinB[73] ,
    input \dinB[74] ,
    input \dinB[75] ,
    input \dinB[76] ,
    input \dinB[77] ,
    input \dinB[78] ,
    input \dinB[79] ,
    input \dinB[80] ,
    input \dinB[81] ,
    input \dinB[82] ,
    input \dinB[83] ,
    input \dinB[84] ,
    input \dinB[85] ,
    input \dinB[86] ,
    input \dinB[87] ,
    input \dinB[88] ,
    input \dinB[89] ,
    input \dinB[90] ,
    input \dinB[91] ,
    input \dinB[92] ,
    input \dinB[93] ,
    input \dinB[94] ,
    input \dinB[95] ,
    input \dinB[96] ,
    input \dinB[97] ,
    input \dinB[98] ,
    input \dinB[99] ,
    input \dinB[100] ,
    input \dinB[101] ,
    input \dinB[102] ,
    input \dinB[103] ,
    input \dinB[104] ,
    input \dinB[105] ,
    input \dinB[106] ,
    input \dinB[107] ,
    input \dinB[108] ,
    input \dinB[109] ,
    input \dinB[110] ,
    input \dinB[111] ,
    input \dinB[112] ,
    input \dinB[113] ,
    input \dinB[114] ,
    input \dinB[115] ,
    input \dinB[116] ,
    input \dinB[117] ,
    input \dinB[118] ,
    input \dinB[119] ,
    input \dinB[120] ,
    input \dinB[121] ,
    input \dinB[122] ,
    input \dinB[123] ,
    input \dinB[124] ,
    input \dinB[125] ,
    input \dinB[126] ,
    input \dinB[127] ,
    input \dinB[128] ,
    input \dinB[129] ,
    input \dinB[130] ,
    input \dinB[131] ,
    input \dinB[132] ,
    input \dinB[133] ,
    input \dinB[134] ,
    input \dinB[135] ,
    input \dinB[136] ,
    input \dinB[137] ,
    input \dinB[138] ,
    input \dinB[139] ,
    input \dinB[140] ,
    input \dinB[141] ,
    input \dinB[142] ,
    input \dinB[143] ,
    input \dinB[144] ,
    input \dinB[145] ,
    input \dinB[146] ,
    input \dinB[147] ,
    input \dinB[148] ,
    input \dinB[149] ,
    input \dinB[150] ,
    input \dinB[151] ,
    input \dinB[152] ,
    input \dinB[153] ,
    input \dinB[154] ,
    input \dinB[155] ,
    input \dinB[156] ,
    input \dinB[157] ,
    input \dinB[158] ,
    input \dinB[159] ,
    input \dinB[160] ,
    input \dinB[161] ,
    input \dinB[162] ,
    input \dinB[163] ,
    input \dinB[164] ,
    input \dinB[165] ,
    input \dinB[166] ,
    input \dinB[167] ,
    input \dinB[168] ,
    input \dinB[169] ,
    input \dinB[170] ,
    input \dinB[171] ,
    input \dinB[172] ,
    input \dinB[173] ,
    input \dinB[174] ,
    input \dinB[175] ,
    input \dinB[176] ,
    input \dinB[177] ,
    input \dinB[178] ,
    input \dinB[179] ,
    input \dinB[180] ,
    input \dinB[181] ,
    input \dinB[182] ,
    input \dinB[183] ,
    input \dinB[184] ,
    input \dinB[185] ,
    input \dinB[186] ,
    input \dinB[187] ,
    input \dinB[188] ,
    input \dinB[189] ,
    input \dinB[190] ,
    input \dinB[191] ,
    input \dinB[192] ,
    input \dinB[193] ,
    input \dinB[194] ,
    input \dinB[195] ,
    input \dinB[196] ,
    input \dinB[197] ,
    input \dinB[198] ,
    input \dinB[199] ,
    input \dinB[200] ,
    input \dinB[201] ,
    input \dinB[202] ,
    input \dinB[203] ,
    input \dinB[204] ,
    input \dinB[205] ,
    input \dinB[206] ,
    input \dinB[207] ,
    input \dinB[208] ,
    input \dinB[209] ,
    input \dinB[210] ,
    input \dinB[211] ,
    input \dinB[212] ,
    input \dinB[213] ,
    input \dinB[214] ,
    input \dinB[215] ,
    input \dinB[216] ,
    input \dinB[217] ,
    input \dinB[218] ,
    input \dinB[219] ,
    input \dinB[220] ,
    input \dinB[221] ,
    input \dinB[222] ,
    input \dinB[223] ,
    input \dinB[224] ,
    input \dinB[225] ,
    input \dinB[226] ,
    input \dinB[227] ,
    input \dinB[228] ,
    input \dinB[229] ,
    input \dinB[230] ,
    input \dinB[231] ,
    input \dinB[232] ,
    input \dinB[233] ,
    input \dinB[234] ,
    input \dinB[235] ,
    input \dinB[236] ,
    input \dinB[237] ,
    input \dinB[238] ,
    input \dinB[239] ,
    input \dinB[240] ,
    input \dinB[241] ,
    input \dinB[242] ,
    input \dinB[243] ,
    input \dinB[244] ,
    input \dinB[245] ,
    input \dinB[246] ,
    input \dinB[247] ,
    input \dinB[248] ,
    input \dinB[249] ,
    input \dinB[250] ,
    input \dinB[251] ,
    input \dinB[252] ,
    input \dinB[253] ,
    input \dinB[254] ,
    input \dinB[255] ,
    input \dinB[256] ,
    input \dinB[257] ,
    input \dinB[258] ,
    input \dinB[259] ,
    input \dinB[260] ,
    input \dinB[261] ,
    input \dinB[262] ,
    input \dinB[263] ,
    input \dinB[264] ,
    input \dinB[265] ,
    input \dinB[266] ,
    input \dinB[267] ,
    input \dinB[268] ,
    input \dinB[269] ,
    input \dinB[270] ,
    input \dinB[271] ,
    input \dinB[272] ,
    input \dinB[273] ,
    input \dinB[274] ,
    input \dinB[275] ,
    input \dinB[276] ,
    input \dinB[277] ,
    input \dinB[278] ,
    input \dinB[279] ,
    input \dinB[280] ,
    input \dinB[281] ,
    input \dinB[282] ,
    input \dinB[283] ,
    input \dinB[284] ,
    input \dinB[285] ,
    input \dinB[286] ,
    input \dinB[287] ,
    input \dinB[288] ,
    input \dinB[289] ,
    input \dinB[290] ,
    input \dinB[291] ,
    input \dinB[292] ,
    input \dinB[293] ,
    input \dinB[294] ,
    input \dinB[295] ,
    input \dinB[296] ,
    input \dinB[297] ,
    input \dinB[298] ,
    input \dinB[299] ,
    input \dinB[300] ,
    input \dinB[301] ,
    input \dinB[302] ,
    input \dinB[303] ,
    input \dinB[304] ,
    input \dinB[305] ,
    input \dinB[306] ,
    input \dinB[307] ,
    input \dinB[308] ,
    input \dinB[309] ,
    input \dinB[310] ,
    input \dinB[311] ,
    input \dinB[312] ,
    input \dinB[313] ,
    input \dinB[314] ,
    input \dinB[315] ,
    input \dinB[316] ,
    input \dinB[317] ,
    input \dinB[318] ,
    input \dinB[319] ,
    input \dinB[320] ,
    input \dinB[321] ,
    input \dinB[322] ,
    input \dinB[323] ,
    input \dinB[324] ,
    input \dinB[325] ,
    input \dinB[326] ,
    input \dinB[327] ,
    input \dinB[328] ,
    input \dinB[329] ,
    input \dinB[330] ,
    input \dinB[331] ,
    input \dinB[332] ,
    input \dinB[333] ,
    input \dinB[334] ,
    input \dinB[335] ,
    input \dinB[336] ,
    input \dinB[337] ,
    input \dinB[338] ,
    input \dinB[339] ,
    input \dinB[340] ,
    input \dinB[341] ,
    input \dinB[342] ,
    input \dinB[343] ,
    input \dinB[344] ,
    input \dinB[345] ,
    input \dinB[346] ,
    input \dinB[347] ,
    input \dinB[348] ,
    input \dinB[349] ,
    input \dinB[350] ,
    input \dinB[351] ,
    input \dinB[352] ,
    input \dinB[353] ,
    input \dinB[354] ,
    input \dinB[355] ,
    input \dinB[356] ,
    input \dinB[357] ,
    input \dinB[358] ,
    input \dinB[359] ,
    input \dinB[360] ,
    input \dinB[361] ,
    input \dinB[362] ,
    input \dinB[363] ,
    input \dinB[364] ,
    input \dinB[365] ,
    input \dinB[366] ,
    input \dinB[367] ,
    input \dinB[368] ,
    input \dinB[369] ,
    input \dinB[370] ,
    input \dinB[371] ,
    input \dinB[372] ,
    input \dinB[373] ,
    input \dinB[374] ,
    input \dinB[375] ,
    input \dinB[376] ,
    input \dinB[377] ,
    input \dinB[378] ,
    input \dinB[379] ,
    input \dinB[380] ,
    input \dinB[381] ,
    input \dinB[382] ,
    input \dinB[383] ,
    input \dinB[384] ,
    input \dinB[385] ,
    input \dinB[386] ,
    input \dinB[387] ,
    input \dinB[388] ,
    input \dinB[389] ,
    input \dinB[390] ,
    input \dinB[391] ,
    input \dinB[392] ,
    input \dinB[393] ,
    input \dinB[394] ,
    input \dinB[395] ,
    input \dinB[396] ,
    input \dinB[397] ,
    input \dinB[398] ,
    input \dinB[399] ,
    input \dinB[400] ,
    input \dinB[401] ,
    input \dinB[402] ,
    input \dinB[403] ,
    input \dinB[404] ,
    input \dinB[405] ,
    input \dinB[406] ,
    input \dinB[407] ,
    input \dinB[408] ,
    input \dinB[409] ,
    input \dinB[410] ,
    input \dinB[411] ,
    input \dinB[412] ,
    input \dinB[413] ,
    input \dinB[414] ,
    input \dinB[415] ,
    input \dinB[416] ,
    input \dinB[417] ,
    input \dinB[418] ,
    input \dinB[419] ,
    input \dinB[420] ,
    input \dinB[421] ,
    input \dinB[422] ,
    input \dinB[423] ,
    input \dinB[424] ,
    input \dinB[425] ,
    input \dinB[426] ,
    input \dinB[427] ,
    input \dinB[428] ,
    input \dinB[429] ,
    input \dinB[430] ,
    input \dinB[431] ,
    input \dinB[432] ,
    input \dinB[433] ,
    input \dinB[434] ,
    input \dinB[435] ,
    input \dinB[436] ,
    input \dinB[437] ,
    input \dinB[438] ,
    input \dinB[439] ,
    input \dinB[440] ,
    input \dinB[441] ,
    input \dinB[442] ,
    input \dinB[443] ,
    input \dinB[444] ,
    input \dinB[445] ,
    input \dinB[446] ,
    input \dinB[447] ,
    input \dinB[448] ,
    input \dinB[449] ,
    input \dinB[450] ,
    input \dinB[451] ,
    input \dinB[452] ,
    input \dinB[453] ,
    input \dinB[454] ,
    input \dinB[455] ,
    input \dinB[456] ,
    input \dinB[457] ,
    input \dinB[458] ,
    input \dinB[459] ,
    input \dinB[460] ,
    input \dinB[461] ,
    input \dinB[462] ,
    input \dinB[463] ,
    input \dinB[464] ,
    input \dinB[465] ,
    input \dinB[466] ,
    input \dinB[467] ,
    input \dinB[468] ,
    input \dinB[469] ,
    input \dinB[470] ,
    input \dinB[471] ,
    input \dinB[472] ,
    input \dinB[473] ,
    input \dinB[474] ,
    input \dinB[475] ,
    input \dinB[476] ,
    input \dinB[477] ,
    input \dinB[478] ,
    input \dinB[479] ,
    input \dinB[480] ,
    input \dinB[481] ,
    input \dinB[482] ,
    input \dinB[483] ,
    input \dinB[484] ,
    input \dinB[485] ,
    input \dinB[486] ,
    input \dinB[487] ,
    input \dinB[488] ,
    input \dinB[489] ,
    input \dinB[490] ,
    input \dinB[491] ,
    input \dinB[492] ,
    input \dinB[493] ,
    input \dinB[494] ,
    input \dinB[495] ,
    input \dinB[496] ,
    input \dinB[497] ,
    input \dinB[498] ,
    input \dinB[499] ,
    input \dinB[500] ,
    input \dinB[501] ,
    input \dinB[502] ,
    input \dinB[503] ,
    input \dinB[504] ,
    input \dinB[505] ,
    input \dinB[506] ,
    input \dinB[507] ,
    input \dinB[508] ,
    input \dinB[509] ,
    input \dinB[510] ,
    input \dinB[511] ,
    doutA_net[45] ,
    doutB_net[401] ,
    doutA_net[0] ,
    doutA_net[1] ,
    doutA_net[2] ,
    doutA_net[3] ,
    doutA_net[4] ,
    doutA_net[5] ,
    doutA_net[6] ,
    doutA_net[7] ,
    doutA_net[8] ,
    doutA_net[9] ,
    doutA_net[10] ,
    doutA_net[11] ,
    doutA_net[12] ,
    doutA_net[13] ,
    doutA_net[14] ,
    doutA_net[15] ,
    doutA_net[16] ,
    doutA_net[17] ,
    doutA_net[36] ,
    doutA_net[37] ,
    doutA_net[38] ,
    doutA_net[39] ,
    doutA_net[40] ,
    doutA_net[41] ,
    doutA_net[42] ,
    doutA_net[43] ,
    doutA_net[44] ,
    doutA_net[46] ,
    doutA_net[47] ,
    doutA_net[48] ,
    doutA_net[49] ,
    doutA_net[50] ,
    doutA_net[51] ,
    doutA_net[52] ,
    doutA_net[53] ,
    doutA_net[72] ,
    doutA_net[73] ,
    doutA_net[74] ,
    doutA_net[75] ,
    doutA_net[76] ,
    doutA_net[77] ,
    doutA_net[78] ,
    doutA_net[79] ,
    doutA_net[80] ,
    doutA_net[81] ,
    doutA_net[82] ,
    doutA_net[83] ,
    doutA_net[84] ,
    doutA_net[85] ,
    doutA_net[86] ,
    doutA_net[87] ,
    doutA_net[88] ,
    doutA_net[89] ,
    doutA_net[108] ,
    doutA_net[109] ,
    doutA_net[110] ,
    doutA_net[111] ,
    doutA_net[112] ,
    doutA_net[113] ,
    doutA_net[114] ,
    doutA_net[115] ,
    doutA_net[116] ,
    doutA_net[117] ,
    doutA_net[118] ,
    doutA_net[119] ,
    doutA_net[120] ,
    doutA_net[121] ,
    doutA_net[122] ,
    doutA_net[123] ,
    doutA_net[124] ,
    doutA_net[125] ,
    doutA_net[144] ,
    doutA_net[145] ,
    doutA_net[146] ,
    doutA_net[147] ,
    doutA_net[148] ,
    doutA_net[149] ,
    doutA_net[150] ,
    doutA_net[151] ,
    doutA_net[152] ,
    doutA_net[153] ,
    doutA_net[154] ,
    doutA_net[155] ,
    doutA_net[156] ,
    doutA_net[157] ,
    doutA_net[158] ,
    doutA_net[159] ,
    doutA_net[160] ,
    doutA_net[161] ,
    doutA_net[180] ,
    doutA_net[181] ,
    doutA_net[182] ,
    doutA_net[183] ,
    doutA_net[184] ,
    doutA_net[185] ,
    doutA_net[186] ,
    doutA_net[187] ,
    doutA_net[188] ,
    doutA_net[189] ,
    doutA_net[190] ,
    doutA_net[191] ,
    doutA_net[192] ,
    doutA_net[193] ,
    doutA_net[194] ,
    doutA_net[195] ,
    doutA_net[196] ,
    doutA_net[197] ,
    doutA_net[216] ,
    doutA_net[217] ,
    doutA_net[218] ,
    doutA_net[219] ,
    doutA_net[220] ,
    doutA_net[221] ,
    doutA_net[222] ,
    doutA_net[223] ,
    doutA_net[224] ,
    doutA_net[225] ,
    doutA_net[226] ,
    doutA_net[227] ,
    doutA_net[228] ,
    doutA_net[229] ,
    doutA_net[230] ,
    doutA_net[231] ,
    doutA_net[232] ,
    doutA_net[233] ,
    doutA_net[252] ,
    doutA_net[253] ,
    doutA_net[254] ,
    doutA_net[255] ,
    doutA_net[256] ,
    doutA_net[257] ,
    doutA_net[258] ,
    doutA_net[259] ,
    doutA_net[260] ,
    doutA_net[261] ,
    doutA_net[262] ,
    doutA_net[263] ,
    doutA_net[264] ,
    doutA_net[265] ,
    doutA_net[266] ,
    doutA_net[267] ,
    doutA_net[268] ,
    doutA_net[269] ,
    doutA_net[288] ,
    doutA_net[289] ,
    doutA_net[290] ,
    doutA_net[291] ,
    doutA_net[292] ,
    doutA_net[293] ,
    doutA_net[294] ,
    doutA_net[295] ,
    doutA_net[296] ,
    doutA_net[297] ,
    doutA_net[298] ,
    doutA_net[299] ,
    doutA_net[300] ,
    doutA_net[301] ,
    doutA_net[302] ,
    doutA_net[303] ,
    doutA_net[304] ,
    doutA_net[305] ,
    doutA_net[324] ,
    doutA_net[325] ,
    doutA_net[326] ,
    doutA_net[327] ,
    doutA_net[328] ,
    doutA_net[329] ,
    doutA_net[330] ,
    doutA_net[331] ,
    doutA_net[332] ,
    doutA_net[333] ,
    doutA_net[334] ,
    doutA_net[335] ,
    doutA_net[336] ,
    doutA_net[337] ,
    doutA_net[338] ,
    doutA_net[339] ,
    doutA_net[340] ,
    doutA_net[341] ,
    doutA_net[360] ,
    doutA_net[361] ,
    doutA_net[362] ,
    doutA_net[363] ,
    doutA_net[364] ,
    doutA_net[365] ,
    doutA_net[366] ,
    doutA_net[367] ,
    doutA_net[368] ,
    doutA_net[369] ,
    doutA_net[370] ,
    doutA_net[371] ,
    doutA_net[372] ,
    doutA_net[373] ,
    doutA_net[374] ,
    doutA_net[375] ,
    doutA_net[376] ,
    doutA_net[377] ,
    doutA_net[396] ,
    doutA_net[397] ,
    doutA_net[398] ,
    doutA_net[399] ,
    doutA_net[400] ,
    doutA_net[401] ,
    doutA_net[402] ,
    doutA_net[403] ,
    doutA_net[404] ,
    doutA_net[405] ,
    doutA_net[406] ,
    doutA_net[407] ,
    doutA_net[408] ,
    doutA_net[409] ,
    doutA_net[410] ,
    doutA_net[411] ,
    doutA_net[412] ,
    doutA_net[413] ,
    doutA_net[432] ,
    doutA_net[433] ,
    doutA_net[434] ,
    doutA_net[435] ,
    doutA_net[436] ,
    doutA_net[437] ,
    doutA_net[438] ,
    doutA_net[439] ,
    doutA_net[440] ,
    doutA_net[441] ,
    doutA_net[442] ,
    doutA_net[443] ,
    doutA_net[444] ,
    doutA_net[445] ,
    doutA_net[446] ,
    doutA_net[447] ,
    doutA_net[448] ,
    doutA_net[449] ,
    doutA_net[468] ,
    doutA_net[469] ,
    doutA_net[470] ,
    doutA_net[471] ,
    doutA_net[472] ,
    doutA_net[473] ,
    doutA_net[474] ,
    doutA_net[475] ,
    doutA_net[476] ,
    doutA_net[477] ,
    doutA_net[478] ,
    doutA_net[479] ,
    doutA_net[480] ,
    doutA_net[481] ,
    doutA_net[482] ,
    doutA_net[483] ,
    doutA_net[484] ,
    doutA_net[485] ,
    doutA_net[504] ,
    doutA_net[505] ,
    doutA_net[506] ,
    doutA_net[507] ,
    doutA_net[508] ,
    doutA_net[509] ,
    doutA_net[510] ,
    doutA_net[511] ,
    doutB_net[0] ,
    doutB_net[1] ,
    doutB_net[2] ,
    doutB_net[3] ,
    doutB_net[4] ,
    doutB_net[5] ,
    doutB_net[6] ,
    doutB_net[7] ,
    doutB_net[8] ,
    doutB_net[9] ,
    doutB_net[10] ,
    doutB_net[11] ,
    doutB_net[12] ,
    doutB_net[13] ,
    doutB_net[14] ,
    doutB_net[15] ,
    doutB_net[16] ,
    doutB_net[17] ,
    doutB_net[36] ,
    doutB_net[37] ,
    doutB_net[38] ,
    doutB_net[39] ,
    doutB_net[40] ,
    doutB_net[41] ,
    doutB_net[42] ,
    doutB_net[43] ,
    doutB_net[44] ,
    doutB_net[45] ,
    doutB_net[46] ,
    doutB_net[47] ,
    doutB_net[48] ,
    doutB_net[49] ,
    doutB_net[50] ,
    doutB_net[51] ,
    doutB_net[52] ,
    doutB_net[53] ,
    doutB_net[72] ,
    doutB_net[73] ,
    doutB_net[74] ,
    doutB_net[75] ,
    doutB_net[76] ,
    doutB_net[77] ,
    doutB_net[78] ,
    doutB_net[79] ,
    doutB_net[80] ,
    doutB_net[81] ,
    doutB_net[82] ,
    doutB_net[83] ,
    doutB_net[84] ,
    doutB_net[85] ,
    doutB_net[86] ,
    doutB_net[87] ,
    doutB_net[88] ,
    doutB_net[89] ,
    doutB_net[108] ,
    doutB_net[109] ,
    doutB_net[110] ,
    doutB_net[111] ,
    doutB_net[112] ,
    doutB_net[113] ,
    doutB_net[114] ,
    doutB_net[115] ,
    doutB_net[116] ,
    doutB_net[117] ,
    doutB_net[118] ,
    doutB_net[119] ,
    doutB_net[120] ,
    doutB_net[121] ,
    doutB_net[122] ,
    doutB_net[123] ,
    doutB_net[124] ,
    doutB_net[125] ,
    doutB_net[144] ,
    doutB_net[145] ,
    doutB_net[146] ,
    doutB_net[147] ,
    doutB_net[148] ,
    doutB_net[149] ,
    doutB_net[150] ,
    doutB_net[151] ,
    doutB_net[152] ,
    doutB_net[153] ,
    doutB_net[154] ,
    doutB_net[155] ,
    doutB_net[156] ,
    doutB_net[157] ,
    doutB_net[158] ,
    doutB_net[159] ,
    doutB_net[160] ,
    doutB_net[161] ,
    doutB_net[180] ,
    doutB_net[181] ,
    doutB_net[182] ,
    doutB_net[183] ,
    doutB_net[184] ,
    doutB_net[185] ,
    doutB_net[186] ,
    doutB_net[187] ,
    doutB_net[188] ,
    doutB_net[189] ,
    doutB_net[190] ,
    doutB_net[191] ,
    doutB_net[192] ,
    doutB_net[193] ,
    doutB_net[194] ,
    doutB_net[195] ,
    doutB_net[196] ,
    doutB_net[197] ,
    doutB_net[216] ,
    doutB_net[217] ,
    doutB_net[218] ,
    doutB_net[219] ,
    doutB_net[220] ,
    doutB_net[221] ,
    doutB_net[222] ,
    doutB_net[223] ,
    doutB_net[224] ,
    doutB_net[225] ,
    doutB_net[226] ,
    doutB_net[227] ,
    doutB_net[228] ,
    doutB_net[229] ,
    doutB_net[230] ,
    doutB_net[231] ,
    doutB_net[232] ,
    doutB_net[233] ,
    doutB_net[252] ,
    doutB_net[253] ,
    doutB_net[254] ,
    doutB_net[255] ,
    doutB_net[256] ,
    doutB_net[257] ,
    doutB_net[258] ,
    doutB_net[259] ,
    doutB_net[260] ,
    doutB_net[261] ,
    doutB_net[262] ,
    doutB_net[263] ,
    doutB_net[264] ,
    doutB_net[265] ,
    doutB_net[266] ,
    doutB_net[267] ,
    doutB_net[268] ,
    doutB_net[269] ,
    doutB_net[288] ,
    doutB_net[289] ,
    doutB_net[290] ,
    doutB_net[291] ,
    doutB_net[292] ,
    doutB_net[293] ,
    doutB_net[294] ,
    doutB_net[295] ,
    doutB_net[296] ,
    doutB_net[297] ,
    doutB_net[298] ,
    doutB_net[299] ,
    doutB_net[300] ,
    doutB_net[301] ,
    doutB_net[302] ,
    doutB_net[303] ,
    doutB_net[304] ,
    doutB_net[305] ,
    doutB_net[324] ,
    doutB_net[325] ,
    doutB_net[326] ,
    doutB_net[327] ,
    doutB_net[328] ,
    doutB_net[329] ,
    doutB_net[330] ,
    doutB_net[331] ,
    doutB_net[332] ,
    doutB_net[333] ,
    doutB_net[334] ,
    doutB_net[335] ,
    doutB_net[336] ,
    doutB_net[337] ,
    doutB_net[338] ,
    doutB_net[339] ,
    doutB_net[340] ,
    doutB_net[341] ,
    doutB_net[360] ,
    doutB_net[361] ,
    doutB_net[362] ,
    doutB_net[363] ,
    doutB_net[364] ,
    doutB_net[365] ,
    doutB_net[366] ,
    doutB_net[367] ,
    doutB_net[368] ,
    doutB_net[369] ,
    doutB_net[370] ,
    doutB_net[371] ,
    doutB_net[372] ,
    doutB_net[373] ,
    doutB_net[374] ,
    doutB_net[375] ,
    doutB_net[376] ,
    doutB_net[377] ,
    doutB_net[396] ,
    doutB_net[397] ,
    doutB_net[398] ,
    doutB_net[399] ,
    doutB_net[400] ,
    doutB_net[402] ,
    doutB_net[403] ,
    doutB_net[404] ,
    doutB_net[405] ,
    doutB_net[406] ,
    doutB_net[407] ,
    doutB_net[408] ,
    doutB_net[409] ,
    doutB_net[410] ,
    doutB_net[411] ,
    doutB_net[412] ,
    doutB_net[413] ,
    doutB_net[432] ,
    doutB_net[433] ,
    doutB_net[434] ,
    doutB_net[435] ,
    doutB_net[436] ,
    doutB_net[437] ,
    doutB_net[438] ,
    doutB_net[439] ,
    doutB_net[440] ,
    doutB_net[441] ,
    doutB_net[442] ,
    doutB_net[443] ,
    doutB_net[444] ,
    doutB_net[445] ,
    doutB_net[446] ,
    doutB_net[447] ,
    doutB_net[448] ,
    doutB_net[449] ,
    doutB_net[468] ,
    doutB_net[469] ,
    doutB_net[470] ,
    doutB_net[471] ,
    doutB_net[472] ,
    doutB_net[473] ,
    doutB_net[474] ,
    doutB_net[475] ,
    doutB_net[476] ,
    doutB_net[477] ,
    doutB_net[478] ,
    doutB_net[479] ,
    doutB_net[480] ,
    doutB_net[481] ,
    doutB_net[482] ,
    doutB_net[483] ,
    doutB_net[484] ,
    doutB_net[485] ,
    doutB_net[504] ,
    doutB_net[505] ,
    doutB_net[506] ,
    doutB_net[507] ,
    doutB_net[508] ,
    doutB_net[509] ,
    doutB_net[510] ,
    doutB_net[511] ,
    doutA_net[18] ,
    doutA_net[19] ,
    doutA_net[20] ,
    doutA_net[21] ,
    doutA_net[22] ,
    doutA_net[23] ,
    doutA_net[24] ,
    doutA_net[25] ,
    doutA_net[26] ,
    doutA_net[27] ,
    doutA_net[28] ,
    doutA_net[29] ,
    doutA_net[30] ,
    doutA_net[31] ,
    doutA_net[32] ,
    doutA_net[33] ,
    doutA_net[34] ,
    doutA_net[35] ,
    doutA_net[54] ,
    doutA_net[55] ,
    doutA_net[56] ,
    doutA_net[57] ,
    doutA_net[58] ,
    doutA_net[59] ,
    doutA_net[60] ,
    doutA_net[61] ,
    doutA_net[62] ,
    doutA_net[63] ,
    doutA_net[64] ,
    doutA_net[65] ,
    doutA_net[66] ,
    doutA_net[67] ,
    doutA_net[68] ,
    doutA_net[69] ,
    doutA_net[70] ,
    doutA_net[71] ,
    doutA_net[90] ,
    doutA_net[91] ,
    doutA_net[92] ,
    doutA_net[93] ,
    doutA_net[94] ,
    doutA_net[95] ,
    doutA_net[96] ,
    doutA_net[97] ,
    doutA_net[98] ,
    doutA_net[99] ,
    doutA_net[100] ,
    doutA_net[101] ,
    doutA_net[102] ,
    doutA_net[103] ,
    doutA_net[104] ,
    doutA_net[105] ,
    doutA_net[106] ,
    doutA_net[107] ,
    doutA_net[126] ,
    doutA_net[127] ,
    doutA_net[128] ,
    doutA_net[129] ,
    doutA_net[130] ,
    doutA_net[131] ,
    doutA_net[132] ,
    doutA_net[133] ,
    doutA_net[134] ,
    doutA_net[135] ,
    doutA_net[136] ,
    doutA_net[137] ,
    doutA_net[138] ,
    doutA_net[139] ,
    doutA_net[140] ,
    doutA_net[141] ,
    doutA_net[142] ,
    doutA_net[143] ,
    doutA_net[162] ,
    doutA_net[163] ,
    doutA_net[164] ,
    doutA_net[165] ,
    doutA_net[166] ,
    doutA_net[167] ,
    doutA_net[168] ,
    doutA_net[169] ,
    doutA_net[170] ,
    doutA_net[171] ,
    doutA_net[172] ,
    doutA_net[173] ,
    doutA_net[174] ,
    doutA_net[175] ,
    doutA_net[176] ,
    doutA_net[177] ,
    doutA_net[178] ,
    doutA_net[179] ,
    doutA_net[198] ,
    doutA_net[199] ,
    doutA_net[200] ,
    doutA_net[201] ,
    doutA_net[202] ,
    doutA_net[203] ,
    doutA_net[204] ,
    doutA_net[205] ,
    doutA_net[206] ,
    doutA_net[207] ,
    doutA_net[208] ,
    doutA_net[209] ,
    doutA_net[210] ,
    doutA_net[211] ,
    doutA_net[212] ,
    doutA_net[213] ,
    doutA_net[214] ,
    doutA_net[215] ,
    doutA_net[234] ,
    doutA_net[235] ,
    doutA_net[236] ,
    doutA_net[237] ,
    doutA_net[238] ,
    doutA_net[239] ,
    doutA_net[240] ,
    doutA_net[241] ,
    doutA_net[242] ,
    doutA_net[243] ,
    doutA_net[244] ,
    doutA_net[245] ,
    doutA_net[246] ,
    doutA_net[247] ,
    doutA_net[248] ,
    doutA_net[249] ,
    doutA_net[250] ,
    doutA_net[251] ,
    doutA_net[270] ,
    doutA_net[271] ,
    doutA_net[272] ,
    doutA_net[273] ,
    doutA_net[274] ,
    doutA_net[275] ,
    doutA_net[276] ,
    doutA_net[277] ,
    doutA_net[278] ,
    doutA_net[279] ,
    doutA_net[280] ,
    doutA_net[281] ,
    doutA_net[282] ,
    doutA_net[283] ,
    doutA_net[284] ,
    doutA_net[285] ,
    doutA_net[286] ,
    doutA_net[287] ,
    doutA_net[306] ,
    doutA_net[307] ,
    doutA_net[308] ,
    doutA_net[309] ,
    doutA_net[310] ,
    doutA_net[311] ,
    doutA_net[312] ,
    doutA_net[313] ,
    doutA_net[314] ,
    doutA_net[315] ,
    doutA_net[316] ,
    doutA_net[317] ,
    doutA_net[318] ,
    doutA_net[319] ,
    doutA_net[320] ,
    doutA_net[321] ,
    doutA_net[322] ,
    doutA_net[323] ,
    doutA_net[342] ,
    doutA_net[343] ,
    doutA_net[344] ,
    doutA_net[345] ,
    doutA_net[346] ,
    doutA_net[347] ,
    doutA_net[348] ,
    doutA_net[349] ,
    doutA_net[350] ,
    doutA_net[351] ,
    doutA_net[352] ,
    doutA_net[353] ,
    doutA_net[354] ,
    doutA_net[355] ,
    doutA_net[356] ,
    doutA_net[357] ,
    doutA_net[358] ,
    doutA_net[359] ,
    doutA_net[378] ,
    doutA_net[379] ,
    doutA_net[380] ,
    doutA_net[381] ,
    doutA_net[382] ,
    doutA_net[383] ,
    doutA_net[384] ,
    doutA_net[385] ,
    doutA_net[386] ,
    doutA_net[387] ,
    doutA_net[388] ,
    doutA_net[389] ,
    doutA_net[390] ,
    doutA_net[391] ,
    doutA_net[392] ,
    doutA_net[393] ,
    doutA_net[394] ,
    doutA_net[395] ,
    doutA_net[414] ,
    doutA_net[415] ,
    doutA_net[416] ,
    doutA_net[417] ,
    doutA_net[418] ,
    doutA_net[419] ,
    doutA_net[420] ,
    doutA_net[421] ,
    doutA_net[422] ,
    doutA_net[423] ,
    doutA_net[424] ,
    doutA_net[425] ,
    doutA_net[426] ,
    doutA_net[427] ,
    doutA_net[428] ,
    doutA_net[429] ,
    doutA_net[430] ,
    doutA_net[431] ,
    doutA_net[450] ,
    doutA_net[451] ,
    doutA_net[452] ,
    doutA_net[453] ,
    doutA_net[454] ,
    doutA_net[455] ,
    doutA_net[456] ,
    doutA_net[457] ,
    doutA_net[458] ,
    doutA_net[459] ,
    doutA_net[460] ,
    doutA_net[461] ,
    doutA_net[462] ,
    doutA_net[463] ,
    doutA_net[464] ,
    doutA_net[465] ,
    doutA_net[466] ,
    doutA_net[467] ,
    doutA_net[486] ,
    doutA_net[487] ,
    doutA_net[488] ,
    doutA_net[489] ,
    doutA_net[490] ,
    doutA_net[491] ,
    doutA_net[492] ,
    doutA_net[493] ,
    doutA_net[494] ,
    doutA_net[495] ,
    doutA_net[496] ,
    doutA_net[497] ,
    doutA_net[498] ,
    doutA_net[499] ,
    doutA_net[500] ,
    doutA_net[501] ,
    doutA_net[502] ,
    doutA_net[503] ,
    doutB_net[18] ,
    doutB_net[19] ,
    doutB_net[20] ,
    doutB_net[21] ,
    doutB_net[22] ,
    doutB_net[23] ,
    doutB_net[24] ,
    doutB_net[25] ,
    doutB_net[26] ,
    doutB_net[27] ,
    doutB_net[28] ,
    doutB_net[29] ,
    doutB_net[30] ,
    doutB_net[31] ,
    doutB_net[32] ,
    doutB_net[33] ,
    doutB_net[34] ,
    doutB_net[35] ,
    doutB_net[54] ,
    doutB_net[55] ,
    doutB_net[56] ,
    doutB_net[57] ,
    doutB_net[58] ,
    doutB_net[59] ,
    doutB_net[60] ,
    doutB_net[61] ,
    doutB_net[62] ,
    doutB_net[63] ,
    doutB_net[64] ,
    doutB_net[65] ,
    doutB_net[66] ,
    doutB_net[67] ,
    doutB_net[68] ,
    doutB_net[69] ,
    doutB_net[70] ,
    doutB_net[71] ,
    doutB_net[90] ,
    doutB_net[91] ,
    doutB_net[92] ,
    doutB_net[93] ,
    doutB_net[94] ,
    doutB_net[95] ,
    doutB_net[96] ,
    doutB_net[97] ,
    doutB_net[98] ,
    doutB_net[99] ,
    doutB_net[100] ,
    doutB_net[101] ,
    doutB_net[102] ,
    doutB_net[103] ,
    doutB_net[104] ,
    doutB_net[105] ,
    doutB_net[106] ,
    doutB_net[107] ,
    doutB_net[126] ,
    doutB_net[127] ,
    doutB_net[128] ,
    doutB_net[129] ,
    doutB_net[130] ,
    doutB_net[131] ,
    doutB_net[132] ,
    doutB_net[133] ,
    doutB_net[134] ,
    doutB_net[135] ,
    doutB_net[136] ,
    doutB_net[137] ,
    doutB_net[138] ,
    doutB_net[139] ,
    doutB_net[140] ,
    doutB_net[141] ,
    doutB_net[142] ,
    doutB_net[143] ,
    doutB_net[162] ,
    doutB_net[163] ,
    doutB_net[164] ,
    doutB_net[165] ,
    doutB_net[166] ,
    doutB_net[167] ,
    doutB_net[168] ,
    doutB_net[169] ,
    doutB_net[170] ,
    doutB_net[171] ,
    doutB_net[172] ,
    doutB_net[173] ,
    doutB_net[174] ,
    doutB_net[175] ,
    doutB_net[176] ,
    doutB_net[177] ,
    doutB_net[178] ,
    doutB_net[179] ,
    doutB_net[198] ,
    doutB_net[199] ,
    doutB_net[200] ,
    doutB_net[201] ,
    doutB_net[202] ,
    doutB_net[203] ,
    doutB_net[204] ,
    doutB_net[205] ,
    doutB_net[206] ,
    doutB_net[207] ,
    doutB_net[208] ,
    doutB_net[209] ,
    doutB_net[210] ,
    doutB_net[211] ,
    doutB_net[212] ,
    doutB_net[213] ,
    doutB_net[214] ,
    doutB_net[215] ,
    doutB_net[234] ,
    doutB_net[235] ,
    doutB_net[236] ,
    doutB_net[237] ,
    doutB_net[238] ,
    doutB_net[239] ,
    doutB_net[240] ,
    doutB_net[241] ,
    doutB_net[242] ,
    doutB_net[243] ,
    doutB_net[244] ,
    doutB_net[245] ,
    doutB_net[246] ,
    doutB_net[247] ,
    doutB_net[248] ,
    doutB_net[249] ,
    doutB_net[250] ,
    doutB_net[251] ,
    doutB_net[270] ,
    doutB_net[271] ,
    doutB_net[272] ,
    doutB_net[273] ,
    doutB_net[274] ,
    doutB_net[275] ,
    doutB_net[276] ,
    doutB_net[277] ,
    doutB_net[278] ,
    doutB_net[279] ,
    doutB_net[280] ,
    doutB_net[281] ,
    doutB_net[282] ,
    doutB_net[283] ,
    doutB_net[284] ,
    doutB_net[285] ,
    doutB_net[286] ,
    doutB_net[287] ,
    doutB_net[306] ,
    doutB_net[307] ,
    doutB_net[308] ,
    doutB_net[309] ,
    doutB_net[310] ,
    doutB_net[311] ,
    doutB_net[312] ,
    doutB_net[313] ,
    doutB_net[314] ,
    doutB_net[315] ,
    doutB_net[316] ,
    doutB_net[317] ,
    doutB_net[318] ,
    doutB_net[319] ,
    doutB_net[320] ,
    doutB_net[321] ,
    doutB_net[322] ,
    doutB_net[323] ,
    doutB_net[342] ,
    doutB_net[343] ,
    doutB_net[344] ,
    doutB_net[345] ,
    doutB_net[346] ,
    doutB_net[347] ,
    doutB_net[348] ,
    doutB_net[349] ,
    doutB_net[350] ,
    doutB_net[351] ,
    doutB_net[352] ,
    doutB_net[353] ,
    doutB_net[354] ,
    doutB_net[355] ,
    doutB_net[356] ,
    doutB_net[357] ,
    doutB_net[358] ,
    doutB_net[359] ,
    doutB_net[378] ,
    doutB_net[379] ,
    doutB_net[380] ,
    doutB_net[381] ,
    doutB_net[382] ,
    doutB_net[383] ,
    doutB_net[384] ,
    doutB_net[385] ,
    doutB_net[386] ,
    doutB_net[387] ,
    doutB_net[388] ,
    doutB_net[389] ,
    doutB_net[390] ,
    doutB_net[391] ,
    doutB_net[392] ,
    doutB_net[393] ,
    doutB_net[394] ,
    doutB_net[395] ,
    doutB_net[414] ,
    doutB_net[415] ,
    doutB_net[416] ,
    doutB_net[417] ,
    doutB_net[418] ,
    doutB_net[419] ,
    doutB_net[420] ,
    doutB_net[421] ,
    doutB_net[422] ,
    doutB_net[423] ,
    doutB_net[424] ,
    doutB_net[425] ,
    doutB_net[426] ,
    doutB_net[427] ,
    doutB_net[428] ,
    doutB_net[429] ,
    doutB_net[430] ,
    doutB_net[431] ,
    doutB_net[450] ,
    doutB_net[451] ,
    doutB_net[452] ,
    doutB_net[453] ,
    doutB_net[454] ,
    doutB_net[455] ,
    doutB_net[456] ,
    doutB_net[457] ,
    doutB_net[458] ,
    doutB_net[459] ,
    doutB_net[460] ,
    doutB_net[461] ,
    doutB_net[462] ,
    doutB_net[463] ,
    doutB_net[464] ,
    doutB_net[465] ,
    doutB_net[466] ,
    doutB_net[467] ,
    doutB_net[486] ,
    doutB_net[487] ,
    doutB_net[488] ,
    doutB_net[489] ,
    doutB_net[490] ,
    doutB_net[491] ,
    doutB_net[492] ,
    doutB_net[493] ,
    doutB_net[494] ,
    doutB_net[495] ,
    doutB_net[496] ,
    doutB_net[497] ,
    doutB_net[498] ,
    doutB_net[499] ,
    doutB_net[500] ,
    doutB_net[501] ,
    doutB_net[502] ,
    doutB_net[503] );
    `else
        tdp_512x10_post_synth netlist(.*, .doutA(doutA_net), .doutB(doutB_net));
    `endif

    
    //clock//
    initial begin
        clkA = 1'b0;
        forever #10 clkA = ~clkA;
    end
    initial begin
        clkB = 1'b0;
        forever #5 clkB = ~clkB;
    end

    initial begin
        for(integer i = 0; i<10; i=i+1) begin 
            golden.ram[i] ='b0;
        end 
    end
    initial begin
    {weA,weB, addrA,addrB, dinA, dinB, cycle, i} = 0;
 
 
    repeat (1) @ (negedge clkA);
    addrA <= 'd1; addrB <= 'd2; weA <=1'b1; weB <=1'b1; dinA<= {$random}; dinB<= {$random};
    compare(cycle);
    repeat (1) @ (negedge clkA);
    addrA <= 'd1; addrB <= 'd2; weA <=1'b0; weB <=1'b0; dinA<= {$random}; dinB<= {$random};
    compare(cycle);

    for (integer i=0; i<512; i=i+1)begin
        repeat (1) @ (negedge clkA)

        addrA <= $urandom_range(0,4); addrB <= $urandom_range(5,9); weA <=1'b1; weB <=1'b1; dinA<= {$random}; dinB<= {$random};
        cycle = cycle +1;
     
        compare(cycle);

    end

    for (integer i=0; i<512; i=i+1)begin
        repeat (1) @ (negedge clkB)

        addrA <= $urandom_range(0,4); addrB <= $urandom_range(5,9); weA <=1'b0; weB <=1'b0; dinA<= {$random}; dinB<= {$random};
        cycle = cycle +1;
     
        compare(cycle);

    end

    for (integer i=0; i<512; i=i+1)begin
        repeat (1) @ (negedge clkA)

        addrA <= $urandom_range(0,4); addrB <= $urandom_range(5,9); weA <=1'b0; weB <=1'b1; dinA<= {$random}; dinB<= {$random};
        cycle = cycle +1;
     
        compare(cycle);

    end

    for (integer i=0; i<512; i=i+1)begin
        repeat (1) @ (negedge clkB)

        addrA <= $urandom_range(0,4); addrB <= $urandom_range(5,9); weA <=1'b1; weB <=1'b0; dinA<= {$random}; dinB<= {$random};
        cycle = cycle +1;
     
        compare(cycle);

    end
    
    //random
    for (integer i=0; i<512; i=i+1)begin
        repeat (1) @ (negedge clkA)
        addrA <= $urandom_range(0,4); addrB <= $urandom_range(5,9); weA <={$random};  weB <={$random};  dinA<= {$random}; dinB<= {$random};
        cycle = cycle +1;
       
        compare(cycle);
    end
    if(mismatch == 0)
        $display("\n**** All Comparison Matched ***\nSimulation Passed");
    else
        $display("%0d comparison(s) mismatched\nERROR: SIM: Simulation Failed", mismatch);
    

    repeat (10) @(negedge clkA); $finish;
    end

    task compare(input integer cycle);
    //$display("\n Comparison at cycle %0d", cycle);
    if(doutA !== doutA_net) begin
        $display("doutA mismatch. Golden: %0h, Netlist: %0h, Time: %0t", doutA, doutA_net,$time);
        mismatch = mismatch+1;
    end

     if(doutB !== doutB_net) begin
        $display("doutB mismatch. Golden: %0h, Netlist: %0h, Time: %0t", doutB, doutB_net,$time);
        mismatch = mismatch+1;
    end
    
    
    endtask


initial begin
    $dumpfile("tb.vcd");
    $dumpvars;
end
endmodule