module LATCHN_primitive_inst_old(D, G, Q);
  input D;
  input G;
  output Q;

LATCHN inst (.*);

endmodule
