// `include "encoder.v"
// `include "invertion.v"
// `include "large_mux.v"
// `include "register.v"
module design26_30_50_top #(parameter WIDTH=32,CHANNEL=30) (clk, rst, in, out);

	localparam OUT_BUS=CHANNEL*WIDTH;
	input clk,rst;
	input [WIDTH-1:0] in;
	output [WIDTH-1:0] out;

	reg [WIDTH-1:0] d_in0;
	reg [WIDTH-1:0] d_in1;
	reg [WIDTH-1:0] d_in2;
	reg [WIDTH-1:0] d_in3;
	reg [WIDTH-1:0] d_in4;
	reg [WIDTH-1:0] d_in5;
	reg [WIDTH-1:0] d_in6;
	reg [WIDTH-1:0] d_in7;
	reg [WIDTH-1:0] d_in8;
	reg [WIDTH-1:0] d_in9;
	reg [WIDTH-1:0] d_in10;
	reg [WIDTH-1:0] d_in11;
	reg [WIDTH-1:0] d_in12;
	reg [WIDTH-1:0] d_in13;
	reg [WIDTH-1:0] d_in14;
	reg [WIDTH-1:0] d_in15;
	reg [WIDTH-1:0] d_in16;
	reg [WIDTH-1:0] d_in17;
	reg [WIDTH-1:0] d_in18;
	reg [WIDTH-1:0] d_in19;
	reg [WIDTH-1:0] d_in20;
	reg [WIDTH-1:0] d_in21;
	reg [WIDTH-1:0] d_in22;
	reg [WIDTH-1:0] d_in23;
	reg [WIDTH-1:0] d_in24;
	reg [WIDTH-1:0] d_in25;
	reg [WIDTH-1:0] d_in26;
	reg [WIDTH-1:0] d_in27;
	reg [WIDTH-1:0] d_in28;
	reg [WIDTH-1:0] d_in29;
	wire [WIDTH-1:0] d_out0;
	wire [WIDTH-1:0] d_out1;
	wire [WIDTH-1:0] d_out2;
	wire [WIDTH-1:0] d_out3;
	wire [WIDTH-1:0] d_out4;
	wire [WIDTH-1:0] d_out5;
	wire [WIDTH-1:0] d_out6;
	wire [WIDTH-1:0] d_out7;
	wire [WIDTH-1:0] d_out8;
	wire [WIDTH-1:0] d_out9;
	wire [WIDTH-1:0] d_out10;
	wire [WIDTH-1:0] d_out11;
	wire [WIDTH-1:0] d_out12;
	wire [WIDTH-1:0] d_out13;
	wire [WIDTH-1:0] d_out14;
	wire [WIDTH-1:0] d_out15;
	wire [WIDTH-1:0] d_out16;
	wire [WIDTH-1:0] d_out17;
	wire [WIDTH-1:0] d_out18;
	wire [WIDTH-1:0] d_out19;
	wire [WIDTH-1:0] d_out20;
	wire [WIDTH-1:0] d_out21;
	wire [WIDTH-1:0] d_out22;
	wire [WIDTH-1:0] d_out23;
	wire [WIDTH-1:0] d_out24;
	wire [WIDTH-1:0] d_out25;
	wire [WIDTH-1:0] d_out26;
	wire [WIDTH-1:0] d_out27;
	wire [WIDTH-1:0] d_out28;
	wire [WIDTH-1:0] d_out29;

	reg [OUT_BUS-1:0] tmp;

	always @ (posedge clk or posedge rst) begin
		if (rst)
			tmp <= 0;
		else
			tmp <= {tmp[OUT_BUS-(WIDTH-1):0],in};
	end

	always @ (posedge clk) begin
		d_in0 <= tmp[WIDTH-1:0];
		d_in1 <= tmp[(WIDTH*2)-1:WIDTH*1];
		d_in2 <= tmp[(WIDTH*3)-1:WIDTH*2];
		d_in3 <= tmp[(WIDTH*4)-1:WIDTH*3];
		d_in4 <= tmp[(WIDTH*5)-1:WIDTH*4];
		d_in5 <= tmp[(WIDTH*6)-1:WIDTH*5];
		d_in6 <= tmp[(WIDTH*7)-1:WIDTH*6];
		d_in7 <= tmp[(WIDTH*8)-1:WIDTH*7];
		d_in8 <= tmp[(WIDTH*9)-1:WIDTH*8];
		d_in9 <= tmp[(WIDTH*10)-1:WIDTH*9];
		d_in10 <= tmp[(WIDTH*11)-1:WIDTH*10];
		d_in11 <= tmp[(WIDTH*12)-1:WIDTH*11];
		d_in12 <= tmp[(WIDTH*13)-1:WIDTH*12];
		d_in13 <= tmp[(WIDTH*14)-1:WIDTH*13];
		d_in14 <= tmp[(WIDTH*15)-1:WIDTH*14];
		d_in15 <= tmp[(WIDTH*16)-1:WIDTH*15];
		d_in16 <= tmp[(WIDTH*17)-1:WIDTH*16];
		d_in17 <= tmp[(WIDTH*18)-1:WIDTH*17];
		d_in18 <= tmp[(WIDTH*19)-1:WIDTH*18];
		d_in19 <= tmp[(WIDTH*20)-1:WIDTH*19];
		d_in20 <= tmp[(WIDTH*21)-1:WIDTH*20];
		d_in21 <= tmp[(WIDTH*22)-1:WIDTH*21];
		d_in22 <= tmp[(WIDTH*23)-1:WIDTH*22];
		d_in23 <= tmp[(WIDTH*24)-1:WIDTH*23];
		d_in24 <= tmp[(WIDTH*25)-1:WIDTH*24];
		d_in25 <= tmp[(WIDTH*26)-1:WIDTH*25];
		d_in26 <= tmp[(WIDTH*27)-1:WIDTH*26];
		d_in27 <= tmp[(WIDTH*28)-1:WIDTH*27];
		d_in28 <= tmp[(WIDTH*29)-1:WIDTH*28];
		d_in29 <= tmp[(WIDTH*30)-1:WIDTH*29];
	end

	design26_30_50 #(.WIDTH(WIDTH)) design26_30_50_inst(.d_in0(d_in0),.d_in1(d_in1),.d_in2(d_in2),.d_in3(d_in3),.d_in4(d_in4),.d_in5(d_in5),.d_in6(d_in6),.d_in7(d_in7),.d_in8(d_in8),.d_in9(d_in9),.d_in10(d_in10),.d_in11(d_in11),.d_in12(d_in12),.d_in13(d_in13),.d_in14(d_in14),.d_in15(d_in15),.d_in16(d_in16),.d_in17(d_in17),.d_in18(d_in18),.d_in19(d_in19),.d_in20(d_in20),.d_in21(d_in21),.d_in22(d_in22),.d_in23(d_in23),.d_in24(d_in24),.d_in25(d_in25),.d_in26(d_in26),.d_in27(d_in27),.d_in28(d_in28),.d_in29(d_in29),.d_out0(d_out0),.d_out1(d_out1),.d_out2(d_out2),.d_out3(d_out3),.d_out4(d_out4),.d_out5(d_out5),.d_out6(d_out6),.d_out7(d_out7),.d_out8(d_out8),.d_out9(d_out9),.d_out10(d_out10),.d_out11(d_out11),.d_out12(d_out12),.d_out13(d_out13),.d_out14(d_out14),.d_out15(d_out15),.d_out16(d_out16),.d_out17(d_out17),.d_out18(d_out18),.d_out19(d_out19),.d_out20(d_out20),.d_out21(d_out21),.d_out22(d_out22),.d_out23(d_out23),.d_out24(d_out24),.d_out25(d_out25),.d_out26(d_out26),.d_out27(d_out27),.d_out28(d_out28),.d_out29(d_out29),.clk(clk),.rst(rst));

	assign out = d_out0^d_out1^d_out2^d_out3^d_out4^d_out5^d_out6^d_out7^d_out8^d_out9^d_out10^d_out11^d_out12^d_out13^d_out14^d_out15^d_out16^d_out17^d_out18^d_out19^d_out20^d_out21^d_out22^d_out23^d_out24^d_out25^d_out26^d_out27^d_out28^d_out29;

endmodule

module design26_30_50 #(parameter WIDTH=32) (d_in0, d_in1, d_in2, d_in3, d_in4, d_in5, d_in6, d_in7, d_in8, d_in9, d_in10, d_in11, d_in12, d_in13, d_in14, d_in15, d_in16, d_in17, d_in18, d_in19, d_in20, d_in21, d_in22, d_in23, d_in24, d_in25, d_in26, d_in27, d_in28, d_in29, d_out0, d_out1, d_out2, d_out3, d_out4, d_out5, d_out6, d_out7, d_out8, d_out9, d_out10, d_out11, d_out12, d_out13, d_out14, d_out15, d_out16, d_out17, d_out18, d_out19, d_out20, d_out21, d_out22, d_out23, d_out24, d_out25, d_out26, d_out27, d_out28, d_out29, clk, rst);
	input clk;
	input rst;
	input [WIDTH-1:0] d_in0; 
	input [WIDTH-1:0] d_in1; 
	input [WIDTH-1:0] d_in2; 
	input [WIDTH-1:0] d_in3; 
	input [WIDTH-1:0] d_in4; 
	input [WIDTH-1:0] d_in5; 
	input [WIDTH-1:0] d_in6; 
	input [WIDTH-1:0] d_in7; 
	input [WIDTH-1:0] d_in8; 
	input [WIDTH-1:0] d_in9; 
	input [WIDTH-1:0] d_in10; 
	input [WIDTH-1:0] d_in11; 
	input [WIDTH-1:0] d_in12; 
	input [WIDTH-1:0] d_in13; 
	input [WIDTH-1:0] d_in14; 
	input [WIDTH-1:0] d_in15; 
	input [WIDTH-1:0] d_in16; 
	input [WIDTH-1:0] d_in17; 
	input [WIDTH-1:0] d_in18; 
	input [WIDTH-1:0] d_in19; 
	input [WIDTH-1:0] d_in20; 
	input [WIDTH-1:0] d_in21; 
	input [WIDTH-1:0] d_in22; 
	input [WIDTH-1:0] d_in23; 
	input [WIDTH-1:0] d_in24; 
	input [WIDTH-1:0] d_in25; 
	input [WIDTH-1:0] d_in26; 
	input [WIDTH-1:0] d_in27; 
	input [WIDTH-1:0] d_in28; 
	input [WIDTH-1:0] d_in29; 
	output [WIDTH-1:0] d_out0; 
	output [WIDTH-1:0] d_out1; 
	output [WIDTH-1:0] d_out2; 
	output [WIDTH-1:0] d_out3; 
	output [WIDTH-1:0] d_out4; 
	output [WIDTH-1:0] d_out5; 
	output [WIDTH-1:0] d_out6; 
	output [WIDTH-1:0] d_out7; 
	output [WIDTH-1:0] d_out8; 
	output [WIDTH-1:0] d_out9; 
	output [WIDTH-1:0] d_out10; 
	output [WIDTH-1:0] d_out11; 
	output [WIDTH-1:0] d_out12; 
	output [WIDTH-1:0] d_out13; 
	output [WIDTH-1:0] d_out14; 
	output [WIDTH-1:0] d_out15; 
	output [WIDTH-1:0] d_out16; 
	output [WIDTH-1:0] d_out17; 
	output [WIDTH-1:0] d_out18; 
	output [WIDTH-1:0] d_out19; 
	output [WIDTH-1:0] d_out20; 
	output [WIDTH-1:0] d_out21; 
	output [WIDTH-1:0] d_out22; 
	output [WIDTH-1:0] d_out23; 
	output [WIDTH-1:0] d_out24; 
	output [WIDTH-1:0] d_out25; 
	output [WIDTH-1:0] d_out26; 
	output [WIDTH-1:0] d_out27; 
	output [WIDTH-1:0] d_out28; 
	output [WIDTH-1:0] d_out29; 

	wire [WIDTH-1:0] wire_d0_0;
	wire [WIDTH-1:0] wire_d0_1;
	wire [WIDTH-1:0] wire_d0_2;
	wire [WIDTH-1:0] wire_d0_3;
	wire [WIDTH-1:0] wire_d0_4;
	wire [WIDTH-1:0] wire_d0_5;
	wire [WIDTH-1:0] wire_d0_6;
	wire [WIDTH-1:0] wire_d0_7;
	wire [WIDTH-1:0] wire_d0_8;
	wire [WIDTH-1:0] wire_d0_9;
	wire [WIDTH-1:0] wire_d0_10;
	wire [WIDTH-1:0] wire_d0_11;
	wire [WIDTH-1:0] wire_d0_12;
	wire [WIDTH-1:0] wire_d0_13;
	wire [WIDTH-1:0] wire_d0_14;
	wire [WIDTH-1:0] wire_d0_15;
	wire [WIDTH-1:0] wire_d0_16;
	wire [WIDTH-1:0] wire_d0_17;
	wire [WIDTH-1:0] wire_d0_18;
	wire [WIDTH-1:0] wire_d0_19;
	wire [WIDTH-1:0] wire_d0_20;
	wire [WIDTH-1:0] wire_d0_21;
	wire [WIDTH-1:0] wire_d0_22;
	wire [WIDTH-1:0] wire_d0_23;
	wire [WIDTH-1:0] wire_d0_24;
	wire [WIDTH-1:0] wire_d0_25;
	wire [WIDTH-1:0] wire_d0_26;
	wire [WIDTH-1:0] wire_d0_27;
	wire [WIDTH-1:0] wire_d0_28;
	wire [WIDTH-1:0] wire_d0_29;
	wire [WIDTH-1:0] wire_d0_30;
	wire [WIDTH-1:0] wire_d0_31;
	wire [WIDTH-1:0] wire_d0_32;
	wire [WIDTH-1:0] wire_d0_33;
	wire [WIDTH-1:0] wire_d0_34;
	wire [WIDTH-1:0] wire_d0_35;
	wire [WIDTH-1:0] wire_d0_36;
	wire [WIDTH-1:0] wire_d0_37;
	wire [WIDTH-1:0] wire_d0_38;
	wire [WIDTH-1:0] wire_d0_39;
	wire [WIDTH-1:0] wire_d0_40;
	wire [WIDTH-1:0] wire_d0_41;
	wire [WIDTH-1:0] wire_d0_42;
	wire [WIDTH-1:0] wire_d0_43;
	wire [WIDTH-1:0] wire_d0_44;
	wire [WIDTH-1:0] wire_d0_45;
	wire [WIDTH-1:0] wire_d0_46;
	wire [WIDTH-1:0] wire_d0_47;
	wire [WIDTH-1:0] wire_d0_48;
	wire [WIDTH-1:0] wire_d1_0;
	wire [WIDTH-1:0] wire_d1_1;
	wire [WIDTH-1:0] wire_d1_2;
	wire [WIDTH-1:0] wire_d1_3;
	wire [WIDTH-1:0] wire_d1_4;
	wire [WIDTH-1:0] wire_d1_5;
	wire [WIDTH-1:0] wire_d1_6;
	wire [WIDTH-1:0] wire_d1_7;
	wire [WIDTH-1:0] wire_d1_8;
	wire [WIDTH-1:0] wire_d1_9;
	wire [WIDTH-1:0] wire_d1_10;
	wire [WIDTH-1:0] wire_d1_11;
	wire [WIDTH-1:0] wire_d1_12;
	wire [WIDTH-1:0] wire_d1_13;
	wire [WIDTH-1:0] wire_d1_14;
	wire [WIDTH-1:0] wire_d1_15;
	wire [WIDTH-1:0] wire_d1_16;
	wire [WIDTH-1:0] wire_d1_17;
	wire [WIDTH-1:0] wire_d1_18;
	wire [WIDTH-1:0] wire_d1_19;
	wire [WIDTH-1:0] wire_d1_20;
	wire [WIDTH-1:0] wire_d1_21;
	wire [WIDTH-1:0] wire_d1_22;
	wire [WIDTH-1:0] wire_d1_23;
	wire [WIDTH-1:0] wire_d1_24;
	wire [WIDTH-1:0] wire_d1_25;
	wire [WIDTH-1:0] wire_d1_26;
	wire [WIDTH-1:0] wire_d1_27;
	wire [WIDTH-1:0] wire_d1_28;
	wire [WIDTH-1:0] wire_d1_29;
	wire [WIDTH-1:0] wire_d1_30;
	wire [WIDTH-1:0] wire_d1_31;
	wire [WIDTH-1:0] wire_d1_32;
	wire [WIDTH-1:0] wire_d1_33;
	wire [WIDTH-1:0] wire_d1_34;
	wire [WIDTH-1:0] wire_d1_35;
	wire [WIDTH-1:0] wire_d1_36;
	wire [WIDTH-1:0] wire_d1_37;
	wire [WIDTH-1:0] wire_d1_38;
	wire [WIDTH-1:0] wire_d1_39;
	wire [WIDTH-1:0] wire_d1_40;
	wire [WIDTH-1:0] wire_d1_41;
	wire [WIDTH-1:0] wire_d1_42;
	wire [WIDTH-1:0] wire_d1_43;
	wire [WIDTH-1:0] wire_d1_44;
	wire [WIDTH-1:0] wire_d1_45;
	wire [WIDTH-1:0] wire_d1_46;
	wire [WIDTH-1:0] wire_d1_47;
	wire [WIDTH-1:0] wire_d1_48;
	wire [WIDTH-1:0] wire_d2_0;
	wire [WIDTH-1:0] wire_d2_1;
	wire [WIDTH-1:0] wire_d2_2;
	wire [WIDTH-1:0] wire_d2_3;
	wire [WIDTH-1:0] wire_d2_4;
	wire [WIDTH-1:0] wire_d2_5;
	wire [WIDTH-1:0] wire_d2_6;
	wire [WIDTH-1:0] wire_d2_7;
	wire [WIDTH-1:0] wire_d2_8;
	wire [WIDTH-1:0] wire_d2_9;
	wire [WIDTH-1:0] wire_d2_10;
	wire [WIDTH-1:0] wire_d2_11;
	wire [WIDTH-1:0] wire_d2_12;
	wire [WIDTH-1:0] wire_d2_13;
	wire [WIDTH-1:0] wire_d2_14;
	wire [WIDTH-1:0] wire_d2_15;
	wire [WIDTH-1:0] wire_d2_16;
	wire [WIDTH-1:0] wire_d2_17;
	wire [WIDTH-1:0] wire_d2_18;
	wire [WIDTH-1:0] wire_d2_19;
	wire [WIDTH-1:0] wire_d2_20;
	wire [WIDTH-1:0] wire_d2_21;
	wire [WIDTH-1:0] wire_d2_22;
	wire [WIDTH-1:0] wire_d2_23;
	wire [WIDTH-1:0] wire_d2_24;
	wire [WIDTH-1:0] wire_d2_25;
	wire [WIDTH-1:0] wire_d2_26;
	wire [WIDTH-1:0] wire_d2_27;
	wire [WIDTH-1:0] wire_d2_28;
	wire [WIDTH-1:0] wire_d2_29;
	wire [WIDTH-1:0] wire_d2_30;
	wire [WIDTH-1:0] wire_d2_31;
	wire [WIDTH-1:0] wire_d2_32;
	wire [WIDTH-1:0] wire_d2_33;
	wire [WIDTH-1:0] wire_d2_34;
	wire [WIDTH-1:0] wire_d2_35;
	wire [WIDTH-1:0] wire_d2_36;
	wire [WIDTH-1:0] wire_d2_37;
	wire [WIDTH-1:0] wire_d2_38;
	wire [WIDTH-1:0] wire_d2_39;
	wire [WIDTH-1:0] wire_d2_40;
	wire [WIDTH-1:0] wire_d2_41;
	wire [WIDTH-1:0] wire_d2_42;
	wire [WIDTH-1:0] wire_d2_43;
	wire [WIDTH-1:0] wire_d2_44;
	wire [WIDTH-1:0] wire_d2_45;
	wire [WIDTH-1:0] wire_d2_46;
	wire [WIDTH-1:0] wire_d2_47;
	wire [WIDTH-1:0] wire_d2_48;
	wire [WIDTH-1:0] wire_d3_0;
	wire [WIDTH-1:0] wire_d3_1;
	wire [WIDTH-1:0] wire_d3_2;
	wire [WIDTH-1:0] wire_d3_3;
	wire [WIDTH-1:0] wire_d3_4;
	wire [WIDTH-1:0] wire_d3_5;
	wire [WIDTH-1:0] wire_d3_6;
	wire [WIDTH-1:0] wire_d3_7;
	wire [WIDTH-1:0] wire_d3_8;
	wire [WIDTH-1:0] wire_d3_9;
	wire [WIDTH-1:0] wire_d3_10;
	wire [WIDTH-1:0] wire_d3_11;
	wire [WIDTH-1:0] wire_d3_12;
	wire [WIDTH-1:0] wire_d3_13;
	wire [WIDTH-1:0] wire_d3_14;
	wire [WIDTH-1:0] wire_d3_15;
	wire [WIDTH-1:0] wire_d3_16;
	wire [WIDTH-1:0] wire_d3_17;
	wire [WIDTH-1:0] wire_d3_18;
	wire [WIDTH-1:0] wire_d3_19;
	wire [WIDTH-1:0] wire_d3_20;
	wire [WIDTH-1:0] wire_d3_21;
	wire [WIDTH-1:0] wire_d3_22;
	wire [WIDTH-1:0] wire_d3_23;
	wire [WIDTH-1:0] wire_d3_24;
	wire [WIDTH-1:0] wire_d3_25;
	wire [WIDTH-1:0] wire_d3_26;
	wire [WIDTH-1:0] wire_d3_27;
	wire [WIDTH-1:0] wire_d3_28;
	wire [WIDTH-1:0] wire_d3_29;
	wire [WIDTH-1:0] wire_d3_30;
	wire [WIDTH-1:0] wire_d3_31;
	wire [WIDTH-1:0] wire_d3_32;
	wire [WIDTH-1:0] wire_d3_33;
	wire [WIDTH-1:0] wire_d3_34;
	wire [WIDTH-1:0] wire_d3_35;
	wire [WIDTH-1:0] wire_d3_36;
	wire [WIDTH-1:0] wire_d3_37;
	wire [WIDTH-1:0] wire_d3_38;
	wire [WIDTH-1:0] wire_d3_39;
	wire [WIDTH-1:0] wire_d3_40;
	wire [WIDTH-1:0] wire_d3_41;
	wire [WIDTH-1:0] wire_d3_42;
	wire [WIDTH-1:0] wire_d3_43;
	wire [WIDTH-1:0] wire_d3_44;
	wire [WIDTH-1:0] wire_d3_45;
	wire [WIDTH-1:0] wire_d3_46;
	wire [WIDTH-1:0] wire_d3_47;
	wire [WIDTH-1:0] wire_d3_48;
	wire [WIDTH-1:0] wire_d4_0;
	wire [WIDTH-1:0] wire_d4_1;
	wire [WIDTH-1:0] wire_d4_2;
	wire [WIDTH-1:0] wire_d4_3;
	wire [WIDTH-1:0] wire_d4_4;
	wire [WIDTH-1:0] wire_d4_5;
	wire [WIDTH-1:0] wire_d4_6;
	wire [WIDTH-1:0] wire_d4_7;
	wire [WIDTH-1:0] wire_d4_8;
	wire [WIDTH-1:0] wire_d4_9;
	wire [WIDTH-1:0] wire_d4_10;
	wire [WIDTH-1:0] wire_d4_11;
	wire [WIDTH-1:0] wire_d4_12;
	wire [WIDTH-1:0] wire_d4_13;
	wire [WIDTH-1:0] wire_d4_14;
	wire [WIDTH-1:0] wire_d4_15;
	wire [WIDTH-1:0] wire_d4_16;
	wire [WIDTH-1:0] wire_d4_17;
	wire [WIDTH-1:0] wire_d4_18;
	wire [WIDTH-1:0] wire_d4_19;
	wire [WIDTH-1:0] wire_d4_20;
	wire [WIDTH-1:0] wire_d4_21;
	wire [WIDTH-1:0] wire_d4_22;
	wire [WIDTH-1:0] wire_d4_23;
	wire [WIDTH-1:0] wire_d4_24;
	wire [WIDTH-1:0] wire_d4_25;
	wire [WIDTH-1:0] wire_d4_26;
	wire [WIDTH-1:0] wire_d4_27;
	wire [WIDTH-1:0] wire_d4_28;
	wire [WIDTH-1:0] wire_d4_29;
	wire [WIDTH-1:0] wire_d4_30;
	wire [WIDTH-1:0] wire_d4_31;
	wire [WIDTH-1:0] wire_d4_32;
	wire [WIDTH-1:0] wire_d4_33;
	wire [WIDTH-1:0] wire_d4_34;
	wire [WIDTH-1:0] wire_d4_35;
	wire [WIDTH-1:0] wire_d4_36;
	wire [WIDTH-1:0] wire_d4_37;
	wire [WIDTH-1:0] wire_d4_38;
	wire [WIDTH-1:0] wire_d4_39;
	wire [WIDTH-1:0] wire_d4_40;
	wire [WIDTH-1:0] wire_d4_41;
	wire [WIDTH-1:0] wire_d4_42;
	wire [WIDTH-1:0] wire_d4_43;
	wire [WIDTH-1:0] wire_d4_44;
	wire [WIDTH-1:0] wire_d4_45;
	wire [WIDTH-1:0] wire_d4_46;
	wire [WIDTH-1:0] wire_d4_47;
	wire [WIDTH-1:0] wire_d4_48;
	wire [WIDTH-1:0] wire_d5_0;
	wire [WIDTH-1:0] wire_d5_1;
	wire [WIDTH-1:0] wire_d5_2;
	wire [WIDTH-1:0] wire_d5_3;
	wire [WIDTH-1:0] wire_d5_4;
	wire [WIDTH-1:0] wire_d5_5;
	wire [WIDTH-1:0] wire_d5_6;
	wire [WIDTH-1:0] wire_d5_7;
	wire [WIDTH-1:0] wire_d5_8;
	wire [WIDTH-1:0] wire_d5_9;
	wire [WIDTH-1:0] wire_d5_10;
	wire [WIDTH-1:0] wire_d5_11;
	wire [WIDTH-1:0] wire_d5_12;
	wire [WIDTH-1:0] wire_d5_13;
	wire [WIDTH-1:0] wire_d5_14;
	wire [WIDTH-1:0] wire_d5_15;
	wire [WIDTH-1:0] wire_d5_16;
	wire [WIDTH-1:0] wire_d5_17;
	wire [WIDTH-1:0] wire_d5_18;
	wire [WIDTH-1:0] wire_d5_19;
	wire [WIDTH-1:0] wire_d5_20;
	wire [WIDTH-1:0] wire_d5_21;
	wire [WIDTH-1:0] wire_d5_22;
	wire [WIDTH-1:0] wire_d5_23;
	wire [WIDTH-1:0] wire_d5_24;
	wire [WIDTH-1:0] wire_d5_25;
	wire [WIDTH-1:0] wire_d5_26;
	wire [WIDTH-1:0] wire_d5_27;
	wire [WIDTH-1:0] wire_d5_28;
	wire [WIDTH-1:0] wire_d5_29;
	wire [WIDTH-1:0] wire_d5_30;
	wire [WIDTH-1:0] wire_d5_31;
	wire [WIDTH-1:0] wire_d5_32;
	wire [WIDTH-1:0] wire_d5_33;
	wire [WIDTH-1:0] wire_d5_34;
	wire [WIDTH-1:0] wire_d5_35;
	wire [WIDTH-1:0] wire_d5_36;
	wire [WIDTH-1:0] wire_d5_37;
	wire [WIDTH-1:0] wire_d5_38;
	wire [WIDTH-1:0] wire_d5_39;
	wire [WIDTH-1:0] wire_d5_40;
	wire [WIDTH-1:0] wire_d5_41;
	wire [WIDTH-1:0] wire_d5_42;
	wire [WIDTH-1:0] wire_d5_43;
	wire [WIDTH-1:0] wire_d5_44;
	wire [WIDTH-1:0] wire_d5_45;
	wire [WIDTH-1:0] wire_d5_46;
	wire [WIDTH-1:0] wire_d5_47;
	wire [WIDTH-1:0] wire_d5_48;
	wire [WIDTH-1:0] wire_d6_0;
	wire [WIDTH-1:0] wire_d6_1;
	wire [WIDTH-1:0] wire_d6_2;
	wire [WIDTH-1:0] wire_d6_3;
	wire [WIDTH-1:0] wire_d6_4;
	wire [WIDTH-1:0] wire_d6_5;
	wire [WIDTH-1:0] wire_d6_6;
	wire [WIDTH-1:0] wire_d6_7;
	wire [WIDTH-1:0] wire_d6_8;
	wire [WIDTH-1:0] wire_d6_9;
	wire [WIDTH-1:0] wire_d6_10;
	wire [WIDTH-1:0] wire_d6_11;
	wire [WIDTH-1:0] wire_d6_12;
	wire [WIDTH-1:0] wire_d6_13;
	wire [WIDTH-1:0] wire_d6_14;
	wire [WIDTH-1:0] wire_d6_15;
	wire [WIDTH-1:0] wire_d6_16;
	wire [WIDTH-1:0] wire_d6_17;
	wire [WIDTH-1:0] wire_d6_18;
	wire [WIDTH-1:0] wire_d6_19;
	wire [WIDTH-1:0] wire_d6_20;
	wire [WIDTH-1:0] wire_d6_21;
	wire [WIDTH-1:0] wire_d6_22;
	wire [WIDTH-1:0] wire_d6_23;
	wire [WIDTH-1:0] wire_d6_24;
	wire [WIDTH-1:0] wire_d6_25;
	wire [WIDTH-1:0] wire_d6_26;
	wire [WIDTH-1:0] wire_d6_27;
	wire [WIDTH-1:0] wire_d6_28;
	wire [WIDTH-1:0] wire_d6_29;
	wire [WIDTH-1:0] wire_d6_30;
	wire [WIDTH-1:0] wire_d6_31;
	wire [WIDTH-1:0] wire_d6_32;
	wire [WIDTH-1:0] wire_d6_33;
	wire [WIDTH-1:0] wire_d6_34;
	wire [WIDTH-1:0] wire_d6_35;
	wire [WIDTH-1:0] wire_d6_36;
	wire [WIDTH-1:0] wire_d6_37;
	wire [WIDTH-1:0] wire_d6_38;
	wire [WIDTH-1:0] wire_d6_39;
	wire [WIDTH-1:0] wire_d6_40;
	wire [WIDTH-1:0] wire_d6_41;
	wire [WIDTH-1:0] wire_d6_42;
	wire [WIDTH-1:0] wire_d6_43;
	wire [WIDTH-1:0] wire_d6_44;
	wire [WIDTH-1:0] wire_d6_45;
	wire [WIDTH-1:0] wire_d6_46;
	wire [WIDTH-1:0] wire_d6_47;
	wire [WIDTH-1:0] wire_d6_48;
	wire [WIDTH-1:0] wire_d7_0;
	wire [WIDTH-1:0] wire_d7_1;
	wire [WIDTH-1:0] wire_d7_2;
	wire [WIDTH-1:0] wire_d7_3;
	wire [WIDTH-1:0] wire_d7_4;
	wire [WIDTH-1:0] wire_d7_5;
	wire [WIDTH-1:0] wire_d7_6;
	wire [WIDTH-1:0] wire_d7_7;
	wire [WIDTH-1:0] wire_d7_8;
	wire [WIDTH-1:0] wire_d7_9;
	wire [WIDTH-1:0] wire_d7_10;
	wire [WIDTH-1:0] wire_d7_11;
	wire [WIDTH-1:0] wire_d7_12;
	wire [WIDTH-1:0] wire_d7_13;
	wire [WIDTH-1:0] wire_d7_14;
	wire [WIDTH-1:0] wire_d7_15;
	wire [WIDTH-1:0] wire_d7_16;
	wire [WIDTH-1:0] wire_d7_17;
	wire [WIDTH-1:0] wire_d7_18;
	wire [WIDTH-1:0] wire_d7_19;
	wire [WIDTH-1:0] wire_d7_20;
	wire [WIDTH-1:0] wire_d7_21;
	wire [WIDTH-1:0] wire_d7_22;
	wire [WIDTH-1:0] wire_d7_23;
	wire [WIDTH-1:0] wire_d7_24;
	wire [WIDTH-1:0] wire_d7_25;
	wire [WIDTH-1:0] wire_d7_26;
	wire [WIDTH-1:0] wire_d7_27;
	wire [WIDTH-1:0] wire_d7_28;
	wire [WIDTH-1:0] wire_d7_29;
	wire [WIDTH-1:0] wire_d7_30;
	wire [WIDTH-1:0] wire_d7_31;
	wire [WIDTH-1:0] wire_d7_32;
	wire [WIDTH-1:0] wire_d7_33;
	wire [WIDTH-1:0] wire_d7_34;
	wire [WIDTH-1:0] wire_d7_35;
	wire [WIDTH-1:0] wire_d7_36;
	wire [WIDTH-1:0] wire_d7_37;
	wire [WIDTH-1:0] wire_d7_38;
	wire [WIDTH-1:0] wire_d7_39;
	wire [WIDTH-1:0] wire_d7_40;
	wire [WIDTH-1:0] wire_d7_41;
	wire [WIDTH-1:0] wire_d7_42;
	wire [WIDTH-1:0] wire_d7_43;
	wire [WIDTH-1:0] wire_d7_44;
	wire [WIDTH-1:0] wire_d7_45;
	wire [WIDTH-1:0] wire_d7_46;
	wire [WIDTH-1:0] wire_d7_47;
	wire [WIDTH-1:0] wire_d7_48;
	wire [WIDTH-1:0] wire_d8_0;
	wire [WIDTH-1:0] wire_d8_1;
	wire [WIDTH-1:0] wire_d8_2;
	wire [WIDTH-1:0] wire_d8_3;
	wire [WIDTH-1:0] wire_d8_4;
	wire [WIDTH-1:0] wire_d8_5;
	wire [WIDTH-1:0] wire_d8_6;
	wire [WIDTH-1:0] wire_d8_7;
	wire [WIDTH-1:0] wire_d8_8;
	wire [WIDTH-1:0] wire_d8_9;
	wire [WIDTH-1:0] wire_d8_10;
	wire [WIDTH-1:0] wire_d8_11;
	wire [WIDTH-1:0] wire_d8_12;
	wire [WIDTH-1:0] wire_d8_13;
	wire [WIDTH-1:0] wire_d8_14;
	wire [WIDTH-1:0] wire_d8_15;
	wire [WIDTH-1:0] wire_d8_16;
	wire [WIDTH-1:0] wire_d8_17;
	wire [WIDTH-1:0] wire_d8_18;
	wire [WIDTH-1:0] wire_d8_19;
	wire [WIDTH-1:0] wire_d8_20;
	wire [WIDTH-1:0] wire_d8_21;
	wire [WIDTH-1:0] wire_d8_22;
	wire [WIDTH-1:0] wire_d8_23;
	wire [WIDTH-1:0] wire_d8_24;
	wire [WIDTH-1:0] wire_d8_25;
	wire [WIDTH-1:0] wire_d8_26;
	wire [WIDTH-1:0] wire_d8_27;
	wire [WIDTH-1:0] wire_d8_28;
	wire [WIDTH-1:0] wire_d8_29;
	wire [WIDTH-1:0] wire_d8_30;
	wire [WIDTH-1:0] wire_d8_31;
	wire [WIDTH-1:0] wire_d8_32;
	wire [WIDTH-1:0] wire_d8_33;
	wire [WIDTH-1:0] wire_d8_34;
	wire [WIDTH-1:0] wire_d8_35;
	wire [WIDTH-1:0] wire_d8_36;
	wire [WIDTH-1:0] wire_d8_37;
	wire [WIDTH-1:0] wire_d8_38;
	wire [WIDTH-1:0] wire_d8_39;
	wire [WIDTH-1:0] wire_d8_40;
	wire [WIDTH-1:0] wire_d8_41;
	wire [WIDTH-1:0] wire_d8_42;
	wire [WIDTH-1:0] wire_d8_43;
	wire [WIDTH-1:0] wire_d8_44;
	wire [WIDTH-1:0] wire_d8_45;
	wire [WIDTH-1:0] wire_d8_46;
	wire [WIDTH-1:0] wire_d8_47;
	wire [WIDTH-1:0] wire_d8_48;
	wire [WIDTH-1:0] wire_d9_0;
	wire [WIDTH-1:0] wire_d9_1;
	wire [WIDTH-1:0] wire_d9_2;
	wire [WIDTH-1:0] wire_d9_3;
	wire [WIDTH-1:0] wire_d9_4;
	wire [WIDTH-1:0] wire_d9_5;
	wire [WIDTH-1:0] wire_d9_6;
	wire [WIDTH-1:0] wire_d9_7;
	wire [WIDTH-1:0] wire_d9_8;
	wire [WIDTH-1:0] wire_d9_9;
	wire [WIDTH-1:0] wire_d9_10;
	wire [WIDTH-1:0] wire_d9_11;
	wire [WIDTH-1:0] wire_d9_12;
	wire [WIDTH-1:0] wire_d9_13;
	wire [WIDTH-1:0] wire_d9_14;
	wire [WIDTH-1:0] wire_d9_15;
	wire [WIDTH-1:0] wire_d9_16;
	wire [WIDTH-1:0] wire_d9_17;
	wire [WIDTH-1:0] wire_d9_18;
	wire [WIDTH-1:0] wire_d9_19;
	wire [WIDTH-1:0] wire_d9_20;
	wire [WIDTH-1:0] wire_d9_21;
	wire [WIDTH-1:0] wire_d9_22;
	wire [WIDTH-1:0] wire_d9_23;
	wire [WIDTH-1:0] wire_d9_24;
	wire [WIDTH-1:0] wire_d9_25;
	wire [WIDTH-1:0] wire_d9_26;
	wire [WIDTH-1:0] wire_d9_27;
	wire [WIDTH-1:0] wire_d9_28;
	wire [WIDTH-1:0] wire_d9_29;
	wire [WIDTH-1:0] wire_d9_30;
	wire [WIDTH-1:0] wire_d9_31;
	wire [WIDTH-1:0] wire_d9_32;
	wire [WIDTH-1:0] wire_d9_33;
	wire [WIDTH-1:0] wire_d9_34;
	wire [WIDTH-1:0] wire_d9_35;
	wire [WIDTH-1:0] wire_d9_36;
	wire [WIDTH-1:0] wire_d9_37;
	wire [WIDTH-1:0] wire_d9_38;
	wire [WIDTH-1:0] wire_d9_39;
	wire [WIDTH-1:0] wire_d9_40;
	wire [WIDTH-1:0] wire_d9_41;
	wire [WIDTH-1:0] wire_d9_42;
	wire [WIDTH-1:0] wire_d9_43;
	wire [WIDTH-1:0] wire_d9_44;
	wire [WIDTH-1:0] wire_d9_45;
	wire [WIDTH-1:0] wire_d9_46;
	wire [WIDTH-1:0] wire_d9_47;
	wire [WIDTH-1:0] wire_d9_48;
	wire [WIDTH-1:0] wire_d10_0;
	wire [WIDTH-1:0] wire_d10_1;
	wire [WIDTH-1:0] wire_d10_2;
	wire [WIDTH-1:0] wire_d10_3;
	wire [WIDTH-1:0] wire_d10_4;
	wire [WIDTH-1:0] wire_d10_5;
	wire [WIDTH-1:0] wire_d10_6;
	wire [WIDTH-1:0] wire_d10_7;
	wire [WIDTH-1:0] wire_d10_8;
	wire [WIDTH-1:0] wire_d10_9;
	wire [WIDTH-1:0] wire_d10_10;
	wire [WIDTH-1:0] wire_d10_11;
	wire [WIDTH-1:0] wire_d10_12;
	wire [WIDTH-1:0] wire_d10_13;
	wire [WIDTH-1:0] wire_d10_14;
	wire [WIDTH-1:0] wire_d10_15;
	wire [WIDTH-1:0] wire_d10_16;
	wire [WIDTH-1:0] wire_d10_17;
	wire [WIDTH-1:0] wire_d10_18;
	wire [WIDTH-1:0] wire_d10_19;
	wire [WIDTH-1:0] wire_d10_20;
	wire [WIDTH-1:0] wire_d10_21;
	wire [WIDTH-1:0] wire_d10_22;
	wire [WIDTH-1:0] wire_d10_23;
	wire [WIDTH-1:0] wire_d10_24;
	wire [WIDTH-1:0] wire_d10_25;
	wire [WIDTH-1:0] wire_d10_26;
	wire [WIDTH-1:0] wire_d10_27;
	wire [WIDTH-1:0] wire_d10_28;
	wire [WIDTH-1:0] wire_d10_29;
	wire [WIDTH-1:0] wire_d10_30;
	wire [WIDTH-1:0] wire_d10_31;
	wire [WIDTH-1:0] wire_d10_32;
	wire [WIDTH-1:0] wire_d10_33;
	wire [WIDTH-1:0] wire_d10_34;
	wire [WIDTH-1:0] wire_d10_35;
	wire [WIDTH-1:0] wire_d10_36;
	wire [WIDTH-1:0] wire_d10_37;
	wire [WIDTH-1:0] wire_d10_38;
	wire [WIDTH-1:0] wire_d10_39;
	wire [WIDTH-1:0] wire_d10_40;
	wire [WIDTH-1:0] wire_d10_41;
	wire [WIDTH-1:0] wire_d10_42;
	wire [WIDTH-1:0] wire_d10_43;
	wire [WIDTH-1:0] wire_d10_44;
	wire [WIDTH-1:0] wire_d10_45;
	wire [WIDTH-1:0] wire_d10_46;
	wire [WIDTH-1:0] wire_d10_47;
	wire [WIDTH-1:0] wire_d10_48;
	wire [WIDTH-1:0] wire_d11_0;
	wire [WIDTH-1:0] wire_d11_1;
	wire [WIDTH-1:0] wire_d11_2;
	wire [WIDTH-1:0] wire_d11_3;
	wire [WIDTH-1:0] wire_d11_4;
	wire [WIDTH-1:0] wire_d11_5;
	wire [WIDTH-1:0] wire_d11_6;
	wire [WIDTH-1:0] wire_d11_7;
	wire [WIDTH-1:0] wire_d11_8;
	wire [WIDTH-1:0] wire_d11_9;
	wire [WIDTH-1:0] wire_d11_10;
	wire [WIDTH-1:0] wire_d11_11;
	wire [WIDTH-1:0] wire_d11_12;
	wire [WIDTH-1:0] wire_d11_13;
	wire [WIDTH-1:0] wire_d11_14;
	wire [WIDTH-1:0] wire_d11_15;
	wire [WIDTH-1:0] wire_d11_16;
	wire [WIDTH-1:0] wire_d11_17;
	wire [WIDTH-1:0] wire_d11_18;
	wire [WIDTH-1:0] wire_d11_19;
	wire [WIDTH-1:0] wire_d11_20;
	wire [WIDTH-1:0] wire_d11_21;
	wire [WIDTH-1:0] wire_d11_22;
	wire [WIDTH-1:0] wire_d11_23;
	wire [WIDTH-1:0] wire_d11_24;
	wire [WIDTH-1:0] wire_d11_25;
	wire [WIDTH-1:0] wire_d11_26;
	wire [WIDTH-1:0] wire_d11_27;
	wire [WIDTH-1:0] wire_d11_28;
	wire [WIDTH-1:0] wire_d11_29;
	wire [WIDTH-1:0] wire_d11_30;
	wire [WIDTH-1:0] wire_d11_31;
	wire [WIDTH-1:0] wire_d11_32;
	wire [WIDTH-1:0] wire_d11_33;
	wire [WIDTH-1:0] wire_d11_34;
	wire [WIDTH-1:0] wire_d11_35;
	wire [WIDTH-1:0] wire_d11_36;
	wire [WIDTH-1:0] wire_d11_37;
	wire [WIDTH-1:0] wire_d11_38;
	wire [WIDTH-1:0] wire_d11_39;
	wire [WIDTH-1:0] wire_d11_40;
	wire [WIDTH-1:0] wire_d11_41;
	wire [WIDTH-1:0] wire_d11_42;
	wire [WIDTH-1:0] wire_d11_43;
	wire [WIDTH-1:0] wire_d11_44;
	wire [WIDTH-1:0] wire_d11_45;
	wire [WIDTH-1:0] wire_d11_46;
	wire [WIDTH-1:0] wire_d11_47;
	wire [WIDTH-1:0] wire_d11_48;
	wire [WIDTH-1:0] wire_d12_0;
	wire [WIDTH-1:0] wire_d12_1;
	wire [WIDTH-1:0] wire_d12_2;
	wire [WIDTH-1:0] wire_d12_3;
	wire [WIDTH-1:0] wire_d12_4;
	wire [WIDTH-1:0] wire_d12_5;
	wire [WIDTH-1:0] wire_d12_6;
	wire [WIDTH-1:0] wire_d12_7;
	wire [WIDTH-1:0] wire_d12_8;
	wire [WIDTH-1:0] wire_d12_9;
	wire [WIDTH-1:0] wire_d12_10;
	wire [WIDTH-1:0] wire_d12_11;
	wire [WIDTH-1:0] wire_d12_12;
	wire [WIDTH-1:0] wire_d12_13;
	wire [WIDTH-1:0] wire_d12_14;
	wire [WIDTH-1:0] wire_d12_15;
	wire [WIDTH-1:0] wire_d12_16;
	wire [WIDTH-1:0] wire_d12_17;
	wire [WIDTH-1:0] wire_d12_18;
	wire [WIDTH-1:0] wire_d12_19;
	wire [WIDTH-1:0] wire_d12_20;
	wire [WIDTH-1:0] wire_d12_21;
	wire [WIDTH-1:0] wire_d12_22;
	wire [WIDTH-1:0] wire_d12_23;
	wire [WIDTH-1:0] wire_d12_24;
	wire [WIDTH-1:0] wire_d12_25;
	wire [WIDTH-1:0] wire_d12_26;
	wire [WIDTH-1:0] wire_d12_27;
	wire [WIDTH-1:0] wire_d12_28;
	wire [WIDTH-1:0] wire_d12_29;
	wire [WIDTH-1:0] wire_d12_30;
	wire [WIDTH-1:0] wire_d12_31;
	wire [WIDTH-1:0] wire_d12_32;
	wire [WIDTH-1:0] wire_d12_33;
	wire [WIDTH-1:0] wire_d12_34;
	wire [WIDTH-1:0] wire_d12_35;
	wire [WIDTH-1:0] wire_d12_36;
	wire [WIDTH-1:0] wire_d12_37;
	wire [WIDTH-1:0] wire_d12_38;
	wire [WIDTH-1:0] wire_d12_39;
	wire [WIDTH-1:0] wire_d12_40;
	wire [WIDTH-1:0] wire_d12_41;
	wire [WIDTH-1:0] wire_d12_42;
	wire [WIDTH-1:0] wire_d12_43;
	wire [WIDTH-1:0] wire_d12_44;
	wire [WIDTH-1:0] wire_d12_45;
	wire [WIDTH-1:0] wire_d12_46;
	wire [WIDTH-1:0] wire_d12_47;
	wire [WIDTH-1:0] wire_d12_48;
	wire [WIDTH-1:0] wire_d13_0;
	wire [WIDTH-1:0] wire_d13_1;
	wire [WIDTH-1:0] wire_d13_2;
	wire [WIDTH-1:0] wire_d13_3;
	wire [WIDTH-1:0] wire_d13_4;
	wire [WIDTH-1:0] wire_d13_5;
	wire [WIDTH-1:0] wire_d13_6;
	wire [WIDTH-1:0] wire_d13_7;
	wire [WIDTH-1:0] wire_d13_8;
	wire [WIDTH-1:0] wire_d13_9;
	wire [WIDTH-1:0] wire_d13_10;
	wire [WIDTH-1:0] wire_d13_11;
	wire [WIDTH-1:0] wire_d13_12;
	wire [WIDTH-1:0] wire_d13_13;
	wire [WIDTH-1:0] wire_d13_14;
	wire [WIDTH-1:0] wire_d13_15;
	wire [WIDTH-1:0] wire_d13_16;
	wire [WIDTH-1:0] wire_d13_17;
	wire [WIDTH-1:0] wire_d13_18;
	wire [WIDTH-1:0] wire_d13_19;
	wire [WIDTH-1:0] wire_d13_20;
	wire [WIDTH-1:0] wire_d13_21;
	wire [WIDTH-1:0] wire_d13_22;
	wire [WIDTH-1:0] wire_d13_23;
	wire [WIDTH-1:0] wire_d13_24;
	wire [WIDTH-1:0] wire_d13_25;
	wire [WIDTH-1:0] wire_d13_26;
	wire [WIDTH-1:0] wire_d13_27;
	wire [WIDTH-1:0] wire_d13_28;
	wire [WIDTH-1:0] wire_d13_29;
	wire [WIDTH-1:0] wire_d13_30;
	wire [WIDTH-1:0] wire_d13_31;
	wire [WIDTH-1:0] wire_d13_32;
	wire [WIDTH-1:0] wire_d13_33;
	wire [WIDTH-1:0] wire_d13_34;
	wire [WIDTH-1:0] wire_d13_35;
	wire [WIDTH-1:0] wire_d13_36;
	wire [WIDTH-1:0] wire_d13_37;
	wire [WIDTH-1:0] wire_d13_38;
	wire [WIDTH-1:0] wire_d13_39;
	wire [WIDTH-1:0] wire_d13_40;
	wire [WIDTH-1:0] wire_d13_41;
	wire [WIDTH-1:0] wire_d13_42;
	wire [WIDTH-1:0] wire_d13_43;
	wire [WIDTH-1:0] wire_d13_44;
	wire [WIDTH-1:0] wire_d13_45;
	wire [WIDTH-1:0] wire_d13_46;
	wire [WIDTH-1:0] wire_d13_47;
	wire [WIDTH-1:0] wire_d13_48;
	wire [WIDTH-1:0] wire_d14_0;
	wire [WIDTH-1:0] wire_d14_1;
	wire [WIDTH-1:0] wire_d14_2;
	wire [WIDTH-1:0] wire_d14_3;
	wire [WIDTH-1:0] wire_d14_4;
	wire [WIDTH-1:0] wire_d14_5;
	wire [WIDTH-1:0] wire_d14_6;
	wire [WIDTH-1:0] wire_d14_7;
	wire [WIDTH-1:0] wire_d14_8;
	wire [WIDTH-1:0] wire_d14_9;
	wire [WIDTH-1:0] wire_d14_10;
	wire [WIDTH-1:0] wire_d14_11;
	wire [WIDTH-1:0] wire_d14_12;
	wire [WIDTH-1:0] wire_d14_13;
	wire [WIDTH-1:0] wire_d14_14;
	wire [WIDTH-1:0] wire_d14_15;
	wire [WIDTH-1:0] wire_d14_16;
	wire [WIDTH-1:0] wire_d14_17;
	wire [WIDTH-1:0] wire_d14_18;
	wire [WIDTH-1:0] wire_d14_19;
	wire [WIDTH-1:0] wire_d14_20;
	wire [WIDTH-1:0] wire_d14_21;
	wire [WIDTH-1:0] wire_d14_22;
	wire [WIDTH-1:0] wire_d14_23;
	wire [WIDTH-1:0] wire_d14_24;
	wire [WIDTH-1:0] wire_d14_25;
	wire [WIDTH-1:0] wire_d14_26;
	wire [WIDTH-1:0] wire_d14_27;
	wire [WIDTH-1:0] wire_d14_28;
	wire [WIDTH-1:0] wire_d14_29;
	wire [WIDTH-1:0] wire_d14_30;
	wire [WIDTH-1:0] wire_d14_31;
	wire [WIDTH-1:0] wire_d14_32;
	wire [WIDTH-1:0] wire_d14_33;
	wire [WIDTH-1:0] wire_d14_34;
	wire [WIDTH-1:0] wire_d14_35;
	wire [WIDTH-1:0] wire_d14_36;
	wire [WIDTH-1:0] wire_d14_37;
	wire [WIDTH-1:0] wire_d14_38;
	wire [WIDTH-1:0] wire_d14_39;
	wire [WIDTH-1:0] wire_d14_40;
	wire [WIDTH-1:0] wire_d14_41;
	wire [WIDTH-1:0] wire_d14_42;
	wire [WIDTH-1:0] wire_d14_43;
	wire [WIDTH-1:0] wire_d14_44;
	wire [WIDTH-1:0] wire_d14_45;
	wire [WIDTH-1:0] wire_d14_46;
	wire [WIDTH-1:0] wire_d14_47;
	wire [WIDTH-1:0] wire_d14_48;
	wire [WIDTH-1:0] wire_d15_0;
	wire [WIDTH-1:0] wire_d15_1;
	wire [WIDTH-1:0] wire_d15_2;
	wire [WIDTH-1:0] wire_d15_3;
	wire [WIDTH-1:0] wire_d15_4;
	wire [WIDTH-1:0] wire_d15_5;
	wire [WIDTH-1:0] wire_d15_6;
	wire [WIDTH-1:0] wire_d15_7;
	wire [WIDTH-1:0] wire_d15_8;
	wire [WIDTH-1:0] wire_d15_9;
	wire [WIDTH-1:0] wire_d15_10;
	wire [WIDTH-1:0] wire_d15_11;
	wire [WIDTH-1:0] wire_d15_12;
	wire [WIDTH-1:0] wire_d15_13;
	wire [WIDTH-1:0] wire_d15_14;
	wire [WIDTH-1:0] wire_d15_15;
	wire [WIDTH-1:0] wire_d15_16;
	wire [WIDTH-1:0] wire_d15_17;
	wire [WIDTH-1:0] wire_d15_18;
	wire [WIDTH-1:0] wire_d15_19;
	wire [WIDTH-1:0] wire_d15_20;
	wire [WIDTH-1:0] wire_d15_21;
	wire [WIDTH-1:0] wire_d15_22;
	wire [WIDTH-1:0] wire_d15_23;
	wire [WIDTH-1:0] wire_d15_24;
	wire [WIDTH-1:0] wire_d15_25;
	wire [WIDTH-1:0] wire_d15_26;
	wire [WIDTH-1:0] wire_d15_27;
	wire [WIDTH-1:0] wire_d15_28;
	wire [WIDTH-1:0] wire_d15_29;
	wire [WIDTH-1:0] wire_d15_30;
	wire [WIDTH-1:0] wire_d15_31;
	wire [WIDTH-1:0] wire_d15_32;
	wire [WIDTH-1:0] wire_d15_33;
	wire [WIDTH-1:0] wire_d15_34;
	wire [WIDTH-1:0] wire_d15_35;
	wire [WIDTH-1:0] wire_d15_36;
	wire [WIDTH-1:0] wire_d15_37;
	wire [WIDTH-1:0] wire_d15_38;
	wire [WIDTH-1:0] wire_d15_39;
	wire [WIDTH-1:0] wire_d15_40;
	wire [WIDTH-1:0] wire_d15_41;
	wire [WIDTH-1:0] wire_d15_42;
	wire [WIDTH-1:0] wire_d15_43;
	wire [WIDTH-1:0] wire_d15_44;
	wire [WIDTH-1:0] wire_d15_45;
	wire [WIDTH-1:0] wire_d15_46;
	wire [WIDTH-1:0] wire_d15_47;
	wire [WIDTH-1:0] wire_d15_48;
	wire [WIDTH-1:0] wire_d16_0;
	wire [WIDTH-1:0] wire_d16_1;
	wire [WIDTH-1:0] wire_d16_2;
	wire [WIDTH-1:0] wire_d16_3;
	wire [WIDTH-1:0] wire_d16_4;
	wire [WIDTH-1:0] wire_d16_5;
	wire [WIDTH-1:0] wire_d16_6;
	wire [WIDTH-1:0] wire_d16_7;
	wire [WIDTH-1:0] wire_d16_8;
	wire [WIDTH-1:0] wire_d16_9;
	wire [WIDTH-1:0] wire_d16_10;
	wire [WIDTH-1:0] wire_d16_11;
	wire [WIDTH-1:0] wire_d16_12;
	wire [WIDTH-1:0] wire_d16_13;
	wire [WIDTH-1:0] wire_d16_14;
	wire [WIDTH-1:0] wire_d16_15;
	wire [WIDTH-1:0] wire_d16_16;
	wire [WIDTH-1:0] wire_d16_17;
	wire [WIDTH-1:0] wire_d16_18;
	wire [WIDTH-1:0] wire_d16_19;
	wire [WIDTH-1:0] wire_d16_20;
	wire [WIDTH-1:0] wire_d16_21;
	wire [WIDTH-1:0] wire_d16_22;
	wire [WIDTH-1:0] wire_d16_23;
	wire [WIDTH-1:0] wire_d16_24;
	wire [WIDTH-1:0] wire_d16_25;
	wire [WIDTH-1:0] wire_d16_26;
	wire [WIDTH-1:0] wire_d16_27;
	wire [WIDTH-1:0] wire_d16_28;
	wire [WIDTH-1:0] wire_d16_29;
	wire [WIDTH-1:0] wire_d16_30;
	wire [WIDTH-1:0] wire_d16_31;
	wire [WIDTH-1:0] wire_d16_32;
	wire [WIDTH-1:0] wire_d16_33;
	wire [WIDTH-1:0] wire_d16_34;
	wire [WIDTH-1:0] wire_d16_35;
	wire [WIDTH-1:0] wire_d16_36;
	wire [WIDTH-1:0] wire_d16_37;
	wire [WIDTH-1:0] wire_d16_38;
	wire [WIDTH-1:0] wire_d16_39;
	wire [WIDTH-1:0] wire_d16_40;
	wire [WIDTH-1:0] wire_d16_41;
	wire [WIDTH-1:0] wire_d16_42;
	wire [WIDTH-1:0] wire_d16_43;
	wire [WIDTH-1:0] wire_d16_44;
	wire [WIDTH-1:0] wire_d16_45;
	wire [WIDTH-1:0] wire_d16_46;
	wire [WIDTH-1:0] wire_d16_47;
	wire [WIDTH-1:0] wire_d16_48;
	wire [WIDTH-1:0] wire_d17_0;
	wire [WIDTH-1:0] wire_d17_1;
	wire [WIDTH-1:0] wire_d17_2;
	wire [WIDTH-1:0] wire_d17_3;
	wire [WIDTH-1:0] wire_d17_4;
	wire [WIDTH-1:0] wire_d17_5;
	wire [WIDTH-1:0] wire_d17_6;
	wire [WIDTH-1:0] wire_d17_7;
	wire [WIDTH-1:0] wire_d17_8;
	wire [WIDTH-1:0] wire_d17_9;
	wire [WIDTH-1:0] wire_d17_10;
	wire [WIDTH-1:0] wire_d17_11;
	wire [WIDTH-1:0] wire_d17_12;
	wire [WIDTH-1:0] wire_d17_13;
	wire [WIDTH-1:0] wire_d17_14;
	wire [WIDTH-1:0] wire_d17_15;
	wire [WIDTH-1:0] wire_d17_16;
	wire [WIDTH-1:0] wire_d17_17;
	wire [WIDTH-1:0] wire_d17_18;
	wire [WIDTH-1:0] wire_d17_19;
	wire [WIDTH-1:0] wire_d17_20;
	wire [WIDTH-1:0] wire_d17_21;
	wire [WIDTH-1:0] wire_d17_22;
	wire [WIDTH-1:0] wire_d17_23;
	wire [WIDTH-1:0] wire_d17_24;
	wire [WIDTH-1:0] wire_d17_25;
	wire [WIDTH-1:0] wire_d17_26;
	wire [WIDTH-1:0] wire_d17_27;
	wire [WIDTH-1:0] wire_d17_28;
	wire [WIDTH-1:0] wire_d17_29;
	wire [WIDTH-1:0] wire_d17_30;
	wire [WIDTH-1:0] wire_d17_31;
	wire [WIDTH-1:0] wire_d17_32;
	wire [WIDTH-1:0] wire_d17_33;
	wire [WIDTH-1:0] wire_d17_34;
	wire [WIDTH-1:0] wire_d17_35;
	wire [WIDTH-1:0] wire_d17_36;
	wire [WIDTH-1:0] wire_d17_37;
	wire [WIDTH-1:0] wire_d17_38;
	wire [WIDTH-1:0] wire_d17_39;
	wire [WIDTH-1:0] wire_d17_40;
	wire [WIDTH-1:0] wire_d17_41;
	wire [WIDTH-1:0] wire_d17_42;
	wire [WIDTH-1:0] wire_d17_43;
	wire [WIDTH-1:0] wire_d17_44;
	wire [WIDTH-1:0] wire_d17_45;
	wire [WIDTH-1:0] wire_d17_46;
	wire [WIDTH-1:0] wire_d17_47;
	wire [WIDTH-1:0] wire_d17_48;
	wire [WIDTH-1:0] wire_d18_0;
	wire [WIDTH-1:0] wire_d18_1;
	wire [WIDTH-1:0] wire_d18_2;
	wire [WIDTH-1:0] wire_d18_3;
	wire [WIDTH-1:0] wire_d18_4;
	wire [WIDTH-1:0] wire_d18_5;
	wire [WIDTH-1:0] wire_d18_6;
	wire [WIDTH-1:0] wire_d18_7;
	wire [WIDTH-1:0] wire_d18_8;
	wire [WIDTH-1:0] wire_d18_9;
	wire [WIDTH-1:0] wire_d18_10;
	wire [WIDTH-1:0] wire_d18_11;
	wire [WIDTH-1:0] wire_d18_12;
	wire [WIDTH-1:0] wire_d18_13;
	wire [WIDTH-1:0] wire_d18_14;
	wire [WIDTH-1:0] wire_d18_15;
	wire [WIDTH-1:0] wire_d18_16;
	wire [WIDTH-1:0] wire_d18_17;
	wire [WIDTH-1:0] wire_d18_18;
	wire [WIDTH-1:0] wire_d18_19;
	wire [WIDTH-1:0] wire_d18_20;
	wire [WIDTH-1:0] wire_d18_21;
	wire [WIDTH-1:0] wire_d18_22;
	wire [WIDTH-1:0] wire_d18_23;
	wire [WIDTH-1:0] wire_d18_24;
	wire [WIDTH-1:0] wire_d18_25;
	wire [WIDTH-1:0] wire_d18_26;
	wire [WIDTH-1:0] wire_d18_27;
	wire [WIDTH-1:0] wire_d18_28;
	wire [WIDTH-1:0] wire_d18_29;
	wire [WIDTH-1:0] wire_d18_30;
	wire [WIDTH-1:0] wire_d18_31;
	wire [WIDTH-1:0] wire_d18_32;
	wire [WIDTH-1:0] wire_d18_33;
	wire [WIDTH-1:0] wire_d18_34;
	wire [WIDTH-1:0] wire_d18_35;
	wire [WIDTH-1:0] wire_d18_36;
	wire [WIDTH-1:0] wire_d18_37;
	wire [WIDTH-1:0] wire_d18_38;
	wire [WIDTH-1:0] wire_d18_39;
	wire [WIDTH-1:0] wire_d18_40;
	wire [WIDTH-1:0] wire_d18_41;
	wire [WIDTH-1:0] wire_d18_42;
	wire [WIDTH-1:0] wire_d18_43;
	wire [WIDTH-1:0] wire_d18_44;
	wire [WIDTH-1:0] wire_d18_45;
	wire [WIDTH-1:0] wire_d18_46;
	wire [WIDTH-1:0] wire_d18_47;
	wire [WIDTH-1:0] wire_d18_48;
	wire [WIDTH-1:0] wire_d19_0;
	wire [WIDTH-1:0] wire_d19_1;
	wire [WIDTH-1:0] wire_d19_2;
	wire [WIDTH-1:0] wire_d19_3;
	wire [WIDTH-1:0] wire_d19_4;
	wire [WIDTH-1:0] wire_d19_5;
	wire [WIDTH-1:0] wire_d19_6;
	wire [WIDTH-1:0] wire_d19_7;
	wire [WIDTH-1:0] wire_d19_8;
	wire [WIDTH-1:0] wire_d19_9;
	wire [WIDTH-1:0] wire_d19_10;
	wire [WIDTH-1:0] wire_d19_11;
	wire [WIDTH-1:0] wire_d19_12;
	wire [WIDTH-1:0] wire_d19_13;
	wire [WIDTH-1:0] wire_d19_14;
	wire [WIDTH-1:0] wire_d19_15;
	wire [WIDTH-1:0] wire_d19_16;
	wire [WIDTH-1:0] wire_d19_17;
	wire [WIDTH-1:0] wire_d19_18;
	wire [WIDTH-1:0] wire_d19_19;
	wire [WIDTH-1:0] wire_d19_20;
	wire [WIDTH-1:0] wire_d19_21;
	wire [WIDTH-1:0] wire_d19_22;
	wire [WIDTH-1:0] wire_d19_23;
	wire [WIDTH-1:0] wire_d19_24;
	wire [WIDTH-1:0] wire_d19_25;
	wire [WIDTH-1:0] wire_d19_26;
	wire [WIDTH-1:0] wire_d19_27;
	wire [WIDTH-1:0] wire_d19_28;
	wire [WIDTH-1:0] wire_d19_29;
	wire [WIDTH-1:0] wire_d19_30;
	wire [WIDTH-1:0] wire_d19_31;
	wire [WIDTH-1:0] wire_d19_32;
	wire [WIDTH-1:0] wire_d19_33;
	wire [WIDTH-1:0] wire_d19_34;
	wire [WIDTH-1:0] wire_d19_35;
	wire [WIDTH-1:0] wire_d19_36;
	wire [WIDTH-1:0] wire_d19_37;
	wire [WIDTH-1:0] wire_d19_38;
	wire [WIDTH-1:0] wire_d19_39;
	wire [WIDTH-1:0] wire_d19_40;
	wire [WIDTH-1:0] wire_d19_41;
	wire [WIDTH-1:0] wire_d19_42;
	wire [WIDTH-1:0] wire_d19_43;
	wire [WIDTH-1:0] wire_d19_44;
	wire [WIDTH-1:0] wire_d19_45;
	wire [WIDTH-1:0] wire_d19_46;
	wire [WIDTH-1:0] wire_d19_47;
	wire [WIDTH-1:0] wire_d19_48;
	wire [WIDTH-1:0] wire_d20_0;
	wire [WIDTH-1:0] wire_d20_1;
	wire [WIDTH-1:0] wire_d20_2;
	wire [WIDTH-1:0] wire_d20_3;
	wire [WIDTH-1:0] wire_d20_4;
	wire [WIDTH-1:0] wire_d20_5;
	wire [WIDTH-1:0] wire_d20_6;
	wire [WIDTH-1:0] wire_d20_7;
	wire [WIDTH-1:0] wire_d20_8;
	wire [WIDTH-1:0] wire_d20_9;
	wire [WIDTH-1:0] wire_d20_10;
	wire [WIDTH-1:0] wire_d20_11;
	wire [WIDTH-1:0] wire_d20_12;
	wire [WIDTH-1:0] wire_d20_13;
	wire [WIDTH-1:0] wire_d20_14;
	wire [WIDTH-1:0] wire_d20_15;
	wire [WIDTH-1:0] wire_d20_16;
	wire [WIDTH-1:0] wire_d20_17;
	wire [WIDTH-1:0] wire_d20_18;
	wire [WIDTH-1:0] wire_d20_19;
	wire [WIDTH-1:0] wire_d20_20;
	wire [WIDTH-1:0] wire_d20_21;
	wire [WIDTH-1:0] wire_d20_22;
	wire [WIDTH-1:0] wire_d20_23;
	wire [WIDTH-1:0] wire_d20_24;
	wire [WIDTH-1:0] wire_d20_25;
	wire [WIDTH-1:0] wire_d20_26;
	wire [WIDTH-1:0] wire_d20_27;
	wire [WIDTH-1:0] wire_d20_28;
	wire [WIDTH-1:0] wire_d20_29;
	wire [WIDTH-1:0] wire_d20_30;
	wire [WIDTH-1:0] wire_d20_31;
	wire [WIDTH-1:0] wire_d20_32;
	wire [WIDTH-1:0] wire_d20_33;
	wire [WIDTH-1:0] wire_d20_34;
	wire [WIDTH-1:0] wire_d20_35;
	wire [WIDTH-1:0] wire_d20_36;
	wire [WIDTH-1:0] wire_d20_37;
	wire [WIDTH-1:0] wire_d20_38;
	wire [WIDTH-1:0] wire_d20_39;
	wire [WIDTH-1:0] wire_d20_40;
	wire [WIDTH-1:0] wire_d20_41;
	wire [WIDTH-1:0] wire_d20_42;
	wire [WIDTH-1:0] wire_d20_43;
	wire [WIDTH-1:0] wire_d20_44;
	wire [WIDTH-1:0] wire_d20_45;
	wire [WIDTH-1:0] wire_d20_46;
	wire [WIDTH-1:0] wire_d20_47;
	wire [WIDTH-1:0] wire_d20_48;
	wire [WIDTH-1:0] wire_d21_0;
	wire [WIDTH-1:0] wire_d21_1;
	wire [WIDTH-1:0] wire_d21_2;
	wire [WIDTH-1:0] wire_d21_3;
	wire [WIDTH-1:0] wire_d21_4;
	wire [WIDTH-1:0] wire_d21_5;
	wire [WIDTH-1:0] wire_d21_6;
	wire [WIDTH-1:0] wire_d21_7;
	wire [WIDTH-1:0] wire_d21_8;
	wire [WIDTH-1:0] wire_d21_9;
	wire [WIDTH-1:0] wire_d21_10;
	wire [WIDTH-1:0] wire_d21_11;
	wire [WIDTH-1:0] wire_d21_12;
	wire [WIDTH-1:0] wire_d21_13;
	wire [WIDTH-1:0] wire_d21_14;
	wire [WIDTH-1:0] wire_d21_15;
	wire [WIDTH-1:0] wire_d21_16;
	wire [WIDTH-1:0] wire_d21_17;
	wire [WIDTH-1:0] wire_d21_18;
	wire [WIDTH-1:0] wire_d21_19;
	wire [WIDTH-1:0] wire_d21_20;
	wire [WIDTH-1:0] wire_d21_21;
	wire [WIDTH-1:0] wire_d21_22;
	wire [WIDTH-1:0] wire_d21_23;
	wire [WIDTH-1:0] wire_d21_24;
	wire [WIDTH-1:0] wire_d21_25;
	wire [WIDTH-1:0] wire_d21_26;
	wire [WIDTH-1:0] wire_d21_27;
	wire [WIDTH-1:0] wire_d21_28;
	wire [WIDTH-1:0] wire_d21_29;
	wire [WIDTH-1:0] wire_d21_30;
	wire [WIDTH-1:0] wire_d21_31;
	wire [WIDTH-1:0] wire_d21_32;
	wire [WIDTH-1:0] wire_d21_33;
	wire [WIDTH-1:0] wire_d21_34;
	wire [WIDTH-1:0] wire_d21_35;
	wire [WIDTH-1:0] wire_d21_36;
	wire [WIDTH-1:0] wire_d21_37;
	wire [WIDTH-1:0] wire_d21_38;
	wire [WIDTH-1:0] wire_d21_39;
	wire [WIDTH-1:0] wire_d21_40;
	wire [WIDTH-1:0] wire_d21_41;
	wire [WIDTH-1:0] wire_d21_42;
	wire [WIDTH-1:0] wire_d21_43;
	wire [WIDTH-1:0] wire_d21_44;
	wire [WIDTH-1:0] wire_d21_45;
	wire [WIDTH-1:0] wire_d21_46;
	wire [WIDTH-1:0] wire_d21_47;
	wire [WIDTH-1:0] wire_d21_48;
	wire [WIDTH-1:0] wire_d22_0;
	wire [WIDTH-1:0] wire_d22_1;
	wire [WIDTH-1:0] wire_d22_2;
	wire [WIDTH-1:0] wire_d22_3;
	wire [WIDTH-1:0] wire_d22_4;
	wire [WIDTH-1:0] wire_d22_5;
	wire [WIDTH-1:0] wire_d22_6;
	wire [WIDTH-1:0] wire_d22_7;
	wire [WIDTH-1:0] wire_d22_8;
	wire [WIDTH-1:0] wire_d22_9;
	wire [WIDTH-1:0] wire_d22_10;
	wire [WIDTH-1:0] wire_d22_11;
	wire [WIDTH-1:0] wire_d22_12;
	wire [WIDTH-1:0] wire_d22_13;
	wire [WIDTH-1:0] wire_d22_14;
	wire [WIDTH-1:0] wire_d22_15;
	wire [WIDTH-1:0] wire_d22_16;
	wire [WIDTH-1:0] wire_d22_17;
	wire [WIDTH-1:0] wire_d22_18;
	wire [WIDTH-1:0] wire_d22_19;
	wire [WIDTH-1:0] wire_d22_20;
	wire [WIDTH-1:0] wire_d22_21;
	wire [WIDTH-1:0] wire_d22_22;
	wire [WIDTH-1:0] wire_d22_23;
	wire [WIDTH-1:0] wire_d22_24;
	wire [WIDTH-1:0] wire_d22_25;
	wire [WIDTH-1:0] wire_d22_26;
	wire [WIDTH-1:0] wire_d22_27;
	wire [WIDTH-1:0] wire_d22_28;
	wire [WIDTH-1:0] wire_d22_29;
	wire [WIDTH-1:0] wire_d22_30;
	wire [WIDTH-1:0] wire_d22_31;
	wire [WIDTH-1:0] wire_d22_32;
	wire [WIDTH-1:0] wire_d22_33;
	wire [WIDTH-1:0] wire_d22_34;
	wire [WIDTH-1:0] wire_d22_35;
	wire [WIDTH-1:0] wire_d22_36;
	wire [WIDTH-1:0] wire_d22_37;
	wire [WIDTH-1:0] wire_d22_38;
	wire [WIDTH-1:0] wire_d22_39;
	wire [WIDTH-1:0] wire_d22_40;
	wire [WIDTH-1:0] wire_d22_41;
	wire [WIDTH-1:0] wire_d22_42;
	wire [WIDTH-1:0] wire_d22_43;
	wire [WIDTH-1:0] wire_d22_44;
	wire [WIDTH-1:0] wire_d22_45;
	wire [WIDTH-1:0] wire_d22_46;
	wire [WIDTH-1:0] wire_d22_47;
	wire [WIDTH-1:0] wire_d22_48;
	wire [WIDTH-1:0] wire_d23_0;
	wire [WIDTH-1:0] wire_d23_1;
	wire [WIDTH-1:0] wire_d23_2;
	wire [WIDTH-1:0] wire_d23_3;
	wire [WIDTH-1:0] wire_d23_4;
	wire [WIDTH-1:0] wire_d23_5;
	wire [WIDTH-1:0] wire_d23_6;
	wire [WIDTH-1:0] wire_d23_7;
	wire [WIDTH-1:0] wire_d23_8;
	wire [WIDTH-1:0] wire_d23_9;
	wire [WIDTH-1:0] wire_d23_10;
	wire [WIDTH-1:0] wire_d23_11;
	wire [WIDTH-1:0] wire_d23_12;
	wire [WIDTH-1:0] wire_d23_13;
	wire [WIDTH-1:0] wire_d23_14;
	wire [WIDTH-1:0] wire_d23_15;
	wire [WIDTH-1:0] wire_d23_16;
	wire [WIDTH-1:0] wire_d23_17;
	wire [WIDTH-1:0] wire_d23_18;
	wire [WIDTH-1:0] wire_d23_19;
	wire [WIDTH-1:0] wire_d23_20;
	wire [WIDTH-1:0] wire_d23_21;
	wire [WIDTH-1:0] wire_d23_22;
	wire [WIDTH-1:0] wire_d23_23;
	wire [WIDTH-1:0] wire_d23_24;
	wire [WIDTH-1:0] wire_d23_25;
	wire [WIDTH-1:0] wire_d23_26;
	wire [WIDTH-1:0] wire_d23_27;
	wire [WIDTH-1:0] wire_d23_28;
	wire [WIDTH-1:0] wire_d23_29;
	wire [WIDTH-1:0] wire_d23_30;
	wire [WIDTH-1:0] wire_d23_31;
	wire [WIDTH-1:0] wire_d23_32;
	wire [WIDTH-1:0] wire_d23_33;
	wire [WIDTH-1:0] wire_d23_34;
	wire [WIDTH-1:0] wire_d23_35;
	wire [WIDTH-1:0] wire_d23_36;
	wire [WIDTH-1:0] wire_d23_37;
	wire [WIDTH-1:0] wire_d23_38;
	wire [WIDTH-1:0] wire_d23_39;
	wire [WIDTH-1:0] wire_d23_40;
	wire [WIDTH-1:0] wire_d23_41;
	wire [WIDTH-1:0] wire_d23_42;
	wire [WIDTH-1:0] wire_d23_43;
	wire [WIDTH-1:0] wire_d23_44;
	wire [WIDTH-1:0] wire_d23_45;
	wire [WIDTH-1:0] wire_d23_46;
	wire [WIDTH-1:0] wire_d23_47;
	wire [WIDTH-1:0] wire_d23_48;
	wire [WIDTH-1:0] wire_d24_0;
	wire [WIDTH-1:0] wire_d24_1;
	wire [WIDTH-1:0] wire_d24_2;
	wire [WIDTH-1:0] wire_d24_3;
	wire [WIDTH-1:0] wire_d24_4;
	wire [WIDTH-1:0] wire_d24_5;
	wire [WIDTH-1:0] wire_d24_6;
	wire [WIDTH-1:0] wire_d24_7;
	wire [WIDTH-1:0] wire_d24_8;
	wire [WIDTH-1:0] wire_d24_9;
	wire [WIDTH-1:0] wire_d24_10;
	wire [WIDTH-1:0] wire_d24_11;
	wire [WIDTH-1:0] wire_d24_12;
	wire [WIDTH-1:0] wire_d24_13;
	wire [WIDTH-1:0] wire_d24_14;
	wire [WIDTH-1:0] wire_d24_15;
	wire [WIDTH-1:0] wire_d24_16;
	wire [WIDTH-1:0] wire_d24_17;
	wire [WIDTH-1:0] wire_d24_18;
	wire [WIDTH-1:0] wire_d24_19;
	wire [WIDTH-1:0] wire_d24_20;
	wire [WIDTH-1:0] wire_d24_21;
	wire [WIDTH-1:0] wire_d24_22;
	wire [WIDTH-1:0] wire_d24_23;
	wire [WIDTH-1:0] wire_d24_24;
	wire [WIDTH-1:0] wire_d24_25;
	wire [WIDTH-1:0] wire_d24_26;
	wire [WIDTH-1:0] wire_d24_27;
	wire [WIDTH-1:0] wire_d24_28;
	wire [WIDTH-1:0] wire_d24_29;
	wire [WIDTH-1:0] wire_d24_30;
	wire [WIDTH-1:0] wire_d24_31;
	wire [WIDTH-1:0] wire_d24_32;
	wire [WIDTH-1:0] wire_d24_33;
	wire [WIDTH-1:0] wire_d24_34;
	wire [WIDTH-1:0] wire_d24_35;
	wire [WIDTH-1:0] wire_d24_36;
	wire [WIDTH-1:0] wire_d24_37;
	wire [WIDTH-1:0] wire_d24_38;
	wire [WIDTH-1:0] wire_d24_39;
	wire [WIDTH-1:0] wire_d24_40;
	wire [WIDTH-1:0] wire_d24_41;
	wire [WIDTH-1:0] wire_d24_42;
	wire [WIDTH-1:0] wire_d24_43;
	wire [WIDTH-1:0] wire_d24_44;
	wire [WIDTH-1:0] wire_d24_45;
	wire [WIDTH-1:0] wire_d24_46;
	wire [WIDTH-1:0] wire_d24_47;
	wire [WIDTH-1:0] wire_d24_48;
	wire [WIDTH-1:0] wire_d25_0;
	wire [WIDTH-1:0] wire_d25_1;
	wire [WIDTH-1:0] wire_d25_2;
	wire [WIDTH-1:0] wire_d25_3;
	wire [WIDTH-1:0] wire_d25_4;
	wire [WIDTH-1:0] wire_d25_5;
	wire [WIDTH-1:0] wire_d25_6;
	wire [WIDTH-1:0] wire_d25_7;
	wire [WIDTH-1:0] wire_d25_8;
	wire [WIDTH-1:0] wire_d25_9;
	wire [WIDTH-1:0] wire_d25_10;
	wire [WIDTH-1:0] wire_d25_11;
	wire [WIDTH-1:0] wire_d25_12;
	wire [WIDTH-1:0] wire_d25_13;
	wire [WIDTH-1:0] wire_d25_14;
	wire [WIDTH-1:0] wire_d25_15;
	wire [WIDTH-1:0] wire_d25_16;
	wire [WIDTH-1:0] wire_d25_17;
	wire [WIDTH-1:0] wire_d25_18;
	wire [WIDTH-1:0] wire_d25_19;
	wire [WIDTH-1:0] wire_d25_20;
	wire [WIDTH-1:0] wire_d25_21;
	wire [WIDTH-1:0] wire_d25_22;
	wire [WIDTH-1:0] wire_d25_23;
	wire [WIDTH-1:0] wire_d25_24;
	wire [WIDTH-1:0] wire_d25_25;
	wire [WIDTH-1:0] wire_d25_26;
	wire [WIDTH-1:0] wire_d25_27;
	wire [WIDTH-1:0] wire_d25_28;
	wire [WIDTH-1:0] wire_d25_29;
	wire [WIDTH-1:0] wire_d25_30;
	wire [WIDTH-1:0] wire_d25_31;
	wire [WIDTH-1:0] wire_d25_32;
	wire [WIDTH-1:0] wire_d25_33;
	wire [WIDTH-1:0] wire_d25_34;
	wire [WIDTH-1:0] wire_d25_35;
	wire [WIDTH-1:0] wire_d25_36;
	wire [WIDTH-1:0] wire_d25_37;
	wire [WIDTH-1:0] wire_d25_38;
	wire [WIDTH-1:0] wire_d25_39;
	wire [WIDTH-1:0] wire_d25_40;
	wire [WIDTH-1:0] wire_d25_41;
	wire [WIDTH-1:0] wire_d25_42;
	wire [WIDTH-1:0] wire_d25_43;
	wire [WIDTH-1:0] wire_d25_44;
	wire [WIDTH-1:0] wire_d25_45;
	wire [WIDTH-1:0] wire_d25_46;
	wire [WIDTH-1:0] wire_d25_47;
	wire [WIDTH-1:0] wire_d25_48;
	wire [WIDTH-1:0] wire_d26_0;
	wire [WIDTH-1:0] wire_d26_1;
	wire [WIDTH-1:0] wire_d26_2;
	wire [WIDTH-1:0] wire_d26_3;
	wire [WIDTH-1:0] wire_d26_4;
	wire [WIDTH-1:0] wire_d26_5;
	wire [WIDTH-1:0] wire_d26_6;
	wire [WIDTH-1:0] wire_d26_7;
	wire [WIDTH-1:0] wire_d26_8;
	wire [WIDTH-1:0] wire_d26_9;
	wire [WIDTH-1:0] wire_d26_10;
	wire [WIDTH-1:0] wire_d26_11;
	wire [WIDTH-1:0] wire_d26_12;
	wire [WIDTH-1:0] wire_d26_13;
	wire [WIDTH-1:0] wire_d26_14;
	wire [WIDTH-1:0] wire_d26_15;
	wire [WIDTH-1:0] wire_d26_16;
	wire [WIDTH-1:0] wire_d26_17;
	wire [WIDTH-1:0] wire_d26_18;
	wire [WIDTH-1:0] wire_d26_19;
	wire [WIDTH-1:0] wire_d26_20;
	wire [WIDTH-1:0] wire_d26_21;
	wire [WIDTH-1:0] wire_d26_22;
	wire [WIDTH-1:0] wire_d26_23;
	wire [WIDTH-1:0] wire_d26_24;
	wire [WIDTH-1:0] wire_d26_25;
	wire [WIDTH-1:0] wire_d26_26;
	wire [WIDTH-1:0] wire_d26_27;
	wire [WIDTH-1:0] wire_d26_28;
	wire [WIDTH-1:0] wire_d26_29;
	wire [WIDTH-1:0] wire_d26_30;
	wire [WIDTH-1:0] wire_d26_31;
	wire [WIDTH-1:0] wire_d26_32;
	wire [WIDTH-1:0] wire_d26_33;
	wire [WIDTH-1:0] wire_d26_34;
	wire [WIDTH-1:0] wire_d26_35;
	wire [WIDTH-1:0] wire_d26_36;
	wire [WIDTH-1:0] wire_d26_37;
	wire [WIDTH-1:0] wire_d26_38;
	wire [WIDTH-1:0] wire_d26_39;
	wire [WIDTH-1:0] wire_d26_40;
	wire [WIDTH-1:0] wire_d26_41;
	wire [WIDTH-1:0] wire_d26_42;
	wire [WIDTH-1:0] wire_d26_43;
	wire [WIDTH-1:0] wire_d26_44;
	wire [WIDTH-1:0] wire_d26_45;
	wire [WIDTH-1:0] wire_d26_46;
	wire [WIDTH-1:0] wire_d26_47;
	wire [WIDTH-1:0] wire_d26_48;
	wire [WIDTH-1:0] wire_d27_0;
	wire [WIDTH-1:0] wire_d27_1;
	wire [WIDTH-1:0] wire_d27_2;
	wire [WIDTH-1:0] wire_d27_3;
	wire [WIDTH-1:0] wire_d27_4;
	wire [WIDTH-1:0] wire_d27_5;
	wire [WIDTH-1:0] wire_d27_6;
	wire [WIDTH-1:0] wire_d27_7;
	wire [WIDTH-1:0] wire_d27_8;
	wire [WIDTH-1:0] wire_d27_9;
	wire [WIDTH-1:0] wire_d27_10;
	wire [WIDTH-1:0] wire_d27_11;
	wire [WIDTH-1:0] wire_d27_12;
	wire [WIDTH-1:0] wire_d27_13;
	wire [WIDTH-1:0] wire_d27_14;
	wire [WIDTH-1:0] wire_d27_15;
	wire [WIDTH-1:0] wire_d27_16;
	wire [WIDTH-1:0] wire_d27_17;
	wire [WIDTH-1:0] wire_d27_18;
	wire [WIDTH-1:0] wire_d27_19;
	wire [WIDTH-1:0] wire_d27_20;
	wire [WIDTH-1:0] wire_d27_21;
	wire [WIDTH-1:0] wire_d27_22;
	wire [WIDTH-1:0] wire_d27_23;
	wire [WIDTH-1:0] wire_d27_24;
	wire [WIDTH-1:0] wire_d27_25;
	wire [WIDTH-1:0] wire_d27_26;
	wire [WIDTH-1:0] wire_d27_27;
	wire [WIDTH-1:0] wire_d27_28;
	wire [WIDTH-1:0] wire_d27_29;
	wire [WIDTH-1:0] wire_d27_30;
	wire [WIDTH-1:0] wire_d27_31;
	wire [WIDTH-1:0] wire_d27_32;
	wire [WIDTH-1:0] wire_d27_33;
	wire [WIDTH-1:0] wire_d27_34;
	wire [WIDTH-1:0] wire_d27_35;
	wire [WIDTH-1:0] wire_d27_36;
	wire [WIDTH-1:0] wire_d27_37;
	wire [WIDTH-1:0] wire_d27_38;
	wire [WIDTH-1:0] wire_d27_39;
	wire [WIDTH-1:0] wire_d27_40;
	wire [WIDTH-1:0] wire_d27_41;
	wire [WIDTH-1:0] wire_d27_42;
	wire [WIDTH-1:0] wire_d27_43;
	wire [WIDTH-1:0] wire_d27_44;
	wire [WIDTH-1:0] wire_d27_45;
	wire [WIDTH-1:0] wire_d27_46;
	wire [WIDTH-1:0] wire_d27_47;
	wire [WIDTH-1:0] wire_d27_48;
	wire [WIDTH-1:0] wire_d28_0;
	wire [WIDTH-1:0] wire_d28_1;
	wire [WIDTH-1:0] wire_d28_2;
	wire [WIDTH-1:0] wire_d28_3;
	wire [WIDTH-1:0] wire_d28_4;
	wire [WIDTH-1:0] wire_d28_5;
	wire [WIDTH-1:0] wire_d28_6;
	wire [WIDTH-1:0] wire_d28_7;
	wire [WIDTH-1:0] wire_d28_8;
	wire [WIDTH-1:0] wire_d28_9;
	wire [WIDTH-1:0] wire_d28_10;
	wire [WIDTH-1:0] wire_d28_11;
	wire [WIDTH-1:0] wire_d28_12;
	wire [WIDTH-1:0] wire_d28_13;
	wire [WIDTH-1:0] wire_d28_14;
	wire [WIDTH-1:0] wire_d28_15;
	wire [WIDTH-1:0] wire_d28_16;
	wire [WIDTH-1:0] wire_d28_17;
	wire [WIDTH-1:0] wire_d28_18;
	wire [WIDTH-1:0] wire_d28_19;
	wire [WIDTH-1:0] wire_d28_20;
	wire [WIDTH-1:0] wire_d28_21;
	wire [WIDTH-1:0] wire_d28_22;
	wire [WIDTH-1:0] wire_d28_23;
	wire [WIDTH-1:0] wire_d28_24;
	wire [WIDTH-1:0] wire_d28_25;
	wire [WIDTH-1:0] wire_d28_26;
	wire [WIDTH-1:0] wire_d28_27;
	wire [WIDTH-1:0] wire_d28_28;
	wire [WIDTH-1:0] wire_d28_29;
	wire [WIDTH-1:0] wire_d28_30;
	wire [WIDTH-1:0] wire_d28_31;
	wire [WIDTH-1:0] wire_d28_32;
	wire [WIDTH-1:0] wire_d28_33;
	wire [WIDTH-1:0] wire_d28_34;
	wire [WIDTH-1:0] wire_d28_35;
	wire [WIDTH-1:0] wire_d28_36;
	wire [WIDTH-1:0] wire_d28_37;
	wire [WIDTH-1:0] wire_d28_38;
	wire [WIDTH-1:0] wire_d28_39;
	wire [WIDTH-1:0] wire_d28_40;
	wire [WIDTH-1:0] wire_d28_41;
	wire [WIDTH-1:0] wire_d28_42;
	wire [WIDTH-1:0] wire_d28_43;
	wire [WIDTH-1:0] wire_d28_44;
	wire [WIDTH-1:0] wire_d28_45;
	wire [WIDTH-1:0] wire_d28_46;
	wire [WIDTH-1:0] wire_d28_47;
	wire [WIDTH-1:0] wire_d28_48;
	wire [WIDTH-1:0] wire_d29_0;
	wire [WIDTH-1:0] wire_d29_1;
	wire [WIDTH-1:0] wire_d29_2;
	wire [WIDTH-1:0] wire_d29_3;
	wire [WIDTH-1:0] wire_d29_4;
	wire [WIDTH-1:0] wire_d29_5;
	wire [WIDTH-1:0] wire_d29_6;
	wire [WIDTH-1:0] wire_d29_7;
	wire [WIDTH-1:0] wire_d29_8;
	wire [WIDTH-1:0] wire_d29_9;
	wire [WIDTH-1:0] wire_d29_10;
	wire [WIDTH-1:0] wire_d29_11;
	wire [WIDTH-1:0] wire_d29_12;
	wire [WIDTH-1:0] wire_d29_13;
	wire [WIDTH-1:0] wire_d29_14;
	wire [WIDTH-1:0] wire_d29_15;
	wire [WIDTH-1:0] wire_d29_16;
	wire [WIDTH-1:0] wire_d29_17;
	wire [WIDTH-1:0] wire_d29_18;
	wire [WIDTH-1:0] wire_d29_19;
	wire [WIDTH-1:0] wire_d29_20;
	wire [WIDTH-1:0] wire_d29_21;
	wire [WIDTH-1:0] wire_d29_22;
	wire [WIDTH-1:0] wire_d29_23;
	wire [WIDTH-1:0] wire_d29_24;
	wire [WIDTH-1:0] wire_d29_25;
	wire [WIDTH-1:0] wire_d29_26;
	wire [WIDTH-1:0] wire_d29_27;
	wire [WIDTH-1:0] wire_d29_28;
	wire [WIDTH-1:0] wire_d29_29;
	wire [WIDTH-1:0] wire_d29_30;
	wire [WIDTH-1:0] wire_d29_31;
	wire [WIDTH-1:0] wire_d29_32;
	wire [WIDTH-1:0] wire_d29_33;
	wire [WIDTH-1:0] wire_d29_34;
	wire [WIDTH-1:0] wire_d29_35;
	wire [WIDTH-1:0] wire_d29_36;
	wire [WIDTH-1:0] wire_d29_37;
	wire [WIDTH-1:0] wire_d29_38;
	wire [WIDTH-1:0] wire_d29_39;
	wire [WIDTH-1:0] wire_d29_40;
	wire [WIDTH-1:0] wire_d29_41;
	wire [WIDTH-1:0] wire_d29_42;
	wire [WIDTH-1:0] wire_d29_43;
	wire [WIDTH-1:0] wire_d29_44;
	wire [WIDTH-1:0] wire_d29_45;
	wire [WIDTH-1:0] wire_d29_46;
	wire [WIDTH-1:0] wire_d29_47;
	wire [WIDTH-1:0] wire_d29_48;

	invertion #(.WIDTH(WIDTH)) invertion_instance100(.data_in(d_in0),.data_out(wire_d0_0),.clk(clk),.rst(rst));            //channel 1
	large_mux #(.WIDTH(WIDTH)) large_mux_instance101(.data_in(wire_d0_0),.data_out(wire_d0_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance102(.data_in(wire_d0_1),.data_out(wire_d0_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance103(.data_in(wire_d0_2),.data_out(wire_d0_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance104(.data_in(wire_d0_3),.data_out(wire_d0_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance105(.data_in(wire_d0_4),.data_out(wire_d0_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance106(.data_in(wire_d0_5),.data_out(wire_d0_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance107(.data_in(wire_d0_6),.data_out(wire_d0_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance108(.data_in(wire_d0_7),.data_out(wire_d0_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance109(.data_in(wire_d0_8),.data_out(wire_d0_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1010(.data_in(wire_d0_9),.data_out(wire_d0_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1011(.data_in(wire_d0_10),.data_out(wire_d0_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1012(.data_in(wire_d0_11),.data_out(wire_d0_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1013(.data_in(wire_d0_12),.data_out(wire_d0_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1014(.data_in(wire_d0_13),.data_out(wire_d0_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1015(.data_in(wire_d0_14),.data_out(wire_d0_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1016(.data_in(wire_d0_15),.data_out(wire_d0_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1017(.data_in(wire_d0_16),.data_out(wire_d0_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1018(.data_in(wire_d0_17),.data_out(wire_d0_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1019(.data_in(wire_d0_18),.data_out(wire_d0_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1020(.data_in(wire_d0_19),.data_out(wire_d0_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1021(.data_in(wire_d0_20),.data_out(wire_d0_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1022(.data_in(wire_d0_21),.data_out(wire_d0_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1023(.data_in(wire_d0_22),.data_out(wire_d0_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1024(.data_in(wire_d0_23),.data_out(wire_d0_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1025(.data_in(wire_d0_24),.data_out(wire_d0_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1026(.data_in(wire_d0_25),.data_out(wire_d0_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1027(.data_in(wire_d0_26),.data_out(wire_d0_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1028(.data_in(wire_d0_27),.data_out(wire_d0_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1029(.data_in(wire_d0_28),.data_out(wire_d0_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1030(.data_in(wire_d0_29),.data_out(wire_d0_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1031(.data_in(wire_d0_30),.data_out(wire_d0_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1032(.data_in(wire_d0_31),.data_out(wire_d0_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1033(.data_in(wire_d0_32),.data_out(wire_d0_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1034(.data_in(wire_d0_33),.data_out(wire_d0_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1035(.data_in(wire_d0_34),.data_out(wire_d0_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1036(.data_in(wire_d0_35),.data_out(wire_d0_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1037(.data_in(wire_d0_36),.data_out(wire_d0_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1038(.data_in(wire_d0_37),.data_out(wire_d0_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1039(.data_in(wire_d0_38),.data_out(wire_d0_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1040(.data_in(wire_d0_39),.data_out(wire_d0_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1041(.data_in(wire_d0_40),.data_out(wire_d0_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1042(.data_in(wire_d0_41),.data_out(wire_d0_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1043(.data_in(wire_d0_42),.data_out(wire_d0_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1044(.data_in(wire_d0_43),.data_out(wire_d0_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1045(.data_in(wire_d0_44),.data_out(wire_d0_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1046(.data_in(wire_d0_45),.data_out(wire_d0_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1047(.data_in(wire_d0_46),.data_out(wire_d0_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1048(.data_in(wire_d0_47),.data_out(wire_d0_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1049(.data_in(wire_d0_48),.data_out(d_out0),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance210(.data_in(d_in1),.data_out(wire_d1_0),.clk(clk),.rst(rst));            //channel 2
	encoder #(.WIDTH(WIDTH)) encoder_instance211(.data_in(wire_d1_0),.data_out(wire_d1_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212(.data_in(wire_d1_1),.data_out(wire_d1_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance213(.data_in(wire_d1_2),.data_out(wire_d1_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance214(.data_in(wire_d1_3),.data_out(wire_d1_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance215(.data_in(wire_d1_4),.data_out(wire_d1_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance216(.data_in(wire_d1_5),.data_out(wire_d1_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance217(.data_in(wire_d1_6),.data_out(wire_d1_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance218(.data_in(wire_d1_7),.data_out(wire_d1_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance219(.data_in(wire_d1_8),.data_out(wire_d1_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2110(.data_in(wire_d1_9),.data_out(wire_d1_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2111(.data_in(wire_d1_10),.data_out(wire_d1_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2112(.data_in(wire_d1_11),.data_out(wire_d1_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2113(.data_in(wire_d1_12),.data_out(wire_d1_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2114(.data_in(wire_d1_13),.data_out(wire_d1_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2115(.data_in(wire_d1_14),.data_out(wire_d1_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2116(.data_in(wire_d1_15),.data_out(wire_d1_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2117(.data_in(wire_d1_16),.data_out(wire_d1_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2118(.data_in(wire_d1_17),.data_out(wire_d1_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2119(.data_in(wire_d1_18),.data_out(wire_d1_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2120(.data_in(wire_d1_19),.data_out(wire_d1_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2121(.data_in(wire_d1_20),.data_out(wire_d1_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2122(.data_in(wire_d1_21),.data_out(wire_d1_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2123(.data_in(wire_d1_22),.data_out(wire_d1_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2124(.data_in(wire_d1_23),.data_out(wire_d1_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2125(.data_in(wire_d1_24),.data_out(wire_d1_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2126(.data_in(wire_d1_25),.data_out(wire_d1_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2127(.data_in(wire_d1_26),.data_out(wire_d1_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2128(.data_in(wire_d1_27),.data_out(wire_d1_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2129(.data_in(wire_d1_28),.data_out(wire_d1_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2130(.data_in(wire_d1_29),.data_out(wire_d1_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2131(.data_in(wire_d1_30),.data_out(wire_d1_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2132(.data_in(wire_d1_31),.data_out(wire_d1_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2133(.data_in(wire_d1_32),.data_out(wire_d1_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2134(.data_in(wire_d1_33),.data_out(wire_d1_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2135(.data_in(wire_d1_34),.data_out(wire_d1_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2136(.data_in(wire_d1_35),.data_out(wire_d1_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2137(.data_in(wire_d1_36),.data_out(wire_d1_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2138(.data_in(wire_d1_37),.data_out(wire_d1_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2139(.data_in(wire_d1_38),.data_out(wire_d1_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2140(.data_in(wire_d1_39),.data_out(wire_d1_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2141(.data_in(wire_d1_40),.data_out(wire_d1_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2142(.data_in(wire_d1_41),.data_out(wire_d1_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2143(.data_in(wire_d1_42),.data_out(wire_d1_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2144(.data_in(wire_d1_43),.data_out(wire_d1_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2145(.data_in(wire_d1_44),.data_out(wire_d1_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2146(.data_in(wire_d1_45),.data_out(wire_d1_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2147(.data_in(wire_d1_46),.data_out(wire_d1_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2148(.data_in(wire_d1_47),.data_out(wire_d1_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2149(.data_in(wire_d1_48),.data_out(d_out1),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance320(.data_in(d_in2),.data_out(wire_d2_0),.clk(clk),.rst(rst));            //channel 3
	large_mux #(.WIDTH(WIDTH)) large_mux_instance321(.data_in(wire_d2_0),.data_out(wire_d2_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance322(.data_in(wire_d2_1),.data_out(wire_d2_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance323(.data_in(wire_d2_2),.data_out(wire_d2_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance324(.data_in(wire_d2_3),.data_out(wire_d2_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance325(.data_in(wire_d2_4),.data_out(wire_d2_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance326(.data_in(wire_d2_5),.data_out(wire_d2_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance327(.data_in(wire_d2_6),.data_out(wire_d2_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance328(.data_in(wire_d2_7),.data_out(wire_d2_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance329(.data_in(wire_d2_8),.data_out(wire_d2_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3210(.data_in(wire_d2_9),.data_out(wire_d2_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3211(.data_in(wire_d2_10),.data_out(wire_d2_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3212(.data_in(wire_d2_11),.data_out(wire_d2_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3213(.data_in(wire_d2_12),.data_out(wire_d2_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3214(.data_in(wire_d2_13),.data_out(wire_d2_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3215(.data_in(wire_d2_14),.data_out(wire_d2_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3216(.data_in(wire_d2_15),.data_out(wire_d2_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3217(.data_in(wire_d2_16),.data_out(wire_d2_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3218(.data_in(wire_d2_17),.data_out(wire_d2_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3219(.data_in(wire_d2_18),.data_out(wire_d2_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3220(.data_in(wire_d2_19),.data_out(wire_d2_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3221(.data_in(wire_d2_20),.data_out(wire_d2_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3222(.data_in(wire_d2_21),.data_out(wire_d2_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3223(.data_in(wire_d2_22),.data_out(wire_d2_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3224(.data_in(wire_d2_23),.data_out(wire_d2_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3225(.data_in(wire_d2_24),.data_out(wire_d2_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3226(.data_in(wire_d2_25),.data_out(wire_d2_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3227(.data_in(wire_d2_26),.data_out(wire_d2_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3228(.data_in(wire_d2_27),.data_out(wire_d2_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3229(.data_in(wire_d2_28),.data_out(wire_d2_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3230(.data_in(wire_d2_29),.data_out(wire_d2_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3231(.data_in(wire_d2_30),.data_out(wire_d2_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3232(.data_in(wire_d2_31),.data_out(wire_d2_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3233(.data_in(wire_d2_32),.data_out(wire_d2_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3234(.data_in(wire_d2_33),.data_out(wire_d2_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3235(.data_in(wire_d2_34),.data_out(wire_d2_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3236(.data_in(wire_d2_35),.data_out(wire_d2_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3237(.data_in(wire_d2_36),.data_out(wire_d2_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3238(.data_in(wire_d2_37),.data_out(wire_d2_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3239(.data_in(wire_d2_38),.data_out(wire_d2_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3240(.data_in(wire_d2_39),.data_out(wire_d2_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3241(.data_in(wire_d2_40),.data_out(wire_d2_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3242(.data_in(wire_d2_41),.data_out(wire_d2_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3243(.data_in(wire_d2_42),.data_out(wire_d2_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3244(.data_in(wire_d2_43),.data_out(wire_d2_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3245(.data_in(wire_d2_44),.data_out(wire_d2_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3246(.data_in(wire_d2_45),.data_out(wire_d2_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3247(.data_in(wire_d2_46),.data_out(wire_d2_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3248(.data_in(wire_d2_47),.data_out(wire_d2_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3249(.data_in(wire_d2_48),.data_out(d_out2),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance430(.data_in(d_in3),.data_out(wire_d3_0),.clk(clk),.rst(rst));            //channel 4
	encoder #(.WIDTH(WIDTH)) encoder_instance431(.data_in(wire_d3_0),.data_out(wire_d3_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance432(.data_in(wire_d3_1),.data_out(wire_d3_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance433(.data_in(wire_d3_2),.data_out(wire_d3_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance434(.data_in(wire_d3_3),.data_out(wire_d3_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance435(.data_in(wire_d3_4),.data_out(wire_d3_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance436(.data_in(wire_d3_5),.data_out(wire_d3_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance437(.data_in(wire_d3_6),.data_out(wire_d3_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance438(.data_in(wire_d3_7),.data_out(wire_d3_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance439(.data_in(wire_d3_8),.data_out(wire_d3_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4310(.data_in(wire_d3_9),.data_out(wire_d3_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4311(.data_in(wire_d3_10),.data_out(wire_d3_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4312(.data_in(wire_d3_11),.data_out(wire_d3_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4313(.data_in(wire_d3_12),.data_out(wire_d3_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4314(.data_in(wire_d3_13),.data_out(wire_d3_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4315(.data_in(wire_d3_14),.data_out(wire_d3_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4316(.data_in(wire_d3_15),.data_out(wire_d3_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4317(.data_in(wire_d3_16),.data_out(wire_d3_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4318(.data_in(wire_d3_17),.data_out(wire_d3_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4319(.data_in(wire_d3_18),.data_out(wire_d3_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4320(.data_in(wire_d3_19),.data_out(wire_d3_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4321(.data_in(wire_d3_20),.data_out(wire_d3_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4322(.data_in(wire_d3_21),.data_out(wire_d3_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4323(.data_in(wire_d3_22),.data_out(wire_d3_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4324(.data_in(wire_d3_23),.data_out(wire_d3_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4325(.data_in(wire_d3_24),.data_out(wire_d3_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4326(.data_in(wire_d3_25),.data_out(wire_d3_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4327(.data_in(wire_d3_26),.data_out(wire_d3_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4328(.data_in(wire_d3_27),.data_out(wire_d3_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4329(.data_in(wire_d3_28),.data_out(wire_d3_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4330(.data_in(wire_d3_29),.data_out(wire_d3_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4331(.data_in(wire_d3_30),.data_out(wire_d3_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4332(.data_in(wire_d3_31),.data_out(wire_d3_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4333(.data_in(wire_d3_32),.data_out(wire_d3_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4334(.data_in(wire_d3_33),.data_out(wire_d3_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4335(.data_in(wire_d3_34),.data_out(wire_d3_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4336(.data_in(wire_d3_35),.data_out(wire_d3_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4337(.data_in(wire_d3_36),.data_out(wire_d3_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4338(.data_in(wire_d3_37),.data_out(wire_d3_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4339(.data_in(wire_d3_38),.data_out(wire_d3_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4340(.data_in(wire_d3_39),.data_out(wire_d3_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4341(.data_in(wire_d3_40),.data_out(wire_d3_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4342(.data_in(wire_d3_41),.data_out(wire_d3_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4343(.data_in(wire_d3_42),.data_out(wire_d3_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4344(.data_in(wire_d3_43),.data_out(wire_d3_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4345(.data_in(wire_d3_44),.data_out(wire_d3_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4346(.data_in(wire_d3_45),.data_out(wire_d3_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4347(.data_in(wire_d3_46),.data_out(wire_d3_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4348(.data_in(wire_d3_47),.data_out(wire_d3_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4349(.data_in(wire_d3_48),.data_out(d_out3),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance540(.data_in(d_in4),.data_out(wire_d4_0),.clk(clk),.rst(rst));            //channel 5
	invertion #(.WIDTH(WIDTH)) invertion_instance541(.data_in(wire_d4_0),.data_out(wire_d4_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance542(.data_in(wire_d4_1),.data_out(wire_d4_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance543(.data_in(wire_d4_2),.data_out(wire_d4_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance544(.data_in(wire_d4_3),.data_out(wire_d4_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance545(.data_in(wire_d4_4),.data_out(wire_d4_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance546(.data_in(wire_d4_5),.data_out(wire_d4_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance547(.data_in(wire_d4_6),.data_out(wire_d4_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance548(.data_in(wire_d4_7),.data_out(wire_d4_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance549(.data_in(wire_d4_8),.data_out(wire_d4_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5410(.data_in(wire_d4_9),.data_out(wire_d4_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5411(.data_in(wire_d4_10),.data_out(wire_d4_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5412(.data_in(wire_d4_11),.data_out(wire_d4_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5413(.data_in(wire_d4_12),.data_out(wire_d4_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5414(.data_in(wire_d4_13),.data_out(wire_d4_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5415(.data_in(wire_d4_14),.data_out(wire_d4_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5416(.data_in(wire_d4_15),.data_out(wire_d4_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5417(.data_in(wire_d4_16),.data_out(wire_d4_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5418(.data_in(wire_d4_17),.data_out(wire_d4_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5419(.data_in(wire_d4_18),.data_out(wire_d4_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5420(.data_in(wire_d4_19),.data_out(wire_d4_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5421(.data_in(wire_d4_20),.data_out(wire_d4_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5422(.data_in(wire_d4_21),.data_out(wire_d4_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5423(.data_in(wire_d4_22),.data_out(wire_d4_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5424(.data_in(wire_d4_23),.data_out(wire_d4_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5425(.data_in(wire_d4_24),.data_out(wire_d4_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5426(.data_in(wire_d4_25),.data_out(wire_d4_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5427(.data_in(wire_d4_26),.data_out(wire_d4_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5428(.data_in(wire_d4_27),.data_out(wire_d4_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5429(.data_in(wire_d4_28),.data_out(wire_d4_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5430(.data_in(wire_d4_29),.data_out(wire_d4_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5431(.data_in(wire_d4_30),.data_out(wire_d4_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5432(.data_in(wire_d4_31),.data_out(wire_d4_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5433(.data_in(wire_d4_32),.data_out(wire_d4_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5434(.data_in(wire_d4_33),.data_out(wire_d4_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5435(.data_in(wire_d4_34),.data_out(wire_d4_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5436(.data_in(wire_d4_35),.data_out(wire_d4_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5437(.data_in(wire_d4_36),.data_out(wire_d4_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5438(.data_in(wire_d4_37),.data_out(wire_d4_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5439(.data_in(wire_d4_38),.data_out(wire_d4_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5440(.data_in(wire_d4_39),.data_out(wire_d4_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5441(.data_in(wire_d4_40),.data_out(wire_d4_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5442(.data_in(wire_d4_41),.data_out(wire_d4_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5443(.data_in(wire_d4_42),.data_out(wire_d4_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5444(.data_in(wire_d4_43),.data_out(wire_d4_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5445(.data_in(wire_d4_44),.data_out(wire_d4_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5446(.data_in(wire_d4_45),.data_out(wire_d4_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5447(.data_in(wire_d4_46),.data_out(wire_d4_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5448(.data_in(wire_d4_47),.data_out(wire_d4_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5449(.data_in(wire_d4_48),.data_out(d_out4),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance650(.data_in(d_in5),.data_out(wire_d5_0),.clk(clk),.rst(rst));            //channel 6
	invertion #(.WIDTH(WIDTH)) invertion_instance651(.data_in(wire_d5_0),.data_out(wire_d5_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance652(.data_in(wire_d5_1),.data_out(wire_d5_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance653(.data_in(wire_d5_2),.data_out(wire_d5_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance654(.data_in(wire_d5_3),.data_out(wire_d5_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance655(.data_in(wire_d5_4),.data_out(wire_d5_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance656(.data_in(wire_d5_5),.data_out(wire_d5_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance657(.data_in(wire_d5_6),.data_out(wire_d5_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance658(.data_in(wire_d5_7),.data_out(wire_d5_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance659(.data_in(wire_d5_8),.data_out(wire_d5_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6510(.data_in(wire_d5_9),.data_out(wire_d5_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6511(.data_in(wire_d5_10),.data_out(wire_d5_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6512(.data_in(wire_d5_11),.data_out(wire_d5_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6513(.data_in(wire_d5_12),.data_out(wire_d5_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6514(.data_in(wire_d5_13),.data_out(wire_d5_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6515(.data_in(wire_d5_14),.data_out(wire_d5_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6516(.data_in(wire_d5_15),.data_out(wire_d5_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6517(.data_in(wire_d5_16),.data_out(wire_d5_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6518(.data_in(wire_d5_17),.data_out(wire_d5_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6519(.data_in(wire_d5_18),.data_out(wire_d5_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6520(.data_in(wire_d5_19),.data_out(wire_d5_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6521(.data_in(wire_d5_20),.data_out(wire_d5_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6522(.data_in(wire_d5_21),.data_out(wire_d5_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6523(.data_in(wire_d5_22),.data_out(wire_d5_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6524(.data_in(wire_d5_23),.data_out(wire_d5_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6525(.data_in(wire_d5_24),.data_out(wire_d5_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6526(.data_in(wire_d5_25),.data_out(wire_d5_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6527(.data_in(wire_d5_26),.data_out(wire_d5_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6528(.data_in(wire_d5_27),.data_out(wire_d5_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6529(.data_in(wire_d5_28),.data_out(wire_d5_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6530(.data_in(wire_d5_29),.data_out(wire_d5_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6531(.data_in(wire_d5_30),.data_out(wire_d5_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6532(.data_in(wire_d5_31),.data_out(wire_d5_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6533(.data_in(wire_d5_32),.data_out(wire_d5_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6534(.data_in(wire_d5_33),.data_out(wire_d5_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6535(.data_in(wire_d5_34),.data_out(wire_d5_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6536(.data_in(wire_d5_35),.data_out(wire_d5_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6537(.data_in(wire_d5_36),.data_out(wire_d5_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6538(.data_in(wire_d5_37),.data_out(wire_d5_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6539(.data_in(wire_d5_38),.data_out(wire_d5_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6540(.data_in(wire_d5_39),.data_out(wire_d5_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6541(.data_in(wire_d5_40),.data_out(wire_d5_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6542(.data_in(wire_d5_41),.data_out(wire_d5_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6543(.data_in(wire_d5_42),.data_out(wire_d5_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6544(.data_in(wire_d5_43),.data_out(wire_d5_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6545(.data_in(wire_d5_44),.data_out(wire_d5_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6546(.data_in(wire_d5_45),.data_out(wire_d5_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6547(.data_in(wire_d5_46),.data_out(wire_d5_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6548(.data_in(wire_d5_47),.data_out(wire_d5_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6549(.data_in(wire_d5_48),.data_out(d_out5),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance760(.data_in(d_in6),.data_out(wire_d6_0),.clk(clk),.rst(rst));            //channel 7
	invertion #(.WIDTH(WIDTH)) invertion_instance761(.data_in(wire_d6_0),.data_out(wire_d6_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance762(.data_in(wire_d6_1),.data_out(wire_d6_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance763(.data_in(wire_d6_2),.data_out(wire_d6_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance764(.data_in(wire_d6_3),.data_out(wire_d6_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance765(.data_in(wire_d6_4),.data_out(wire_d6_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance766(.data_in(wire_d6_5),.data_out(wire_d6_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance767(.data_in(wire_d6_6),.data_out(wire_d6_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance768(.data_in(wire_d6_7),.data_out(wire_d6_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance769(.data_in(wire_d6_8),.data_out(wire_d6_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7610(.data_in(wire_d6_9),.data_out(wire_d6_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7611(.data_in(wire_d6_10),.data_out(wire_d6_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7612(.data_in(wire_d6_11),.data_out(wire_d6_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7613(.data_in(wire_d6_12),.data_out(wire_d6_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7614(.data_in(wire_d6_13),.data_out(wire_d6_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7615(.data_in(wire_d6_14),.data_out(wire_d6_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7616(.data_in(wire_d6_15),.data_out(wire_d6_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7617(.data_in(wire_d6_16),.data_out(wire_d6_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7618(.data_in(wire_d6_17),.data_out(wire_d6_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7619(.data_in(wire_d6_18),.data_out(wire_d6_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7620(.data_in(wire_d6_19),.data_out(wire_d6_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7621(.data_in(wire_d6_20),.data_out(wire_d6_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7622(.data_in(wire_d6_21),.data_out(wire_d6_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7623(.data_in(wire_d6_22),.data_out(wire_d6_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7624(.data_in(wire_d6_23),.data_out(wire_d6_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7625(.data_in(wire_d6_24),.data_out(wire_d6_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7626(.data_in(wire_d6_25),.data_out(wire_d6_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7627(.data_in(wire_d6_26),.data_out(wire_d6_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7628(.data_in(wire_d6_27),.data_out(wire_d6_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7629(.data_in(wire_d6_28),.data_out(wire_d6_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7630(.data_in(wire_d6_29),.data_out(wire_d6_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7631(.data_in(wire_d6_30),.data_out(wire_d6_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7632(.data_in(wire_d6_31),.data_out(wire_d6_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7633(.data_in(wire_d6_32),.data_out(wire_d6_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7634(.data_in(wire_d6_33),.data_out(wire_d6_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7635(.data_in(wire_d6_34),.data_out(wire_d6_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7636(.data_in(wire_d6_35),.data_out(wire_d6_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7637(.data_in(wire_d6_36),.data_out(wire_d6_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7638(.data_in(wire_d6_37),.data_out(wire_d6_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7639(.data_in(wire_d6_38),.data_out(wire_d6_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7640(.data_in(wire_d6_39),.data_out(wire_d6_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7641(.data_in(wire_d6_40),.data_out(wire_d6_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7642(.data_in(wire_d6_41),.data_out(wire_d6_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7643(.data_in(wire_d6_42),.data_out(wire_d6_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7644(.data_in(wire_d6_43),.data_out(wire_d6_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7645(.data_in(wire_d6_44),.data_out(wire_d6_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7646(.data_in(wire_d6_45),.data_out(wire_d6_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7647(.data_in(wire_d6_46),.data_out(wire_d6_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7648(.data_in(wire_d6_47),.data_out(wire_d6_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7649(.data_in(wire_d6_48),.data_out(d_out6),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance870(.data_in(d_in7),.data_out(wire_d7_0),.clk(clk),.rst(rst));            //channel 8
	register #(.WIDTH(WIDTH)) register_instance871(.data_in(wire_d7_0),.data_out(wire_d7_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance872(.data_in(wire_d7_1),.data_out(wire_d7_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance873(.data_in(wire_d7_2),.data_out(wire_d7_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance874(.data_in(wire_d7_3),.data_out(wire_d7_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance875(.data_in(wire_d7_4),.data_out(wire_d7_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance876(.data_in(wire_d7_5),.data_out(wire_d7_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance877(.data_in(wire_d7_6),.data_out(wire_d7_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance878(.data_in(wire_d7_7),.data_out(wire_d7_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance879(.data_in(wire_d7_8),.data_out(wire_d7_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8710(.data_in(wire_d7_9),.data_out(wire_d7_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8711(.data_in(wire_d7_10),.data_out(wire_d7_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8712(.data_in(wire_d7_11),.data_out(wire_d7_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8713(.data_in(wire_d7_12),.data_out(wire_d7_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8714(.data_in(wire_d7_13),.data_out(wire_d7_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8715(.data_in(wire_d7_14),.data_out(wire_d7_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8716(.data_in(wire_d7_15),.data_out(wire_d7_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8717(.data_in(wire_d7_16),.data_out(wire_d7_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8718(.data_in(wire_d7_17),.data_out(wire_d7_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8719(.data_in(wire_d7_18),.data_out(wire_d7_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8720(.data_in(wire_d7_19),.data_out(wire_d7_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8721(.data_in(wire_d7_20),.data_out(wire_d7_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8722(.data_in(wire_d7_21),.data_out(wire_d7_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8723(.data_in(wire_d7_22),.data_out(wire_d7_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8724(.data_in(wire_d7_23),.data_out(wire_d7_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8725(.data_in(wire_d7_24),.data_out(wire_d7_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8726(.data_in(wire_d7_25),.data_out(wire_d7_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8727(.data_in(wire_d7_26),.data_out(wire_d7_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8728(.data_in(wire_d7_27),.data_out(wire_d7_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8729(.data_in(wire_d7_28),.data_out(wire_d7_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8730(.data_in(wire_d7_29),.data_out(wire_d7_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8731(.data_in(wire_d7_30),.data_out(wire_d7_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8732(.data_in(wire_d7_31),.data_out(wire_d7_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8733(.data_in(wire_d7_32),.data_out(wire_d7_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8734(.data_in(wire_d7_33),.data_out(wire_d7_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8735(.data_in(wire_d7_34),.data_out(wire_d7_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8736(.data_in(wire_d7_35),.data_out(wire_d7_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8737(.data_in(wire_d7_36),.data_out(wire_d7_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8738(.data_in(wire_d7_37),.data_out(wire_d7_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8739(.data_in(wire_d7_38),.data_out(wire_d7_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8740(.data_in(wire_d7_39),.data_out(wire_d7_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8741(.data_in(wire_d7_40),.data_out(wire_d7_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8742(.data_in(wire_d7_41),.data_out(wire_d7_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8743(.data_in(wire_d7_42),.data_out(wire_d7_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8744(.data_in(wire_d7_43),.data_out(wire_d7_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8745(.data_in(wire_d7_44),.data_out(wire_d7_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8746(.data_in(wire_d7_45),.data_out(wire_d7_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8747(.data_in(wire_d7_46),.data_out(wire_d7_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8748(.data_in(wire_d7_47),.data_out(wire_d7_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8749(.data_in(wire_d7_48),.data_out(d_out7),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance980(.data_in(d_in8),.data_out(wire_d8_0),.clk(clk),.rst(rst));            //channel 9
	encoder #(.WIDTH(WIDTH)) encoder_instance981(.data_in(wire_d8_0),.data_out(wire_d8_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance982(.data_in(wire_d8_1),.data_out(wire_d8_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance983(.data_in(wire_d8_2),.data_out(wire_d8_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance984(.data_in(wire_d8_3),.data_out(wire_d8_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance985(.data_in(wire_d8_4),.data_out(wire_d8_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance986(.data_in(wire_d8_5),.data_out(wire_d8_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance987(.data_in(wire_d8_6),.data_out(wire_d8_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance988(.data_in(wire_d8_7),.data_out(wire_d8_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance989(.data_in(wire_d8_8),.data_out(wire_d8_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9810(.data_in(wire_d8_9),.data_out(wire_d8_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9811(.data_in(wire_d8_10),.data_out(wire_d8_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9812(.data_in(wire_d8_11),.data_out(wire_d8_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9813(.data_in(wire_d8_12),.data_out(wire_d8_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9814(.data_in(wire_d8_13),.data_out(wire_d8_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9815(.data_in(wire_d8_14),.data_out(wire_d8_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9816(.data_in(wire_d8_15),.data_out(wire_d8_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9817(.data_in(wire_d8_16),.data_out(wire_d8_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9818(.data_in(wire_d8_17),.data_out(wire_d8_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9819(.data_in(wire_d8_18),.data_out(wire_d8_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9820(.data_in(wire_d8_19),.data_out(wire_d8_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9821(.data_in(wire_d8_20),.data_out(wire_d8_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9822(.data_in(wire_d8_21),.data_out(wire_d8_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9823(.data_in(wire_d8_22),.data_out(wire_d8_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9824(.data_in(wire_d8_23),.data_out(wire_d8_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9825(.data_in(wire_d8_24),.data_out(wire_d8_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9826(.data_in(wire_d8_25),.data_out(wire_d8_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9827(.data_in(wire_d8_26),.data_out(wire_d8_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9828(.data_in(wire_d8_27),.data_out(wire_d8_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9829(.data_in(wire_d8_28),.data_out(wire_d8_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9830(.data_in(wire_d8_29),.data_out(wire_d8_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9831(.data_in(wire_d8_30),.data_out(wire_d8_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9832(.data_in(wire_d8_31),.data_out(wire_d8_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9833(.data_in(wire_d8_32),.data_out(wire_d8_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9834(.data_in(wire_d8_33),.data_out(wire_d8_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9835(.data_in(wire_d8_34),.data_out(wire_d8_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9836(.data_in(wire_d8_35),.data_out(wire_d8_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9837(.data_in(wire_d8_36),.data_out(wire_d8_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9838(.data_in(wire_d8_37),.data_out(wire_d8_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9839(.data_in(wire_d8_38),.data_out(wire_d8_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9840(.data_in(wire_d8_39),.data_out(wire_d8_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9841(.data_in(wire_d8_40),.data_out(wire_d8_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9842(.data_in(wire_d8_41),.data_out(wire_d8_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9843(.data_in(wire_d8_42),.data_out(wire_d8_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9844(.data_in(wire_d8_43),.data_out(wire_d8_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9845(.data_in(wire_d8_44),.data_out(wire_d8_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9846(.data_in(wire_d8_45),.data_out(wire_d8_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9847(.data_in(wire_d8_46),.data_out(wire_d8_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9848(.data_in(wire_d8_47),.data_out(wire_d8_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9849(.data_in(wire_d8_48),.data_out(d_out8),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance1090(.data_in(d_in9),.data_out(wire_d9_0),.clk(clk),.rst(rst));            //channel 10
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1091(.data_in(wire_d9_0),.data_out(wire_d9_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1092(.data_in(wire_d9_1),.data_out(wire_d9_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1093(.data_in(wire_d9_2),.data_out(wire_d9_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1094(.data_in(wire_d9_3),.data_out(wire_d9_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1095(.data_in(wire_d9_4),.data_out(wire_d9_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1096(.data_in(wire_d9_5),.data_out(wire_d9_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1097(.data_in(wire_d9_6),.data_out(wire_d9_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1098(.data_in(wire_d9_7),.data_out(wire_d9_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1099(.data_in(wire_d9_8),.data_out(wire_d9_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10910(.data_in(wire_d9_9),.data_out(wire_d9_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10911(.data_in(wire_d9_10),.data_out(wire_d9_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10912(.data_in(wire_d9_11),.data_out(wire_d9_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10913(.data_in(wire_d9_12),.data_out(wire_d9_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10914(.data_in(wire_d9_13),.data_out(wire_d9_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10915(.data_in(wire_d9_14),.data_out(wire_d9_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10916(.data_in(wire_d9_15),.data_out(wire_d9_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10917(.data_in(wire_d9_16),.data_out(wire_d9_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10918(.data_in(wire_d9_17),.data_out(wire_d9_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10919(.data_in(wire_d9_18),.data_out(wire_d9_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10920(.data_in(wire_d9_19),.data_out(wire_d9_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10921(.data_in(wire_d9_20),.data_out(wire_d9_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10922(.data_in(wire_d9_21),.data_out(wire_d9_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10923(.data_in(wire_d9_22),.data_out(wire_d9_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10924(.data_in(wire_d9_23),.data_out(wire_d9_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10925(.data_in(wire_d9_24),.data_out(wire_d9_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10926(.data_in(wire_d9_25),.data_out(wire_d9_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10927(.data_in(wire_d9_26),.data_out(wire_d9_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10928(.data_in(wire_d9_27),.data_out(wire_d9_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10929(.data_in(wire_d9_28),.data_out(wire_d9_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10930(.data_in(wire_d9_29),.data_out(wire_d9_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10931(.data_in(wire_d9_30),.data_out(wire_d9_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10932(.data_in(wire_d9_31),.data_out(wire_d9_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10933(.data_in(wire_d9_32),.data_out(wire_d9_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10934(.data_in(wire_d9_33),.data_out(wire_d9_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10935(.data_in(wire_d9_34),.data_out(wire_d9_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10936(.data_in(wire_d9_35),.data_out(wire_d9_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10937(.data_in(wire_d9_36),.data_out(wire_d9_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10938(.data_in(wire_d9_37),.data_out(wire_d9_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10939(.data_in(wire_d9_38),.data_out(wire_d9_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10940(.data_in(wire_d9_39),.data_out(wire_d9_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance10941(.data_in(wire_d9_40),.data_out(wire_d9_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10942(.data_in(wire_d9_41),.data_out(wire_d9_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10943(.data_in(wire_d9_42),.data_out(wire_d9_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10944(.data_in(wire_d9_43),.data_out(wire_d9_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10945(.data_in(wire_d9_44),.data_out(wire_d9_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10946(.data_in(wire_d9_45),.data_out(wire_d9_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10947(.data_in(wire_d9_46),.data_out(wire_d9_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance10948(.data_in(wire_d9_47),.data_out(wire_d9_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10949(.data_in(wire_d9_48),.data_out(d_out9),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance11100(.data_in(d_in10),.data_out(wire_d10_0),.clk(clk),.rst(rst));            //channel 11
	large_mux #(.WIDTH(WIDTH)) large_mux_instance11101(.data_in(wire_d10_0),.data_out(wire_d10_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance11102(.data_in(wire_d10_1),.data_out(wire_d10_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance11103(.data_in(wire_d10_2),.data_out(wire_d10_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance11104(.data_in(wire_d10_3),.data_out(wire_d10_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance11105(.data_in(wire_d10_4),.data_out(wire_d10_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance11106(.data_in(wire_d10_5),.data_out(wire_d10_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance11107(.data_in(wire_d10_6),.data_out(wire_d10_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance11108(.data_in(wire_d10_7),.data_out(wire_d10_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance11109(.data_in(wire_d10_8),.data_out(wire_d10_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111010(.data_in(wire_d10_9),.data_out(wire_d10_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111011(.data_in(wire_d10_10),.data_out(wire_d10_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111012(.data_in(wire_d10_11),.data_out(wire_d10_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111013(.data_in(wire_d10_12),.data_out(wire_d10_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111014(.data_in(wire_d10_13),.data_out(wire_d10_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111015(.data_in(wire_d10_14),.data_out(wire_d10_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111016(.data_in(wire_d10_15),.data_out(wire_d10_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111017(.data_in(wire_d10_16),.data_out(wire_d10_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111018(.data_in(wire_d10_17),.data_out(wire_d10_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111019(.data_in(wire_d10_18),.data_out(wire_d10_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111020(.data_in(wire_d10_19),.data_out(wire_d10_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111021(.data_in(wire_d10_20),.data_out(wire_d10_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111022(.data_in(wire_d10_21),.data_out(wire_d10_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111023(.data_in(wire_d10_22),.data_out(wire_d10_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111024(.data_in(wire_d10_23),.data_out(wire_d10_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111025(.data_in(wire_d10_24),.data_out(wire_d10_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111026(.data_in(wire_d10_25),.data_out(wire_d10_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111027(.data_in(wire_d10_26),.data_out(wire_d10_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111028(.data_in(wire_d10_27),.data_out(wire_d10_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111029(.data_in(wire_d10_28),.data_out(wire_d10_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111030(.data_in(wire_d10_29),.data_out(wire_d10_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111031(.data_in(wire_d10_30),.data_out(wire_d10_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111032(.data_in(wire_d10_31),.data_out(wire_d10_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111033(.data_in(wire_d10_32),.data_out(wire_d10_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111034(.data_in(wire_d10_33),.data_out(wire_d10_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111035(.data_in(wire_d10_34),.data_out(wire_d10_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111036(.data_in(wire_d10_35),.data_out(wire_d10_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111037(.data_in(wire_d10_36),.data_out(wire_d10_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111038(.data_in(wire_d10_37),.data_out(wire_d10_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111039(.data_in(wire_d10_38),.data_out(wire_d10_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111040(.data_in(wire_d10_39),.data_out(wire_d10_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111041(.data_in(wire_d10_40),.data_out(wire_d10_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111042(.data_in(wire_d10_41),.data_out(wire_d10_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111043(.data_in(wire_d10_42),.data_out(wire_d10_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111044(.data_in(wire_d10_43),.data_out(wire_d10_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111045(.data_in(wire_d10_44),.data_out(wire_d10_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance111046(.data_in(wire_d10_45),.data_out(wire_d10_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance111047(.data_in(wire_d10_46),.data_out(wire_d10_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance111048(.data_in(wire_d10_47),.data_out(wire_d10_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance111049(.data_in(wire_d10_48),.data_out(d_out10),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance12110(.data_in(d_in11),.data_out(wire_d11_0),.clk(clk),.rst(rst));            //channel 12
	invertion #(.WIDTH(WIDTH)) invertion_instance12111(.data_in(wire_d11_0),.data_out(wire_d11_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance12112(.data_in(wire_d11_1),.data_out(wire_d11_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance12113(.data_in(wire_d11_2),.data_out(wire_d11_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance12114(.data_in(wire_d11_3),.data_out(wire_d11_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance12115(.data_in(wire_d11_4),.data_out(wire_d11_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance12116(.data_in(wire_d11_5),.data_out(wire_d11_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance12117(.data_in(wire_d11_6),.data_out(wire_d11_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance12118(.data_in(wire_d11_7),.data_out(wire_d11_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance12119(.data_in(wire_d11_8),.data_out(wire_d11_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121110(.data_in(wire_d11_9),.data_out(wire_d11_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121111(.data_in(wire_d11_10),.data_out(wire_d11_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121112(.data_in(wire_d11_11),.data_out(wire_d11_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121113(.data_in(wire_d11_12),.data_out(wire_d11_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121114(.data_in(wire_d11_13),.data_out(wire_d11_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121115(.data_in(wire_d11_14),.data_out(wire_d11_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121116(.data_in(wire_d11_15),.data_out(wire_d11_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121117(.data_in(wire_d11_16),.data_out(wire_d11_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121118(.data_in(wire_d11_17),.data_out(wire_d11_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121119(.data_in(wire_d11_18),.data_out(wire_d11_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121120(.data_in(wire_d11_19),.data_out(wire_d11_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121121(.data_in(wire_d11_20),.data_out(wire_d11_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121122(.data_in(wire_d11_21),.data_out(wire_d11_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121123(.data_in(wire_d11_22),.data_out(wire_d11_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121124(.data_in(wire_d11_23),.data_out(wire_d11_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121125(.data_in(wire_d11_24),.data_out(wire_d11_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121126(.data_in(wire_d11_25),.data_out(wire_d11_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121127(.data_in(wire_d11_26),.data_out(wire_d11_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121128(.data_in(wire_d11_27),.data_out(wire_d11_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121129(.data_in(wire_d11_28),.data_out(wire_d11_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121130(.data_in(wire_d11_29),.data_out(wire_d11_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121131(.data_in(wire_d11_30),.data_out(wire_d11_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121132(.data_in(wire_d11_31),.data_out(wire_d11_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121133(.data_in(wire_d11_32),.data_out(wire_d11_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121134(.data_in(wire_d11_33),.data_out(wire_d11_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121135(.data_in(wire_d11_34),.data_out(wire_d11_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121136(.data_in(wire_d11_35),.data_out(wire_d11_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121137(.data_in(wire_d11_36),.data_out(wire_d11_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121138(.data_in(wire_d11_37),.data_out(wire_d11_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121139(.data_in(wire_d11_38),.data_out(wire_d11_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121140(.data_in(wire_d11_39),.data_out(wire_d11_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121141(.data_in(wire_d11_40),.data_out(wire_d11_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121142(.data_in(wire_d11_41),.data_out(wire_d11_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121143(.data_in(wire_d11_42),.data_out(wire_d11_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121144(.data_in(wire_d11_43),.data_out(wire_d11_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121145(.data_in(wire_d11_44),.data_out(wire_d11_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance121146(.data_in(wire_d11_45),.data_out(wire_d11_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance121147(.data_in(wire_d11_46),.data_out(wire_d11_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance121148(.data_in(wire_d11_47),.data_out(wire_d11_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance121149(.data_in(wire_d11_48),.data_out(d_out11),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance13120(.data_in(d_in12),.data_out(wire_d12_0),.clk(clk),.rst(rst));            //channel 13
	large_mux #(.WIDTH(WIDTH)) large_mux_instance13121(.data_in(wire_d12_0),.data_out(wire_d12_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance13122(.data_in(wire_d12_1),.data_out(wire_d12_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance13123(.data_in(wire_d12_2),.data_out(wire_d12_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance13124(.data_in(wire_d12_3),.data_out(wire_d12_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance13125(.data_in(wire_d12_4),.data_out(wire_d12_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance13126(.data_in(wire_d12_5),.data_out(wire_d12_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance13127(.data_in(wire_d12_6),.data_out(wire_d12_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance13128(.data_in(wire_d12_7),.data_out(wire_d12_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance13129(.data_in(wire_d12_8),.data_out(wire_d12_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131210(.data_in(wire_d12_9),.data_out(wire_d12_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131211(.data_in(wire_d12_10),.data_out(wire_d12_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131212(.data_in(wire_d12_11),.data_out(wire_d12_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131213(.data_in(wire_d12_12),.data_out(wire_d12_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131214(.data_in(wire_d12_13),.data_out(wire_d12_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131215(.data_in(wire_d12_14),.data_out(wire_d12_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131216(.data_in(wire_d12_15),.data_out(wire_d12_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131217(.data_in(wire_d12_16),.data_out(wire_d12_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131218(.data_in(wire_d12_17),.data_out(wire_d12_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131219(.data_in(wire_d12_18),.data_out(wire_d12_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131220(.data_in(wire_d12_19),.data_out(wire_d12_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131221(.data_in(wire_d12_20),.data_out(wire_d12_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131222(.data_in(wire_d12_21),.data_out(wire_d12_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131223(.data_in(wire_d12_22),.data_out(wire_d12_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131224(.data_in(wire_d12_23),.data_out(wire_d12_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131225(.data_in(wire_d12_24),.data_out(wire_d12_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131226(.data_in(wire_d12_25),.data_out(wire_d12_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131227(.data_in(wire_d12_26),.data_out(wire_d12_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131228(.data_in(wire_d12_27),.data_out(wire_d12_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131229(.data_in(wire_d12_28),.data_out(wire_d12_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131230(.data_in(wire_d12_29),.data_out(wire_d12_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131231(.data_in(wire_d12_30),.data_out(wire_d12_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131232(.data_in(wire_d12_31),.data_out(wire_d12_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131233(.data_in(wire_d12_32),.data_out(wire_d12_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131234(.data_in(wire_d12_33),.data_out(wire_d12_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131235(.data_in(wire_d12_34),.data_out(wire_d12_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131236(.data_in(wire_d12_35),.data_out(wire_d12_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131237(.data_in(wire_d12_36),.data_out(wire_d12_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131238(.data_in(wire_d12_37),.data_out(wire_d12_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131239(.data_in(wire_d12_38),.data_out(wire_d12_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131240(.data_in(wire_d12_39),.data_out(wire_d12_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131241(.data_in(wire_d12_40),.data_out(wire_d12_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131242(.data_in(wire_d12_41),.data_out(wire_d12_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131243(.data_in(wire_d12_42),.data_out(wire_d12_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131244(.data_in(wire_d12_43),.data_out(wire_d12_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131245(.data_in(wire_d12_44),.data_out(wire_d12_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance131246(.data_in(wire_d12_45),.data_out(wire_d12_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance131247(.data_in(wire_d12_46),.data_out(wire_d12_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance131248(.data_in(wire_d12_47),.data_out(wire_d12_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance131249(.data_in(wire_d12_48),.data_out(d_out12),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance14130(.data_in(d_in13),.data_out(wire_d13_0),.clk(clk),.rst(rst));            //channel 14
	encoder #(.WIDTH(WIDTH)) encoder_instance14131(.data_in(wire_d13_0),.data_out(wire_d13_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance14132(.data_in(wire_d13_1),.data_out(wire_d13_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance14133(.data_in(wire_d13_2),.data_out(wire_d13_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance14134(.data_in(wire_d13_3),.data_out(wire_d13_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance14135(.data_in(wire_d13_4),.data_out(wire_d13_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance14136(.data_in(wire_d13_5),.data_out(wire_d13_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance14137(.data_in(wire_d13_6),.data_out(wire_d13_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance14138(.data_in(wire_d13_7),.data_out(wire_d13_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance14139(.data_in(wire_d13_8),.data_out(wire_d13_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141310(.data_in(wire_d13_9),.data_out(wire_d13_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141311(.data_in(wire_d13_10),.data_out(wire_d13_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141312(.data_in(wire_d13_11),.data_out(wire_d13_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141313(.data_in(wire_d13_12),.data_out(wire_d13_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141314(.data_in(wire_d13_13),.data_out(wire_d13_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141315(.data_in(wire_d13_14),.data_out(wire_d13_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141316(.data_in(wire_d13_15),.data_out(wire_d13_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141317(.data_in(wire_d13_16),.data_out(wire_d13_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141318(.data_in(wire_d13_17),.data_out(wire_d13_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141319(.data_in(wire_d13_18),.data_out(wire_d13_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141320(.data_in(wire_d13_19),.data_out(wire_d13_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141321(.data_in(wire_d13_20),.data_out(wire_d13_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141322(.data_in(wire_d13_21),.data_out(wire_d13_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141323(.data_in(wire_d13_22),.data_out(wire_d13_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141324(.data_in(wire_d13_23),.data_out(wire_d13_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141325(.data_in(wire_d13_24),.data_out(wire_d13_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141326(.data_in(wire_d13_25),.data_out(wire_d13_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141327(.data_in(wire_d13_26),.data_out(wire_d13_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141328(.data_in(wire_d13_27),.data_out(wire_d13_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141329(.data_in(wire_d13_28),.data_out(wire_d13_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141330(.data_in(wire_d13_29),.data_out(wire_d13_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141331(.data_in(wire_d13_30),.data_out(wire_d13_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141332(.data_in(wire_d13_31),.data_out(wire_d13_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141333(.data_in(wire_d13_32),.data_out(wire_d13_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141334(.data_in(wire_d13_33),.data_out(wire_d13_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141335(.data_in(wire_d13_34),.data_out(wire_d13_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141336(.data_in(wire_d13_35),.data_out(wire_d13_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141337(.data_in(wire_d13_36),.data_out(wire_d13_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141338(.data_in(wire_d13_37),.data_out(wire_d13_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141339(.data_in(wire_d13_38),.data_out(wire_d13_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141340(.data_in(wire_d13_39),.data_out(wire_d13_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance141341(.data_in(wire_d13_40),.data_out(wire_d13_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141342(.data_in(wire_d13_41),.data_out(wire_d13_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141343(.data_in(wire_d13_42),.data_out(wire_d13_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141344(.data_in(wire_d13_43),.data_out(wire_d13_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141345(.data_in(wire_d13_44),.data_out(wire_d13_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141346(.data_in(wire_d13_45),.data_out(wire_d13_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance141347(.data_in(wire_d13_46),.data_out(wire_d13_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance141348(.data_in(wire_d13_47),.data_out(wire_d13_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance141349(.data_in(wire_d13_48),.data_out(d_out13),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance15140(.data_in(d_in14),.data_out(wire_d14_0),.clk(clk),.rst(rst));            //channel 15
	invertion #(.WIDTH(WIDTH)) invertion_instance15141(.data_in(wire_d14_0),.data_out(wire_d14_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance15142(.data_in(wire_d14_1),.data_out(wire_d14_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance15143(.data_in(wire_d14_2),.data_out(wire_d14_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance15144(.data_in(wire_d14_3),.data_out(wire_d14_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance15145(.data_in(wire_d14_4),.data_out(wire_d14_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance15146(.data_in(wire_d14_5),.data_out(wire_d14_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance15147(.data_in(wire_d14_6),.data_out(wire_d14_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance15148(.data_in(wire_d14_7),.data_out(wire_d14_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance15149(.data_in(wire_d14_8),.data_out(wire_d14_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151410(.data_in(wire_d14_9),.data_out(wire_d14_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151411(.data_in(wire_d14_10),.data_out(wire_d14_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151412(.data_in(wire_d14_11),.data_out(wire_d14_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151413(.data_in(wire_d14_12),.data_out(wire_d14_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151414(.data_in(wire_d14_13),.data_out(wire_d14_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151415(.data_in(wire_d14_14),.data_out(wire_d14_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151416(.data_in(wire_d14_15),.data_out(wire_d14_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151417(.data_in(wire_d14_16),.data_out(wire_d14_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151418(.data_in(wire_d14_17),.data_out(wire_d14_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151419(.data_in(wire_d14_18),.data_out(wire_d14_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151420(.data_in(wire_d14_19),.data_out(wire_d14_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151421(.data_in(wire_d14_20),.data_out(wire_d14_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151422(.data_in(wire_d14_21),.data_out(wire_d14_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151423(.data_in(wire_d14_22),.data_out(wire_d14_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151424(.data_in(wire_d14_23),.data_out(wire_d14_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151425(.data_in(wire_d14_24),.data_out(wire_d14_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151426(.data_in(wire_d14_25),.data_out(wire_d14_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151427(.data_in(wire_d14_26),.data_out(wire_d14_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151428(.data_in(wire_d14_27),.data_out(wire_d14_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151429(.data_in(wire_d14_28),.data_out(wire_d14_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151430(.data_in(wire_d14_29),.data_out(wire_d14_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151431(.data_in(wire_d14_30),.data_out(wire_d14_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151432(.data_in(wire_d14_31),.data_out(wire_d14_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151433(.data_in(wire_d14_32),.data_out(wire_d14_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151434(.data_in(wire_d14_33),.data_out(wire_d14_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151435(.data_in(wire_d14_34),.data_out(wire_d14_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151436(.data_in(wire_d14_35),.data_out(wire_d14_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151437(.data_in(wire_d14_36),.data_out(wire_d14_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151438(.data_in(wire_d14_37),.data_out(wire_d14_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151439(.data_in(wire_d14_38),.data_out(wire_d14_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151440(.data_in(wire_d14_39),.data_out(wire_d14_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151441(.data_in(wire_d14_40),.data_out(wire_d14_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151442(.data_in(wire_d14_41),.data_out(wire_d14_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151443(.data_in(wire_d14_42),.data_out(wire_d14_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151444(.data_in(wire_d14_43),.data_out(wire_d14_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance151445(.data_in(wire_d14_44),.data_out(wire_d14_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151446(.data_in(wire_d14_45),.data_out(wire_d14_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance151447(.data_in(wire_d14_46),.data_out(wire_d14_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance151448(.data_in(wire_d14_47),.data_out(wire_d14_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance151449(.data_in(wire_d14_48),.data_out(d_out14),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance16150(.data_in(d_in15),.data_out(wire_d15_0),.clk(clk),.rst(rst));            //channel 16
	large_mux #(.WIDTH(WIDTH)) large_mux_instance16151(.data_in(wire_d15_0),.data_out(wire_d15_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance16152(.data_in(wire_d15_1),.data_out(wire_d15_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance16153(.data_in(wire_d15_2),.data_out(wire_d15_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance16154(.data_in(wire_d15_3),.data_out(wire_d15_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance16155(.data_in(wire_d15_4),.data_out(wire_d15_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance16156(.data_in(wire_d15_5),.data_out(wire_d15_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance16157(.data_in(wire_d15_6),.data_out(wire_d15_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance16158(.data_in(wire_d15_7),.data_out(wire_d15_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance16159(.data_in(wire_d15_8),.data_out(wire_d15_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161510(.data_in(wire_d15_9),.data_out(wire_d15_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161511(.data_in(wire_d15_10),.data_out(wire_d15_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161512(.data_in(wire_d15_11),.data_out(wire_d15_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161513(.data_in(wire_d15_12),.data_out(wire_d15_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161514(.data_in(wire_d15_13),.data_out(wire_d15_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161515(.data_in(wire_d15_14),.data_out(wire_d15_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161516(.data_in(wire_d15_15),.data_out(wire_d15_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161517(.data_in(wire_d15_16),.data_out(wire_d15_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161518(.data_in(wire_d15_17),.data_out(wire_d15_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161519(.data_in(wire_d15_18),.data_out(wire_d15_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161520(.data_in(wire_d15_19),.data_out(wire_d15_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161521(.data_in(wire_d15_20),.data_out(wire_d15_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161522(.data_in(wire_d15_21),.data_out(wire_d15_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161523(.data_in(wire_d15_22),.data_out(wire_d15_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161524(.data_in(wire_d15_23),.data_out(wire_d15_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161525(.data_in(wire_d15_24),.data_out(wire_d15_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161526(.data_in(wire_d15_25),.data_out(wire_d15_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161527(.data_in(wire_d15_26),.data_out(wire_d15_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161528(.data_in(wire_d15_27),.data_out(wire_d15_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161529(.data_in(wire_d15_28),.data_out(wire_d15_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161530(.data_in(wire_d15_29),.data_out(wire_d15_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161531(.data_in(wire_d15_30),.data_out(wire_d15_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161532(.data_in(wire_d15_31),.data_out(wire_d15_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161533(.data_in(wire_d15_32),.data_out(wire_d15_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161534(.data_in(wire_d15_33),.data_out(wire_d15_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161535(.data_in(wire_d15_34),.data_out(wire_d15_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161536(.data_in(wire_d15_35),.data_out(wire_d15_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161537(.data_in(wire_d15_36),.data_out(wire_d15_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161538(.data_in(wire_d15_37),.data_out(wire_d15_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance161539(.data_in(wire_d15_38),.data_out(wire_d15_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161540(.data_in(wire_d15_39),.data_out(wire_d15_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161541(.data_in(wire_d15_40),.data_out(wire_d15_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161542(.data_in(wire_d15_41),.data_out(wire_d15_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161543(.data_in(wire_d15_42),.data_out(wire_d15_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161544(.data_in(wire_d15_43),.data_out(wire_d15_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance161545(.data_in(wire_d15_44),.data_out(wire_d15_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161546(.data_in(wire_d15_45),.data_out(wire_d15_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161547(.data_in(wire_d15_46),.data_out(wire_d15_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance161548(.data_in(wire_d15_47),.data_out(wire_d15_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance161549(.data_in(wire_d15_48),.data_out(d_out15),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance17160(.data_in(d_in16),.data_out(wire_d16_0),.clk(clk),.rst(rst));            //channel 17
	encoder #(.WIDTH(WIDTH)) encoder_instance17161(.data_in(wire_d16_0),.data_out(wire_d16_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance17162(.data_in(wire_d16_1),.data_out(wire_d16_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance17163(.data_in(wire_d16_2),.data_out(wire_d16_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance17164(.data_in(wire_d16_3),.data_out(wire_d16_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance17165(.data_in(wire_d16_4),.data_out(wire_d16_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance17166(.data_in(wire_d16_5),.data_out(wire_d16_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance17167(.data_in(wire_d16_6),.data_out(wire_d16_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance17168(.data_in(wire_d16_7),.data_out(wire_d16_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance17169(.data_in(wire_d16_8),.data_out(wire_d16_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171610(.data_in(wire_d16_9),.data_out(wire_d16_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171611(.data_in(wire_d16_10),.data_out(wire_d16_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171612(.data_in(wire_d16_11),.data_out(wire_d16_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171613(.data_in(wire_d16_12),.data_out(wire_d16_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171614(.data_in(wire_d16_13),.data_out(wire_d16_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171615(.data_in(wire_d16_14),.data_out(wire_d16_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171616(.data_in(wire_d16_15),.data_out(wire_d16_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171617(.data_in(wire_d16_16),.data_out(wire_d16_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171618(.data_in(wire_d16_17),.data_out(wire_d16_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171619(.data_in(wire_d16_18),.data_out(wire_d16_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171620(.data_in(wire_d16_19),.data_out(wire_d16_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171621(.data_in(wire_d16_20),.data_out(wire_d16_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171622(.data_in(wire_d16_21),.data_out(wire_d16_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171623(.data_in(wire_d16_22),.data_out(wire_d16_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171624(.data_in(wire_d16_23),.data_out(wire_d16_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171625(.data_in(wire_d16_24),.data_out(wire_d16_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171626(.data_in(wire_d16_25),.data_out(wire_d16_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171627(.data_in(wire_d16_26),.data_out(wire_d16_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171628(.data_in(wire_d16_27),.data_out(wire_d16_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171629(.data_in(wire_d16_28),.data_out(wire_d16_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171630(.data_in(wire_d16_29),.data_out(wire_d16_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171631(.data_in(wire_d16_30),.data_out(wire_d16_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171632(.data_in(wire_d16_31),.data_out(wire_d16_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171633(.data_in(wire_d16_32),.data_out(wire_d16_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171634(.data_in(wire_d16_33),.data_out(wire_d16_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171635(.data_in(wire_d16_34),.data_out(wire_d16_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171636(.data_in(wire_d16_35),.data_out(wire_d16_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171637(.data_in(wire_d16_36),.data_out(wire_d16_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171638(.data_in(wire_d16_37),.data_out(wire_d16_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance171639(.data_in(wire_d16_38),.data_out(wire_d16_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171640(.data_in(wire_d16_39),.data_out(wire_d16_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171641(.data_in(wire_d16_40),.data_out(wire_d16_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171642(.data_in(wire_d16_41),.data_out(wire_d16_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171643(.data_in(wire_d16_42),.data_out(wire_d16_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171644(.data_in(wire_d16_43),.data_out(wire_d16_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171645(.data_in(wire_d16_44),.data_out(wire_d16_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171646(.data_in(wire_d16_45),.data_out(wire_d16_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance171647(.data_in(wire_d16_46),.data_out(wire_d16_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance171648(.data_in(wire_d16_47),.data_out(wire_d16_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance171649(.data_in(wire_d16_48),.data_out(d_out16),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance18170(.data_in(d_in17),.data_out(wire_d17_0),.clk(clk),.rst(rst));            //channel 18
	register #(.WIDTH(WIDTH)) register_instance18171(.data_in(wire_d17_0),.data_out(wire_d17_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance18172(.data_in(wire_d17_1),.data_out(wire_d17_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance18173(.data_in(wire_d17_2),.data_out(wire_d17_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance18174(.data_in(wire_d17_3),.data_out(wire_d17_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance18175(.data_in(wire_d17_4),.data_out(wire_d17_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance18176(.data_in(wire_d17_5),.data_out(wire_d17_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance18177(.data_in(wire_d17_6),.data_out(wire_d17_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance18178(.data_in(wire_d17_7),.data_out(wire_d17_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance18179(.data_in(wire_d17_8),.data_out(wire_d17_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181710(.data_in(wire_d17_9),.data_out(wire_d17_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181711(.data_in(wire_d17_10),.data_out(wire_d17_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181712(.data_in(wire_d17_11),.data_out(wire_d17_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181713(.data_in(wire_d17_12),.data_out(wire_d17_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181714(.data_in(wire_d17_13),.data_out(wire_d17_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181715(.data_in(wire_d17_14),.data_out(wire_d17_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181716(.data_in(wire_d17_15),.data_out(wire_d17_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181717(.data_in(wire_d17_16),.data_out(wire_d17_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181718(.data_in(wire_d17_17),.data_out(wire_d17_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181719(.data_in(wire_d17_18),.data_out(wire_d17_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181720(.data_in(wire_d17_19),.data_out(wire_d17_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181721(.data_in(wire_d17_20),.data_out(wire_d17_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181722(.data_in(wire_d17_21),.data_out(wire_d17_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181723(.data_in(wire_d17_22),.data_out(wire_d17_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181724(.data_in(wire_d17_23),.data_out(wire_d17_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181725(.data_in(wire_d17_24),.data_out(wire_d17_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181726(.data_in(wire_d17_25),.data_out(wire_d17_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181727(.data_in(wire_d17_26),.data_out(wire_d17_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181728(.data_in(wire_d17_27),.data_out(wire_d17_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181729(.data_in(wire_d17_28),.data_out(wire_d17_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181730(.data_in(wire_d17_29),.data_out(wire_d17_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181731(.data_in(wire_d17_30),.data_out(wire_d17_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181732(.data_in(wire_d17_31),.data_out(wire_d17_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181733(.data_in(wire_d17_32),.data_out(wire_d17_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181734(.data_in(wire_d17_33),.data_out(wire_d17_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181735(.data_in(wire_d17_34),.data_out(wire_d17_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181736(.data_in(wire_d17_35),.data_out(wire_d17_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181737(.data_in(wire_d17_36),.data_out(wire_d17_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181738(.data_in(wire_d17_37),.data_out(wire_d17_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181739(.data_in(wire_d17_38),.data_out(wire_d17_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance181740(.data_in(wire_d17_39),.data_out(wire_d17_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181741(.data_in(wire_d17_40),.data_out(wire_d17_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181742(.data_in(wire_d17_41),.data_out(wire_d17_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181743(.data_in(wire_d17_42),.data_out(wire_d17_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance181744(.data_in(wire_d17_43),.data_out(wire_d17_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181745(.data_in(wire_d17_44),.data_out(wire_d17_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181746(.data_in(wire_d17_45),.data_out(wire_d17_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181747(.data_in(wire_d17_46),.data_out(wire_d17_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance181748(.data_in(wire_d17_47),.data_out(wire_d17_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance181749(.data_in(wire_d17_48),.data_out(d_out17),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance19180(.data_in(d_in18),.data_out(wire_d18_0),.clk(clk),.rst(rst));            //channel 19
	large_mux #(.WIDTH(WIDTH)) large_mux_instance19181(.data_in(wire_d18_0),.data_out(wire_d18_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance19182(.data_in(wire_d18_1),.data_out(wire_d18_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance19183(.data_in(wire_d18_2),.data_out(wire_d18_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance19184(.data_in(wire_d18_3),.data_out(wire_d18_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance19185(.data_in(wire_d18_4),.data_out(wire_d18_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance19186(.data_in(wire_d18_5),.data_out(wire_d18_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance19187(.data_in(wire_d18_6),.data_out(wire_d18_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance19188(.data_in(wire_d18_7),.data_out(wire_d18_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance19189(.data_in(wire_d18_8),.data_out(wire_d18_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191810(.data_in(wire_d18_9),.data_out(wire_d18_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191811(.data_in(wire_d18_10),.data_out(wire_d18_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191812(.data_in(wire_d18_11),.data_out(wire_d18_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191813(.data_in(wire_d18_12),.data_out(wire_d18_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191814(.data_in(wire_d18_13),.data_out(wire_d18_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191815(.data_in(wire_d18_14),.data_out(wire_d18_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191816(.data_in(wire_d18_15),.data_out(wire_d18_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191817(.data_in(wire_d18_16),.data_out(wire_d18_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191818(.data_in(wire_d18_17),.data_out(wire_d18_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191819(.data_in(wire_d18_18),.data_out(wire_d18_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191820(.data_in(wire_d18_19),.data_out(wire_d18_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191821(.data_in(wire_d18_20),.data_out(wire_d18_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191822(.data_in(wire_d18_21),.data_out(wire_d18_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191823(.data_in(wire_d18_22),.data_out(wire_d18_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191824(.data_in(wire_d18_23),.data_out(wire_d18_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191825(.data_in(wire_d18_24),.data_out(wire_d18_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191826(.data_in(wire_d18_25),.data_out(wire_d18_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191827(.data_in(wire_d18_26),.data_out(wire_d18_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191828(.data_in(wire_d18_27),.data_out(wire_d18_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191829(.data_in(wire_d18_28),.data_out(wire_d18_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191830(.data_in(wire_d18_29),.data_out(wire_d18_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191831(.data_in(wire_d18_30),.data_out(wire_d18_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191832(.data_in(wire_d18_31),.data_out(wire_d18_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191833(.data_in(wire_d18_32),.data_out(wire_d18_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191834(.data_in(wire_d18_33),.data_out(wire_d18_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191835(.data_in(wire_d18_34),.data_out(wire_d18_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191836(.data_in(wire_d18_35),.data_out(wire_d18_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191837(.data_in(wire_d18_36),.data_out(wire_d18_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191838(.data_in(wire_d18_37),.data_out(wire_d18_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191839(.data_in(wire_d18_38),.data_out(wire_d18_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191840(.data_in(wire_d18_39),.data_out(wire_d18_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191841(.data_in(wire_d18_40),.data_out(wire_d18_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191842(.data_in(wire_d18_41),.data_out(wire_d18_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191843(.data_in(wire_d18_42),.data_out(wire_d18_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance191844(.data_in(wire_d18_43),.data_out(wire_d18_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance191845(.data_in(wire_d18_44),.data_out(wire_d18_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191846(.data_in(wire_d18_45),.data_out(wire_d18_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191847(.data_in(wire_d18_46),.data_out(wire_d18_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance191848(.data_in(wire_d18_47),.data_out(wire_d18_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance191849(.data_in(wire_d18_48),.data_out(d_out18),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance20190(.data_in(d_in19),.data_out(wire_d19_0),.clk(clk),.rst(rst));            //channel 20
	register #(.WIDTH(WIDTH)) register_instance20191(.data_in(wire_d19_0),.data_out(wire_d19_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance20192(.data_in(wire_d19_1),.data_out(wire_d19_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance20193(.data_in(wire_d19_2),.data_out(wire_d19_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance20194(.data_in(wire_d19_3),.data_out(wire_d19_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance20195(.data_in(wire_d19_4),.data_out(wire_d19_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance20196(.data_in(wire_d19_5),.data_out(wire_d19_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance20197(.data_in(wire_d19_6),.data_out(wire_d19_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance20198(.data_in(wire_d19_7),.data_out(wire_d19_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance20199(.data_in(wire_d19_8),.data_out(wire_d19_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201910(.data_in(wire_d19_9),.data_out(wire_d19_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201911(.data_in(wire_d19_10),.data_out(wire_d19_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201912(.data_in(wire_d19_11),.data_out(wire_d19_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201913(.data_in(wire_d19_12),.data_out(wire_d19_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201914(.data_in(wire_d19_13),.data_out(wire_d19_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201915(.data_in(wire_d19_14),.data_out(wire_d19_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201916(.data_in(wire_d19_15),.data_out(wire_d19_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201917(.data_in(wire_d19_16),.data_out(wire_d19_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201918(.data_in(wire_d19_17),.data_out(wire_d19_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201919(.data_in(wire_d19_18),.data_out(wire_d19_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201920(.data_in(wire_d19_19),.data_out(wire_d19_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201921(.data_in(wire_d19_20),.data_out(wire_d19_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201922(.data_in(wire_d19_21),.data_out(wire_d19_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201923(.data_in(wire_d19_22),.data_out(wire_d19_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201924(.data_in(wire_d19_23),.data_out(wire_d19_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201925(.data_in(wire_d19_24),.data_out(wire_d19_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201926(.data_in(wire_d19_25),.data_out(wire_d19_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201927(.data_in(wire_d19_26),.data_out(wire_d19_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201928(.data_in(wire_d19_27),.data_out(wire_d19_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201929(.data_in(wire_d19_28),.data_out(wire_d19_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201930(.data_in(wire_d19_29),.data_out(wire_d19_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201931(.data_in(wire_d19_30),.data_out(wire_d19_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201932(.data_in(wire_d19_31),.data_out(wire_d19_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201933(.data_in(wire_d19_32),.data_out(wire_d19_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201934(.data_in(wire_d19_33),.data_out(wire_d19_34),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201935(.data_in(wire_d19_34),.data_out(wire_d19_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201936(.data_in(wire_d19_35),.data_out(wire_d19_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201937(.data_in(wire_d19_36),.data_out(wire_d19_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201938(.data_in(wire_d19_37),.data_out(wire_d19_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201939(.data_in(wire_d19_38),.data_out(wire_d19_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201940(.data_in(wire_d19_39),.data_out(wire_d19_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201941(.data_in(wire_d19_40),.data_out(wire_d19_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201942(.data_in(wire_d19_41),.data_out(wire_d19_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201943(.data_in(wire_d19_42),.data_out(wire_d19_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201944(.data_in(wire_d19_43),.data_out(wire_d19_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201945(.data_in(wire_d19_44),.data_out(wire_d19_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance201946(.data_in(wire_d19_45),.data_out(wire_d19_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance201947(.data_in(wire_d19_46),.data_out(wire_d19_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance201948(.data_in(wire_d19_47),.data_out(wire_d19_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance201949(.data_in(wire_d19_48),.data_out(d_out19),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance21200(.data_in(d_in20),.data_out(wire_d20_0),.clk(clk),.rst(rst));            //channel 21
	register #(.WIDTH(WIDTH)) register_instance21201(.data_in(wire_d20_0),.data_out(wire_d20_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance21202(.data_in(wire_d20_1),.data_out(wire_d20_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance21203(.data_in(wire_d20_2),.data_out(wire_d20_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance21204(.data_in(wire_d20_3),.data_out(wire_d20_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance21205(.data_in(wire_d20_4),.data_out(wire_d20_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance21206(.data_in(wire_d20_5),.data_out(wire_d20_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance21207(.data_in(wire_d20_6),.data_out(wire_d20_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance21208(.data_in(wire_d20_7),.data_out(wire_d20_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance21209(.data_in(wire_d20_8),.data_out(wire_d20_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212010(.data_in(wire_d20_9),.data_out(wire_d20_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212011(.data_in(wire_d20_10),.data_out(wire_d20_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212012(.data_in(wire_d20_11),.data_out(wire_d20_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212013(.data_in(wire_d20_12),.data_out(wire_d20_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212014(.data_in(wire_d20_13),.data_out(wire_d20_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212015(.data_in(wire_d20_14),.data_out(wire_d20_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212016(.data_in(wire_d20_15),.data_out(wire_d20_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212017(.data_in(wire_d20_16),.data_out(wire_d20_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212018(.data_in(wire_d20_17),.data_out(wire_d20_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212019(.data_in(wire_d20_18),.data_out(wire_d20_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212020(.data_in(wire_d20_19),.data_out(wire_d20_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212021(.data_in(wire_d20_20),.data_out(wire_d20_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212022(.data_in(wire_d20_21),.data_out(wire_d20_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212023(.data_in(wire_d20_22),.data_out(wire_d20_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212024(.data_in(wire_d20_23),.data_out(wire_d20_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212025(.data_in(wire_d20_24),.data_out(wire_d20_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212026(.data_in(wire_d20_25),.data_out(wire_d20_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212027(.data_in(wire_d20_26),.data_out(wire_d20_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212028(.data_in(wire_d20_27),.data_out(wire_d20_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212029(.data_in(wire_d20_28),.data_out(wire_d20_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212030(.data_in(wire_d20_29),.data_out(wire_d20_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212031(.data_in(wire_d20_30),.data_out(wire_d20_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212032(.data_in(wire_d20_31),.data_out(wire_d20_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212033(.data_in(wire_d20_32),.data_out(wire_d20_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212034(.data_in(wire_d20_33),.data_out(wire_d20_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212035(.data_in(wire_d20_34),.data_out(wire_d20_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212036(.data_in(wire_d20_35),.data_out(wire_d20_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212037(.data_in(wire_d20_36),.data_out(wire_d20_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212038(.data_in(wire_d20_37),.data_out(wire_d20_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212039(.data_in(wire_d20_38),.data_out(wire_d20_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212040(.data_in(wire_d20_39),.data_out(wire_d20_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212041(.data_in(wire_d20_40),.data_out(wire_d20_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212042(.data_in(wire_d20_41),.data_out(wire_d20_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212043(.data_in(wire_d20_42),.data_out(wire_d20_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212044(.data_in(wire_d20_43),.data_out(wire_d20_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212045(.data_in(wire_d20_44),.data_out(wire_d20_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance212046(.data_in(wire_d20_45),.data_out(wire_d20_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance212047(.data_in(wire_d20_46),.data_out(wire_d20_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212048(.data_in(wire_d20_47),.data_out(wire_d20_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance212049(.data_in(wire_d20_48),.data_out(d_out20),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance22210(.data_in(d_in21),.data_out(wire_d21_0),.clk(clk),.rst(rst));            //channel 22
	register #(.WIDTH(WIDTH)) register_instance22211(.data_in(wire_d21_0),.data_out(wire_d21_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance22212(.data_in(wire_d21_1),.data_out(wire_d21_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance22213(.data_in(wire_d21_2),.data_out(wire_d21_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance22214(.data_in(wire_d21_3),.data_out(wire_d21_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance22215(.data_in(wire_d21_4),.data_out(wire_d21_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance22216(.data_in(wire_d21_5),.data_out(wire_d21_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance22217(.data_in(wire_d21_6),.data_out(wire_d21_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance22218(.data_in(wire_d21_7),.data_out(wire_d21_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance22219(.data_in(wire_d21_8),.data_out(wire_d21_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222110(.data_in(wire_d21_9),.data_out(wire_d21_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222111(.data_in(wire_d21_10),.data_out(wire_d21_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222112(.data_in(wire_d21_11),.data_out(wire_d21_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222113(.data_in(wire_d21_12),.data_out(wire_d21_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222114(.data_in(wire_d21_13),.data_out(wire_d21_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222115(.data_in(wire_d21_14),.data_out(wire_d21_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222116(.data_in(wire_d21_15),.data_out(wire_d21_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222117(.data_in(wire_d21_16),.data_out(wire_d21_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222118(.data_in(wire_d21_17),.data_out(wire_d21_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222119(.data_in(wire_d21_18),.data_out(wire_d21_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222120(.data_in(wire_d21_19),.data_out(wire_d21_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222121(.data_in(wire_d21_20),.data_out(wire_d21_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222122(.data_in(wire_d21_21),.data_out(wire_d21_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222123(.data_in(wire_d21_22),.data_out(wire_d21_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222124(.data_in(wire_d21_23),.data_out(wire_d21_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222125(.data_in(wire_d21_24),.data_out(wire_d21_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222126(.data_in(wire_d21_25),.data_out(wire_d21_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222127(.data_in(wire_d21_26),.data_out(wire_d21_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222128(.data_in(wire_d21_27),.data_out(wire_d21_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222129(.data_in(wire_d21_28),.data_out(wire_d21_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222130(.data_in(wire_d21_29),.data_out(wire_d21_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222131(.data_in(wire_d21_30),.data_out(wire_d21_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222132(.data_in(wire_d21_31),.data_out(wire_d21_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222133(.data_in(wire_d21_32),.data_out(wire_d21_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222134(.data_in(wire_d21_33),.data_out(wire_d21_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222135(.data_in(wire_d21_34),.data_out(wire_d21_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222136(.data_in(wire_d21_35),.data_out(wire_d21_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222137(.data_in(wire_d21_36),.data_out(wire_d21_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222138(.data_in(wire_d21_37),.data_out(wire_d21_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222139(.data_in(wire_d21_38),.data_out(wire_d21_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222140(.data_in(wire_d21_39),.data_out(wire_d21_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222141(.data_in(wire_d21_40),.data_out(wire_d21_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222142(.data_in(wire_d21_41),.data_out(wire_d21_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222143(.data_in(wire_d21_42),.data_out(wire_d21_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance222144(.data_in(wire_d21_43),.data_out(wire_d21_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222145(.data_in(wire_d21_44),.data_out(wire_d21_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance222146(.data_in(wire_d21_45),.data_out(wire_d21_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222147(.data_in(wire_d21_46),.data_out(wire_d21_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance222148(.data_in(wire_d21_47),.data_out(wire_d21_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance222149(.data_in(wire_d21_48),.data_out(d_out21),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance23220(.data_in(d_in22),.data_out(wire_d22_0),.clk(clk),.rst(rst));            //channel 23
	large_mux #(.WIDTH(WIDTH)) large_mux_instance23221(.data_in(wire_d22_0),.data_out(wire_d22_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance23222(.data_in(wire_d22_1),.data_out(wire_d22_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance23223(.data_in(wire_d22_2),.data_out(wire_d22_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance23224(.data_in(wire_d22_3),.data_out(wire_d22_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance23225(.data_in(wire_d22_4),.data_out(wire_d22_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance23226(.data_in(wire_d22_5),.data_out(wire_d22_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance23227(.data_in(wire_d22_6),.data_out(wire_d22_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance23228(.data_in(wire_d22_7),.data_out(wire_d22_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance23229(.data_in(wire_d22_8),.data_out(wire_d22_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232210(.data_in(wire_d22_9),.data_out(wire_d22_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232211(.data_in(wire_d22_10),.data_out(wire_d22_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232212(.data_in(wire_d22_11),.data_out(wire_d22_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232213(.data_in(wire_d22_12),.data_out(wire_d22_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232214(.data_in(wire_d22_13),.data_out(wire_d22_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232215(.data_in(wire_d22_14),.data_out(wire_d22_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232216(.data_in(wire_d22_15),.data_out(wire_d22_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232217(.data_in(wire_d22_16),.data_out(wire_d22_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232218(.data_in(wire_d22_17),.data_out(wire_d22_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232219(.data_in(wire_d22_18),.data_out(wire_d22_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232220(.data_in(wire_d22_19),.data_out(wire_d22_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232221(.data_in(wire_d22_20),.data_out(wire_d22_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232222(.data_in(wire_d22_21),.data_out(wire_d22_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232223(.data_in(wire_d22_22),.data_out(wire_d22_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232224(.data_in(wire_d22_23),.data_out(wire_d22_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232225(.data_in(wire_d22_24),.data_out(wire_d22_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232226(.data_in(wire_d22_25),.data_out(wire_d22_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232227(.data_in(wire_d22_26),.data_out(wire_d22_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232228(.data_in(wire_d22_27),.data_out(wire_d22_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232229(.data_in(wire_d22_28),.data_out(wire_d22_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232230(.data_in(wire_d22_29),.data_out(wire_d22_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232231(.data_in(wire_d22_30),.data_out(wire_d22_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232232(.data_in(wire_d22_31),.data_out(wire_d22_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232233(.data_in(wire_d22_32),.data_out(wire_d22_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232234(.data_in(wire_d22_33),.data_out(wire_d22_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232235(.data_in(wire_d22_34),.data_out(wire_d22_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232236(.data_in(wire_d22_35),.data_out(wire_d22_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232237(.data_in(wire_d22_36),.data_out(wire_d22_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232238(.data_in(wire_d22_37),.data_out(wire_d22_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232239(.data_in(wire_d22_38),.data_out(wire_d22_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232240(.data_in(wire_d22_39),.data_out(wire_d22_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232241(.data_in(wire_d22_40),.data_out(wire_d22_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232242(.data_in(wire_d22_41),.data_out(wire_d22_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232243(.data_in(wire_d22_42),.data_out(wire_d22_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232244(.data_in(wire_d22_43),.data_out(wire_d22_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance232245(.data_in(wire_d22_44),.data_out(wire_d22_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance232246(.data_in(wire_d22_45),.data_out(wire_d22_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232247(.data_in(wire_d22_46),.data_out(wire_d22_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance232248(.data_in(wire_d22_47),.data_out(wire_d22_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance232249(.data_in(wire_d22_48),.data_out(d_out22),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance24230(.data_in(d_in23),.data_out(wire_d23_0),.clk(clk),.rst(rst));            //channel 24
	encoder #(.WIDTH(WIDTH)) encoder_instance24231(.data_in(wire_d23_0),.data_out(wire_d23_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance24232(.data_in(wire_d23_1),.data_out(wire_d23_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance24233(.data_in(wire_d23_2),.data_out(wire_d23_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance24234(.data_in(wire_d23_3),.data_out(wire_d23_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance24235(.data_in(wire_d23_4),.data_out(wire_d23_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance24236(.data_in(wire_d23_5),.data_out(wire_d23_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance24237(.data_in(wire_d23_6),.data_out(wire_d23_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance24238(.data_in(wire_d23_7),.data_out(wire_d23_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance24239(.data_in(wire_d23_8),.data_out(wire_d23_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242310(.data_in(wire_d23_9),.data_out(wire_d23_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242311(.data_in(wire_d23_10),.data_out(wire_d23_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242312(.data_in(wire_d23_11),.data_out(wire_d23_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242313(.data_in(wire_d23_12),.data_out(wire_d23_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242314(.data_in(wire_d23_13),.data_out(wire_d23_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242315(.data_in(wire_d23_14),.data_out(wire_d23_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242316(.data_in(wire_d23_15),.data_out(wire_d23_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242317(.data_in(wire_d23_16),.data_out(wire_d23_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242318(.data_in(wire_d23_17),.data_out(wire_d23_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242319(.data_in(wire_d23_18),.data_out(wire_d23_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242320(.data_in(wire_d23_19),.data_out(wire_d23_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242321(.data_in(wire_d23_20),.data_out(wire_d23_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242322(.data_in(wire_d23_21),.data_out(wire_d23_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242323(.data_in(wire_d23_22),.data_out(wire_d23_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242324(.data_in(wire_d23_23),.data_out(wire_d23_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242325(.data_in(wire_d23_24),.data_out(wire_d23_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242326(.data_in(wire_d23_25),.data_out(wire_d23_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242327(.data_in(wire_d23_26),.data_out(wire_d23_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242328(.data_in(wire_d23_27),.data_out(wire_d23_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242329(.data_in(wire_d23_28),.data_out(wire_d23_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242330(.data_in(wire_d23_29),.data_out(wire_d23_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242331(.data_in(wire_d23_30),.data_out(wire_d23_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242332(.data_in(wire_d23_31),.data_out(wire_d23_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242333(.data_in(wire_d23_32),.data_out(wire_d23_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242334(.data_in(wire_d23_33),.data_out(wire_d23_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242335(.data_in(wire_d23_34),.data_out(wire_d23_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242336(.data_in(wire_d23_35),.data_out(wire_d23_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242337(.data_in(wire_d23_36),.data_out(wire_d23_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242338(.data_in(wire_d23_37),.data_out(wire_d23_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242339(.data_in(wire_d23_38),.data_out(wire_d23_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242340(.data_in(wire_d23_39),.data_out(wire_d23_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242341(.data_in(wire_d23_40),.data_out(wire_d23_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242342(.data_in(wire_d23_41),.data_out(wire_d23_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance242343(.data_in(wire_d23_42),.data_out(wire_d23_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242344(.data_in(wire_d23_43),.data_out(wire_d23_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242345(.data_in(wire_d23_44),.data_out(wire_d23_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242346(.data_in(wire_d23_45),.data_out(wire_d23_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance242347(.data_in(wire_d23_46),.data_out(wire_d23_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance242348(.data_in(wire_d23_47),.data_out(wire_d23_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance242349(.data_in(wire_d23_48),.data_out(d_out23),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance25240(.data_in(d_in24),.data_out(wire_d24_0),.clk(clk),.rst(rst));            //channel 25
	invertion #(.WIDTH(WIDTH)) invertion_instance25241(.data_in(wire_d24_0),.data_out(wire_d24_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance25242(.data_in(wire_d24_1),.data_out(wire_d24_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance25243(.data_in(wire_d24_2),.data_out(wire_d24_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance25244(.data_in(wire_d24_3),.data_out(wire_d24_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance25245(.data_in(wire_d24_4),.data_out(wire_d24_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance25246(.data_in(wire_d24_5),.data_out(wire_d24_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance25247(.data_in(wire_d24_6),.data_out(wire_d24_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance25248(.data_in(wire_d24_7),.data_out(wire_d24_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance25249(.data_in(wire_d24_8),.data_out(wire_d24_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252410(.data_in(wire_d24_9),.data_out(wire_d24_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252411(.data_in(wire_d24_10),.data_out(wire_d24_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252412(.data_in(wire_d24_11),.data_out(wire_d24_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252413(.data_in(wire_d24_12),.data_out(wire_d24_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252414(.data_in(wire_d24_13),.data_out(wire_d24_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252415(.data_in(wire_d24_14),.data_out(wire_d24_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252416(.data_in(wire_d24_15),.data_out(wire_d24_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252417(.data_in(wire_d24_16),.data_out(wire_d24_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252418(.data_in(wire_d24_17),.data_out(wire_d24_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252419(.data_in(wire_d24_18),.data_out(wire_d24_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252420(.data_in(wire_d24_19),.data_out(wire_d24_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252421(.data_in(wire_d24_20),.data_out(wire_d24_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252422(.data_in(wire_d24_21),.data_out(wire_d24_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252423(.data_in(wire_d24_22),.data_out(wire_d24_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252424(.data_in(wire_d24_23),.data_out(wire_d24_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252425(.data_in(wire_d24_24),.data_out(wire_d24_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252426(.data_in(wire_d24_25),.data_out(wire_d24_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance252427(.data_in(wire_d24_26),.data_out(wire_d24_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252428(.data_in(wire_d24_27),.data_out(wire_d24_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252429(.data_in(wire_d24_28),.data_out(wire_d24_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252430(.data_in(wire_d24_29),.data_out(wire_d24_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252431(.data_in(wire_d24_30),.data_out(wire_d24_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252432(.data_in(wire_d24_31),.data_out(wire_d24_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252433(.data_in(wire_d24_32),.data_out(wire_d24_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252434(.data_in(wire_d24_33),.data_out(wire_d24_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252435(.data_in(wire_d24_34),.data_out(wire_d24_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252436(.data_in(wire_d24_35),.data_out(wire_d24_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252437(.data_in(wire_d24_36),.data_out(wire_d24_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252438(.data_in(wire_d24_37),.data_out(wire_d24_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252439(.data_in(wire_d24_38),.data_out(wire_d24_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252440(.data_in(wire_d24_39),.data_out(wire_d24_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252441(.data_in(wire_d24_40),.data_out(wire_d24_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252442(.data_in(wire_d24_41),.data_out(wire_d24_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252443(.data_in(wire_d24_42),.data_out(wire_d24_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252444(.data_in(wire_d24_43),.data_out(wire_d24_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252445(.data_in(wire_d24_44),.data_out(wire_d24_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance252446(.data_in(wire_d24_45),.data_out(wire_d24_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252447(.data_in(wire_d24_46),.data_out(wire_d24_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance252448(.data_in(wire_d24_47),.data_out(wire_d24_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance252449(.data_in(wire_d24_48),.data_out(d_out24),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance26250(.data_in(d_in25),.data_out(wire_d25_0),.clk(clk),.rst(rst));            //channel 26
	invertion #(.WIDTH(WIDTH)) invertion_instance26251(.data_in(wire_d25_0),.data_out(wire_d25_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance26252(.data_in(wire_d25_1),.data_out(wire_d25_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance26253(.data_in(wire_d25_2),.data_out(wire_d25_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance26254(.data_in(wire_d25_3),.data_out(wire_d25_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance26255(.data_in(wire_d25_4),.data_out(wire_d25_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance26256(.data_in(wire_d25_5),.data_out(wire_d25_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance26257(.data_in(wire_d25_6),.data_out(wire_d25_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance26258(.data_in(wire_d25_7),.data_out(wire_d25_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance26259(.data_in(wire_d25_8),.data_out(wire_d25_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262510(.data_in(wire_d25_9),.data_out(wire_d25_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262511(.data_in(wire_d25_10),.data_out(wire_d25_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262512(.data_in(wire_d25_11),.data_out(wire_d25_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262513(.data_in(wire_d25_12),.data_out(wire_d25_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262514(.data_in(wire_d25_13),.data_out(wire_d25_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262515(.data_in(wire_d25_14),.data_out(wire_d25_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262516(.data_in(wire_d25_15),.data_out(wire_d25_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262517(.data_in(wire_d25_16),.data_out(wire_d25_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262518(.data_in(wire_d25_17),.data_out(wire_d25_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262519(.data_in(wire_d25_18),.data_out(wire_d25_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262520(.data_in(wire_d25_19),.data_out(wire_d25_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262521(.data_in(wire_d25_20),.data_out(wire_d25_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262522(.data_in(wire_d25_21),.data_out(wire_d25_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262523(.data_in(wire_d25_22),.data_out(wire_d25_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262524(.data_in(wire_d25_23),.data_out(wire_d25_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262525(.data_in(wire_d25_24),.data_out(wire_d25_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262526(.data_in(wire_d25_25),.data_out(wire_d25_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262527(.data_in(wire_d25_26),.data_out(wire_d25_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262528(.data_in(wire_d25_27),.data_out(wire_d25_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262529(.data_in(wire_d25_28),.data_out(wire_d25_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262530(.data_in(wire_d25_29),.data_out(wire_d25_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262531(.data_in(wire_d25_30),.data_out(wire_d25_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262532(.data_in(wire_d25_31),.data_out(wire_d25_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance262533(.data_in(wire_d25_32),.data_out(wire_d25_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262534(.data_in(wire_d25_33),.data_out(wire_d25_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262535(.data_in(wire_d25_34),.data_out(wire_d25_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262536(.data_in(wire_d25_35),.data_out(wire_d25_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262537(.data_in(wire_d25_36),.data_out(wire_d25_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262538(.data_in(wire_d25_37),.data_out(wire_d25_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262539(.data_in(wire_d25_38),.data_out(wire_d25_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262540(.data_in(wire_d25_39),.data_out(wire_d25_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262541(.data_in(wire_d25_40),.data_out(wire_d25_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262542(.data_in(wire_d25_41),.data_out(wire_d25_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262543(.data_in(wire_d25_42),.data_out(wire_d25_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262544(.data_in(wire_d25_43),.data_out(wire_d25_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262545(.data_in(wire_d25_44),.data_out(wire_d25_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance262546(.data_in(wire_d25_45),.data_out(wire_d25_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262547(.data_in(wire_d25_46),.data_out(wire_d25_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance262548(.data_in(wire_d25_47),.data_out(wire_d25_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance262549(.data_in(wire_d25_48),.data_out(d_out25),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance27260(.data_in(d_in26),.data_out(wire_d26_0),.clk(clk),.rst(rst));            //channel 27
	register #(.WIDTH(WIDTH)) register_instance27261(.data_in(wire_d26_0),.data_out(wire_d26_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance27262(.data_in(wire_d26_1),.data_out(wire_d26_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance27263(.data_in(wire_d26_2),.data_out(wire_d26_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance27264(.data_in(wire_d26_3),.data_out(wire_d26_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance27265(.data_in(wire_d26_4),.data_out(wire_d26_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance27266(.data_in(wire_d26_5),.data_out(wire_d26_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance27267(.data_in(wire_d26_6),.data_out(wire_d26_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance27268(.data_in(wire_d26_7),.data_out(wire_d26_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance27269(.data_in(wire_d26_8),.data_out(wire_d26_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272610(.data_in(wire_d26_9),.data_out(wire_d26_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272611(.data_in(wire_d26_10),.data_out(wire_d26_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272612(.data_in(wire_d26_11),.data_out(wire_d26_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272613(.data_in(wire_d26_12),.data_out(wire_d26_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272614(.data_in(wire_d26_13),.data_out(wire_d26_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272615(.data_in(wire_d26_14),.data_out(wire_d26_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272616(.data_in(wire_d26_15),.data_out(wire_d26_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272617(.data_in(wire_d26_16),.data_out(wire_d26_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272618(.data_in(wire_d26_17),.data_out(wire_d26_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272619(.data_in(wire_d26_18),.data_out(wire_d26_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272620(.data_in(wire_d26_19),.data_out(wire_d26_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272621(.data_in(wire_d26_20),.data_out(wire_d26_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272622(.data_in(wire_d26_21),.data_out(wire_d26_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272623(.data_in(wire_d26_22),.data_out(wire_d26_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272624(.data_in(wire_d26_23),.data_out(wire_d26_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272625(.data_in(wire_d26_24),.data_out(wire_d26_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272626(.data_in(wire_d26_25),.data_out(wire_d26_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272627(.data_in(wire_d26_26),.data_out(wire_d26_27),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272628(.data_in(wire_d26_27),.data_out(wire_d26_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272629(.data_in(wire_d26_28),.data_out(wire_d26_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272630(.data_in(wire_d26_29),.data_out(wire_d26_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272631(.data_in(wire_d26_30),.data_out(wire_d26_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272632(.data_in(wire_d26_31),.data_out(wire_d26_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272633(.data_in(wire_d26_32),.data_out(wire_d26_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272634(.data_in(wire_d26_33),.data_out(wire_d26_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272635(.data_in(wire_d26_34),.data_out(wire_d26_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272636(.data_in(wire_d26_35),.data_out(wire_d26_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272637(.data_in(wire_d26_36),.data_out(wire_d26_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272638(.data_in(wire_d26_37),.data_out(wire_d26_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272639(.data_in(wire_d26_38),.data_out(wire_d26_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272640(.data_in(wire_d26_39),.data_out(wire_d26_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272641(.data_in(wire_d26_40),.data_out(wire_d26_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance272642(.data_in(wire_d26_41),.data_out(wire_d26_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272643(.data_in(wire_d26_42),.data_out(wire_d26_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272644(.data_in(wire_d26_43),.data_out(wire_d26_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272645(.data_in(wire_d26_44),.data_out(wire_d26_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272646(.data_in(wire_d26_45),.data_out(wire_d26_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance272647(.data_in(wire_d26_46),.data_out(wire_d26_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance272648(.data_in(wire_d26_47),.data_out(wire_d26_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance272649(.data_in(wire_d26_48),.data_out(d_out26),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance28270(.data_in(d_in27),.data_out(wire_d27_0),.clk(clk),.rst(rst));            //channel 28
	register #(.WIDTH(WIDTH)) register_instance28271(.data_in(wire_d27_0),.data_out(wire_d27_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance28272(.data_in(wire_d27_1),.data_out(wire_d27_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance28273(.data_in(wire_d27_2),.data_out(wire_d27_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance28274(.data_in(wire_d27_3),.data_out(wire_d27_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance28275(.data_in(wire_d27_4),.data_out(wire_d27_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance28276(.data_in(wire_d27_5),.data_out(wire_d27_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance28277(.data_in(wire_d27_6),.data_out(wire_d27_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance28278(.data_in(wire_d27_7),.data_out(wire_d27_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance28279(.data_in(wire_d27_8),.data_out(wire_d27_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282710(.data_in(wire_d27_9),.data_out(wire_d27_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282711(.data_in(wire_d27_10),.data_out(wire_d27_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282712(.data_in(wire_d27_11),.data_out(wire_d27_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282713(.data_in(wire_d27_12),.data_out(wire_d27_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282714(.data_in(wire_d27_13),.data_out(wire_d27_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282715(.data_in(wire_d27_14),.data_out(wire_d27_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282716(.data_in(wire_d27_15),.data_out(wire_d27_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282717(.data_in(wire_d27_16),.data_out(wire_d27_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282718(.data_in(wire_d27_17),.data_out(wire_d27_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282719(.data_in(wire_d27_18),.data_out(wire_d27_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282720(.data_in(wire_d27_19),.data_out(wire_d27_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282721(.data_in(wire_d27_20),.data_out(wire_d27_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282722(.data_in(wire_d27_21),.data_out(wire_d27_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282723(.data_in(wire_d27_22),.data_out(wire_d27_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282724(.data_in(wire_d27_23),.data_out(wire_d27_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282725(.data_in(wire_d27_24),.data_out(wire_d27_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282726(.data_in(wire_d27_25),.data_out(wire_d27_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282727(.data_in(wire_d27_26),.data_out(wire_d27_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282728(.data_in(wire_d27_27),.data_out(wire_d27_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282729(.data_in(wire_d27_28),.data_out(wire_d27_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282730(.data_in(wire_d27_29),.data_out(wire_d27_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282731(.data_in(wire_d27_30),.data_out(wire_d27_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282732(.data_in(wire_d27_31),.data_out(wire_d27_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282733(.data_in(wire_d27_32),.data_out(wire_d27_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282734(.data_in(wire_d27_33),.data_out(wire_d27_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282735(.data_in(wire_d27_34),.data_out(wire_d27_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282736(.data_in(wire_d27_35),.data_out(wire_d27_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282737(.data_in(wire_d27_36),.data_out(wire_d27_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282738(.data_in(wire_d27_37),.data_out(wire_d27_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282739(.data_in(wire_d27_38),.data_out(wire_d27_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282740(.data_in(wire_d27_39),.data_out(wire_d27_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282741(.data_in(wire_d27_40),.data_out(wire_d27_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282742(.data_in(wire_d27_41),.data_out(wire_d27_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282743(.data_in(wire_d27_42),.data_out(wire_d27_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282744(.data_in(wire_d27_43),.data_out(wire_d27_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282745(.data_in(wire_d27_44),.data_out(wire_d27_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance282746(.data_in(wire_d27_45),.data_out(wire_d27_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance282747(.data_in(wire_d27_46),.data_out(wire_d27_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance282748(.data_in(wire_d27_47),.data_out(wire_d27_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance282749(.data_in(wire_d27_48),.data_out(d_out27),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance29280(.data_in(d_in28),.data_out(wire_d28_0),.clk(clk),.rst(rst));            //channel 29
	encoder #(.WIDTH(WIDTH)) encoder_instance29281(.data_in(wire_d28_0),.data_out(wire_d28_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance29282(.data_in(wire_d28_1),.data_out(wire_d28_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance29283(.data_in(wire_d28_2),.data_out(wire_d28_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance29284(.data_in(wire_d28_3),.data_out(wire_d28_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance29285(.data_in(wire_d28_4),.data_out(wire_d28_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance29286(.data_in(wire_d28_5),.data_out(wire_d28_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance29287(.data_in(wire_d28_6),.data_out(wire_d28_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance29288(.data_in(wire_d28_7),.data_out(wire_d28_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance29289(.data_in(wire_d28_8),.data_out(wire_d28_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292810(.data_in(wire_d28_9),.data_out(wire_d28_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292811(.data_in(wire_d28_10),.data_out(wire_d28_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292812(.data_in(wire_d28_11),.data_out(wire_d28_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292813(.data_in(wire_d28_12),.data_out(wire_d28_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292814(.data_in(wire_d28_13),.data_out(wire_d28_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292815(.data_in(wire_d28_14),.data_out(wire_d28_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292816(.data_in(wire_d28_15),.data_out(wire_d28_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292817(.data_in(wire_d28_16),.data_out(wire_d28_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292818(.data_in(wire_d28_17),.data_out(wire_d28_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292819(.data_in(wire_d28_18),.data_out(wire_d28_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292820(.data_in(wire_d28_19),.data_out(wire_d28_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292821(.data_in(wire_d28_20),.data_out(wire_d28_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292822(.data_in(wire_d28_21),.data_out(wire_d28_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292823(.data_in(wire_d28_22),.data_out(wire_d28_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292824(.data_in(wire_d28_23),.data_out(wire_d28_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292825(.data_in(wire_d28_24),.data_out(wire_d28_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292826(.data_in(wire_d28_25),.data_out(wire_d28_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292827(.data_in(wire_d28_26),.data_out(wire_d28_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292828(.data_in(wire_d28_27),.data_out(wire_d28_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292829(.data_in(wire_d28_28),.data_out(wire_d28_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292830(.data_in(wire_d28_29),.data_out(wire_d28_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292831(.data_in(wire_d28_30),.data_out(wire_d28_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292832(.data_in(wire_d28_31),.data_out(wire_d28_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292833(.data_in(wire_d28_32),.data_out(wire_d28_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292834(.data_in(wire_d28_33),.data_out(wire_d28_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292835(.data_in(wire_d28_34),.data_out(wire_d28_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292836(.data_in(wire_d28_35),.data_out(wire_d28_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292837(.data_in(wire_d28_36),.data_out(wire_d28_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292838(.data_in(wire_d28_37),.data_out(wire_d28_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292839(.data_in(wire_d28_38),.data_out(wire_d28_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292840(.data_in(wire_d28_39),.data_out(wire_d28_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance292841(.data_in(wire_d28_40),.data_out(wire_d28_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292842(.data_in(wire_d28_41),.data_out(wire_d28_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292843(.data_in(wire_d28_42),.data_out(wire_d28_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292844(.data_in(wire_d28_43),.data_out(wire_d28_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292845(.data_in(wire_d28_44),.data_out(wire_d28_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance292846(.data_in(wire_d28_45),.data_out(wire_d28_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance292847(.data_in(wire_d28_46),.data_out(wire_d28_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292848(.data_in(wire_d28_47),.data_out(wire_d28_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance292849(.data_in(wire_d28_48),.data_out(d_out28),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance30290(.data_in(d_in29),.data_out(wire_d29_0),.clk(clk),.rst(rst));            //channel 30
	encoder #(.WIDTH(WIDTH)) encoder_instance30291(.data_in(wire_d29_0),.data_out(wire_d29_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance30292(.data_in(wire_d29_1),.data_out(wire_d29_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance30293(.data_in(wire_d29_2),.data_out(wire_d29_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance30294(.data_in(wire_d29_3),.data_out(wire_d29_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance30295(.data_in(wire_d29_4),.data_out(wire_d29_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance30296(.data_in(wire_d29_5),.data_out(wire_d29_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance30297(.data_in(wire_d29_6),.data_out(wire_d29_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance30298(.data_in(wire_d29_7),.data_out(wire_d29_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance30299(.data_in(wire_d29_8),.data_out(wire_d29_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302910(.data_in(wire_d29_9),.data_out(wire_d29_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302911(.data_in(wire_d29_10),.data_out(wire_d29_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302912(.data_in(wire_d29_11),.data_out(wire_d29_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302913(.data_in(wire_d29_12),.data_out(wire_d29_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302914(.data_in(wire_d29_13),.data_out(wire_d29_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302915(.data_in(wire_d29_14),.data_out(wire_d29_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302916(.data_in(wire_d29_15),.data_out(wire_d29_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302917(.data_in(wire_d29_16),.data_out(wire_d29_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302918(.data_in(wire_d29_17),.data_out(wire_d29_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302919(.data_in(wire_d29_18),.data_out(wire_d29_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302920(.data_in(wire_d29_19),.data_out(wire_d29_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302921(.data_in(wire_d29_20),.data_out(wire_d29_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302922(.data_in(wire_d29_21),.data_out(wire_d29_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302923(.data_in(wire_d29_22),.data_out(wire_d29_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302924(.data_in(wire_d29_23),.data_out(wire_d29_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302925(.data_in(wire_d29_24),.data_out(wire_d29_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302926(.data_in(wire_d29_25),.data_out(wire_d29_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302927(.data_in(wire_d29_26),.data_out(wire_d29_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302928(.data_in(wire_d29_27),.data_out(wire_d29_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302929(.data_in(wire_d29_28),.data_out(wire_d29_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302930(.data_in(wire_d29_29),.data_out(wire_d29_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302931(.data_in(wire_d29_30),.data_out(wire_d29_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302932(.data_in(wire_d29_31),.data_out(wire_d29_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302933(.data_in(wire_d29_32),.data_out(wire_d29_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance302934(.data_in(wire_d29_33),.data_out(wire_d29_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302935(.data_in(wire_d29_34),.data_out(wire_d29_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302936(.data_in(wire_d29_35),.data_out(wire_d29_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302937(.data_in(wire_d29_36),.data_out(wire_d29_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302938(.data_in(wire_d29_37),.data_out(wire_d29_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302939(.data_in(wire_d29_38),.data_out(wire_d29_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302940(.data_in(wire_d29_39),.data_out(wire_d29_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302941(.data_in(wire_d29_40),.data_out(wire_d29_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302942(.data_in(wire_d29_41),.data_out(wire_d29_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302943(.data_in(wire_d29_42),.data_out(wire_d29_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance302944(.data_in(wire_d29_43),.data_out(wire_d29_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302945(.data_in(wire_d29_44),.data_out(wire_d29_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302946(.data_in(wire_d29_45),.data_out(wire_d29_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance302947(.data_in(wire_d29_46),.data_out(wire_d29_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302948(.data_in(wire_d29_47),.data_out(wire_d29_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance302949(.data_in(wire_d29_48),.data_out(d_out29),.clk(clk),.rst(rst));


endmodule