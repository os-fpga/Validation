`include "encoder.v"
`include "invertion.v"
`include "large_adder.v"
`include "large_mux.v"
`include "memory_cntrl.v"
`include "register.v"
`include "full_adder.v"
`include "d_latch.v"
`include "shift_reg.v"
`include "mod_n_counter.v"
`include "decoder.v"
`include "parity_generator.v"

module design205_55_50_top #(parameter WIDTH=32,CHANNEL=55) (clk, rst, in, out);

	localparam OUT_BUS=CHANNEL*WIDTH;
	input clk,rst;
	input [WIDTH-1:0] in;
	output [WIDTH-1:0] out;

	reg [WIDTH-1:0] d_in0;
	reg [WIDTH-1:0] d_in1;
	reg [WIDTH-1:0] d_in2;
	reg [WIDTH-1:0] d_in3;
	reg [WIDTH-1:0] d_in4;
	reg [WIDTH-1:0] d_in5;
	reg [WIDTH-1:0] d_in6;
	reg [WIDTH-1:0] d_in7;
	reg [WIDTH-1:0] d_in8;
	reg [WIDTH-1:0] d_in9;
	reg [WIDTH-1:0] d_in10;
	reg [WIDTH-1:0] d_in11;
	reg [WIDTH-1:0] d_in12;
	reg [WIDTH-1:0] d_in13;
	reg [WIDTH-1:0] d_in14;
	reg [WIDTH-1:0] d_in15;
	reg [WIDTH-1:0] d_in16;
	reg [WIDTH-1:0] d_in17;
	reg [WIDTH-1:0] d_in18;
	reg [WIDTH-1:0] d_in19;
	reg [WIDTH-1:0] d_in20;
	reg [WIDTH-1:0] d_in21;
	reg [WIDTH-1:0] d_in22;
	reg [WIDTH-1:0] d_in23;
	reg [WIDTH-1:0] d_in24;
	reg [WIDTH-1:0] d_in25;
	reg [WIDTH-1:0] d_in26;
	reg [WIDTH-1:0] d_in27;
	reg [WIDTH-1:0] d_in28;
	reg [WIDTH-1:0] d_in29;
	reg [WIDTH-1:0] d_in30;
	reg [WIDTH-1:0] d_in31;
	reg [WIDTH-1:0] d_in32;
	reg [WIDTH-1:0] d_in33;
	reg [WIDTH-1:0] d_in34;
	reg [WIDTH-1:0] d_in35;
	reg [WIDTH-1:0] d_in36;
	reg [WIDTH-1:0] d_in37;
	reg [WIDTH-1:0] d_in38;
	reg [WIDTH-1:0] d_in39;
	reg [WIDTH-1:0] d_in40;
	reg [WIDTH-1:0] d_in41;
	reg [WIDTH-1:0] d_in42;
	reg [WIDTH-1:0] d_in43;
	reg [WIDTH-1:0] d_in44;
	reg [WIDTH-1:0] d_in45;
	reg [WIDTH-1:0] d_in46;
	reg [WIDTH-1:0] d_in47;
	reg [WIDTH-1:0] d_in48;
	reg [WIDTH-1:0] d_in49;
	reg [WIDTH-1:0] d_in50;
	reg [WIDTH-1:0] d_in51;
	reg [WIDTH-1:0] d_in52;
	reg [WIDTH-1:0] d_in53;
	reg [WIDTH-1:0] d_in54;
	wire [WIDTH-1:0] d_out0;
	wire [WIDTH-1:0] d_out1;
	wire [WIDTH-1:0] d_out2;
	wire [WIDTH-1:0] d_out3;
	wire [WIDTH-1:0] d_out4;
	wire [WIDTH-1:0] d_out5;
	wire [WIDTH-1:0] d_out6;
	wire [WIDTH-1:0] d_out7;
	wire [WIDTH-1:0] d_out8;
	wire [WIDTH-1:0] d_out9;
	wire [WIDTH-1:0] d_out10;
	wire [WIDTH-1:0] d_out11;
	wire [WIDTH-1:0] d_out12;
	wire [WIDTH-1:0] d_out13;
	wire [WIDTH-1:0] d_out14;
	wire [WIDTH-1:0] d_out15;
	wire [WIDTH-1:0] d_out16;
	wire [WIDTH-1:0] d_out17;
	wire [WIDTH-1:0] d_out18;
	wire [WIDTH-1:0] d_out19;
	wire [WIDTH-1:0] d_out20;
	wire [WIDTH-1:0] d_out21;
	wire [WIDTH-1:0] d_out22;
	wire [WIDTH-1:0] d_out23;
	wire [WIDTH-1:0] d_out24;
	wire [WIDTH-1:0] d_out25;
	wire [WIDTH-1:0] d_out26;
	wire [WIDTH-1:0] d_out27;
	wire [WIDTH-1:0] d_out28;
	wire [WIDTH-1:0] d_out29;
	wire [WIDTH-1:0] d_out30;
	wire [WIDTH-1:0] d_out31;
	wire [WIDTH-1:0] d_out32;
	wire [WIDTH-1:0] d_out33;
	wire [WIDTH-1:0] d_out34;
	wire [WIDTH-1:0] d_out35;
	wire [WIDTH-1:0] d_out36;
	wire [WIDTH-1:0] d_out37;
	wire [WIDTH-1:0] d_out38;
	wire [WIDTH-1:0] d_out39;
	wire [WIDTH-1:0] d_out40;
	wire [WIDTH-1:0] d_out41;
	wire [WIDTH-1:0] d_out42;
	wire [WIDTH-1:0] d_out43;
	wire [WIDTH-1:0] d_out44;
	wire [WIDTH-1:0] d_out45;
	wire [WIDTH-1:0] d_out46;
	wire [WIDTH-1:0] d_out47;
	wire [WIDTH-1:0] d_out48;
	wire [WIDTH-1:0] d_out49;
	wire [WIDTH-1:0] d_out50;
	wire [WIDTH-1:0] d_out51;
	wire [WIDTH-1:0] d_out52;
	wire [WIDTH-1:0] d_out53;
	wire [WIDTH-1:0] d_out54;

	reg [OUT_BUS-1:0] tmp;

	always @ (posedge clk or posedge rst) begin
		if (rst)
			tmp <= 0;
		else
			tmp <= {tmp[OUT_BUS-(WIDTH-1):0],in};
	end

	always @ (posedge clk) begin
		d_in0 <= tmp[WIDTH-1:0];
		d_in1 <= tmp[(WIDTH*2)-1:WIDTH*1];
		d_in2 <= tmp[(WIDTH*3)-1:WIDTH*2];
		d_in3 <= tmp[(WIDTH*4)-1:WIDTH*3];
		d_in4 <= tmp[(WIDTH*5)-1:WIDTH*4];
		d_in5 <= tmp[(WIDTH*6)-1:WIDTH*5];
		d_in6 <= tmp[(WIDTH*7)-1:WIDTH*6];
		d_in7 <= tmp[(WIDTH*8)-1:WIDTH*7];
		d_in8 <= tmp[(WIDTH*9)-1:WIDTH*8];
		d_in9 <= tmp[(WIDTH*10)-1:WIDTH*9];
		d_in10 <= tmp[(WIDTH*11)-1:WIDTH*10];
		d_in11 <= tmp[(WIDTH*12)-1:WIDTH*11];
		d_in12 <= tmp[(WIDTH*13)-1:WIDTH*12];
		d_in13 <= tmp[(WIDTH*14)-1:WIDTH*13];
		d_in14 <= tmp[(WIDTH*15)-1:WIDTH*14];
		d_in15 <= tmp[(WIDTH*16)-1:WIDTH*15];
		d_in16 <= tmp[(WIDTH*17)-1:WIDTH*16];
		d_in17 <= tmp[(WIDTH*18)-1:WIDTH*17];
		d_in18 <= tmp[(WIDTH*19)-1:WIDTH*18];
		d_in19 <= tmp[(WIDTH*20)-1:WIDTH*19];
		d_in20 <= tmp[(WIDTH*21)-1:WIDTH*20];
		d_in21 <= tmp[(WIDTH*22)-1:WIDTH*21];
		d_in22 <= tmp[(WIDTH*23)-1:WIDTH*22];
		d_in23 <= tmp[(WIDTH*24)-1:WIDTH*23];
		d_in24 <= tmp[(WIDTH*25)-1:WIDTH*24];
		d_in25 <= tmp[(WIDTH*26)-1:WIDTH*25];
		d_in26 <= tmp[(WIDTH*27)-1:WIDTH*26];
		d_in27 <= tmp[(WIDTH*28)-1:WIDTH*27];
		d_in28 <= tmp[(WIDTH*29)-1:WIDTH*28];
		d_in29 <= tmp[(WIDTH*30)-1:WIDTH*29];
		d_in30 <= tmp[(WIDTH*31)-1:WIDTH*30];
		d_in31 <= tmp[(WIDTH*32)-1:WIDTH*31];
		d_in32 <= tmp[(WIDTH*33)-1:WIDTH*32];
		d_in33 <= tmp[(WIDTH*34)-1:WIDTH*33];
		d_in34 <= tmp[(WIDTH*35)-1:WIDTH*34];
		d_in35 <= tmp[(WIDTH*36)-1:WIDTH*35];
		d_in36 <= tmp[(WIDTH*37)-1:WIDTH*36];
		d_in37 <= tmp[(WIDTH*38)-1:WIDTH*37];
		d_in38 <= tmp[(WIDTH*39)-1:WIDTH*38];
		d_in39 <= tmp[(WIDTH*40)-1:WIDTH*39];
		d_in40 <= tmp[(WIDTH*41)-1:WIDTH*40];
		d_in41 <= tmp[(WIDTH*42)-1:WIDTH*41];
		d_in42 <= tmp[(WIDTH*43)-1:WIDTH*42];
		d_in43 <= tmp[(WIDTH*44)-1:WIDTH*43];
		d_in44 <= tmp[(WIDTH*45)-1:WIDTH*44];
		d_in45 <= tmp[(WIDTH*46)-1:WIDTH*45];
		d_in46 <= tmp[(WIDTH*47)-1:WIDTH*46];
		d_in47 <= tmp[(WIDTH*48)-1:WIDTH*47];
		d_in48 <= tmp[(WIDTH*49)-1:WIDTH*48];
		d_in49 <= tmp[(WIDTH*50)-1:WIDTH*49];
		d_in50 <= tmp[(WIDTH*51)-1:WIDTH*50];
		d_in51 <= tmp[(WIDTH*52)-1:WIDTH*51];
		d_in52 <= tmp[(WIDTH*53)-1:WIDTH*52];
		d_in53 <= tmp[(WIDTH*54)-1:WIDTH*53];
		d_in54 <= tmp[(WIDTH*55)-1:WIDTH*54];
	end

	design205_55_50 #(.WIDTH(WIDTH)) design205_55_50_inst(.d_in0(d_in0),.d_in1(d_in1),.d_in2(d_in2),.d_in3(d_in3),.d_in4(d_in4),.d_in5(d_in5),.d_in6(d_in6),.d_in7(d_in7),.d_in8(d_in8),.d_in9(d_in9),.d_in10(d_in10),.d_in11(d_in11),.d_in12(d_in12),.d_in13(d_in13),.d_in14(d_in14),.d_in15(d_in15),.d_in16(d_in16),.d_in17(d_in17),.d_in18(d_in18),.d_in19(d_in19),.d_in20(d_in20),.d_in21(d_in21),.d_in22(d_in22),.d_in23(d_in23),.d_in24(d_in24),.d_in25(d_in25),.d_in26(d_in26),.d_in27(d_in27),.d_in28(d_in28),.d_in29(d_in29),.d_in30(d_in30),.d_in31(d_in31),.d_in32(d_in32),.d_in33(d_in33),.d_in34(d_in34),.d_in35(d_in35),.d_in36(d_in36),.d_in37(d_in37),.d_in38(d_in38),.d_in39(d_in39),.d_in40(d_in40),.d_in41(d_in41),.d_in42(d_in42),.d_in43(d_in43),.d_in44(d_in44),.d_in45(d_in45),.d_in46(d_in46),.d_in47(d_in47),.d_in48(d_in48),.d_in49(d_in49),.d_in50(d_in50),.d_in51(d_in51),.d_in52(d_in52),.d_in53(d_in53),.d_in54(d_in54),.d_out0(d_out0),.d_out1(d_out1),.d_out2(d_out2),.d_out3(d_out3),.d_out4(d_out4),.d_out5(d_out5),.d_out6(d_out6),.d_out7(d_out7),.d_out8(d_out8),.d_out9(d_out9),.d_out10(d_out10),.d_out11(d_out11),.d_out12(d_out12),.d_out13(d_out13),.d_out14(d_out14),.d_out15(d_out15),.d_out16(d_out16),.d_out17(d_out17),.d_out18(d_out18),.d_out19(d_out19),.d_out20(d_out20),.d_out21(d_out21),.d_out22(d_out22),.d_out23(d_out23),.d_out24(d_out24),.d_out25(d_out25),.d_out26(d_out26),.d_out27(d_out27),.d_out28(d_out28),.d_out29(d_out29),.d_out30(d_out30),.d_out31(d_out31),.d_out32(d_out32),.d_out33(d_out33),.d_out34(d_out34),.d_out35(d_out35),.d_out36(d_out36),.d_out37(d_out37),.d_out38(d_out38),.d_out39(d_out39),.d_out40(d_out40),.d_out41(d_out41),.d_out42(d_out42),.d_out43(d_out43),.d_out44(d_out44),.d_out45(d_out45),.d_out46(d_out46),.d_out47(d_out47),.d_out48(d_out48),.d_out49(d_out49),.d_out50(d_out50),.d_out51(d_out51),.d_out52(d_out52),.d_out53(d_out53),.d_out54(d_out54),.clk(clk),.rst(rst));

	assign out = d_out0^d_out1^d_out2^d_out3^d_out4^d_out5^d_out6^d_out7^d_out8^d_out9^d_out10^d_out11^d_out12^d_out13^d_out14^d_out15^d_out16^d_out17^d_out18^d_out19^d_out20^d_out21^d_out22^d_out23^d_out24^d_out25^d_out26^d_out27^d_out28^d_out29^d_out30^d_out31^d_out32^d_out33^d_out34^d_out35^d_out36^d_out37^d_out38^d_out39^d_out40^d_out41^d_out42^d_out43^d_out44^d_out45^d_out46^d_out47^d_out48^d_out49^d_out50^d_out51^d_out52^d_out53^d_out54;

endmodule

module design205_55_50 #(parameter WIDTH=32) (d_in0, d_in1, d_in2, d_in3, d_in4, d_in5, d_in6, d_in7, d_in8, d_in9, d_in10, d_in11, d_in12, d_in13, d_in14, d_in15, d_in16, d_in17, d_in18, d_in19, d_in20, d_in21, d_in22, d_in23, d_in24, d_in25, d_in26, d_in27, d_in28, d_in29, d_in30, d_in31, d_in32, d_in33, d_in34, d_in35, d_in36, d_in37, d_in38, d_in39, d_in40, d_in41, d_in42, d_in43, d_in44, d_in45, d_in46, d_in47, d_in48, d_in49, d_in50, d_in51, d_in52, d_in53, d_in54, d_out0, d_out1, d_out2, d_out3, d_out4, d_out5, d_out6, d_out7, d_out8, d_out9, d_out10, d_out11, d_out12, d_out13, d_out14, d_out15, d_out16, d_out17, d_out18, d_out19, d_out20, d_out21, d_out22, d_out23, d_out24, d_out25, d_out26, d_out27, d_out28, d_out29, d_out30, d_out31, d_out32, d_out33, d_out34, d_out35, d_out36, d_out37, d_out38, d_out39, d_out40, d_out41, d_out42, d_out43, d_out44, d_out45, d_out46, d_out47, d_out48, d_out49, d_out50, d_out51, d_out52, d_out53, d_out54, clk, rst);
	input clk;
	input rst;
	input [WIDTH-1:0] d_in0; 
	input [WIDTH-1:0] d_in1; 
	input [WIDTH-1:0] d_in2; 
	input [WIDTH-1:0] d_in3; 
	input [WIDTH-1:0] d_in4; 
	input [WIDTH-1:0] d_in5; 
	input [WIDTH-1:0] d_in6; 
	input [WIDTH-1:0] d_in7; 
	input [WIDTH-1:0] d_in8; 
	input [WIDTH-1:0] d_in9; 
	input [WIDTH-1:0] d_in10; 
	input [WIDTH-1:0] d_in11; 
	input [WIDTH-1:0] d_in12; 
	input [WIDTH-1:0] d_in13; 
	input [WIDTH-1:0] d_in14; 
	input [WIDTH-1:0] d_in15; 
	input [WIDTH-1:0] d_in16; 
	input [WIDTH-1:0] d_in17; 
	input [WIDTH-1:0] d_in18; 
	input [WIDTH-1:0] d_in19; 
	input [WIDTH-1:0] d_in20; 
	input [WIDTH-1:0] d_in21; 
	input [WIDTH-1:0] d_in22; 
	input [WIDTH-1:0] d_in23; 
	input [WIDTH-1:0] d_in24; 
	input [WIDTH-1:0] d_in25; 
	input [WIDTH-1:0] d_in26; 
	input [WIDTH-1:0] d_in27; 
	input [WIDTH-1:0] d_in28; 
	input [WIDTH-1:0] d_in29; 
	input [WIDTH-1:0] d_in30; 
	input [WIDTH-1:0] d_in31; 
	input [WIDTH-1:0] d_in32; 
	input [WIDTH-1:0] d_in33; 
	input [WIDTH-1:0] d_in34; 
	input [WIDTH-1:0] d_in35; 
	input [WIDTH-1:0] d_in36; 
	input [WIDTH-1:0] d_in37; 
	input [WIDTH-1:0] d_in38; 
	input [WIDTH-1:0] d_in39; 
	input [WIDTH-1:0] d_in40; 
	input [WIDTH-1:0] d_in41; 
	input [WIDTH-1:0] d_in42; 
	input [WIDTH-1:0] d_in43; 
	input [WIDTH-1:0] d_in44; 
	input [WIDTH-1:0] d_in45; 
	input [WIDTH-1:0] d_in46; 
	input [WIDTH-1:0] d_in47; 
	input [WIDTH-1:0] d_in48; 
	input [WIDTH-1:0] d_in49; 
	input [WIDTH-1:0] d_in50; 
	input [WIDTH-1:0] d_in51; 
	input [WIDTH-1:0] d_in52; 
	input [WIDTH-1:0] d_in53; 
	input [WIDTH-1:0] d_in54; 
	output [WIDTH-1:0] d_out0; 
	output [WIDTH-1:0] d_out1; 
	output [WIDTH-1:0] d_out2; 
	output [WIDTH-1:0] d_out3; 
	output [WIDTH-1:0] d_out4; 
	output [WIDTH-1:0] d_out5; 
	output [WIDTH-1:0] d_out6; 
	output [WIDTH-1:0] d_out7; 
	output [WIDTH-1:0] d_out8; 
	output [WIDTH-1:0] d_out9; 
	output [WIDTH-1:0] d_out10; 
	output [WIDTH-1:0] d_out11; 
	output [WIDTH-1:0] d_out12; 
	output [WIDTH-1:0] d_out13; 
	output [WIDTH-1:0] d_out14; 
	output [WIDTH-1:0] d_out15; 
	output [WIDTH-1:0] d_out16; 
	output [WIDTH-1:0] d_out17; 
	output [WIDTH-1:0] d_out18; 
	output [WIDTH-1:0] d_out19; 
	output [WIDTH-1:0] d_out20; 
	output [WIDTH-1:0] d_out21; 
	output [WIDTH-1:0] d_out22; 
	output [WIDTH-1:0] d_out23; 
	output [WIDTH-1:0] d_out24; 
	output [WIDTH-1:0] d_out25; 
	output [WIDTH-1:0] d_out26; 
	output [WIDTH-1:0] d_out27; 
	output [WIDTH-1:0] d_out28; 
	output [WIDTH-1:0] d_out29; 
	output [WIDTH-1:0] d_out30; 
	output [WIDTH-1:0] d_out31; 
	output [WIDTH-1:0] d_out32; 
	output [WIDTH-1:0] d_out33; 
	output [WIDTH-1:0] d_out34; 
	output [WIDTH-1:0] d_out35; 
	output [WIDTH-1:0] d_out36; 
	output [WIDTH-1:0] d_out37; 
	output [WIDTH-1:0] d_out38; 
	output [WIDTH-1:0] d_out39; 
	output [WIDTH-1:0] d_out40; 
	output [WIDTH-1:0] d_out41; 
	output [WIDTH-1:0] d_out42; 
	output [WIDTH-1:0] d_out43; 
	output [WIDTH-1:0] d_out44; 
	output [WIDTH-1:0] d_out45; 
	output [WIDTH-1:0] d_out46; 
	output [WIDTH-1:0] d_out47; 
	output [WIDTH-1:0] d_out48; 
	output [WIDTH-1:0] d_out49; 
	output [WIDTH-1:0] d_out50; 
	output [WIDTH-1:0] d_out51; 
	output [WIDTH-1:0] d_out52; 
	output [WIDTH-1:0] d_out53; 
	output [WIDTH-1:0] d_out54; 

	wire [WIDTH-1:0] wire_d0_0;
	wire [WIDTH-1:0] wire_d0_1;
	wire [WIDTH-1:0] wire_d0_2;
	wire [WIDTH-1:0] wire_d0_3;
	wire [WIDTH-1:0] wire_d0_4;
	wire [WIDTH-1:0] wire_d0_5;
	wire [WIDTH-1:0] wire_d0_6;
	wire [WIDTH-1:0] wire_d0_7;
	wire [WIDTH-1:0] wire_d0_8;
	wire [WIDTH-1:0] wire_d0_9;
	wire [WIDTH-1:0] wire_d0_10;
	wire [WIDTH-1:0] wire_d0_11;
	wire [WIDTH-1:0] wire_d0_12;
	wire [WIDTH-1:0] wire_d0_13;
	wire [WIDTH-1:0] wire_d0_14;
	wire [WIDTH-1:0] wire_d0_15;
	wire [WIDTH-1:0] wire_d0_16;
	wire [WIDTH-1:0] wire_d0_17;
	wire [WIDTH-1:0] wire_d0_18;
	wire [WIDTH-1:0] wire_d0_19;
	wire [WIDTH-1:0] wire_d0_20;
	wire [WIDTH-1:0] wire_d0_21;
	wire [WIDTH-1:0] wire_d0_22;
	wire [WIDTH-1:0] wire_d0_23;
	wire [WIDTH-1:0] wire_d0_24;
	wire [WIDTH-1:0] wire_d0_25;
	wire [WIDTH-1:0] wire_d0_26;
	wire [WIDTH-1:0] wire_d0_27;
	wire [WIDTH-1:0] wire_d0_28;
	wire [WIDTH-1:0] wire_d0_29;
	wire [WIDTH-1:0] wire_d0_30;
	wire [WIDTH-1:0] wire_d0_31;
	wire [WIDTH-1:0] wire_d0_32;
	wire [WIDTH-1:0] wire_d0_33;
	wire [WIDTH-1:0] wire_d0_34;
	wire [WIDTH-1:0] wire_d0_35;
	wire [WIDTH-1:0] wire_d0_36;
	wire [WIDTH-1:0] wire_d0_37;
	wire [WIDTH-1:0] wire_d0_38;
	wire [WIDTH-1:0] wire_d0_39;
	wire [WIDTH-1:0] wire_d0_40;
	wire [WIDTH-1:0] wire_d0_41;
	wire [WIDTH-1:0] wire_d0_42;
	wire [WIDTH-1:0] wire_d0_43;
	wire [WIDTH-1:0] wire_d0_44;
	wire [WIDTH-1:0] wire_d0_45;
	wire [WIDTH-1:0] wire_d0_46;
	wire [WIDTH-1:0] wire_d0_47;
	wire [WIDTH-1:0] wire_d0_48;
	wire [WIDTH-1:0] wire_d1_0;
	wire [WIDTH-1:0] wire_d1_1;
	wire [WIDTH-1:0] wire_d1_2;
	wire [WIDTH-1:0] wire_d1_3;
	wire [WIDTH-1:0] wire_d1_4;
	wire [WIDTH-1:0] wire_d1_5;
	wire [WIDTH-1:0] wire_d1_6;
	wire [WIDTH-1:0] wire_d1_7;
	wire [WIDTH-1:0] wire_d1_8;
	wire [WIDTH-1:0] wire_d1_9;
	wire [WIDTH-1:0] wire_d1_10;
	wire [WIDTH-1:0] wire_d1_11;
	wire [WIDTH-1:0] wire_d1_12;
	wire [WIDTH-1:0] wire_d1_13;
	wire [WIDTH-1:0] wire_d1_14;
	wire [WIDTH-1:0] wire_d1_15;
	wire [WIDTH-1:0] wire_d1_16;
	wire [WIDTH-1:0] wire_d1_17;
	wire [WIDTH-1:0] wire_d1_18;
	wire [WIDTH-1:0] wire_d1_19;
	wire [WIDTH-1:0] wire_d1_20;
	wire [WIDTH-1:0] wire_d1_21;
	wire [WIDTH-1:0] wire_d1_22;
	wire [WIDTH-1:0] wire_d1_23;
	wire [WIDTH-1:0] wire_d1_24;
	wire [WIDTH-1:0] wire_d1_25;
	wire [WIDTH-1:0] wire_d1_26;
	wire [WIDTH-1:0] wire_d1_27;
	wire [WIDTH-1:0] wire_d1_28;
	wire [WIDTH-1:0] wire_d1_29;
	wire [WIDTH-1:0] wire_d1_30;
	wire [WIDTH-1:0] wire_d1_31;
	wire [WIDTH-1:0] wire_d1_32;
	wire [WIDTH-1:0] wire_d1_33;
	wire [WIDTH-1:0] wire_d1_34;
	wire [WIDTH-1:0] wire_d1_35;
	wire [WIDTH-1:0] wire_d1_36;
	wire [WIDTH-1:0] wire_d1_37;
	wire [WIDTH-1:0] wire_d1_38;
	wire [WIDTH-1:0] wire_d1_39;
	wire [WIDTH-1:0] wire_d1_40;
	wire [WIDTH-1:0] wire_d1_41;
	wire [WIDTH-1:0] wire_d1_42;
	wire [WIDTH-1:0] wire_d1_43;
	wire [WIDTH-1:0] wire_d1_44;
	wire [WIDTH-1:0] wire_d1_45;
	wire [WIDTH-1:0] wire_d1_46;
	wire [WIDTH-1:0] wire_d1_47;
	wire [WIDTH-1:0] wire_d1_48;
	wire [WIDTH-1:0] wire_d2_0;
	wire [WIDTH-1:0] wire_d2_1;
	wire [WIDTH-1:0] wire_d2_2;
	wire [WIDTH-1:0] wire_d2_3;
	wire [WIDTH-1:0] wire_d2_4;
	wire [WIDTH-1:0] wire_d2_5;
	wire [WIDTH-1:0] wire_d2_6;
	wire [WIDTH-1:0] wire_d2_7;
	wire [WIDTH-1:0] wire_d2_8;
	wire [WIDTH-1:0] wire_d2_9;
	wire [WIDTH-1:0] wire_d2_10;
	wire [WIDTH-1:0] wire_d2_11;
	wire [WIDTH-1:0] wire_d2_12;
	wire [WIDTH-1:0] wire_d2_13;
	wire [WIDTH-1:0] wire_d2_14;
	wire [WIDTH-1:0] wire_d2_15;
	wire [WIDTH-1:0] wire_d2_16;
	wire [WIDTH-1:0] wire_d2_17;
	wire [WIDTH-1:0] wire_d2_18;
	wire [WIDTH-1:0] wire_d2_19;
	wire [WIDTH-1:0] wire_d2_20;
	wire [WIDTH-1:0] wire_d2_21;
	wire [WIDTH-1:0] wire_d2_22;
	wire [WIDTH-1:0] wire_d2_23;
	wire [WIDTH-1:0] wire_d2_24;
	wire [WIDTH-1:0] wire_d2_25;
	wire [WIDTH-1:0] wire_d2_26;
	wire [WIDTH-1:0] wire_d2_27;
	wire [WIDTH-1:0] wire_d2_28;
	wire [WIDTH-1:0] wire_d2_29;
	wire [WIDTH-1:0] wire_d2_30;
	wire [WIDTH-1:0] wire_d2_31;
	wire [WIDTH-1:0] wire_d2_32;
	wire [WIDTH-1:0] wire_d2_33;
	wire [WIDTH-1:0] wire_d2_34;
	wire [WIDTH-1:0] wire_d2_35;
	wire [WIDTH-1:0] wire_d2_36;
	wire [WIDTH-1:0] wire_d2_37;
	wire [WIDTH-1:0] wire_d2_38;
	wire [WIDTH-1:0] wire_d2_39;
	wire [WIDTH-1:0] wire_d2_40;
	wire [WIDTH-1:0] wire_d2_41;
	wire [WIDTH-1:0] wire_d2_42;
	wire [WIDTH-1:0] wire_d2_43;
	wire [WIDTH-1:0] wire_d2_44;
	wire [WIDTH-1:0] wire_d2_45;
	wire [WIDTH-1:0] wire_d2_46;
	wire [WIDTH-1:0] wire_d2_47;
	wire [WIDTH-1:0] wire_d2_48;
	wire [WIDTH-1:0] wire_d3_0;
	wire [WIDTH-1:0] wire_d3_1;
	wire [WIDTH-1:0] wire_d3_2;
	wire [WIDTH-1:0] wire_d3_3;
	wire [WIDTH-1:0] wire_d3_4;
	wire [WIDTH-1:0] wire_d3_5;
	wire [WIDTH-1:0] wire_d3_6;
	wire [WIDTH-1:0] wire_d3_7;
	wire [WIDTH-1:0] wire_d3_8;
	wire [WIDTH-1:0] wire_d3_9;
	wire [WIDTH-1:0] wire_d3_10;
	wire [WIDTH-1:0] wire_d3_11;
	wire [WIDTH-1:0] wire_d3_12;
	wire [WIDTH-1:0] wire_d3_13;
	wire [WIDTH-1:0] wire_d3_14;
	wire [WIDTH-1:0] wire_d3_15;
	wire [WIDTH-1:0] wire_d3_16;
	wire [WIDTH-1:0] wire_d3_17;
	wire [WIDTH-1:0] wire_d3_18;
	wire [WIDTH-1:0] wire_d3_19;
	wire [WIDTH-1:0] wire_d3_20;
	wire [WIDTH-1:0] wire_d3_21;
	wire [WIDTH-1:0] wire_d3_22;
	wire [WIDTH-1:0] wire_d3_23;
	wire [WIDTH-1:0] wire_d3_24;
	wire [WIDTH-1:0] wire_d3_25;
	wire [WIDTH-1:0] wire_d3_26;
	wire [WIDTH-1:0] wire_d3_27;
	wire [WIDTH-1:0] wire_d3_28;
	wire [WIDTH-1:0] wire_d3_29;
	wire [WIDTH-1:0] wire_d3_30;
	wire [WIDTH-1:0] wire_d3_31;
	wire [WIDTH-1:0] wire_d3_32;
	wire [WIDTH-1:0] wire_d3_33;
	wire [WIDTH-1:0] wire_d3_34;
	wire [WIDTH-1:0] wire_d3_35;
	wire [WIDTH-1:0] wire_d3_36;
	wire [WIDTH-1:0] wire_d3_37;
	wire [WIDTH-1:0] wire_d3_38;
	wire [WIDTH-1:0] wire_d3_39;
	wire [WIDTH-1:0] wire_d3_40;
	wire [WIDTH-1:0] wire_d3_41;
	wire [WIDTH-1:0] wire_d3_42;
	wire [WIDTH-1:0] wire_d3_43;
	wire [WIDTH-1:0] wire_d3_44;
	wire [WIDTH-1:0] wire_d3_45;
	wire [WIDTH-1:0] wire_d3_46;
	wire [WIDTH-1:0] wire_d3_47;
	wire [WIDTH-1:0] wire_d3_48;
	wire [WIDTH-1:0] wire_d4_0;
	wire [WIDTH-1:0] wire_d4_1;
	wire [WIDTH-1:0] wire_d4_2;
	wire [WIDTH-1:0] wire_d4_3;
	wire [WIDTH-1:0] wire_d4_4;
	wire [WIDTH-1:0] wire_d4_5;
	wire [WIDTH-1:0] wire_d4_6;
	wire [WIDTH-1:0] wire_d4_7;
	wire [WIDTH-1:0] wire_d4_8;
	wire [WIDTH-1:0] wire_d4_9;
	wire [WIDTH-1:0] wire_d4_10;
	wire [WIDTH-1:0] wire_d4_11;
	wire [WIDTH-1:0] wire_d4_12;
	wire [WIDTH-1:0] wire_d4_13;
	wire [WIDTH-1:0] wire_d4_14;
	wire [WIDTH-1:0] wire_d4_15;
	wire [WIDTH-1:0] wire_d4_16;
	wire [WIDTH-1:0] wire_d4_17;
	wire [WIDTH-1:0] wire_d4_18;
	wire [WIDTH-1:0] wire_d4_19;
	wire [WIDTH-1:0] wire_d4_20;
	wire [WIDTH-1:0] wire_d4_21;
	wire [WIDTH-1:0] wire_d4_22;
	wire [WIDTH-1:0] wire_d4_23;
	wire [WIDTH-1:0] wire_d4_24;
	wire [WIDTH-1:0] wire_d4_25;
	wire [WIDTH-1:0] wire_d4_26;
	wire [WIDTH-1:0] wire_d4_27;
	wire [WIDTH-1:0] wire_d4_28;
	wire [WIDTH-1:0] wire_d4_29;
	wire [WIDTH-1:0] wire_d4_30;
	wire [WIDTH-1:0] wire_d4_31;
	wire [WIDTH-1:0] wire_d4_32;
	wire [WIDTH-1:0] wire_d4_33;
	wire [WIDTH-1:0] wire_d4_34;
	wire [WIDTH-1:0] wire_d4_35;
	wire [WIDTH-1:0] wire_d4_36;
	wire [WIDTH-1:0] wire_d4_37;
	wire [WIDTH-1:0] wire_d4_38;
	wire [WIDTH-1:0] wire_d4_39;
	wire [WIDTH-1:0] wire_d4_40;
	wire [WIDTH-1:0] wire_d4_41;
	wire [WIDTH-1:0] wire_d4_42;
	wire [WIDTH-1:0] wire_d4_43;
	wire [WIDTH-1:0] wire_d4_44;
	wire [WIDTH-1:0] wire_d4_45;
	wire [WIDTH-1:0] wire_d4_46;
	wire [WIDTH-1:0] wire_d4_47;
	wire [WIDTH-1:0] wire_d4_48;
	wire [WIDTH-1:0] wire_d5_0;
	wire [WIDTH-1:0] wire_d5_1;
	wire [WIDTH-1:0] wire_d5_2;
	wire [WIDTH-1:0] wire_d5_3;
	wire [WIDTH-1:0] wire_d5_4;
	wire [WIDTH-1:0] wire_d5_5;
	wire [WIDTH-1:0] wire_d5_6;
	wire [WIDTH-1:0] wire_d5_7;
	wire [WIDTH-1:0] wire_d5_8;
	wire [WIDTH-1:0] wire_d5_9;
	wire [WIDTH-1:0] wire_d5_10;
	wire [WIDTH-1:0] wire_d5_11;
	wire [WIDTH-1:0] wire_d5_12;
	wire [WIDTH-1:0] wire_d5_13;
	wire [WIDTH-1:0] wire_d5_14;
	wire [WIDTH-1:0] wire_d5_15;
	wire [WIDTH-1:0] wire_d5_16;
	wire [WIDTH-1:0] wire_d5_17;
	wire [WIDTH-1:0] wire_d5_18;
	wire [WIDTH-1:0] wire_d5_19;
	wire [WIDTH-1:0] wire_d5_20;
	wire [WIDTH-1:0] wire_d5_21;
	wire [WIDTH-1:0] wire_d5_22;
	wire [WIDTH-1:0] wire_d5_23;
	wire [WIDTH-1:0] wire_d5_24;
	wire [WIDTH-1:0] wire_d5_25;
	wire [WIDTH-1:0] wire_d5_26;
	wire [WIDTH-1:0] wire_d5_27;
	wire [WIDTH-1:0] wire_d5_28;
	wire [WIDTH-1:0] wire_d5_29;
	wire [WIDTH-1:0] wire_d5_30;
	wire [WIDTH-1:0] wire_d5_31;
	wire [WIDTH-1:0] wire_d5_32;
	wire [WIDTH-1:0] wire_d5_33;
	wire [WIDTH-1:0] wire_d5_34;
	wire [WIDTH-1:0] wire_d5_35;
	wire [WIDTH-1:0] wire_d5_36;
	wire [WIDTH-1:0] wire_d5_37;
	wire [WIDTH-1:0] wire_d5_38;
	wire [WIDTH-1:0] wire_d5_39;
	wire [WIDTH-1:0] wire_d5_40;
	wire [WIDTH-1:0] wire_d5_41;
	wire [WIDTH-1:0] wire_d5_42;
	wire [WIDTH-1:0] wire_d5_43;
	wire [WIDTH-1:0] wire_d5_44;
	wire [WIDTH-1:0] wire_d5_45;
	wire [WIDTH-1:0] wire_d5_46;
	wire [WIDTH-1:0] wire_d5_47;
	wire [WIDTH-1:0] wire_d5_48;
	wire [WIDTH-1:0] wire_d6_0;
	wire [WIDTH-1:0] wire_d6_1;
	wire [WIDTH-1:0] wire_d6_2;
	wire [WIDTH-1:0] wire_d6_3;
	wire [WIDTH-1:0] wire_d6_4;
	wire [WIDTH-1:0] wire_d6_5;
	wire [WIDTH-1:0] wire_d6_6;
	wire [WIDTH-1:0] wire_d6_7;
	wire [WIDTH-1:0] wire_d6_8;
	wire [WIDTH-1:0] wire_d6_9;
	wire [WIDTH-1:0] wire_d6_10;
	wire [WIDTH-1:0] wire_d6_11;
	wire [WIDTH-1:0] wire_d6_12;
	wire [WIDTH-1:0] wire_d6_13;
	wire [WIDTH-1:0] wire_d6_14;
	wire [WIDTH-1:0] wire_d6_15;
	wire [WIDTH-1:0] wire_d6_16;
	wire [WIDTH-1:0] wire_d6_17;
	wire [WIDTH-1:0] wire_d6_18;
	wire [WIDTH-1:0] wire_d6_19;
	wire [WIDTH-1:0] wire_d6_20;
	wire [WIDTH-1:0] wire_d6_21;
	wire [WIDTH-1:0] wire_d6_22;
	wire [WIDTH-1:0] wire_d6_23;
	wire [WIDTH-1:0] wire_d6_24;
	wire [WIDTH-1:0] wire_d6_25;
	wire [WIDTH-1:0] wire_d6_26;
	wire [WIDTH-1:0] wire_d6_27;
	wire [WIDTH-1:0] wire_d6_28;
	wire [WIDTH-1:0] wire_d6_29;
	wire [WIDTH-1:0] wire_d6_30;
	wire [WIDTH-1:0] wire_d6_31;
	wire [WIDTH-1:0] wire_d6_32;
	wire [WIDTH-1:0] wire_d6_33;
	wire [WIDTH-1:0] wire_d6_34;
	wire [WIDTH-1:0] wire_d6_35;
	wire [WIDTH-1:0] wire_d6_36;
	wire [WIDTH-1:0] wire_d6_37;
	wire [WIDTH-1:0] wire_d6_38;
	wire [WIDTH-1:0] wire_d6_39;
	wire [WIDTH-1:0] wire_d6_40;
	wire [WIDTH-1:0] wire_d6_41;
	wire [WIDTH-1:0] wire_d6_42;
	wire [WIDTH-1:0] wire_d6_43;
	wire [WIDTH-1:0] wire_d6_44;
	wire [WIDTH-1:0] wire_d6_45;
	wire [WIDTH-1:0] wire_d6_46;
	wire [WIDTH-1:0] wire_d6_47;
	wire [WIDTH-1:0] wire_d6_48;
	wire [WIDTH-1:0] wire_d7_0;
	wire [WIDTH-1:0] wire_d7_1;
	wire [WIDTH-1:0] wire_d7_2;
	wire [WIDTH-1:0] wire_d7_3;
	wire [WIDTH-1:0] wire_d7_4;
	wire [WIDTH-1:0] wire_d7_5;
	wire [WIDTH-1:0] wire_d7_6;
	wire [WIDTH-1:0] wire_d7_7;
	wire [WIDTH-1:0] wire_d7_8;
	wire [WIDTH-1:0] wire_d7_9;
	wire [WIDTH-1:0] wire_d7_10;
	wire [WIDTH-1:0] wire_d7_11;
	wire [WIDTH-1:0] wire_d7_12;
	wire [WIDTH-1:0] wire_d7_13;
	wire [WIDTH-1:0] wire_d7_14;
	wire [WIDTH-1:0] wire_d7_15;
	wire [WIDTH-1:0] wire_d7_16;
	wire [WIDTH-1:0] wire_d7_17;
	wire [WIDTH-1:0] wire_d7_18;
	wire [WIDTH-1:0] wire_d7_19;
	wire [WIDTH-1:0] wire_d7_20;
	wire [WIDTH-1:0] wire_d7_21;
	wire [WIDTH-1:0] wire_d7_22;
	wire [WIDTH-1:0] wire_d7_23;
	wire [WIDTH-1:0] wire_d7_24;
	wire [WIDTH-1:0] wire_d7_25;
	wire [WIDTH-1:0] wire_d7_26;
	wire [WIDTH-1:0] wire_d7_27;
	wire [WIDTH-1:0] wire_d7_28;
	wire [WIDTH-1:0] wire_d7_29;
	wire [WIDTH-1:0] wire_d7_30;
	wire [WIDTH-1:0] wire_d7_31;
	wire [WIDTH-1:0] wire_d7_32;
	wire [WIDTH-1:0] wire_d7_33;
	wire [WIDTH-1:0] wire_d7_34;
	wire [WIDTH-1:0] wire_d7_35;
	wire [WIDTH-1:0] wire_d7_36;
	wire [WIDTH-1:0] wire_d7_37;
	wire [WIDTH-1:0] wire_d7_38;
	wire [WIDTH-1:0] wire_d7_39;
	wire [WIDTH-1:0] wire_d7_40;
	wire [WIDTH-1:0] wire_d7_41;
	wire [WIDTH-1:0] wire_d7_42;
	wire [WIDTH-1:0] wire_d7_43;
	wire [WIDTH-1:0] wire_d7_44;
	wire [WIDTH-1:0] wire_d7_45;
	wire [WIDTH-1:0] wire_d7_46;
	wire [WIDTH-1:0] wire_d7_47;
	wire [WIDTH-1:0] wire_d7_48;
	wire [WIDTH-1:0] wire_d8_0;
	wire [WIDTH-1:0] wire_d8_1;
	wire [WIDTH-1:0] wire_d8_2;
	wire [WIDTH-1:0] wire_d8_3;
	wire [WIDTH-1:0] wire_d8_4;
	wire [WIDTH-1:0] wire_d8_5;
	wire [WIDTH-1:0] wire_d8_6;
	wire [WIDTH-1:0] wire_d8_7;
	wire [WIDTH-1:0] wire_d8_8;
	wire [WIDTH-1:0] wire_d8_9;
	wire [WIDTH-1:0] wire_d8_10;
	wire [WIDTH-1:0] wire_d8_11;
	wire [WIDTH-1:0] wire_d8_12;
	wire [WIDTH-1:0] wire_d8_13;
	wire [WIDTH-1:0] wire_d8_14;
	wire [WIDTH-1:0] wire_d8_15;
	wire [WIDTH-1:0] wire_d8_16;
	wire [WIDTH-1:0] wire_d8_17;
	wire [WIDTH-1:0] wire_d8_18;
	wire [WIDTH-1:0] wire_d8_19;
	wire [WIDTH-1:0] wire_d8_20;
	wire [WIDTH-1:0] wire_d8_21;
	wire [WIDTH-1:0] wire_d8_22;
	wire [WIDTH-1:0] wire_d8_23;
	wire [WIDTH-1:0] wire_d8_24;
	wire [WIDTH-1:0] wire_d8_25;
	wire [WIDTH-1:0] wire_d8_26;
	wire [WIDTH-1:0] wire_d8_27;
	wire [WIDTH-1:0] wire_d8_28;
	wire [WIDTH-1:0] wire_d8_29;
	wire [WIDTH-1:0] wire_d8_30;
	wire [WIDTH-1:0] wire_d8_31;
	wire [WIDTH-1:0] wire_d8_32;
	wire [WIDTH-1:0] wire_d8_33;
	wire [WIDTH-1:0] wire_d8_34;
	wire [WIDTH-1:0] wire_d8_35;
	wire [WIDTH-1:0] wire_d8_36;
	wire [WIDTH-1:0] wire_d8_37;
	wire [WIDTH-1:0] wire_d8_38;
	wire [WIDTH-1:0] wire_d8_39;
	wire [WIDTH-1:0] wire_d8_40;
	wire [WIDTH-1:0] wire_d8_41;
	wire [WIDTH-1:0] wire_d8_42;
	wire [WIDTH-1:0] wire_d8_43;
	wire [WIDTH-1:0] wire_d8_44;
	wire [WIDTH-1:0] wire_d8_45;
	wire [WIDTH-1:0] wire_d8_46;
	wire [WIDTH-1:0] wire_d8_47;
	wire [WIDTH-1:0] wire_d8_48;
	wire [WIDTH-1:0] wire_d9_0;
	wire [WIDTH-1:0] wire_d9_1;
	wire [WIDTH-1:0] wire_d9_2;
	wire [WIDTH-1:0] wire_d9_3;
	wire [WIDTH-1:0] wire_d9_4;
	wire [WIDTH-1:0] wire_d9_5;
	wire [WIDTH-1:0] wire_d9_6;
	wire [WIDTH-1:0] wire_d9_7;
	wire [WIDTH-1:0] wire_d9_8;
	wire [WIDTH-1:0] wire_d9_9;
	wire [WIDTH-1:0] wire_d9_10;
	wire [WIDTH-1:0] wire_d9_11;
	wire [WIDTH-1:0] wire_d9_12;
	wire [WIDTH-1:0] wire_d9_13;
	wire [WIDTH-1:0] wire_d9_14;
	wire [WIDTH-1:0] wire_d9_15;
	wire [WIDTH-1:0] wire_d9_16;
	wire [WIDTH-1:0] wire_d9_17;
	wire [WIDTH-1:0] wire_d9_18;
	wire [WIDTH-1:0] wire_d9_19;
	wire [WIDTH-1:0] wire_d9_20;
	wire [WIDTH-1:0] wire_d9_21;
	wire [WIDTH-1:0] wire_d9_22;
	wire [WIDTH-1:0] wire_d9_23;
	wire [WIDTH-1:0] wire_d9_24;
	wire [WIDTH-1:0] wire_d9_25;
	wire [WIDTH-1:0] wire_d9_26;
	wire [WIDTH-1:0] wire_d9_27;
	wire [WIDTH-1:0] wire_d9_28;
	wire [WIDTH-1:0] wire_d9_29;
	wire [WIDTH-1:0] wire_d9_30;
	wire [WIDTH-1:0] wire_d9_31;
	wire [WIDTH-1:0] wire_d9_32;
	wire [WIDTH-1:0] wire_d9_33;
	wire [WIDTH-1:0] wire_d9_34;
	wire [WIDTH-1:0] wire_d9_35;
	wire [WIDTH-1:0] wire_d9_36;
	wire [WIDTH-1:0] wire_d9_37;
	wire [WIDTH-1:0] wire_d9_38;
	wire [WIDTH-1:0] wire_d9_39;
	wire [WIDTH-1:0] wire_d9_40;
	wire [WIDTH-1:0] wire_d9_41;
	wire [WIDTH-1:0] wire_d9_42;
	wire [WIDTH-1:0] wire_d9_43;
	wire [WIDTH-1:0] wire_d9_44;
	wire [WIDTH-1:0] wire_d9_45;
	wire [WIDTH-1:0] wire_d9_46;
	wire [WIDTH-1:0] wire_d9_47;
	wire [WIDTH-1:0] wire_d9_48;
	wire [WIDTH-1:0] wire_d10_0;
	wire [WIDTH-1:0] wire_d10_1;
	wire [WIDTH-1:0] wire_d10_2;
	wire [WIDTH-1:0] wire_d10_3;
	wire [WIDTH-1:0] wire_d10_4;
	wire [WIDTH-1:0] wire_d10_5;
	wire [WIDTH-1:0] wire_d10_6;
	wire [WIDTH-1:0] wire_d10_7;
	wire [WIDTH-1:0] wire_d10_8;
	wire [WIDTH-1:0] wire_d10_9;
	wire [WIDTH-1:0] wire_d10_10;
	wire [WIDTH-1:0] wire_d10_11;
	wire [WIDTH-1:0] wire_d10_12;
	wire [WIDTH-1:0] wire_d10_13;
	wire [WIDTH-1:0] wire_d10_14;
	wire [WIDTH-1:0] wire_d10_15;
	wire [WIDTH-1:0] wire_d10_16;
	wire [WIDTH-1:0] wire_d10_17;
	wire [WIDTH-1:0] wire_d10_18;
	wire [WIDTH-1:0] wire_d10_19;
	wire [WIDTH-1:0] wire_d10_20;
	wire [WIDTH-1:0] wire_d10_21;
	wire [WIDTH-1:0] wire_d10_22;
	wire [WIDTH-1:0] wire_d10_23;
	wire [WIDTH-1:0] wire_d10_24;
	wire [WIDTH-1:0] wire_d10_25;
	wire [WIDTH-1:0] wire_d10_26;
	wire [WIDTH-1:0] wire_d10_27;
	wire [WIDTH-1:0] wire_d10_28;
	wire [WIDTH-1:0] wire_d10_29;
	wire [WIDTH-1:0] wire_d10_30;
	wire [WIDTH-1:0] wire_d10_31;
	wire [WIDTH-1:0] wire_d10_32;
	wire [WIDTH-1:0] wire_d10_33;
	wire [WIDTH-1:0] wire_d10_34;
	wire [WIDTH-1:0] wire_d10_35;
	wire [WIDTH-1:0] wire_d10_36;
	wire [WIDTH-1:0] wire_d10_37;
	wire [WIDTH-1:0] wire_d10_38;
	wire [WIDTH-1:0] wire_d10_39;
	wire [WIDTH-1:0] wire_d10_40;
	wire [WIDTH-1:0] wire_d10_41;
	wire [WIDTH-1:0] wire_d10_42;
	wire [WIDTH-1:0] wire_d10_43;
	wire [WIDTH-1:0] wire_d10_44;
	wire [WIDTH-1:0] wire_d10_45;
	wire [WIDTH-1:0] wire_d10_46;
	wire [WIDTH-1:0] wire_d10_47;
	wire [WIDTH-1:0] wire_d10_48;
	wire [WIDTH-1:0] wire_d11_0;
	wire [WIDTH-1:0] wire_d11_1;
	wire [WIDTH-1:0] wire_d11_2;
	wire [WIDTH-1:0] wire_d11_3;
	wire [WIDTH-1:0] wire_d11_4;
	wire [WIDTH-1:0] wire_d11_5;
	wire [WIDTH-1:0] wire_d11_6;
	wire [WIDTH-1:0] wire_d11_7;
	wire [WIDTH-1:0] wire_d11_8;
	wire [WIDTH-1:0] wire_d11_9;
	wire [WIDTH-1:0] wire_d11_10;
	wire [WIDTH-1:0] wire_d11_11;
	wire [WIDTH-1:0] wire_d11_12;
	wire [WIDTH-1:0] wire_d11_13;
	wire [WIDTH-1:0] wire_d11_14;
	wire [WIDTH-1:0] wire_d11_15;
	wire [WIDTH-1:0] wire_d11_16;
	wire [WIDTH-1:0] wire_d11_17;
	wire [WIDTH-1:0] wire_d11_18;
	wire [WIDTH-1:0] wire_d11_19;
	wire [WIDTH-1:0] wire_d11_20;
	wire [WIDTH-1:0] wire_d11_21;
	wire [WIDTH-1:0] wire_d11_22;
	wire [WIDTH-1:0] wire_d11_23;
	wire [WIDTH-1:0] wire_d11_24;
	wire [WIDTH-1:0] wire_d11_25;
	wire [WIDTH-1:0] wire_d11_26;
	wire [WIDTH-1:0] wire_d11_27;
	wire [WIDTH-1:0] wire_d11_28;
	wire [WIDTH-1:0] wire_d11_29;
	wire [WIDTH-1:0] wire_d11_30;
	wire [WIDTH-1:0] wire_d11_31;
	wire [WIDTH-1:0] wire_d11_32;
	wire [WIDTH-1:0] wire_d11_33;
	wire [WIDTH-1:0] wire_d11_34;
	wire [WIDTH-1:0] wire_d11_35;
	wire [WIDTH-1:0] wire_d11_36;
	wire [WIDTH-1:0] wire_d11_37;
	wire [WIDTH-1:0] wire_d11_38;
	wire [WIDTH-1:0] wire_d11_39;
	wire [WIDTH-1:0] wire_d11_40;
	wire [WIDTH-1:0] wire_d11_41;
	wire [WIDTH-1:0] wire_d11_42;
	wire [WIDTH-1:0] wire_d11_43;
	wire [WIDTH-1:0] wire_d11_44;
	wire [WIDTH-1:0] wire_d11_45;
	wire [WIDTH-1:0] wire_d11_46;
	wire [WIDTH-1:0] wire_d11_47;
	wire [WIDTH-1:0] wire_d11_48;
	wire [WIDTH-1:0] wire_d12_0;
	wire [WIDTH-1:0] wire_d12_1;
	wire [WIDTH-1:0] wire_d12_2;
	wire [WIDTH-1:0] wire_d12_3;
	wire [WIDTH-1:0] wire_d12_4;
	wire [WIDTH-1:0] wire_d12_5;
	wire [WIDTH-1:0] wire_d12_6;
	wire [WIDTH-1:0] wire_d12_7;
	wire [WIDTH-1:0] wire_d12_8;
	wire [WIDTH-1:0] wire_d12_9;
	wire [WIDTH-1:0] wire_d12_10;
	wire [WIDTH-1:0] wire_d12_11;
	wire [WIDTH-1:0] wire_d12_12;
	wire [WIDTH-1:0] wire_d12_13;
	wire [WIDTH-1:0] wire_d12_14;
	wire [WIDTH-1:0] wire_d12_15;
	wire [WIDTH-1:0] wire_d12_16;
	wire [WIDTH-1:0] wire_d12_17;
	wire [WIDTH-1:0] wire_d12_18;
	wire [WIDTH-1:0] wire_d12_19;
	wire [WIDTH-1:0] wire_d12_20;
	wire [WIDTH-1:0] wire_d12_21;
	wire [WIDTH-1:0] wire_d12_22;
	wire [WIDTH-1:0] wire_d12_23;
	wire [WIDTH-1:0] wire_d12_24;
	wire [WIDTH-1:0] wire_d12_25;
	wire [WIDTH-1:0] wire_d12_26;
	wire [WIDTH-1:0] wire_d12_27;
	wire [WIDTH-1:0] wire_d12_28;
	wire [WIDTH-1:0] wire_d12_29;
	wire [WIDTH-1:0] wire_d12_30;
	wire [WIDTH-1:0] wire_d12_31;
	wire [WIDTH-1:0] wire_d12_32;
	wire [WIDTH-1:0] wire_d12_33;
	wire [WIDTH-1:0] wire_d12_34;
	wire [WIDTH-1:0] wire_d12_35;
	wire [WIDTH-1:0] wire_d12_36;
	wire [WIDTH-1:0] wire_d12_37;
	wire [WIDTH-1:0] wire_d12_38;
	wire [WIDTH-1:0] wire_d12_39;
	wire [WIDTH-1:0] wire_d12_40;
	wire [WIDTH-1:0] wire_d12_41;
	wire [WIDTH-1:0] wire_d12_42;
	wire [WIDTH-1:0] wire_d12_43;
	wire [WIDTH-1:0] wire_d12_44;
	wire [WIDTH-1:0] wire_d12_45;
	wire [WIDTH-1:0] wire_d12_46;
	wire [WIDTH-1:0] wire_d12_47;
	wire [WIDTH-1:0] wire_d12_48;
	wire [WIDTH-1:0] wire_d13_0;
	wire [WIDTH-1:0] wire_d13_1;
	wire [WIDTH-1:0] wire_d13_2;
	wire [WIDTH-1:0] wire_d13_3;
	wire [WIDTH-1:0] wire_d13_4;
	wire [WIDTH-1:0] wire_d13_5;
	wire [WIDTH-1:0] wire_d13_6;
	wire [WIDTH-1:0] wire_d13_7;
	wire [WIDTH-1:0] wire_d13_8;
	wire [WIDTH-1:0] wire_d13_9;
	wire [WIDTH-1:0] wire_d13_10;
	wire [WIDTH-1:0] wire_d13_11;
	wire [WIDTH-1:0] wire_d13_12;
	wire [WIDTH-1:0] wire_d13_13;
	wire [WIDTH-1:0] wire_d13_14;
	wire [WIDTH-1:0] wire_d13_15;
	wire [WIDTH-1:0] wire_d13_16;
	wire [WIDTH-1:0] wire_d13_17;
	wire [WIDTH-1:0] wire_d13_18;
	wire [WIDTH-1:0] wire_d13_19;
	wire [WIDTH-1:0] wire_d13_20;
	wire [WIDTH-1:0] wire_d13_21;
	wire [WIDTH-1:0] wire_d13_22;
	wire [WIDTH-1:0] wire_d13_23;
	wire [WIDTH-1:0] wire_d13_24;
	wire [WIDTH-1:0] wire_d13_25;
	wire [WIDTH-1:0] wire_d13_26;
	wire [WIDTH-1:0] wire_d13_27;
	wire [WIDTH-1:0] wire_d13_28;
	wire [WIDTH-1:0] wire_d13_29;
	wire [WIDTH-1:0] wire_d13_30;
	wire [WIDTH-1:0] wire_d13_31;
	wire [WIDTH-1:0] wire_d13_32;
	wire [WIDTH-1:0] wire_d13_33;
	wire [WIDTH-1:0] wire_d13_34;
	wire [WIDTH-1:0] wire_d13_35;
	wire [WIDTH-1:0] wire_d13_36;
	wire [WIDTH-1:0] wire_d13_37;
	wire [WIDTH-1:0] wire_d13_38;
	wire [WIDTH-1:0] wire_d13_39;
	wire [WIDTH-1:0] wire_d13_40;
	wire [WIDTH-1:0] wire_d13_41;
	wire [WIDTH-1:0] wire_d13_42;
	wire [WIDTH-1:0] wire_d13_43;
	wire [WIDTH-1:0] wire_d13_44;
	wire [WIDTH-1:0] wire_d13_45;
	wire [WIDTH-1:0] wire_d13_46;
	wire [WIDTH-1:0] wire_d13_47;
	wire [WIDTH-1:0] wire_d13_48;
	wire [WIDTH-1:0] wire_d14_0;
	wire [WIDTH-1:0] wire_d14_1;
	wire [WIDTH-1:0] wire_d14_2;
	wire [WIDTH-1:0] wire_d14_3;
	wire [WIDTH-1:0] wire_d14_4;
	wire [WIDTH-1:0] wire_d14_5;
	wire [WIDTH-1:0] wire_d14_6;
	wire [WIDTH-1:0] wire_d14_7;
	wire [WIDTH-1:0] wire_d14_8;
	wire [WIDTH-1:0] wire_d14_9;
	wire [WIDTH-1:0] wire_d14_10;
	wire [WIDTH-1:0] wire_d14_11;
	wire [WIDTH-1:0] wire_d14_12;
	wire [WIDTH-1:0] wire_d14_13;
	wire [WIDTH-1:0] wire_d14_14;
	wire [WIDTH-1:0] wire_d14_15;
	wire [WIDTH-1:0] wire_d14_16;
	wire [WIDTH-1:0] wire_d14_17;
	wire [WIDTH-1:0] wire_d14_18;
	wire [WIDTH-1:0] wire_d14_19;
	wire [WIDTH-1:0] wire_d14_20;
	wire [WIDTH-1:0] wire_d14_21;
	wire [WIDTH-1:0] wire_d14_22;
	wire [WIDTH-1:0] wire_d14_23;
	wire [WIDTH-1:0] wire_d14_24;
	wire [WIDTH-1:0] wire_d14_25;
	wire [WIDTH-1:0] wire_d14_26;
	wire [WIDTH-1:0] wire_d14_27;
	wire [WIDTH-1:0] wire_d14_28;
	wire [WIDTH-1:0] wire_d14_29;
	wire [WIDTH-1:0] wire_d14_30;
	wire [WIDTH-1:0] wire_d14_31;
	wire [WIDTH-1:0] wire_d14_32;
	wire [WIDTH-1:0] wire_d14_33;
	wire [WIDTH-1:0] wire_d14_34;
	wire [WIDTH-1:0] wire_d14_35;
	wire [WIDTH-1:0] wire_d14_36;
	wire [WIDTH-1:0] wire_d14_37;
	wire [WIDTH-1:0] wire_d14_38;
	wire [WIDTH-1:0] wire_d14_39;
	wire [WIDTH-1:0] wire_d14_40;
	wire [WIDTH-1:0] wire_d14_41;
	wire [WIDTH-1:0] wire_d14_42;
	wire [WIDTH-1:0] wire_d14_43;
	wire [WIDTH-1:0] wire_d14_44;
	wire [WIDTH-1:0] wire_d14_45;
	wire [WIDTH-1:0] wire_d14_46;
	wire [WIDTH-1:0] wire_d14_47;
	wire [WIDTH-1:0] wire_d14_48;
	wire [WIDTH-1:0] wire_d15_0;
	wire [WIDTH-1:0] wire_d15_1;
	wire [WIDTH-1:0] wire_d15_2;
	wire [WIDTH-1:0] wire_d15_3;
	wire [WIDTH-1:0] wire_d15_4;
	wire [WIDTH-1:0] wire_d15_5;
	wire [WIDTH-1:0] wire_d15_6;
	wire [WIDTH-1:0] wire_d15_7;
	wire [WIDTH-1:0] wire_d15_8;
	wire [WIDTH-1:0] wire_d15_9;
	wire [WIDTH-1:0] wire_d15_10;
	wire [WIDTH-1:0] wire_d15_11;
	wire [WIDTH-1:0] wire_d15_12;
	wire [WIDTH-1:0] wire_d15_13;
	wire [WIDTH-1:0] wire_d15_14;
	wire [WIDTH-1:0] wire_d15_15;
	wire [WIDTH-1:0] wire_d15_16;
	wire [WIDTH-1:0] wire_d15_17;
	wire [WIDTH-1:0] wire_d15_18;
	wire [WIDTH-1:0] wire_d15_19;
	wire [WIDTH-1:0] wire_d15_20;
	wire [WIDTH-1:0] wire_d15_21;
	wire [WIDTH-1:0] wire_d15_22;
	wire [WIDTH-1:0] wire_d15_23;
	wire [WIDTH-1:0] wire_d15_24;
	wire [WIDTH-1:0] wire_d15_25;
	wire [WIDTH-1:0] wire_d15_26;
	wire [WIDTH-1:0] wire_d15_27;
	wire [WIDTH-1:0] wire_d15_28;
	wire [WIDTH-1:0] wire_d15_29;
	wire [WIDTH-1:0] wire_d15_30;
	wire [WIDTH-1:0] wire_d15_31;
	wire [WIDTH-1:0] wire_d15_32;
	wire [WIDTH-1:0] wire_d15_33;
	wire [WIDTH-1:0] wire_d15_34;
	wire [WIDTH-1:0] wire_d15_35;
	wire [WIDTH-1:0] wire_d15_36;
	wire [WIDTH-1:0] wire_d15_37;
	wire [WIDTH-1:0] wire_d15_38;
	wire [WIDTH-1:0] wire_d15_39;
	wire [WIDTH-1:0] wire_d15_40;
	wire [WIDTH-1:0] wire_d15_41;
	wire [WIDTH-1:0] wire_d15_42;
	wire [WIDTH-1:0] wire_d15_43;
	wire [WIDTH-1:0] wire_d15_44;
	wire [WIDTH-1:0] wire_d15_45;
	wire [WIDTH-1:0] wire_d15_46;
	wire [WIDTH-1:0] wire_d15_47;
	wire [WIDTH-1:0] wire_d15_48;
	wire [WIDTH-1:0] wire_d16_0;
	wire [WIDTH-1:0] wire_d16_1;
	wire [WIDTH-1:0] wire_d16_2;
	wire [WIDTH-1:0] wire_d16_3;
	wire [WIDTH-1:0] wire_d16_4;
	wire [WIDTH-1:0] wire_d16_5;
	wire [WIDTH-1:0] wire_d16_6;
	wire [WIDTH-1:0] wire_d16_7;
	wire [WIDTH-1:0] wire_d16_8;
	wire [WIDTH-1:0] wire_d16_9;
	wire [WIDTH-1:0] wire_d16_10;
	wire [WIDTH-1:0] wire_d16_11;
	wire [WIDTH-1:0] wire_d16_12;
	wire [WIDTH-1:0] wire_d16_13;
	wire [WIDTH-1:0] wire_d16_14;
	wire [WIDTH-1:0] wire_d16_15;
	wire [WIDTH-1:0] wire_d16_16;
	wire [WIDTH-1:0] wire_d16_17;
	wire [WIDTH-1:0] wire_d16_18;
	wire [WIDTH-1:0] wire_d16_19;
	wire [WIDTH-1:0] wire_d16_20;
	wire [WIDTH-1:0] wire_d16_21;
	wire [WIDTH-1:0] wire_d16_22;
	wire [WIDTH-1:0] wire_d16_23;
	wire [WIDTH-1:0] wire_d16_24;
	wire [WIDTH-1:0] wire_d16_25;
	wire [WIDTH-1:0] wire_d16_26;
	wire [WIDTH-1:0] wire_d16_27;
	wire [WIDTH-1:0] wire_d16_28;
	wire [WIDTH-1:0] wire_d16_29;
	wire [WIDTH-1:0] wire_d16_30;
	wire [WIDTH-1:0] wire_d16_31;
	wire [WIDTH-1:0] wire_d16_32;
	wire [WIDTH-1:0] wire_d16_33;
	wire [WIDTH-1:0] wire_d16_34;
	wire [WIDTH-1:0] wire_d16_35;
	wire [WIDTH-1:0] wire_d16_36;
	wire [WIDTH-1:0] wire_d16_37;
	wire [WIDTH-1:0] wire_d16_38;
	wire [WIDTH-1:0] wire_d16_39;
	wire [WIDTH-1:0] wire_d16_40;
	wire [WIDTH-1:0] wire_d16_41;
	wire [WIDTH-1:0] wire_d16_42;
	wire [WIDTH-1:0] wire_d16_43;
	wire [WIDTH-1:0] wire_d16_44;
	wire [WIDTH-1:0] wire_d16_45;
	wire [WIDTH-1:0] wire_d16_46;
	wire [WIDTH-1:0] wire_d16_47;
	wire [WIDTH-1:0] wire_d16_48;
	wire [WIDTH-1:0] wire_d17_0;
	wire [WIDTH-1:0] wire_d17_1;
	wire [WIDTH-1:0] wire_d17_2;
	wire [WIDTH-1:0] wire_d17_3;
	wire [WIDTH-1:0] wire_d17_4;
	wire [WIDTH-1:0] wire_d17_5;
	wire [WIDTH-1:0] wire_d17_6;
	wire [WIDTH-1:0] wire_d17_7;
	wire [WIDTH-1:0] wire_d17_8;
	wire [WIDTH-1:0] wire_d17_9;
	wire [WIDTH-1:0] wire_d17_10;
	wire [WIDTH-1:0] wire_d17_11;
	wire [WIDTH-1:0] wire_d17_12;
	wire [WIDTH-1:0] wire_d17_13;
	wire [WIDTH-1:0] wire_d17_14;
	wire [WIDTH-1:0] wire_d17_15;
	wire [WIDTH-1:0] wire_d17_16;
	wire [WIDTH-1:0] wire_d17_17;
	wire [WIDTH-1:0] wire_d17_18;
	wire [WIDTH-1:0] wire_d17_19;
	wire [WIDTH-1:0] wire_d17_20;
	wire [WIDTH-1:0] wire_d17_21;
	wire [WIDTH-1:0] wire_d17_22;
	wire [WIDTH-1:0] wire_d17_23;
	wire [WIDTH-1:0] wire_d17_24;
	wire [WIDTH-1:0] wire_d17_25;
	wire [WIDTH-1:0] wire_d17_26;
	wire [WIDTH-1:0] wire_d17_27;
	wire [WIDTH-1:0] wire_d17_28;
	wire [WIDTH-1:0] wire_d17_29;
	wire [WIDTH-1:0] wire_d17_30;
	wire [WIDTH-1:0] wire_d17_31;
	wire [WIDTH-1:0] wire_d17_32;
	wire [WIDTH-1:0] wire_d17_33;
	wire [WIDTH-1:0] wire_d17_34;
	wire [WIDTH-1:0] wire_d17_35;
	wire [WIDTH-1:0] wire_d17_36;
	wire [WIDTH-1:0] wire_d17_37;
	wire [WIDTH-1:0] wire_d17_38;
	wire [WIDTH-1:0] wire_d17_39;
	wire [WIDTH-1:0] wire_d17_40;
	wire [WIDTH-1:0] wire_d17_41;
	wire [WIDTH-1:0] wire_d17_42;
	wire [WIDTH-1:0] wire_d17_43;
	wire [WIDTH-1:0] wire_d17_44;
	wire [WIDTH-1:0] wire_d17_45;
	wire [WIDTH-1:0] wire_d17_46;
	wire [WIDTH-1:0] wire_d17_47;
	wire [WIDTH-1:0] wire_d17_48;
	wire [WIDTH-1:0] wire_d18_0;
	wire [WIDTH-1:0] wire_d18_1;
	wire [WIDTH-1:0] wire_d18_2;
	wire [WIDTH-1:0] wire_d18_3;
	wire [WIDTH-1:0] wire_d18_4;
	wire [WIDTH-1:0] wire_d18_5;
	wire [WIDTH-1:0] wire_d18_6;
	wire [WIDTH-1:0] wire_d18_7;
	wire [WIDTH-1:0] wire_d18_8;
	wire [WIDTH-1:0] wire_d18_9;
	wire [WIDTH-1:0] wire_d18_10;
	wire [WIDTH-1:0] wire_d18_11;
	wire [WIDTH-1:0] wire_d18_12;
	wire [WIDTH-1:0] wire_d18_13;
	wire [WIDTH-1:0] wire_d18_14;
	wire [WIDTH-1:0] wire_d18_15;
	wire [WIDTH-1:0] wire_d18_16;
	wire [WIDTH-1:0] wire_d18_17;
	wire [WIDTH-1:0] wire_d18_18;
	wire [WIDTH-1:0] wire_d18_19;
	wire [WIDTH-1:0] wire_d18_20;
	wire [WIDTH-1:0] wire_d18_21;
	wire [WIDTH-1:0] wire_d18_22;
	wire [WIDTH-1:0] wire_d18_23;
	wire [WIDTH-1:0] wire_d18_24;
	wire [WIDTH-1:0] wire_d18_25;
	wire [WIDTH-1:0] wire_d18_26;
	wire [WIDTH-1:0] wire_d18_27;
	wire [WIDTH-1:0] wire_d18_28;
	wire [WIDTH-1:0] wire_d18_29;
	wire [WIDTH-1:0] wire_d18_30;
	wire [WIDTH-1:0] wire_d18_31;
	wire [WIDTH-1:0] wire_d18_32;
	wire [WIDTH-1:0] wire_d18_33;
	wire [WIDTH-1:0] wire_d18_34;
	wire [WIDTH-1:0] wire_d18_35;
	wire [WIDTH-1:0] wire_d18_36;
	wire [WIDTH-1:0] wire_d18_37;
	wire [WIDTH-1:0] wire_d18_38;
	wire [WIDTH-1:0] wire_d18_39;
	wire [WIDTH-1:0] wire_d18_40;
	wire [WIDTH-1:0] wire_d18_41;
	wire [WIDTH-1:0] wire_d18_42;
	wire [WIDTH-1:0] wire_d18_43;
	wire [WIDTH-1:0] wire_d18_44;
	wire [WIDTH-1:0] wire_d18_45;
	wire [WIDTH-1:0] wire_d18_46;
	wire [WIDTH-1:0] wire_d18_47;
	wire [WIDTH-1:0] wire_d18_48;
	wire [WIDTH-1:0] wire_d19_0;
	wire [WIDTH-1:0] wire_d19_1;
	wire [WIDTH-1:0] wire_d19_2;
	wire [WIDTH-1:0] wire_d19_3;
	wire [WIDTH-1:0] wire_d19_4;
	wire [WIDTH-1:0] wire_d19_5;
	wire [WIDTH-1:0] wire_d19_6;
	wire [WIDTH-1:0] wire_d19_7;
	wire [WIDTH-1:0] wire_d19_8;
	wire [WIDTH-1:0] wire_d19_9;
	wire [WIDTH-1:0] wire_d19_10;
	wire [WIDTH-1:0] wire_d19_11;
	wire [WIDTH-1:0] wire_d19_12;
	wire [WIDTH-1:0] wire_d19_13;
	wire [WIDTH-1:0] wire_d19_14;
	wire [WIDTH-1:0] wire_d19_15;
	wire [WIDTH-1:0] wire_d19_16;
	wire [WIDTH-1:0] wire_d19_17;
	wire [WIDTH-1:0] wire_d19_18;
	wire [WIDTH-1:0] wire_d19_19;
	wire [WIDTH-1:0] wire_d19_20;
	wire [WIDTH-1:0] wire_d19_21;
	wire [WIDTH-1:0] wire_d19_22;
	wire [WIDTH-1:0] wire_d19_23;
	wire [WIDTH-1:0] wire_d19_24;
	wire [WIDTH-1:0] wire_d19_25;
	wire [WIDTH-1:0] wire_d19_26;
	wire [WIDTH-1:0] wire_d19_27;
	wire [WIDTH-1:0] wire_d19_28;
	wire [WIDTH-1:0] wire_d19_29;
	wire [WIDTH-1:0] wire_d19_30;
	wire [WIDTH-1:0] wire_d19_31;
	wire [WIDTH-1:0] wire_d19_32;
	wire [WIDTH-1:0] wire_d19_33;
	wire [WIDTH-1:0] wire_d19_34;
	wire [WIDTH-1:0] wire_d19_35;
	wire [WIDTH-1:0] wire_d19_36;
	wire [WIDTH-1:0] wire_d19_37;
	wire [WIDTH-1:0] wire_d19_38;
	wire [WIDTH-1:0] wire_d19_39;
	wire [WIDTH-1:0] wire_d19_40;
	wire [WIDTH-1:0] wire_d19_41;
	wire [WIDTH-1:0] wire_d19_42;
	wire [WIDTH-1:0] wire_d19_43;
	wire [WIDTH-1:0] wire_d19_44;
	wire [WIDTH-1:0] wire_d19_45;
	wire [WIDTH-1:0] wire_d19_46;
	wire [WIDTH-1:0] wire_d19_47;
	wire [WIDTH-1:0] wire_d19_48;
	wire [WIDTH-1:0] wire_d20_0;
	wire [WIDTH-1:0] wire_d20_1;
	wire [WIDTH-1:0] wire_d20_2;
	wire [WIDTH-1:0] wire_d20_3;
	wire [WIDTH-1:0] wire_d20_4;
	wire [WIDTH-1:0] wire_d20_5;
	wire [WIDTH-1:0] wire_d20_6;
	wire [WIDTH-1:0] wire_d20_7;
	wire [WIDTH-1:0] wire_d20_8;
	wire [WIDTH-1:0] wire_d20_9;
	wire [WIDTH-1:0] wire_d20_10;
	wire [WIDTH-1:0] wire_d20_11;
	wire [WIDTH-1:0] wire_d20_12;
	wire [WIDTH-1:0] wire_d20_13;
	wire [WIDTH-1:0] wire_d20_14;
	wire [WIDTH-1:0] wire_d20_15;
	wire [WIDTH-1:0] wire_d20_16;
	wire [WIDTH-1:0] wire_d20_17;
	wire [WIDTH-1:0] wire_d20_18;
	wire [WIDTH-1:0] wire_d20_19;
	wire [WIDTH-1:0] wire_d20_20;
	wire [WIDTH-1:0] wire_d20_21;
	wire [WIDTH-1:0] wire_d20_22;
	wire [WIDTH-1:0] wire_d20_23;
	wire [WIDTH-1:0] wire_d20_24;
	wire [WIDTH-1:0] wire_d20_25;
	wire [WIDTH-1:0] wire_d20_26;
	wire [WIDTH-1:0] wire_d20_27;
	wire [WIDTH-1:0] wire_d20_28;
	wire [WIDTH-1:0] wire_d20_29;
	wire [WIDTH-1:0] wire_d20_30;
	wire [WIDTH-1:0] wire_d20_31;
	wire [WIDTH-1:0] wire_d20_32;
	wire [WIDTH-1:0] wire_d20_33;
	wire [WIDTH-1:0] wire_d20_34;
	wire [WIDTH-1:0] wire_d20_35;
	wire [WIDTH-1:0] wire_d20_36;
	wire [WIDTH-1:0] wire_d20_37;
	wire [WIDTH-1:0] wire_d20_38;
	wire [WIDTH-1:0] wire_d20_39;
	wire [WIDTH-1:0] wire_d20_40;
	wire [WIDTH-1:0] wire_d20_41;
	wire [WIDTH-1:0] wire_d20_42;
	wire [WIDTH-1:0] wire_d20_43;
	wire [WIDTH-1:0] wire_d20_44;
	wire [WIDTH-1:0] wire_d20_45;
	wire [WIDTH-1:0] wire_d20_46;
	wire [WIDTH-1:0] wire_d20_47;
	wire [WIDTH-1:0] wire_d20_48;
	wire [WIDTH-1:0] wire_d21_0;
	wire [WIDTH-1:0] wire_d21_1;
	wire [WIDTH-1:0] wire_d21_2;
	wire [WIDTH-1:0] wire_d21_3;
	wire [WIDTH-1:0] wire_d21_4;
	wire [WIDTH-1:0] wire_d21_5;
	wire [WIDTH-1:0] wire_d21_6;
	wire [WIDTH-1:0] wire_d21_7;
	wire [WIDTH-1:0] wire_d21_8;
	wire [WIDTH-1:0] wire_d21_9;
	wire [WIDTH-1:0] wire_d21_10;
	wire [WIDTH-1:0] wire_d21_11;
	wire [WIDTH-1:0] wire_d21_12;
	wire [WIDTH-1:0] wire_d21_13;
	wire [WIDTH-1:0] wire_d21_14;
	wire [WIDTH-1:0] wire_d21_15;
	wire [WIDTH-1:0] wire_d21_16;
	wire [WIDTH-1:0] wire_d21_17;
	wire [WIDTH-1:0] wire_d21_18;
	wire [WIDTH-1:0] wire_d21_19;
	wire [WIDTH-1:0] wire_d21_20;
	wire [WIDTH-1:0] wire_d21_21;
	wire [WIDTH-1:0] wire_d21_22;
	wire [WIDTH-1:0] wire_d21_23;
	wire [WIDTH-1:0] wire_d21_24;
	wire [WIDTH-1:0] wire_d21_25;
	wire [WIDTH-1:0] wire_d21_26;
	wire [WIDTH-1:0] wire_d21_27;
	wire [WIDTH-1:0] wire_d21_28;
	wire [WIDTH-1:0] wire_d21_29;
	wire [WIDTH-1:0] wire_d21_30;
	wire [WIDTH-1:0] wire_d21_31;
	wire [WIDTH-1:0] wire_d21_32;
	wire [WIDTH-1:0] wire_d21_33;
	wire [WIDTH-1:0] wire_d21_34;
	wire [WIDTH-1:0] wire_d21_35;
	wire [WIDTH-1:0] wire_d21_36;
	wire [WIDTH-1:0] wire_d21_37;
	wire [WIDTH-1:0] wire_d21_38;
	wire [WIDTH-1:0] wire_d21_39;
	wire [WIDTH-1:0] wire_d21_40;
	wire [WIDTH-1:0] wire_d21_41;
	wire [WIDTH-1:0] wire_d21_42;
	wire [WIDTH-1:0] wire_d21_43;
	wire [WIDTH-1:0] wire_d21_44;
	wire [WIDTH-1:0] wire_d21_45;
	wire [WIDTH-1:0] wire_d21_46;
	wire [WIDTH-1:0] wire_d21_47;
	wire [WIDTH-1:0] wire_d21_48;
	wire [WIDTH-1:0] wire_d22_0;
	wire [WIDTH-1:0] wire_d22_1;
	wire [WIDTH-1:0] wire_d22_2;
	wire [WIDTH-1:0] wire_d22_3;
	wire [WIDTH-1:0] wire_d22_4;
	wire [WIDTH-1:0] wire_d22_5;
	wire [WIDTH-1:0] wire_d22_6;
	wire [WIDTH-1:0] wire_d22_7;
	wire [WIDTH-1:0] wire_d22_8;
	wire [WIDTH-1:0] wire_d22_9;
	wire [WIDTH-1:0] wire_d22_10;
	wire [WIDTH-1:0] wire_d22_11;
	wire [WIDTH-1:0] wire_d22_12;
	wire [WIDTH-1:0] wire_d22_13;
	wire [WIDTH-1:0] wire_d22_14;
	wire [WIDTH-1:0] wire_d22_15;
	wire [WIDTH-1:0] wire_d22_16;
	wire [WIDTH-1:0] wire_d22_17;
	wire [WIDTH-1:0] wire_d22_18;
	wire [WIDTH-1:0] wire_d22_19;
	wire [WIDTH-1:0] wire_d22_20;
	wire [WIDTH-1:0] wire_d22_21;
	wire [WIDTH-1:0] wire_d22_22;
	wire [WIDTH-1:0] wire_d22_23;
	wire [WIDTH-1:0] wire_d22_24;
	wire [WIDTH-1:0] wire_d22_25;
	wire [WIDTH-1:0] wire_d22_26;
	wire [WIDTH-1:0] wire_d22_27;
	wire [WIDTH-1:0] wire_d22_28;
	wire [WIDTH-1:0] wire_d22_29;
	wire [WIDTH-1:0] wire_d22_30;
	wire [WIDTH-1:0] wire_d22_31;
	wire [WIDTH-1:0] wire_d22_32;
	wire [WIDTH-1:0] wire_d22_33;
	wire [WIDTH-1:0] wire_d22_34;
	wire [WIDTH-1:0] wire_d22_35;
	wire [WIDTH-1:0] wire_d22_36;
	wire [WIDTH-1:0] wire_d22_37;
	wire [WIDTH-1:0] wire_d22_38;
	wire [WIDTH-1:0] wire_d22_39;
	wire [WIDTH-1:0] wire_d22_40;
	wire [WIDTH-1:0] wire_d22_41;
	wire [WIDTH-1:0] wire_d22_42;
	wire [WIDTH-1:0] wire_d22_43;
	wire [WIDTH-1:0] wire_d22_44;
	wire [WIDTH-1:0] wire_d22_45;
	wire [WIDTH-1:0] wire_d22_46;
	wire [WIDTH-1:0] wire_d22_47;
	wire [WIDTH-1:0] wire_d22_48;
	wire [WIDTH-1:0] wire_d23_0;
	wire [WIDTH-1:0] wire_d23_1;
	wire [WIDTH-1:0] wire_d23_2;
	wire [WIDTH-1:0] wire_d23_3;
	wire [WIDTH-1:0] wire_d23_4;
	wire [WIDTH-1:0] wire_d23_5;
	wire [WIDTH-1:0] wire_d23_6;
	wire [WIDTH-1:0] wire_d23_7;
	wire [WIDTH-1:0] wire_d23_8;
	wire [WIDTH-1:0] wire_d23_9;
	wire [WIDTH-1:0] wire_d23_10;
	wire [WIDTH-1:0] wire_d23_11;
	wire [WIDTH-1:0] wire_d23_12;
	wire [WIDTH-1:0] wire_d23_13;
	wire [WIDTH-1:0] wire_d23_14;
	wire [WIDTH-1:0] wire_d23_15;
	wire [WIDTH-1:0] wire_d23_16;
	wire [WIDTH-1:0] wire_d23_17;
	wire [WIDTH-1:0] wire_d23_18;
	wire [WIDTH-1:0] wire_d23_19;
	wire [WIDTH-1:0] wire_d23_20;
	wire [WIDTH-1:0] wire_d23_21;
	wire [WIDTH-1:0] wire_d23_22;
	wire [WIDTH-1:0] wire_d23_23;
	wire [WIDTH-1:0] wire_d23_24;
	wire [WIDTH-1:0] wire_d23_25;
	wire [WIDTH-1:0] wire_d23_26;
	wire [WIDTH-1:0] wire_d23_27;
	wire [WIDTH-1:0] wire_d23_28;
	wire [WIDTH-1:0] wire_d23_29;
	wire [WIDTH-1:0] wire_d23_30;
	wire [WIDTH-1:0] wire_d23_31;
	wire [WIDTH-1:0] wire_d23_32;
	wire [WIDTH-1:0] wire_d23_33;
	wire [WIDTH-1:0] wire_d23_34;
	wire [WIDTH-1:0] wire_d23_35;
	wire [WIDTH-1:0] wire_d23_36;
	wire [WIDTH-1:0] wire_d23_37;
	wire [WIDTH-1:0] wire_d23_38;
	wire [WIDTH-1:0] wire_d23_39;
	wire [WIDTH-1:0] wire_d23_40;
	wire [WIDTH-1:0] wire_d23_41;
	wire [WIDTH-1:0] wire_d23_42;
	wire [WIDTH-1:0] wire_d23_43;
	wire [WIDTH-1:0] wire_d23_44;
	wire [WIDTH-1:0] wire_d23_45;
	wire [WIDTH-1:0] wire_d23_46;
	wire [WIDTH-1:0] wire_d23_47;
	wire [WIDTH-1:0] wire_d23_48;
	wire [WIDTH-1:0] wire_d24_0;
	wire [WIDTH-1:0] wire_d24_1;
	wire [WIDTH-1:0] wire_d24_2;
	wire [WIDTH-1:0] wire_d24_3;
	wire [WIDTH-1:0] wire_d24_4;
	wire [WIDTH-1:0] wire_d24_5;
	wire [WIDTH-1:0] wire_d24_6;
	wire [WIDTH-1:0] wire_d24_7;
	wire [WIDTH-1:0] wire_d24_8;
	wire [WIDTH-1:0] wire_d24_9;
	wire [WIDTH-1:0] wire_d24_10;
	wire [WIDTH-1:0] wire_d24_11;
	wire [WIDTH-1:0] wire_d24_12;
	wire [WIDTH-1:0] wire_d24_13;
	wire [WIDTH-1:0] wire_d24_14;
	wire [WIDTH-1:0] wire_d24_15;
	wire [WIDTH-1:0] wire_d24_16;
	wire [WIDTH-1:0] wire_d24_17;
	wire [WIDTH-1:0] wire_d24_18;
	wire [WIDTH-1:0] wire_d24_19;
	wire [WIDTH-1:0] wire_d24_20;
	wire [WIDTH-1:0] wire_d24_21;
	wire [WIDTH-1:0] wire_d24_22;
	wire [WIDTH-1:0] wire_d24_23;
	wire [WIDTH-1:0] wire_d24_24;
	wire [WIDTH-1:0] wire_d24_25;
	wire [WIDTH-1:0] wire_d24_26;
	wire [WIDTH-1:0] wire_d24_27;
	wire [WIDTH-1:0] wire_d24_28;
	wire [WIDTH-1:0] wire_d24_29;
	wire [WIDTH-1:0] wire_d24_30;
	wire [WIDTH-1:0] wire_d24_31;
	wire [WIDTH-1:0] wire_d24_32;
	wire [WIDTH-1:0] wire_d24_33;
	wire [WIDTH-1:0] wire_d24_34;
	wire [WIDTH-1:0] wire_d24_35;
	wire [WIDTH-1:0] wire_d24_36;
	wire [WIDTH-1:0] wire_d24_37;
	wire [WIDTH-1:0] wire_d24_38;
	wire [WIDTH-1:0] wire_d24_39;
	wire [WIDTH-1:0] wire_d24_40;
	wire [WIDTH-1:0] wire_d24_41;
	wire [WIDTH-1:0] wire_d24_42;
	wire [WIDTH-1:0] wire_d24_43;
	wire [WIDTH-1:0] wire_d24_44;
	wire [WIDTH-1:0] wire_d24_45;
	wire [WIDTH-1:0] wire_d24_46;
	wire [WIDTH-1:0] wire_d24_47;
	wire [WIDTH-1:0] wire_d24_48;
	wire [WIDTH-1:0] wire_d25_0;
	wire [WIDTH-1:0] wire_d25_1;
	wire [WIDTH-1:0] wire_d25_2;
	wire [WIDTH-1:0] wire_d25_3;
	wire [WIDTH-1:0] wire_d25_4;
	wire [WIDTH-1:0] wire_d25_5;
	wire [WIDTH-1:0] wire_d25_6;
	wire [WIDTH-1:0] wire_d25_7;
	wire [WIDTH-1:0] wire_d25_8;
	wire [WIDTH-1:0] wire_d25_9;
	wire [WIDTH-1:0] wire_d25_10;
	wire [WIDTH-1:0] wire_d25_11;
	wire [WIDTH-1:0] wire_d25_12;
	wire [WIDTH-1:0] wire_d25_13;
	wire [WIDTH-1:0] wire_d25_14;
	wire [WIDTH-1:0] wire_d25_15;
	wire [WIDTH-1:0] wire_d25_16;
	wire [WIDTH-1:0] wire_d25_17;
	wire [WIDTH-1:0] wire_d25_18;
	wire [WIDTH-1:0] wire_d25_19;
	wire [WIDTH-1:0] wire_d25_20;
	wire [WIDTH-1:0] wire_d25_21;
	wire [WIDTH-1:0] wire_d25_22;
	wire [WIDTH-1:0] wire_d25_23;
	wire [WIDTH-1:0] wire_d25_24;
	wire [WIDTH-1:0] wire_d25_25;
	wire [WIDTH-1:0] wire_d25_26;
	wire [WIDTH-1:0] wire_d25_27;
	wire [WIDTH-1:0] wire_d25_28;
	wire [WIDTH-1:0] wire_d25_29;
	wire [WIDTH-1:0] wire_d25_30;
	wire [WIDTH-1:0] wire_d25_31;
	wire [WIDTH-1:0] wire_d25_32;
	wire [WIDTH-1:0] wire_d25_33;
	wire [WIDTH-1:0] wire_d25_34;
	wire [WIDTH-1:0] wire_d25_35;
	wire [WIDTH-1:0] wire_d25_36;
	wire [WIDTH-1:0] wire_d25_37;
	wire [WIDTH-1:0] wire_d25_38;
	wire [WIDTH-1:0] wire_d25_39;
	wire [WIDTH-1:0] wire_d25_40;
	wire [WIDTH-1:0] wire_d25_41;
	wire [WIDTH-1:0] wire_d25_42;
	wire [WIDTH-1:0] wire_d25_43;
	wire [WIDTH-1:0] wire_d25_44;
	wire [WIDTH-1:0] wire_d25_45;
	wire [WIDTH-1:0] wire_d25_46;
	wire [WIDTH-1:0] wire_d25_47;
	wire [WIDTH-1:0] wire_d25_48;
	wire [WIDTH-1:0] wire_d26_0;
	wire [WIDTH-1:0] wire_d26_1;
	wire [WIDTH-1:0] wire_d26_2;
	wire [WIDTH-1:0] wire_d26_3;
	wire [WIDTH-1:0] wire_d26_4;
	wire [WIDTH-1:0] wire_d26_5;
	wire [WIDTH-1:0] wire_d26_6;
	wire [WIDTH-1:0] wire_d26_7;
	wire [WIDTH-1:0] wire_d26_8;
	wire [WIDTH-1:0] wire_d26_9;
	wire [WIDTH-1:0] wire_d26_10;
	wire [WIDTH-1:0] wire_d26_11;
	wire [WIDTH-1:0] wire_d26_12;
	wire [WIDTH-1:0] wire_d26_13;
	wire [WIDTH-1:0] wire_d26_14;
	wire [WIDTH-1:0] wire_d26_15;
	wire [WIDTH-1:0] wire_d26_16;
	wire [WIDTH-1:0] wire_d26_17;
	wire [WIDTH-1:0] wire_d26_18;
	wire [WIDTH-1:0] wire_d26_19;
	wire [WIDTH-1:0] wire_d26_20;
	wire [WIDTH-1:0] wire_d26_21;
	wire [WIDTH-1:0] wire_d26_22;
	wire [WIDTH-1:0] wire_d26_23;
	wire [WIDTH-1:0] wire_d26_24;
	wire [WIDTH-1:0] wire_d26_25;
	wire [WIDTH-1:0] wire_d26_26;
	wire [WIDTH-1:0] wire_d26_27;
	wire [WIDTH-1:0] wire_d26_28;
	wire [WIDTH-1:0] wire_d26_29;
	wire [WIDTH-1:0] wire_d26_30;
	wire [WIDTH-1:0] wire_d26_31;
	wire [WIDTH-1:0] wire_d26_32;
	wire [WIDTH-1:0] wire_d26_33;
	wire [WIDTH-1:0] wire_d26_34;
	wire [WIDTH-1:0] wire_d26_35;
	wire [WIDTH-1:0] wire_d26_36;
	wire [WIDTH-1:0] wire_d26_37;
	wire [WIDTH-1:0] wire_d26_38;
	wire [WIDTH-1:0] wire_d26_39;
	wire [WIDTH-1:0] wire_d26_40;
	wire [WIDTH-1:0] wire_d26_41;
	wire [WIDTH-1:0] wire_d26_42;
	wire [WIDTH-1:0] wire_d26_43;
	wire [WIDTH-1:0] wire_d26_44;
	wire [WIDTH-1:0] wire_d26_45;
	wire [WIDTH-1:0] wire_d26_46;
	wire [WIDTH-1:0] wire_d26_47;
	wire [WIDTH-1:0] wire_d26_48;
	wire [WIDTH-1:0] wire_d27_0;
	wire [WIDTH-1:0] wire_d27_1;
	wire [WIDTH-1:0] wire_d27_2;
	wire [WIDTH-1:0] wire_d27_3;
	wire [WIDTH-1:0] wire_d27_4;
	wire [WIDTH-1:0] wire_d27_5;
	wire [WIDTH-1:0] wire_d27_6;
	wire [WIDTH-1:0] wire_d27_7;
	wire [WIDTH-1:0] wire_d27_8;
	wire [WIDTH-1:0] wire_d27_9;
	wire [WIDTH-1:0] wire_d27_10;
	wire [WIDTH-1:0] wire_d27_11;
	wire [WIDTH-1:0] wire_d27_12;
	wire [WIDTH-1:0] wire_d27_13;
	wire [WIDTH-1:0] wire_d27_14;
	wire [WIDTH-1:0] wire_d27_15;
	wire [WIDTH-1:0] wire_d27_16;
	wire [WIDTH-1:0] wire_d27_17;
	wire [WIDTH-1:0] wire_d27_18;
	wire [WIDTH-1:0] wire_d27_19;
	wire [WIDTH-1:0] wire_d27_20;
	wire [WIDTH-1:0] wire_d27_21;
	wire [WIDTH-1:0] wire_d27_22;
	wire [WIDTH-1:0] wire_d27_23;
	wire [WIDTH-1:0] wire_d27_24;
	wire [WIDTH-1:0] wire_d27_25;
	wire [WIDTH-1:0] wire_d27_26;
	wire [WIDTH-1:0] wire_d27_27;
	wire [WIDTH-1:0] wire_d27_28;
	wire [WIDTH-1:0] wire_d27_29;
	wire [WIDTH-1:0] wire_d27_30;
	wire [WIDTH-1:0] wire_d27_31;
	wire [WIDTH-1:0] wire_d27_32;
	wire [WIDTH-1:0] wire_d27_33;
	wire [WIDTH-1:0] wire_d27_34;
	wire [WIDTH-1:0] wire_d27_35;
	wire [WIDTH-1:0] wire_d27_36;
	wire [WIDTH-1:0] wire_d27_37;
	wire [WIDTH-1:0] wire_d27_38;
	wire [WIDTH-1:0] wire_d27_39;
	wire [WIDTH-1:0] wire_d27_40;
	wire [WIDTH-1:0] wire_d27_41;
	wire [WIDTH-1:0] wire_d27_42;
	wire [WIDTH-1:0] wire_d27_43;
	wire [WIDTH-1:0] wire_d27_44;
	wire [WIDTH-1:0] wire_d27_45;
	wire [WIDTH-1:0] wire_d27_46;
	wire [WIDTH-1:0] wire_d27_47;
	wire [WIDTH-1:0] wire_d27_48;
	wire [WIDTH-1:0] wire_d28_0;
	wire [WIDTH-1:0] wire_d28_1;
	wire [WIDTH-1:0] wire_d28_2;
	wire [WIDTH-1:0] wire_d28_3;
	wire [WIDTH-1:0] wire_d28_4;
	wire [WIDTH-1:0] wire_d28_5;
	wire [WIDTH-1:0] wire_d28_6;
	wire [WIDTH-1:0] wire_d28_7;
	wire [WIDTH-1:0] wire_d28_8;
	wire [WIDTH-1:0] wire_d28_9;
	wire [WIDTH-1:0] wire_d28_10;
	wire [WIDTH-1:0] wire_d28_11;
	wire [WIDTH-1:0] wire_d28_12;
	wire [WIDTH-1:0] wire_d28_13;
	wire [WIDTH-1:0] wire_d28_14;
	wire [WIDTH-1:0] wire_d28_15;
	wire [WIDTH-1:0] wire_d28_16;
	wire [WIDTH-1:0] wire_d28_17;
	wire [WIDTH-1:0] wire_d28_18;
	wire [WIDTH-1:0] wire_d28_19;
	wire [WIDTH-1:0] wire_d28_20;
	wire [WIDTH-1:0] wire_d28_21;
	wire [WIDTH-1:0] wire_d28_22;
	wire [WIDTH-1:0] wire_d28_23;
	wire [WIDTH-1:0] wire_d28_24;
	wire [WIDTH-1:0] wire_d28_25;
	wire [WIDTH-1:0] wire_d28_26;
	wire [WIDTH-1:0] wire_d28_27;
	wire [WIDTH-1:0] wire_d28_28;
	wire [WIDTH-1:0] wire_d28_29;
	wire [WIDTH-1:0] wire_d28_30;
	wire [WIDTH-1:0] wire_d28_31;
	wire [WIDTH-1:0] wire_d28_32;
	wire [WIDTH-1:0] wire_d28_33;
	wire [WIDTH-1:0] wire_d28_34;
	wire [WIDTH-1:0] wire_d28_35;
	wire [WIDTH-1:0] wire_d28_36;
	wire [WIDTH-1:0] wire_d28_37;
	wire [WIDTH-1:0] wire_d28_38;
	wire [WIDTH-1:0] wire_d28_39;
	wire [WIDTH-1:0] wire_d28_40;
	wire [WIDTH-1:0] wire_d28_41;
	wire [WIDTH-1:0] wire_d28_42;
	wire [WIDTH-1:0] wire_d28_43;
	wire [WIDTH-1:0] wire_d28_44;
	wire [WIDTH-1:0] wire_d28_45;
	wire [WIDTH-1:0] wire_d28_46;
	wire [WIDTH-1:0] wire_d28_47;
	wire [WIDTH-1:0] wire_d28_48;
	wire [WIDTH-1:0] wire_d29_0;
	wire [WIDTH-1:0] wire_d29_1;
	wire [WIDTH-1:0] wire_d29_2;
	wire [WIDTH-1:0] wire_d29_3;
	wire [WIDTH-1:0] wire_d29_4;
	wire [WIDTH-1:0] wire_d29_5;
	wire [WIDTH-1:0] wire_d29_6;
	wire [WIDTH-1:0] wire_d29_7;
	wire [WIDTH-1:0] wire_d29_8;
	wire [WIDTH-1:0] wire_d29_9;
	wire [WIDTH-1:0] wire_d29_10;
	wire [WIDTH-1:0] wire_d29_11;
	wire [WIDTH-1:0] wire_d29_12;
	wire [WIDTH-1:0] wire_d29_13;
	wire [WIDTH-1:0] wire_d29_14;
	wire [WIDTH-1:0] wire_d29_15;
	wire [WIDTH-1:0] wire_d29_16;
	wire [WIDTH-1:0] wire_d29_17;
	wire [WIDTH-1:0] wire_d29_18;
	wire [WIDTH-1:0] wire_d29_19;
	wire [WIDTH-1:0] wire_d29_20;
	wire [WIDTH-1:0] wire_d29_21;
	wire [WIDTH-1:0] wire_d29_22;
	wire [WIDTH-1:0] wire_d29_23;
	wire [WIDTH-1:0] wire_d29_24;
	wire [WIDTH-1:0] wire_d29_25;
	wire [WIDTH-1:0] wire_d29_26;
	wire [WIDTH-1:0] wire_d29_27;
	wire [WIDTH-1:0] wire_d29_28;
	wire [WIDTH-1:0] wire_d29_29;
	wire [WIDTH-1:0] wire_d29_30;
	wire [WIDTH-1:0] wire_d29_31;
	wire [WIDTH-1:0] wire_d29_32;
	wire [WIDTH-1:0] wire_d29_33;
	wire [WIDTH-1:0] wire_d29_34;
	wire [WIDTH-1:0] wire_d29_35;
	wire [WIDTH-1:0] wire_d29_36;
	wire [WIDTH-1:0] wire_d29_37;
	wire [WIDTH-1:0] wire_d29_38;
	wire [WIDTH-1:0] wire_d29_39;
	wire [WIDTH-1:0] wire_d29_40;
	wire [WIDTH-1:0] wire_d29_41;
	wire [WIDTH-1:0] wire_d29_42;
	wire [WIDTH-1:0] wire_d29_43;
	wire [WIDTH-1:0] wire_d29_44;
	wire [WIDTH-1:0] wire_d29_45;
	wire [WIDTH-1:0] wire_d29_46;
	wire [WIDTH-1:0] wire_d29_47;
	wire [WIDTH-1:0] wire_d29_48;
	wire [WIDTH-1:0] wire_d30_0;
	wire [WIDTH-1:0] wire_d30_1;
	wire [WIDTH-1:0] wire_d30_2;
	wire [WIDTH-1:0] wire_d30_3;
	wire [WIDTH-1:0] wire_d30_4;
	wire [WIDTH-1:0] wire_d30_5;
	wire [WIDTH-1:0] wire_d30_6;
	wire [WIDTH-1:0] wire_d30_7;
	wire [WIDTH-1:0] wire_d30_8;
	wire [WIDTH-1:0] wire_d30_9;
	wire [WIDTH-1:0] wire_d30_10;
	wire [WIDTH-1:0] wire_d30_11;
	wire [WIDTH-1:0] wire_d30_12;
	wire [WIDTH-1:0] wire_d30_13;
	wire [WIDTH-1:0] wire_d30_14;
	wire [WIDTH-1:0] wire_d30_15;
	wire [WIDTH-1:0] wire_d30_16;
	wire [WIDTH-1:0] wire_d30_17;
	wire [WIDTH-1:0] wire_d30_18;
	wire [WIDTH-1:0] wire_d30_19;
	wire [WIDTH-1:0] wire_d30_20;
	wire [WIDTH-1:0] wire_d30_21;
	wire [WIDTH-1:0] wire_d30_22;
	wire [WIDTH-1:0] wire_d30_23;
	wire [WIDTH-1:0] wire_d30_24;
	wire [WIDTH-1:0] wire_d30_25;
	wire [WIDTH-1:0] wire_d30_26;
	wire [WIDTH-1:0] wire_d30_27;
	wire [WIDTH-1:0] wire_d30_28;
	wire [WIDTH-1:0] wire_d30_29;
	wire [WIDTH-1:0] wire_d30_30;
	wire [WIDTH-1:0] wire_d30_31;
	wire [WIDTH-1:0] wire_d30_32;
	wire [WIDTH-1:0] wire_d30_33;
	wire [WIDTH-1:0] wire_d30_34;
	wire [WIDTH-1:0] wire_d30_35;
	wire [WIDTH-1:0] wire_d30_36;
	wire [WIDTH-1:0] wire_d30_37;
	wire [WIDTH-1:0] wire_d30_38;
	wire [WIDTH-1:0] wire_d30_39;
	wire [WIDTH-1:0] wire_d30_40;
	wire [WIDTH-1:0] wire_d30_41;
	wire [WIDTH-1:0] wire_d30_42;
	wire [WIDTH-1:0] wire_d30_43;
	wire [WIDTH-1:0] wire_d30_44;
	wire [WIDTH-1:0] wire_d30_45;
	wire [WIDTH-1:0] wire_d30_46;
	wire [WIDTH-1:0] wire_d30_47;
	wire [WIDTH-1:0] wire_d30_48;
	wire [WIDTH-1:0] wire_d31_0;
	wire [WIDTH-1:0] wire_d31_1;
	wire [WIDTH-1:0] wire_d31_2;
	wire [WIDTH-1:0] wire_d31_3;
	wire [WIDTH-1:0] wire_d31_4;
	wire [WIDTH-1:0] wire_d31_5;
	wire [WIDTH-1:0] wire_d31_6;
	wire [WIDTH-1:0] wire_d31_7;
	wire [WIDTH-1:0] wire_d31_8;
	wire [WIDTH-1:0] wire_d31_9;
	wire [WIDTH-1:0] wire_d31_10;
	wire [WIDTH-1:0] wire_d31_11;
	wire [WIDTH-1:0] wire_d31_12;
	wire [WIDTH-1:0] wire_d31_13;
	wire [WIDTH-1:0] wire_d31_14;
	wire [WIDTH-1:0] wire_d31_15;
	wire [WIDTH-1:0] wire_d31_16;
	wire [WIDTH-1:0] wire_d31_17;
	wire [WIDTH-1:0] wire_d31_18;
	wire [WIDTH-1:0] wire_d31_19;
	wire [WIDTH-1:0] wire_d31_20;
	wire [WIDTH-1:0] wire_d31_21;
	wire [WIDTH-1:0] wire_d31_22;
	wire [WIDTH-1:0] wire_d31_23;
	wire [WIDTH-1:0] wire_d31_24;
	wire [WIDTH-1:0] wire_d31_25;
	wire [WIDTH-1:0] wire_d31_26;
	wire [WIDTH-1:0] wire_d31_27;
	wire [WIDTH-1:0] wire_d31_28;
	wire [WIDTH-1:0] wire_d31_29;
	wire [WIDTH-1:0] wire_d31_30;
	wire [WIDTH-1:0] wire_d31_31;
	wire [WIDTH-1:0] wire_d31_32;
	wire [WIDTH-1:0] wire_d31_33;
	wire [WIDTH-1:0] wire_d31_34;
	wire [WIDTH-1:0] wire_d31_35;
	wire [WIDTH-1:0] wire_d31_36;
	wire [WIDTH-1:0] wire_d31_37;
	wire [WIDTH-1:0] wire_d31_38;
	wire [WIDTH-1:0] wire_d31_39;
	wire [WIDTH-1:0] wire_d31_40;
	wire [WIDTH-1:0] wire_d31_41;
	wire [WIDTH-1:0] wire_d31_42;
	wire [WIDTH-1:0] wire_d31_43;
	wire [WIDTH-1:0] wire_d31_44;
	wire [WIDTH-1:0] wire_d31_45;
	wire [WIDTH-1:0] wire_d31_46;
	wire [WIDTH-1:0] wire_d31_47;
	wire [WIDTH-1:0] wire_d31_48;
	wire [WIDTH-1:0] wire_d32_0;
	wire [WIDTH-1:0] wire_d32_1;
	wire [WIDTH-1:0] wire_d32_2;
	wire [WIDTH-1:0] wire_d32_3;
	wire [WIDTH-1:0] wire_d32_4;
	wire [WIDTH-1:0] wire_d32_5;
	wire [WIDTH-1:0] wire_d32_6;
	wire [WIDTH-1:0] wire_d32_7;
	wire [WIDTH-1:0] wire_d32_8;
	wire [WIDTH-1:0] wire_d32_9;
	wire [WIDTH-1:0] wire_d32_10;
	wire [WIDTH-1:0] wire_d32_11;
	wire [WIDTH-1:0] wire_d32_12;
	wire [WIDTH-1:0] wire_d32_13;
	wire [WIDTH-1:0] wire_d32_14;
	wire [WIDTH-1:0] wire_d32_15;
	wire [WIDTH-1:0] wire_d32_16;
	wire [WIDTH-1:0] wire_d32_17;
	wire [WIDTH-1:0] wire_d32_18;
	wire [WIDTH-1:0] wire_d32_19;
	wire [WIDTH-1:0] wire_d32_20;
	wire [WIDTH-1:0] wire_d32_21;
	wire [WIDTH-1:0] wire_d32_22;
	wire [WIDTH-1:0] wire_d32_23;
	wire [WIDTH-1:0] wire_d32_24;
	wire [WIDTH-1:0] wire_d32_25;
	wire [WIDTH-1:0] wire_d32_26;
	wire [WIDTH-1:0] wire_d32_27;
	wire [WIDTH-1:0] wire_d32_28;
	wire [WIDTH-1:0] wire_d32_29;
	wire [WIDTH-1:0] wire_d32_30;
	wire [WIDTH-1:0] wire_d32_31;
	wire [WIDTH-1:0] wire_d32_32;
	wire [WIDTH-1:0] wire_d32_33;
	wire [WIDTH-1:0] wire_d32_34;
	wire [WIDTH-1:0] wire_d32_35;
	wire [WIDTH-1:0] wire_d32_36;
	wire [WIDTH-1:0] wire_d32_37;
	wire [WIDTH-1:0] wire_d32_38;
	wire [WIDTH-1:0] wire_d32_39;
	wire [WIDTH-1:0] wire_d32_40;
	wire [WIDTH-1:0] wire_d32_41;
	wire [WIDTH-1:0] wire_d32_42;
	wire [WIDTH-1:0] wire_d32_43;
	wire [WIDTH-1:0] wire_d32_44;
	wire [WIDTH-1:0] wire_d32_45;
	wire [WIDTH-1:0] wire_d32_46;
	wire [WIDTH-1:0] wire_d32_47;
	wire [WIDTH-1:0] wire_d32_48;
	wire [WIDTH-1:0] wire_d33_0;
	wire [WIDTH-1:0] wire_d33_1;
	wire [WIDTH-1:0] wire_d33_2;
	wire [WIDTH-1:0] wire_d33_3;
	wire [WIDTH-1:0] wire_d33_4;
	wire [WIDTH-1:0] wire_d33_5;
	wire [WIDTH-1:0] wire_d33_6;
	wire [WIDTH-1:0] wire_d33_7;
	wire [WIDTH-1:0] wire_d33_8;
	wire [WIDTH-1:0] wire_d33_9;
	wire [WIDTH-1:0] wire_d33_10;
	wire [WIDTH-1:0] wire_d33_11;
	wire [WIDTH-1:0] wire_d33_12;
	wire [WIDTH-1:0] wire_d33_13;
	wire [WIDTH-1:0] wire_d33_14;
	wire [WIDTH-1:0] wire_d33_15;
	wire [WIDTH-1:0] wire_d33_16;
	wire [WIDTH-1:0] wire_d33_17;
	wire [WIDTH-1:0] wire_d33_18;
	wire [WIDTH-1:0] wire_d33_19;
	wire [WIDTH-1:0] wire_d33_20;
	wire [WIDTH-1:0] wire_d33_21;
	wire [WIDTH-1:0] wire_d33_22;
	wire [WIDTH-1:0] wire_d33_23;
	wire [WIDTH-1:0] wire_d33_24;
	wire [WIDTH-1:0] wire_d33_25;
	wire [WIDTH-1:0] wire_d33_26;
	wire [WIDTH-1:0] wire_d33_27;
	wire [WIDTH-1:0] wire_d33_28;
	wire [WIDTH-1:0] wire_d33_29;
	wire [WIDTH-1:0] wire_d33_30;
	wire [WIDTH-1:0] wire_d33_31;
	wire [WIDTH-1:0] wire_d33_32;
	wire [WIDTH-1:0] wire_d33_33;
	wire [WIDTH-1:0] wire_d33_34;
	wire [WIDTH-1:0] wire_d33_35;
	wire [WIDTH-1:0] wire_d33_36;
	wire [WIDTH-1:0] wire_d33_37;
	wire [WIDTH-1:0] wire_d33_38;
	wire [WIDTH-1:0] wire_d33_39;
	wire [WIDTH-1:0] wire_d33_40;
	wire [WIDTH-1:0] wire_d33_41;
	wire [WIDTH-1:0] wire_d33_42;
	wire [WIDTH-1:0] wire_d33_43;
	wire [WIDTH-1:0] wire_d33_44;
	wire [WIDTH-1:0] wire_d33_45;
	wire [WIDTH-1:0] wire_d33_46;
	wire [WIDTH-1:0] wire_d33_47;
	wire [WIDTH-1:0] wire_d33_48;
	wire [WIDTH-1:0] wire_d34_0;
	wire [WIDTH-1:0] wire_d34_1;
	wire [WIDTH-1:0] wire_d34_2;
	wire [WIDTH-1:0] wire_d34_3;
	wire [WIDTH-1:0] wire_d34_4;
	wire [WIDTH-1:0] wire_d34_5;
	wire [WIDTH-1:0] wire_d34_6;
	wire [WIDTH-1:0] wire_d34_7;
	wire [WIDTH-1:0] wire_d34_8;
	wire [WIDTH-1:0] wire_d34_9;
	wire [WIDTH-1:0] wire_d34_10;
	wire [WIDTH-1:0] wire_d34_11;
	wire [WIDTH-1:0] wire_d34_12;
	wire [WIDTH-1:0] wire_d34_13;
	wire [WIDTH-1:0] wire_d34_14;
	wire [WIDTH-1:0] wire_d34_15;
	wire [WIDTH-1:0] wire_d34_16;
	wire [WIDTH-1:0] wire_d34_17;
	wire [WIDTH-1:0] wire_d34_18;
	wire [WIDTH-1:0] wire_d34_19;
	wire [WIDTH-1:0] wire_d34_20;
	wire [WIDTH-1:0] wire_d34_21;
	wire [WIDTH-1:0] wire_d34_22;
	wire [WIDTH-1:0] wire_d34_23;
	wire [WIDTH-1:0] wire_d34_24;
	wire [WIDTH-1:0] wire_d34_25;
	wire [WIDTH-1:0] wire_d34_26;
	wire [WIDTH-1:0] wire_d34_27;
	wire [WIDTH-1:0] wire_d34_28;
	wire [WIDTH-1:0] wire_d34_29;
	wire [WIDTH-1:0] wire_d34_30;
	wire [WIDTH-1:0] wire_d34_31;
	wire [WIDTH-1:0] wire_d34_32;
	wire [WIDTH-1:0] wire_d34_33;
	wire [WIDTH-1:0] wire_d34_34;
	wire [WIDTH-1:0] wire_d34_35;
	wire [WIDTH-1:0] wire_d34_36;
	wire [WIDTH-1:0] wire_d34_37;
	wire [WIDTH-1:0] wire_d34_38;
	wire [WIDTH-1:0] wire_d34_39;
	wire [WIDTH-1:0] wire_d34_40;
	wire [WIDTH-1:0] wire_d34_41;
	wire [WIDTH-1:0] wire_d34_42;
	wire [WIDTH-1:0] wire_d34_43;
	wire [WIDTH-1:0] wire_d34_44;
	wire [WIDTH-1:0] wire_d34_45;
	wire [WIDTH-1:0] wire_d34_46;
	wire [WIDTH-1:0] wire_d34_47;
	wire [WIDTH-1:0] wire_d34_48;
	wire [WIDTH-1:0] wire_d35_0;
	wire [WIDTH-1:0] wire_d35_1;
	wire [WIDTH-1:0] wire_d35_2;
	wire [WIDTH-1:0] wire_d35_3;
	wire [WIDTH-1:0] wire_d35_4;
	wire [WIDTH-1:0] wire_d35_5;
	wire [WIDTH-1:0] wire_d35_6;
	wire [WIDTH-1:0] wire_d35_7;
	wire [WIDTH-1:0] wire_d35_8;
	wire [WIDTH-1:0] wire_d35_9;
	wire [WIDTH-1:0] wire_d35_10;
	wire [WIDTH-1:0] wire_d35_11;
	wire [WIDTH-1:0] wire_d35_12;
	wire [WIDTH-1:0] wire_d35_13;
	wire [WIDTH-1:0] wire_d35_14;
	wire [WIDTH-1:0] wire_d35_15;
	wire [WIDTH-1:0] wire_d35_16;
	wire [WIDTH-1:0] wire_d35_17;
	wire [WIDTH-1:0] wire_d35_18;
	wire [WIDTH-1:0] wire_d35_19;
	wire [WIDTH-1:0] wire_d35_20;
	wire [WIDTH-1:0] wire_d35_21;
	wire [WIDTH-1:0] wire_d35_22;
	wire [WIDTH-1:0] wire_d35_23;
	wire [WIDTH-1:0] wire_d35_24;
	wire [WIDTH-1:0] wire_d35_25;
	wire [WIDTH-1:0] wire_d35_26;
	wire [WIDTH-1:0] wire_d35_27;
	wire [WIDTH-1:0] wire_d35_28;
	wire [WIDTH-1:0] wire_d35_29;
	wire [WIDTH-1:0] wire_d35_30;
	wire [WIDTH-1:0] wire_d35_31;
	wire [WIDTH-1:0] wire_d35_32;
	wire [WIDTH-1:0] wire_d35_33;
	wire [WIDTH-1:0] wire_d35_34;
	wire [WIDTH-1:0] wire_d35_35;
	wire [WIDTH-1:0] wire_d35_36;
	wire [WIDTH-1:0] wire_d35_37;
	wire [WIDTH-1:0] wire_d35_38;
	wire [WIDTH-1:0] wire_d35_39;
	wire [WIDTH-1:0] wire_d35_40;
	wire [WIDTH-1:0] wire_d35_41;
	wire [WIDTH-1:0] wire_d35_42;
	wire [WIDTH-1:0] wire_d35_43;
	wire [WIDTH-1:0] wire_d35_44;
	wire [WIDTH-1:0] wire_d35_45;
	wire [WIDTH-1:0] wire_d35_46;
	wire [WIDTH-1:0] wire_d35_47;
	wire [WIDTH-1:0] wire_d35_48;
	wire [WIDTH-1:0] wire_d36_0;
	wire [WIDTH-1:0] wire_d36_1;
	wire [WIDTH-1:0] wire_d36_2;
	wire [WIDTH-1:0] wire_d36_3;
	wire [WIDTH-1:0] wire_d36_4;
	wire [WIDTH-1:0] wire_d36_5;
	wire [WIDTH-1:0] wire_d36_6;
	wire [WIDTH-1:0] wire_d36_7;
	wire [WIDTH-1:0] wire_d36_8;
	wire [WIDTH-1:0] wire_d36_9;
	wire [WIDTH-1:0] wire_d36_10;
	wire [WIDTH-1:0] wire_d36_11;
	wire [WIDTH-1:0] wire_d36_12;
	wire [WIDTH-1:0] wire_d36_13;
	wire [WIDTH-1:0] wire_d36_14;
	wire [WIDTH-1:0] wire_d36_15;
	wire [WIDTH-1:0] wire_d36_16;
	wire [WIDTH-1:0] wire_d36_17;
	wire [WIDTH-1:0] wire_d36_18;
	wire [WIDTH-1:0] wire_d36_19;
	wire [WIDTH-1:0] wire_d36_20;
	wire [WIDTH-1:0] wire_d36_21;
	wire [WIDTH-1:0] wire_d36_22;
	wire [WIDTH-1:0] wire_d36_23;
	wire [WIDTH-1:0] wire_d36_24;
	wire [WIDTH-1:0] wire_d36_25;
	wire [WIDTH-1:0] wire_d36_26;
	wire [WIDTH-1:0] wire_d36_27;
	wire [WIDTH-1:0] wire_d36_28;
	wire [WIDTH-1:0] wire_d36_29;
	wire [WIDTH-1:0] wire_d36_30;
	wire [WIDTH-1:0] wire_d36_31;
	wire [WIDTH-1:0] wire_d36_32;
	wire [WIDTH-1:0] wire_d36_33;
	wire [WIDTH-1:0] wire_d36_34;
	wire [WIDTH-1:0] wire_d36_35;
	wire [WIDTH-1:0] wire_d36_36;
	wire [WIDTH-1:0] wire_d36_37;
	wire [WIDTH-1:0] wire_d36_38;
	wire [WIDTH-1:0] wire_d36_39;
	wire [WIDTH-1:0] wire_d36_40;
	wire [WIDTH-1:0] wire_d36_41;
	wire [WIDTH-1:0] wire_d36_42;
	wire [WIDTH-1:0] wire_d36_43;
	wire [WIDTH-1:0] wire_d36_44;
	wire [WIDTH-1:0] wire_d36_45;
	wire [WIDTH-1:0] wire_d36_46;
	wire [WIDTH-1:0] wire_d36_47;
	wire [WIDTH-1:0] wire_d36_48;
	wire [WIDTH-1:0] wire_d37_0;
	wire [WIDTH-1:0] wire_d37_1;
	wire [WIDTH-1:0] wire_d37_2;
	wire [WIDTH-1:0] wire_d37_3;
	wire [WIDTH-1:0] wire_d37_4;
	wire [WIDTH-1:0] wire_d37_5;
	wire [WIDTH-1:0] wire_d37_6;
	wire [WIDTH-1:0] wire_d37_7;
	wire [WIDTH-1:0] wire_d37_8;
	wire [WIDTH-1:0] wire_d37_9;
	wire [WIDTH-1:0] wire_d37_10;
	wire [WIDTH-1:0] wire_d37_11;
	wire [WIDTH-1:0] wire_d37_12;
	wire [WIDTH-1:0] wire_d37_13;
	wire [WIDTH-1:0] wire_d37_14;
	wire [WIDTH-1:0] wire_d37_15;
	wire [WIDTH-1:0] wire_d37_16;
	wire [WIDTH-1:0] wire_d37_17;
	wire [WIDTH-1:0] wire_d37_18;
	wire [WIDTH-1:0] wire_d37_19;
	wire [WIDTH-1:0] wire_d37_20;
	wire [WIDTH-1:0] wire_d37_21;
	wire [WIDTH-1:0] wire_d37_22;
	wire [WIDTH-1:0] wire_d37_23;
	wire [WIDTH-1:0] wire_d37_24;
	wire [WIDTH-1:0] wire_d37_25;
	wire [WIDTH-1:0] wire_d37_26;
	wire [WIDTH-1:0] wire_d37_27;
	wire [WIDTH-1:0] wire_d37_28;
	wire [WIDTH-1:0] wire_d37_29;
	wire [WIDTH-1:0] wire_d37_30;
	wire [WIDTH-1:0] wire_d37_31;
	wire [WIDTH-1:0] wire_d37_32;
	wire [WIDTH-1:0] wire_d37_33;
	wire [WIDTH-1:0] wire_d37_34;
	wire [WIDTH-1:0] wire_d37_35;
	wire [WIDTH-1:0] wire_d37_36;
	wire [WIDTH-1:0] wire_d37_37;
	wire [WIDTH-1:0] wire_d37_38;
	wire [WIDTH-1:0] wire_d37_39;
	wire [WIDTH-1:0] wire_d37_40;
	wire [WIDTH-1:0] wire_d37_41;
	wire [WIDTH-1:0] wire_d37_42;
	wire [WIDTH-1:0] wire_d37_43;
	wire [WIDTH-1:0] wire_d37_44;
	wire [WIDTH-1:0] wire_d37_45;
	wire [WIDTH-1:0] wire_d37_46;
	wire [WIDTH-1:0] wire_d37_47;
	wire [WIDTH-1:0] wire_d37_48;
	wire [WIDTH-1:0] wire_d38_0;
	wire [WIDTH-1:0] wire_d38_1;
	wire [WIDTH-1:0] wire_d38_2;
	wire [WIDTH-1:0] wire_d38_3;
	wire [WIDTH-1:0] wire_d38_4;
	wire [WIDTH-1:0] wire_d38_5;
	wire [WIDTH-1:0] wire_d38_6;
	wire [WIDTH-1:0] wire_d38_7;
	wire [WIDTH-1:0] wire_d38_8;
	wire [WIDTH-1:0] wire_d38_9;
	wire [WIDTH-1:0] wire_d38_10;
	wire [WIDTH-1:0] wire_d38_11;
	wire [WIDTH-1:0] wire_d38_12;
	wire [WIDTH-1:0] wire_d38_13;
	wire [WIDTH-1:0] wire_d38_14;
	wire [WIDTH-1:0] wire_d38_15;
	wire [WIDTH-1:0] wire_d38_16;
	wire [WIDTH-1:0] wire_d38_17;
	wire [WIDTH-1:0] wire_d38_18;
	wire [WIDTH-1:0] wire_d38_19;
	wire [WIDTH-1:0] wire_d38_20;
	wire [WIDTH-1:0] wire_d38_21;
	wire [WIDTH-1:0] wire_d38_22;
	wire [WIDTH-1:0] wire_d38_23;
	wire [WIDTH-1:0] wire_d38_24;
	wire [WIDTH-1:0] wire_d38_25;
	wire [WIDTH-1:0] wire_d38_26;
	wire [WIDTH-1:0] wire_d38_27;
	wire [WIDTH-1:0] wire_d38_28;
	wire [WIDTH-1:0] wire_d38_29;
	wire [WIDTH-1:0] wire_d38_30;
	wire [WIDTH-1:0] wire_d38_31;
	wire [WIDTH-1:0] wire_d38_32;
	wire [WIDTH-1:0] wire_d38_33;
	wire [WIDTH-1:0] wire_d38_34;
	wire [WIDTH-1:0] wire_d38_35;
	wire [WIDTH-1:0] wire_d38_36;
	wire [WIDTH-1:0] wire_d38_37;
	wire [WIDTH-1:0] wire_d38_38;
	wire [WIDTH-1:0] wire_d38_39;
	wire [WIDTH-1:0] wire_d38_40;
	wire [WIDTH-1:0] wire_d38_41;
	wire [WIDTH-1:0] wire_d38_42;
	wire [WIDTH-1:0] wire_d38_43;
	wire [WIDTH-1:0] wire_d38_44;
	wire [WIDTH-1:0] wire_d38_45;
	wire [WIDTH-1:0] wire_d38_46;
	wire [WIDTH-1:0] wire_d38_47;
	wire [WIDTH-1:0] wire_d38_48;
	wire [WIDTH-1:0] wire_d39_0;
	wire [WIDTH-1:0] wire_d39_1;
	wire [WIDTH-1:0] wire_d39_2;
	wire [WIDTH-1:0] wire_d39_3;
	wire [WIDTH-1:0] wire_d39_4;
	wire [WIDTH-1:0] wire_d39_5;
	wire [WIDTH-1:0] wire_d39_6;
	wire [WIDTH-1:0] wire_d39_7;
	wire [WIDTH-1:0] wire_d39_8;
	wire [WIDTH-1:0] wire_d39_9;
	wire [WIDTH-1:0] wire_d39_10;
	wire [WIDTH-1:0] wire_d39_11;
	wire [WIDTH-1:0] wire_d39_12;
	wire [WIDTH-1:0] wire_d39_13;
	wire [WIDTH-1:0] wire_d39_14;
	wire [WIDTH-1:0] wire_d39_15;
	wire [WIDTH-1:0] wire_d39_16;
	wire [WIDTH-1:0] wire_d39_17;
	wire [WIDTH-1:0] wire_d39_18;
	wire [WIDTH-1:0] wire_d39_19;
	wire [WIDTH-1:0] wire_d39_20;
	wire [WIDTH-1:0] wire_d39_21;
	wire [WIDTH-1:0] wire_d39_22;
	wire [WIDTH-1:0] wire_d39_23;
	wire [WIDTH-1:0] wire_d39_24;
	wire [WIDTH-1:0] wire_d39_25;
	wire [WIDTH-1:0] wire_d39_26;
	wire [WIDTH-1:0] wire_d39_27;
	wire [WIDTH-1:0] wire_d39_28;
	wire [WIDTH-1:0] wire_d39_29;
	wire [WIDTH-1:0] wire_d39_30;
	wire [WIDTH-1:0] wire_d39_31;
	wire [WIDTH-1:0] wire_d39_32;
	wire [WIDTH-1:0] wire_d39_33;
	wire [WIDTH-1:0] wire_d39_34;
	wire [WIDTH-1:0] wire_d39_35;
	wire [WIDTH-1:0] wire_d39_36;
	wire [WIDTH-1:0] wire_d39_37;
	wire [WIDTH-1:0] wire_d39_38;
	wire [WIDTH-1:0] wire_d39_39;
	wire [WIDTH-1:0] wire_d39_40;
	wire [WIDTH-1:0] wire_d39_41;
	wire [WIDTH-1:0] wire_d39_42;
	wire [WIDTH-1:0] wire_d39_43;
	wire [WIDTH-1:0] wire_d39_44;
	wire [WIDTH-1:0] wire_d39_45;
	wire [WIDTH-1:0] wire_d39_46;
	wire [WIDTH-1:0] wire_d39_47;
	wire [WIDTH-1:0] wire_d39_48;
	wire [WIDTH-1:0] wire_d40_0;
	wire [WIDTH-1:0] wire_d40_1;
	wire [WIDTH-1:0] wire_d40_2;
	wire [WIDTH-1:0] wire_d40_3;
	wire [WIDTH-1:0] wire_d40_4;
	wire [WIDTH-1:0] wire_d40_5;
	wire [WIDTH-1:0] wire_d40_6;
	wire [WIDTH-1:0] wire_d40_7;
	wire [WIDTH-1:0] wire_d40_8;
	wire [WIDTH-1:0] wire_d40_9;
	wire [WIDTH-1:0] wire_d40_10;
	wire [WIDTH-1:0] wire_d40_11;
	wire [WIDTH-1:0] wire_d40_12;
	wire [WIDTH-1:0] wire_d40_13;
	wire [WIDTH-1:0] wire_d40_14;
	wire [WIDTH-1:0] wire_d40_15;
	wire [WIDTH-1:0] wire_d40_16;
	wire [WIDTH-1:0] wire_d40_17;
	wire [WIDTH-1:0] wire_d40_18;
	wire [WIDTH-1:0] wire_d40_19;
	wire [WIDTH-1:0] wire_d40_20;
	wire [WIDTH-1:0] wire_d40_21;
	wire [WIDTH-1:0] wire_d40_22;
	wire [WIDTH-1:0] wire_d40_23;
	wire [WIDTH-1:0] wire_d40_24;
	wire [WIDTH-1:0] wire_d40_25;
	wire [WIDTH-1:0] wire_d40_26;
	wire [WIDTH-1:0] wire_d40_27;
	wire [WIDTH-1:0] wire_d40_28;
	wire [WIDTH-1:0] wire_d40_29;
	wire [WIDTH-1:0] wire_d40_30;
	wire [WIDTH-1:0] wire_d40_31;
	wire [WIDTH-1:0] wire_d40_32;
	wire [WIDTH-1:0] wire_d40_33;
	wire [WIDTH-1:0] wire_d40_34;
	wire [WIDTH-1:0] wire_d40_35;
	wire [WIDTH-1:0] wire_d40_36;
	wire [WIDTH-1:0] wire_d40_37;
	wire [WIDTH-1:0] wire_d40_38;
	wire [WIDTH-1:0] wire_d40_39;
	wire [WIDTH-1:0] wire_d40_40;
	wire [WIDTH-1:0] wire_d40_41;
	wire [WIDTH-1:0] wire_d40_42;
	wire [WIDTH-1:0] wire_d40_43;
	wire [WIDTH-1:0] wire_d40_44;
	wire [WIDTH-1:0] wire_d40_45;
	wire [WIDTH-1:0] wire_d40_46;
	wire [WIDTH-1:0] wire_d40_47;
	wire [WIDTH-1:0] wire_d40_48;
	wire [WIDTH-1:0] wire_d41_0;
	wire [WIDTH-1:0] wire_d41_1;
	wire [WIDTH-1:0] wire_d41_2;
	wire [WIDTH-1:0] wire_d41_3;
	wire [WIDTH-1:0] wire_d41_4;
	wire [WIDTH-1:0] wire_d41_5;
	wire [WIDTH-1:0] wire_d41_6;
	wire [WIDTH-1:0] wire_d41_7;
	wire [WIDTH-1:0] wire_d41_8;
	wire [WIDTH-1:0] wire_d41_9;
	wire [WIDTH-1:0] wire_d41_10;
	wire [WIDTH-1:0] wire_d41_11;
	wire [WIDTH-1:0] wire_d41_12;
	wire [WIDTH-1:0] wire_d41_13;
	wire [WIDTH-1:0] wire_d41_14;
	wire [WIDTH-1:0] wire_d41_15;
	wire [WIDTH-1:0] wire_d41_16;
	wire [WIDTH-1:0] wire_d41_17;
	wire [WIDTH-1:0] wire_d41_18;
	wire [WIDTH-1:0] wire_d41_19;
	wire [WIDTH-1:0] wire_d41_20;
	wire [WIDTH-1:0] wire_d41_21;
	wire [WIDTH-1:0] wire_d41_22;
	wire [WIDTH-1:0] wire_d41_23;
	wire [WIDTH-1:0] wire_d41_24;
	wire [WIDTH-1:0] wire_d41_25;
	wire [WIDTH-1:0] wire_d41_26;
	wire [WIDTH-1:0] wire_d41_27;
	wire [WIDTH-1:0] wire_d41_28;
	wire [WIDTH-1:0] wire_d41_29;
	wire [WIDTH-1:0] wire_d41_30;
	wire [WIDTH-1:0] wire_d41_31;
	wire [WIDTH-1:0] wire_d41_32;
	wire [WIDTH-1:0] wire_d41_33;
	wire [WIDTH-1:0] wire_d41_34;
	wire [WIDTH-1:0] wire_d41_35;
	wire [WIDTH-1:0] wire_d41_36;
	wire [WIDTH-1:0] wire_d41_37;
	wire [WIDTH-1:0] wire_d41_38;
	wire [WIDTH-1:0] wire_d41_39;
	wire [WIDTH-1:0] wire_d41_40;
	wire [WIDTH-1:0] wire_d41_41;
	wire [WIDTH-1:0] wire_d41_42;
	wire [WIDTH-1:0] wire_d41_43;
	wire [WIDTH-1:0] wire_d41_44;
	wire [WIDTH-1:0] wire_d41_45;
	wire [WIDTH-1:0] wire_d41_46;
	wire [WIDTH-1:0] wire_d41_47;
	wire [WIDTH-1:0] wire_d41_48;
	wire [WIDTH-1:0] wire_d42_0;
	wire [WIDTH-1:0] wire_d42_1;
	wire [WIDTH-1:0] wire_d42_2;
	wire [WIDTH-1:0] wire_d42_3;
	wire [WIDTH-1:0] wire_d42_4;
	wire [WIDTH-1:0] wire_d42_5;
	wire [WIDTH-1:0] wire_d42_6;
	wire [WIDTH-1:0] wire_d42_7;
	wire [WIDTH-1:0] wire_d42_8;
	wire [WIDTH-1:0] wire_d42_9;
	wire [WIDTH-1:0] wire_d42_10;
	wire [WIDTH-1:0] wire_d42_11;
	wire [WIDTH-1:0] wire_d42_12;
	wire [WIDTH-1:0] wire_d42_13;
	wire [WIDTH-1:0] wire_d42_14;
	wire [WIDTH-1:0] wire_d42_15;
	wire [WIDTH-1:0] wire_d42_16;
	wire [WIDTH-1:0] wire_d42_17;
	wire [WIDTH-1:0] wire_d42_18;
	wire [WIDTH-1:0] wire_d42_19;
	wire [WIDTH-1:0] wire_d42_20;
	wire [WIDTH-1:0] wire_d42_21;
	wire [WIDTH-1:0] wire_d42_22;
	wire [WIDTH-1:0] wire_d42_23;
	wire [WIDTH-1:0] wire_d42_24;
	wire [WIDTH-1:0] wire_d42_25;
	wire [WIDTH-1:0] wire_d42_26;
	wire [WIDTH-1:0] wire_d42_27;
	wire [WIDTH-1:0] wire_d42_28;
	wire [WIDTH-1:0] wire_d42_29;
	wire [WIDTH-1:0] wire_d42_30;
	wire [WIDTH-1:0] wire_d42_31;
	wire [WIDTH-1:0] wire_d42_32;
	wire [WIDTH-1:0] wire_d42_33;
	wire [WIDTH-1:0] wire_d42_34;
	wire [WIDTH-1:0] wire_d42_35;
	wire [WIDTH-1:0] wire_d42_36;
	wire [WIDTH-1:0] wire_d42_37;
	wire [WIDTH-1:0] wire_d42_38;
	wire [WIDTH-1:0] wire_d42_39;
	wire [WIDTH-1:0] wire_d42_40;
	wire [WIDTH-1:0] wire_d42_41;
	wire [WIDTH-1:0] wire_d42_42;
	wire [WIDTH-1:0] wire_d42_43;
	wire [WIDTH-1:0] wire_d42_44;
	wire [WIDTH-1:0] wire_d42_45;
	wire [WIDTH-1:0] wire_d42_46;
	wire [WIDTH-1:0] wire_d42_47;
	wire [WIDTH-1:0] wire_d42_48;
	wire [WIDTH-1:0] wire_d43_0;
	wire [WIDTH-1:0] wire_d43_1;
	wire [WIDTH-1:0] wire_d43_2;
	wire [WIDTH-1:0] wire_d43_3;
	wire [WIDTH-1:0] wire_d43_4;
	wire [WIDTH-1:0] wire_d43_5;
	wire [WIDTH-1:0] wire_d43_6;
	wire [WIDTH-1:0] wire_d43_7;
	wire [WIDTH-1:0] wire_d43_8;
	wire [WIDTH-1:0] wire_d43_9;
	wire [WIDTH-1:0] wire_d43_10;
	wire [WIDTH-1:0] wire_d43_11;
	wire [WIDTH-1:0] wire_d43_12;
	wire [WIDTH-1:0] wire_d43_13;
	wire [WIDTH-1:0] wire_d43_14;
	wire [WIDTH-1:0] wire_d43_15;
	wire [WIDTH-1:0] wire_d43_16;
	wire [WIDTH-1:0] wire_d43_17;
	wire [WIDTH-1:0] wire_d43_18;
	wire [WIDTH-1:0] wire_d43_19;
	wire [WIDTH-1:0] wire_d43_20;
	wire [WIDTH-1:0] wire_d43_21;
	wire [WIDTH-1:0] wire_d43_22;
	wire [WIDTH-1:0] wire_d43_23;
	wire [WIDTH-1:0] wire_d43_24;
	wire [WIDTH-1:0] wire_d43_25;
	wire [WIDTH-1:0] wire_d43_26;
	wire [WIDTH-1:0] wire_d43_27;
	wire [WIDTH-1:0] wire_d43_28;
	wire [WIDTH-1:0] wire_d43_29;
	wire [WIDTH-1:0] wire_d43_30;
	wire [WIDTH-1:0] wire_d43_31;
	wire [WIDTH-1:0] wire_d43_32;
	wire [WIDTH-1:0] wire_d43_33;
	wire [WIDTH-1:0] wire_d43_34;
	wire [WIDTH-1:0] wire_d43_35;
	wire [WIDTH-1:0] wire_d43_36;
	wire [WIDTH-1:0] wire_d43_37;
	wire [WIDTH-1:0] wire_d43_38;
	wire [WIDTH-1:0] wire_d43_39;
	wire [WIDTH-1:0] wire_d43_40;
	wire [WIDTH-1:0] wire_d43_41;
	wire [WIDTH-1:0] wire_d43_42;
	wire [WIDTH-1:0] wire_d43_43;
	wire [WIDTH-1:0] wire_d43_44;
	wire [WIDTH-1:0] wire_d43_45;
	wire [WIDTH-1:0] wire_d43_46;
	wire [WIDTH-1:0] wire_d43_47;
	wire [WIDTH-1:0] wire_d43_48;
	wire [WIDTH-1:0] wire_d44_0;
	wire [WIDTH-1:0] wire_d44_1;
	wire [WIDTH-1:0] wire_d44_2;
	wire [WIDTH-1:0] wire_d44_3;
	wire [WIDTH-1:0] wire_d44_4;
	wire [WIDTH-1:0] wire_d44_5;
	wire [WIDTH-1:0] wire_d44_6;
	wire [WIDTH-1:0] wire_d44_7;
	wire [WIDTH-1:0] wire_d44_8;
	wire [WIDTH-1:0] wire_d44_9;
	wire [WIDTH-1:0] wire_d44_10;
	wire [WIDTH-1:0] wire_d44_11;
	wire [WIDTH-1:0] wire_d44_12;
	wire [WIDTH-1:0] wire_d44_13;
	wire [WIDTH-1:0] wire_d44_14;
	wire [WIDTH-1:0] wire_d44_15;
	wire [WIDTH-1:0] wire_d44_16;
	wire [WIDTH-1:0] wire_d44_17;
	wire [WIDTH-1:0] wire_d44_18;
	wire [WIDTH-1:0] wire_d44_19;
	wire [WIDTH-1:0] wire_d44_20;
	wire [WIDTH-1:0] wire_d44_21;
	wire [WIDTH-1:0] wire_d44_22;
	wire [WIDTH-1:0] wire_d44_23;
	wire [WIDTH-1:0] wire_d44_24;
	wire [WIDTH-1:0] wire_d44_25;
	wire [WIDTH-1:0] wire_d44_26;
	wire [WIDTH-1:0] wire_d44_27;
	wire [WIDTH-1:0] wire_d44_28;
	wire [WIDTH-1:0] wire_d44_29;
	wire [WIDTH-1:0] wire_d44_30;
	wire [WIDTH-1:0] wire_d44_31;
	wire [WIDTH-1:0] wire_d44_32;
	wire [WIDTH-1:0] wire_d44_33;
	wire [WIDTH-1:0] wire_d44_34;
	wire [WIDTH-1:0] wire_d44_35;
	wire [WIDTH-1:0] wire_d44_36;
	wire [WIDTH-1:0] wire_d44_37;
	wire [WIDTH-1:0] wire_d44_38;
	wire [WIDTH-1:0] wire_d44_39;
	wire [WIDTH-1:0] wire_d44_40;
	wire [WIDTH-1:0] wire_d44_41;
	wire [WIDTH-1:0] wire_d44_42;
	wire [WIDTH-1:0] wire_d44_43;
	wire [WIDTH-1:0] wire_d44_44;
	wire [WIDTH-1:0] wire_d44_45;
	wire [WIDTH-1:0] wire_d44_46;
	wire [WIDTH-1:0] wire_d44_47;
	wire [WIDTH-1:0] wire_d44_48;
	wire [WIDTH-1:0] wire_d45_0;
	wire [WIDTH-1:0] wire_d45_1;
	wire [WIDTH-1:0] wire_d45_2;
	wire [WIDTH-1:0] wire_d45_3;
	wire [WIDTH-1:0] wire_d45_4;
	wire [WIDTH-1:0] wire_d45_5;
	wire [WIDTH-1:0] wire_d45_6;
	wire [WIDTH-1:0] wire_d45_7;
	wire [WIDTH-1:0] wire_d45_8;
	wire [WIDTH-1:0] wire_d45_9;
	wire [WIDTH-1:0] wire_d45_10;
	wire [WIDTH-1:0] wire_d45_11;
	wire [WIDTH-1:0] wire_d45_12;
	wire [WIDTH-1:0] wire_d45_13;
	wire [WIDTH-1:0] wire_d45_14;
	wire [WIDTH-1:0] wire_d45_15;
	wire [WIDTH-1:0] wire_d45_16;
	wire [WIDTH-1:0] wire_d45_17;
	wire [WIDTH-1:0] wire_d45_18;
	wire [WIDTH-1:0] wire_d45_19;
	wire [WIDTH-1:0] wire_d45_20;
	wire [WIDTH-1:0] wire_d45_21;
	wire [WIDTH-1:0] wire_d45_22;
	wire [WIDTH-1:0] wire_d45_23;
	wire [WIDTH-1:0] wire_d45_24;
	wire [WIDTH-1:0] wire_d45_25;
	wire [WIDTH-1:0] wire_d45_26;
	wire [WIDTH-1:0] wire_d45_27;
	wire [WIDTH-1:0] wire_d45_28;
	wire [WIDTH-1:0] wire_d45_29;
	wire [WIDTH-1:0] wire_d45_30;
	wire [WIDTH-1:0] wire_d45_31;
	wire [WIDTH-1:0] wire_d45_32;
	wire [WIDTH-1:0] wire_d45_33;
	wire [WIDTH-1:0] wire_d45_34;
	wire [WIDTH-1:0] wire_d45_35;
	wire [WIDTH-1:0] wire_d45_36;
	wire [WIDTH-1:0] wire_d45_37;
	wire [WIDTH-1:0] wire_d45_38;
	wire [WIDTH-1:0] wire_d45_39;
	wire [WIDTH-1:0] wire_d45_40;
	wire [WIDTH-1:0] wire_d45_41;
	wire [WIDTH-1:0] wire_d45_42;
	wire [WIDTH-1:0] wire_d45_43;
	wire [WIDTH-1:0] wire_d45_44;
	wire [WIDTH-1:0] wire_d45_45;
	wire [WIDTH-1:0] wire_d45_46;
	wire [WIDTH-1:0] wire_d45_47;
	wire [WIDTH-1:0] wire_d45_48;
	wire [WIDTH-1:0] wire_d46_0;
	wire [WIDTH-1:0] wire_d46_1;
	wire [WIDTH-1:0] wire_d46_2;
	wire [WIDTH-1:0] wire_d46_3;
	wire [WIDTH-1:0] wire_d46_4;
	wire [WIDTH-1:0] wire_d46_5;
	wire [WIDTH-1:0] wire_d46_6;
	wire [WIDTH-1:0] wire_d46_7;
	wire [WIDTH-1:0] wire_d46_8;
	wire [WIDTH-1:0] wire_d46_9;
	wire [WIDTH-1:0] wire_d46_10;
	wire [WIDTH-1:0] wire_d46_11;
	wire [WIDTH-1:0] wire_d46_12;
	wire [WIDTH-1:0] wire_d46_13;
	wire [WIDTH-1:0] wire_d46_14;
	wire [WIDTH-1:0] wire_d46_15;
	wire [WIDTH-1:0] wire_d46_16;
	wire [WIDTH-1:0] wire_d46_17;
	wire [WIDTH-1:0] wire_d46_18;
	wire [WIDTH-1:0] wire_d46_19;
	wire [WIDTH-1:0] wire_d46_20;
	wire [WIDTH-1:0] wire_d46_21;
	wire [WIDTH-1:0] wire_d46_22;
	wire [WIDTH-1:0] wire_d46_23;
	wire [WIDTH-1:0] wire_d46_24;
	wire [WIDTH-1:0] wire_d46_25;
	wire [WIDTH-1:0] wire_d46_26;
	wire [WIDTH-1:0] wire_d46_27;
	wire [WIDTH-1:0] wire_d46_28;
	wire [WIDTH-1:0] wire_d46_29;
	wire [WIDTH-1:0] wire_d46_30;
	wire [WIDTH-1:0] wire_d46_31;
	wire [WIDTH-1:0] wire_d46_32;
	wire [WIDTH-1:0] wire_d46_33;
	wire [WIDTH-1:0] wire_d46_34;
	wire [WIDTH-1:0] wire_d46_35;
	wire [WIDTH-1:0] wire_d46_36;
	wire [WIDTH-1:0] wire_d46_37;
	wire [WIDTH-1:0] wire_d46_38;
	wire [WIDTH-1:0] wire_d46_39;
	wire [WIDTH-1:0] wire_d46_40;
	wire [WIDTH-1:0] wire_d46_41;
	wire [WIDTH-1:0] wire_d46_42;
	wire [WIDTH-1:0] wire_d46_43;
	wire [WIDTH-1:0] wire_d46_44;
	wire [WIDTH-1:0] wire_d46_45;
	wire [WIDTH-1:0] wire_d46_46;
	wire [WIDTH-1:0] wire_d46_47;
	wire [WIDTH-1:0] wire_d46_48;
	wire [WIDTH-1:0] wire_d47_0;
	wire [WIDTH-1:0] wire_d47_1;
	wire [WIDTH-1:0] wire_d47_2;
	wire [WIDTH-1:0] wire_d47_3;
	wire [WIDTH-1:0] wire_d47_4;
	wire [WIDTH-1:0] wire_d47_5;
	wire [WIDTH-1:0] wire_d47_6;
	wire [WIDTH-1:0] wire_d47_7;
	wire [WIDTH-1:0] wire_d47_8;
	wire [WIDTH-1:0] wire_d47_9;
	wire [WIDTH-1:0] wire_d47_10;
	wire [WIDTH-1:0] wire_d47_11;
	wire [WIDTH-1:0] wire_d47_12;
	wire [WIDTH-1:0] wire_d47_13;
	wire [WIDTH-1:0] wire_d47_14;
	wire [WIDTH-1:0] wire_d47_15;
	wire [WIDTH-1:0] wire_d47_16;
	wire [WIDTH-1:0] wire_d47_17;
	wire [WIDTH-1:0] wire_d47_18;
	wire [WIDTH-1:0] wire_d47_19;
	wire [WIDTH-1:0] wire_d47_20;
	wire [WIDTH-1:0] wire_d47_21;
	wire [WIDTH-1:0] wire_d47_22;
	wire [WIDTH-1:0] wire_d47_23;
	wire [WIDTH-1:0] wire_d47_24;
	wire [WIDTH-1:0] wire_d47_25;
	wire [WIDTH-1:0] wire_d47_26;
	wire [WIDTH-1:0] wire_d47_27;
	wire [WIDTH-1:0] wire_d47_28;
	wire [WIDTH-1:0] wire_d47_29;
	wire [WIDTH-1:0] wire_d47_30;
	wire [WIDTH-1:0] wire_d47_31;
	wire [WIDTH-1:0] wire_d47_32;
	wire [WIDTH-1:0] wire_d47_33;
	wire [WIDTH-1:0] wire_d47_34;
	wire [WIDTH-1:0] wire_d47_35;
	wire [WIDTH-1:0] wire_d47_36;
	wire [WIDTH-1:0] wire_d47_37;
	wire [WIDTH-1:0] wire_d47_38;
	wire [WIDTH-1:0] wire_d47_39;
	wire [WIDTH-1:0] wire_d47_40;
	wire [WIDTH-1:0] wire_d47_41;
	wire [WIDTH-1:0] wire_d47_42;
	wire [WIDTH-1:0] wire_d47_43;
	wire [WIDTH-1:0] wire_d47_44;
	wire [WIDTH-1:0] wire_d47_45;
	wire [WIDTH-1:0] wire_d47_46;
	wire [WIDTH-1:0] wire_d47_47;
	wire [WIDTH-1:0] wire_d47_48;
	wire [WIDTH-1:0] wire_d48_0;
	wire [WIDTH-1:0] wire_d48_1;
	wire [WIDTH-1:0] wire_d48_2;
	wire [WIDTH-1:0] wire_d48_3;
	wire [WIDTH-1:0] wire_d48_4;
	wire [WIDTH-1:0] wire_d48_5;
	wire [WIDTH-1:0] wire_d48_6;
	wire [WIDTH-1:0] wire_d48_7;
	wire [WIDTH-1:0] wire_d48_8;
	wire [WIDTH-1:0] wire_d48_9;
	wire [WIDTH-1:0] wire_d48_10;
	wire [WIDTH-1:0] wire_d48_11;
	wire [WIDTH-1:0] wire_d48_12;
	wire [WIDTH-1:0] wire_d48_13;
	wire [WIDTH-1:0] wire_d48_14;
	wire [WIDTH-1:0] wire_d48_15;
	wire [WIDTH-1:0] wire_d48_16;
	wire [WIDTH-1:0] wire_d48_17;
	wire [WIDTH-1:0] wire_d48_18;
	wire [WIDTH-1:0] wire_d48_19;
	wire [WIDTH-1:0] wire_d48_20;
	wire [WIDTH-1:0] wire_d48_21;
	wire [WIDTH-1:0] wire_d48_22;
	wire [WIDTH-1:0] wire_d48_23;
	wire [WIDTH-1:0] wire_d48_24;
	wire [WIDTH-1:0] wire_d48_25;
	wire [WIDTH-1:0] wire_d48_26;
	wire [WIDTH-1:0] wire_d48_27;
	wire [WIDTH-1:0] wire_d48_28;
	wire [WIDTH-1:0] wire_d48_29;
	wire [WIDTH-1:0] wire_d48_30;
	wire [WIDTH-1:0] wire_d48_31;
	wire [WIDTH-1:0] wire_d48_32;
	wire [WIDTH-1:0] wire_d48_33;
	wire [WIDTH-1:0] wire_d48_34;
	wire [WIDTH-1:0] wire_d48_35;
	wire [WIDTH-1:0] wire_d48_36;
	wire [WIDTH-1:0] wire_d48_37;
	wire [WIDTH-1:0] wire_d48_38;
	wire [WIDTH-1:0] wire_d48_39;
	wire [WIDTH-1:0] wire_d48_40;
	wire [WIDTH-1:0] wire_d48_41;
	wire [WIDTH-1:0] wire_d48_42;
	wire [WIDTH-1:0] wire_d48_43;
	wire [WIDTH-1:0] wire_d48_44;
	wire [WIDTH-1:0] wire_d48_45;
	wire [WIDTH-1:0] wire_d48_46;
	wire [WIDTH-1:0] wire_d48_47;
	wire [WIDTH-1:0] wire_d48_48;
	wire [WIDTH-1:0] wire_d49_0;
	wire [WIDTH-1:0] wire_d49_1;
	wire [WIDTH-1:0] wire_d49_2;
	wire [WIDTH-1:0] wire_d49_3;
	wire [WIDTH-1:0] wire_d49_4;
	wire [WIDTH-1:0] wire_d49_5;
	wire [WIDTH-1:0] wire_d49_6;
	wire [WIDTH-1:0] wire_d49_7;
	wire [WIDTH-1:0] wire_d49_8;
	wire [WIDTH-1:0] wire_d49_9;
	wire [WIDTH-1:0] wire_d49_10;
	wire [WIDTH-1:0] wire_d49_11;
	wire [WIDTH-1:0] wire_d49_12;
	wire [WIDTH-1:0] wire_d49_13;
	wire [WIDTH-1:0] wire_d49_14;
	wire [WIDTH-1:0] wire_d49_15;
	wire [WIDTH-1:0] wire_d49_16;
	wire [WIDTH-1:0] wire_d49_17;
	wire [WIDTH-1:0] wire_d49_18;
	wire [WIDTH-1:0] wire_d49_19;
	wire [WIDTH-1:0] wire_d49_20;
	wire [WIDTH-1:0] wire_d49_21;
	wire [WIDTH-1:0] wire_d49_22;
	wire [WIDTH-1:0] wire_d49_23;
	wire [WIDTH-1:0] wire_d49_24;
	wire [WIDTH-1:0] wire_d49_25;
	wire [WIDTH-1:0] wire_d49_26;
	wire [WIDTH-1:0] wire_d49_27;
	wire [WIDTH-1:0] wire_d49_28;
	wire [WIDTH-1:0] wire_d49_29;
	wire [WIDTH-1:0] wire_d49_30;
	wire [WIDTH-1:0] wire_d49_31;
	wire [WIDTH-1:0] wire_d49_32;
	wire [WIDTH-1:0] wire_d49_33;
	wire [WIDTH-1:0] wire_d49_34;
	wire [WIDTH-1:0] wire_d49_35;
	wire [WIDTH-1:0] wire_d49_36;
	wire [WIDTH-1:0] wire_d49_37;
	wire [WIDTH-1:0] wire_d49_38;
	wire [WIDTH-1:0] wire_d49_39;
	wire [WIDTH-1:0] wire_d49_40;
	wire [WIDTH-1:0] wire_d49_41;
	wire [WIDTH-1:0] wire_d49_42;
	wire [WIDTH-1:0] wire_d49_43;
	wire [WIDTH-1:0] wire_d49_44;
	wire [WIDTH-1:0] wire_d49_45;
	wire [WIDTH-1:0] wire_d49_46;
	wire [WIDTH-1:0] wire_d49_47;
	wire [WIDTH-1:0] wire_d49_48;
	wire [WIDTH-1:0] wire_d50_0;
	wire [WIDTH-1:0] wire_d50_1;
	wire [WIDTH-1:0] wire_d50_2;
	wire [WIDTH-1:0] wire_d50_3;
	wire [WIDTH-1:0] wire_d50_4;
	wire [WIDTH-1:0] wire_d50_5;
	wire [WIDTH-1:0] wire_d50_6;
	wire [WIDTH-1:0] wire_d50_7;
	wire [WIDTH-1:0] wire_d50_8;
	wire [WIDTH-1:0] wire_d50_9;
	wire [WIDTH-1:0] wire_d50_10;
	wire [WIDTH-1:0] wire_d50_11;
	wire [WIDTH-1:0] wire_d50_12;
	wire [WIDTH-1:0] wire_d50_13;
	wire [WIDTH-1:0] wire_d50_14;
	wire [WIDTH-1:0] wire_d50_15;
	wire [WIDTH-1:0] wire_d50_16;
	wire [WIDTH-1:0] wire_d50_17;
	wire [WIDTH-1:0] wire_d50_18;
	wire [WIDTH-1:0] wire_d50_19;
	wire [WIDTH-1:0] wire_d50_20;
	wire [WIDTH-1:0] wire_d50_21;
	wire [WIDTH-1:0] wire_d50_22;
	wire [WIDTH-1:0] wire_d50_23;
	wire [WIDTH-1:0] wire_d50_24;
	wire [WIDTH-1:0] wire_d50_25;
	wire [WIDTH-1:0] wire_d50_26;
	wire [WIDTH-1:0] wire_d50_27;
	wire [WIDTH-1:0] wire_d50_28;
	wire [WIDTH-1:0] wire_d50_29;
	wire [WIDTH-1:0] wire_d50_30;
	wire [WIDTH-1:0] wire_d50_31;
	wire [WIDTH-1:0] wire_d50_32;
	wire [WIDTH-1:0] wire_d50_33;
	wire [WIDTH-1:0] wire_d50_34;
	wire [WIDTH-1:0] wire_d50_35;
	wire [WIDTH-1:0] wire_d50_36;
	wire [WIDTH-1:0] wire_d50_37;
	wire [WIDTH-1:0] wire_d50_38;
	wire [WIDTH-1:0] wire_d50_39;
	wire [WIDTH-1:0] wire_d50_40;
	wire [WIDTH-1:0] wire_d50_41;
	wire [WIDTH-1:0] wire_d50_42;
	wire [WIDTH-1:0] wire_d50_43;
	wire [WIDTH-1:0] wire_d50_44;
	wire [WIDTH-1:0] wire_d50_45;
	wire [WIDTH-1:0] wire_d50_46;
	wire [WIDTH-1:0] wire_d50_47;
	wire [WIDTH-1:0] wire_d50_48;
	wire [WIDTH-1:0] wire_d51_0;
	wire [WIDTH-1:0] wire_d51_1;
	wire [WIDTH-1:0] wire_d51_2;
	wire [WIDTH-1:0] wire_d51_3;
	wire [WIDTH-1:0] wire_d51_4;
	wire [WIDTH-1:0] wire_d51_5;
	wire [WIDTH-1:0] wire_d51_6;
	wire [WIDTH-1:0] wire_d51_7;
	wire [WIDTH-1:0] wire_d51_8;
	wire [WIDTH-1:0] wire_d51_9;
	wire [WIDTH-1:0] wire_d51_10;
	wire [WIDTH-1:0] wire_d51_11;
	wire [WIDTH-1:0] wire_d51_12;
	wire [WIDTH-1:0] wire_d51_13;
	wire [WIDTH-1:0] wire_d51_14;
	wire [WIDTH-1:0] wire_d51_15;
	wire [WIDTH-1:0] wire_d51_16;
	wire [WIDTH-1:0] wire_d51_17;
	wire [WIDTH-1:0] wire_d51_18;
	wire [WIDTH-1:0] wire_d51_19;
	wire [WIDTH-1:0] wire_d51_20;
	wire [WIDTH-1:0] wire_d51_21;
	wire [WIDTH-1:0] wire_d51_22;
	wire [WIDTH-1:0] wire_d51_23;
	wire [WIDTH-1:0] wire_d51_24;
	wire [WIDTH-1:0] wire_d51_25;
	wire [WIDTH-1:0] wire_d51_26;
	wire [WIDTH-1:0] wire_d51_27;
	wire [WIDTH-1:0] wire_d51_28;
	wire [WIDTH-1:0] wire_d51_29;
	wire [WIDTH-1:0] wire_d51_30;
	wire [WIDTH-1:0] wire_d51_31;
	wire [WIDTH-1:0] wire_d51_32;
	wire [WIDTH-1:0] wire_d51_33;
	wire [WIDTH-1:0] wire_d51_34;
	wire [WIDTH-1:0] wire_d51_35;
	wire [WIDTH-1:0] wire_d51_36;
	wire [WIDTH-1:0] wire_d51_37;
	wire [WIDTH-1:0] wire_d51_38;
	wire [WIDTH-1:0] wire_d51_39;
	wire [WIDTH-1:0] wire_d51_40;
	wire [WIDTH-1:0] wire_d51_41;
	wire [WIDTH-1:0] wire_d51_42;
	wire [WIDTH-1:0] wire_d51_43;
	wire [WIDTH-1:0] wire_d51_44;
	wire [WIDTH-1:0] wire_d51_45;
	wire [WIDTH-1:0] wire_d51_46;
	wire [WIDTH-1:0] wire_d51_47;
	wire [WIDTH-1:0] wire_d51_48;
	wire [WIDTH-1:0] wire_d52_0;
	wire [WIDTH-1:0] wire_d52_1;
	wire [WIDTH-1:0] wire_d52_2;
	wire [WIDTH-1:0] wire_d52_3;
	wire [WIDTH-1:0] wire_d52_4;
	wire [WIDTH-1:0] wire_d52_5;
	wire [WIDTH-1:0] wire_d52_6;
	wire [WIDTH-1:0] wire_d52_7;
	wire [WIDTH-1:0] wire_d52_8;
	wire [WIDTH-1:0] wire_d52_9;
	wire [WIDTH-1:0] wire_d52_10;
	wire [WIDTH-1:0] wire_d52_11;
	wire [WIDTH-1:0] wire_d52_12;
	wire [WIDTH-1:0] wire_d52_13;
	wire [WIDTH-1:0] wire_d52_14;
	wire [WIDTH-1:0] wire_d52_15;
	wire [WIDTH-1:0] wire_d52_16;
	wire [WIDTH-1:0] wire_d52_17;
	wire [WIDTH-1:0] wire_d52_18;
	wire [WIDTH-1:0] wire_d52_19;
	wire [WIDTH-1:0] wire_d52_20;
	wire [WIDTH-1:0] wire_d52_21;
	wire [WIDTH-1:0] wire_d52_22;
	wire [WIDTH-1:0] wire_d52_23;
	wire [WIDTH-1:0] wire_d52_24;
	wire [WIDTH-1:0] wire_d52_25;
	wire [WIDTH-1:0] wire_d52_26;
	wire [WIDTH-1:0] wire_d52_27;
	wire [WIDTH-1:0] wire_d52_28;
	wire [WIDTH-1:0] wire_d52_29;
	wire [WIDTH-1:0] wire_d52_30;
	wire [WIDTH-1:0] wire_d52_31;
	wire [WIDTH-1:0] wire_d52_32;
	wire [WIDTH-1:0] wire_d52_33;
	wire [WIDTH-1:0] wire_d52_34;
	wire [WIDTH-1:0] wire_d52_35;
	wire [WIDTH-1:0] wire_d52_36;
	wire [WIDTH-1:0] wire_d52_37;
	wire [WIDTH-1:0] wire_d52_38;
	wire [WIDTH-1:0] wire_d52_39;
	wire [WIDTH-1:0] wire_d52_40;
	wire [WIDTH-1:0] wire_d52_41;
	wire [WIDTH-1:0] wire_d52_42;
	wire [WIDTH-1:0] wire_d52_43;
	wire [WIDTH-1:0] wire_d52_44;
	wire [WIDTH-1:0] wire_d52_45;
	wire [WIDTH-1:0] wire_d52_46;
	wire [WIDTH-1:0] wire_d52_47;
	wire [WIDTH-1:0] wire_d52_48;
	wire [WIDTH-1:0] wire_d53_0;
	wire [WIDTH-1:0] wire_d53_1;
	wire [WIDTH-1:0] wire_d53_2;
	wire [WIDTH-1:0] wire_d53_3;
	wire [WIDTH-1:0] wire_d53_4;
	wire [WIDTH-1:0] wire_d53_5;
	wire [WIDTH-1:0] wire_d53_6;
	wire [WIDTH-1:0] wire_d53_7;
	wire [WIDTH-1:0] wire_d53_8;
	wire [WIDTH-1:0] wire_d53_9;
	wire [WIDTH-1:0] wire_d53_10;
	wire [WIDTH-1:0] wire_d53_11;
	wire [WIDTH-1:0] wire_d53_12;
	wire [WIDTH-1:0] wire_d53_13;
	wire [WIDTH-1:0] wire_d53_14;
	wire [WIDTH-1:0] wire_d53_15;
	wire [WIDTH-1:0] wire_d53_16;
	wire [WIDTH-1:0] wire_d53_17;
	wire [WIDTH-1:0] wire_d53_18;
	wire [WIDTH-1:0] wire_d53_19;
	wire [WIDTH-1:0] wire_d53_20;
	wire [WIDTH-1:0] wire_d53_21;
	wire [WIDTH-1:0] wire_d53_22;
	wire [WIDTH-1:0] wire_d53_23;
	wire [WIDTH-1:0] wire_d53_24;
	wire [WIDTH-1:0] wire_d53_25;
	wire [WIDTH-1:0] wire_d53_26;
	wire [WIDTH-1:0] wire_d53_27;
	wire [WIDTH-1:0] wire_d53_28;
	wire [WIDTH-1:0] wire_d53_29;
	wire [WIDTH-1:0] wire_d53_30;
	wire [WIDTH-1:0] wire_d53_31;
	wire [WIDTH-1:0] wire_d53_32;
	wire [WIDTH-1:0] wire_d53_33;
	wire [WIDTH-1:0] wire_d53_34;
	wire [WIDTH-1:0] wire_d53_35;
	wire [WIDTH-1:0] wire_d53_36;
	wire [WIDTH-1:0] wire_d53_37;
	wire [WIDTH-1:0] wire_d53_38;
	wire [WIDTH-1:0] wire_d53_39;
	wire [WIDTH-1:0] wire_d53_40;
	wire [WIDTH-1:0] wire_d53_41;
	wire [WIDTH-1:0] wire_d53_42;
	wire [WIDTH-1:0] wire_d53_43;
	wire [WIDTH-1:0] wire_d53_44;
	wire [WIDTH-1:0] wire_d53_45;
	wire [WIDTH-1:0] wire_d53_46;
	wire [WIDTH-1:0] wire_d53_47;
	wire [WIDTH-1:0] wire_d53_48;
	wire [WIDTH-1:0] wire_d54_0;
	wire [WIDTH-1:0] wire_d54_1;
	wire [WIDTH-1:0] wire_d54_2;
	wire [WIDTH-1:0] wire_d54_3;
	wire [WIDTH-1:0] wire_d54_4;
	wire [WIDTH-1:0] wire_d54_5;
	wire [WIDTH-1:0] wire_d54_6;
	wire [WIDTH-1:0] wire_d54_7;
	wire [WIDTH-1:0] wire_d54_8;
	wire [WIDTH-1:0] wire_d54_9;
	wire [WIDTH-1:0] wire_d54_10;
	wire [WIDTH-1:0] wire_d54_11;
	wire [WIDTH-1:0] wire_d54_12;
	wire [WIDTH-1:0] wire_d54_13;
	wire [WIDTH-1:0] wire_d54_14;
	wire [WIDTH-1:0] wire_d54_15;
	wire [WIDTH-1:0] wire_d54_16;
	wire [WIDTH-1:0] wire_d54_17;
	wire [WIDTH-1:0] wire_d54_18;
	wire [WIDTH-1:0] wire_d54_19;
	wire [WIDTH-1:0] wire_d54_20;
	wire [WIDTH-1:0] wire_d54_21;
	wire [WIDTH-1:0] wire_d54_22;
	wire [WIDTH-1:0] wire_d54_23;
	wire [WIDTH-1:0] wire_d54_24;
	wire [WIDTH-1:0] wire_d54_25;
	wire [WIDTH-1:0] wire_d54_26;
	wire [WIDTH-1:0] wire_d54_27;
	wire [WIDTH-1:0] wire_d54_28;
	wire [WIDTH-1:0] wire_d54_29;
	wire [WIDTH-1:0] wire_d54_30;
	wire [WIDTH-1:0] wire_d54_31;
	wire [WIDTH-1:0] wire_d54_32;
	wire [WIDTH-1:0] wire_d54_33;
	wire [WIDTH-1:0] wire_d54_34;
	wire [WIDTH-1:0] wire_d54_35;
	wire [WIDTH-1:0] wire_d54_36;
	wire [WIDTH-1:0] wire_d54_37;
	wire [WIDTH-1:0] wire_d54_38;
	wire [WIDTH-1:0] wire_d54_39;
	wire [WIDTH-1:0] wire_d54_40;
	wire [WIDTH-1:0] wire_d54_41;
	wire [WIDTH-1:0] wire_d54_42;
	wire [WIDTH-1:0] wire_d54_43;
	wire [WIDTH-1:0] wire_d54_44;
	wire [WIDTH-1:0] wire_d54_45;
	wire [WIDTH-1:0] wire_d54_46;
	wire [WIDTH-1:0] wire_d54_47;
	wire [WIDTH-1:0] wire_d54_48;

	large_adder #(.WIDTH(WIDTH)) large_adder_instance100(.data_in(d_in0),.data_out(wire_d0_0),.clk(clk),.rst(rst));            //channel 1
	large_mux #(.WIDTH(WIDTH)) large_mux_instance101(.data_in(wire_d0_0),.data_out(wire_d0_1),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance102(.data_in(wire_d0_1),.data_out(wire_d0_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance103(.data_in(wire_d0_2),.data_out(wire_d0_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance104(.data_in(wire_d0_3),.data_out(wire_d0_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance105(.data_in(wire_d0_4),.data_out(wire_d0_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance106(.data_in(wire_d0_5),.data_out(wire_d0_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance107(.data_in(wire_d0_6),.data_out(wire_d0_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance108(.data_in(wire_d0_7),.data_out(wire_d0_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance109(.data_in(wire_d0_8),.data_out(wire_d0_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1010(.data_in(wire_d0_9),.data_out(wire_d0_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1011(.data_in(wire_d0_10),.data_out(wire_d0_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1012(.data_in(wire_d0_11),.data_out(wire_d0_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1013(.data_in(wire_d0_12),.data_out(wire_d0_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1014(.data_in(wire_d0_13),.data_out(wire_d0_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1015(.data_in(wire_d0_14),.data_out(wire_d0_15),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1016(.data_in(wire_d0_15),.data_out(wire_d0_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1017(.data_in(wire_d0_16),.data_out(wire_d0_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1018(.data_in(wire_d0_17),.data_out(wire_d0_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1019(.data_in(wire_d0_18),.data_out(wire_d0_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1020(.data_in(wire_d0_19),.data_out(wire_d0_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1021(.data_in(wire_d0_20),.data_out(wire_d0_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1022(.data_in(wire_d0_21),.data_out(wire_d0_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1023(.data_in(wire_d0_22),.data_out(wire_d0_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1024(.data_in(wire_d0_23),.data_out(wire_d0_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1025(.data_in(wire_d0_24),.data_out(wire_d0_25),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1026(.data_in(wire_d0_25),.data_out(wire_d0_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1027(.data_in(wire_d0_26),.data_out(wire_d0_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1028(.data_in(wire_d0_27),.data_out(wire_d0_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1029(.data_in(wire_d0_28),.data_out(wire_d0_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1030(.data_in(wire_d0_29),.data_out(wire_d0_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1031(.data_in(wire_d0_30),.data_out(wire_d0_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1032(.data_in(wire_d0_31),.data_out(wire_d0_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1033(.data_in(wire_d0_32),.data_out(wire_d0_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1034(.data_in(wire_d0_33),.data_out(wire_d0_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1035(.data_in(wire_d0_34),.data_out(wire_d0_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1036(.data_in(wire_d0_35),.data_out(wire_d0_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1037(.data_in(wire_d0_36),.data_out(wire_d0_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1038(.data_in(wire_d0_37),.data_out(wire_d0_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1039(.data_in(wire_d0_38),.data_out(wire_d0_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1040(.data_in(wire_d0_39),.data_out(wire_d0_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1041(.data_in(wire_d0_40),.data_out(wire_d0_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1042(.data_in(wire_d0_41),.data_out(wire_d0_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1043(.data_in(wire_d0_42),.data_out(wire_d0_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1044(.data_in(wire_d0_43),.data_out(wire_d0_44),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1045(.data_in(wire_d0_44),.data_out(wire_d0_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1046(.data_in(wire_d0_45),.data_out(wire_d0_46),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1047(.data_in(wire_d0_46),.data_out(wire_d0_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1048(.data_in(wire_d0_47),.data_out(wire_d0_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1049(.data_in(wire_d0_48),.data_out(d_out0),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance210(.data_in(d_in1),.data_out(wire_d1_0),.clk(clk),.rst(rst));            //channel 2
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance211(.data_in(wire_d1_0),.data_out(wire_d1_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance212(.data_in(wire_d1_1),.data_out(wire_d1_2),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance213(.data_in(wire_d1_2),.data_out(wire_d1_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance214(.data_in(wire_d1_3),.data_out(wire_d1_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance215(.data_in(wire_d1_4),.data_out(wire_d1_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance216(.data_in(wire_d1_5),.data_out(wire_d1_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance217(.data_in(wire_d1_6),.data_out(wire_d1_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance218(.data_in(wire_d1_7),.data_out(wire_d1_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance219(.data_in(wire_d1_8),.data_out(wire_d1_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2110(.data_in(wire_d1_9),.data_out(wire_d1_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2111(.data_in(wire_d1_10),.data_out(wire_d1_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2112(.data_in(wire_d1_11),.data_out(wire_d1_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2113(.data_in(wire_d1_12),.data_out(wire_d1_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2114(.data_in(wire_d1_13),.data_out(wire_d1_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2115(.data_in(wire_d1_14),.data_out(wire_d1_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2116(.data_in(wire_d1_15),.data_out(wire_d1_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2117(.data_in(wire_d1_16),.data_out(wire_d1_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2118(.data_in(wire_d1_17),.data_out(wire_d1_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2119(.data_in(wire_d1_18),.data_out(wire_d1_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2120(.data_in(wire_d1_19),.data_out(wire_d1_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2121(.data_in(wire_d1_20),.data_out(wire_d1_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2122(.data_in(wire_d1_21),.data_out(wire_d1_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2123(.data_in(wire_d1_22),.data_out(wire_d1_23),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2124(.data_in(wire_d1_23),.data_out(wire_d1_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2125(.data_in(wire_d1_24),.data_out(wire_d1_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2126(.data_in(wire_d1_25),.data_out(wire_d1_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2127(.data_in(wire_d1_26),.data_out(wire_d1_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2128(.data_in(wire_d1_27),.data_out(wire_d1_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2129(.data_in(wire_d1_28),.data_out(wire_d1_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2130(.data_in(wire_d1_29),.data_out(wire_d1_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2131(.data_in(wire_d1_30),.data_out(wire_d1_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2132(.data_in(wire_d1_31),.data_out(wire_d1_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2133(.data_in(wire_d1_32),.data_out(wire_d1_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2134(.data_in(wire_d1_33),.data_out(wire_d1_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2135(.data_in(wire_d1_34),.data_out(wire_d1_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2136(.data_in(wire_d1_35),.data_out(wire_d1_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2137(.data_in(wire_d1_36),.data_out(wire_d1_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2138(.data_in(wire_d1_37),.data_out(wire_d1_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2139(.data_in(wire_d1_38),.data_out(wire_d1_39),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2140(.data_in(wire_d1_39),.data_out(wire_d1_40),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2141(.data_in(wire_d1_40),.data_out(wire_d1_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2142(.data_in(wire_d1_41),.data_out(wire_d1_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2143(.data_in(wire_d1_42),.data_out(wire_d1_43),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2144(.data_in(wire_d1_43),.data_out(wire_d1_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2145(.data_in(wire_d1_44),.data_out(wire_d1_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2146(.data_in(wire_d1_45),.data_out(wire_d1_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2147(.data_in(wire_d1_46),.data_out(wire_d1_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2148(.data_in(wire_d1_47),.data_out(wire_d1_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2149(.data_in(wire_d1_48),.data_out(d_out1),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance320(.data_in(d_in2),.data_out(wire_d2_0),.clk(clk),.rst(rst));            //channel 3
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance321(.data_in(wire_d2_0),.data_out(wire_d2_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance322(.data_in(wire_d2_1),.data_out(wire_d2_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance323(.data_in(wire_d2_2),.data_out(wire_d2_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance324(.data_in(wire_d2_3),.data_out(wire_d2_4),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance325(.data_in(wire_d2_4),.data_out(wire_d2_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance326(.data_in(wire_d2_5),.data_out(wire_d2_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance327(.data_in(wire_d2_6),.data_out(wire_d2_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance328(.data_in(wire_d2_7),.data_out(wire_d2_8),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance329(.data_in(wire_d2_8),.data_out(wire_d2_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3210(.data_in(wire_d2_9),.data_out(wire_d2_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3211(.data_in(wire_d2_10),.data_out(wire_d2_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3212(.data_in(wire_d2_11),.data_out(wire_d2_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3213(.data_in(wire_d2_12),.data_out(wire_d2_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3214(.data_in(wire_d2_13),.data_out(wire_d2_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3215(.data_in(wire_d2_14),.data_out(wire_d2_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3216(.data_in(wire_d2_15),.data_out(wire_d2_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3217(.data_in(wire_d2_16),.data_out(wire_d2_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3218(.data_in(wire_d2_17),.data_out(wire_d2_18),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3219(.data_in(wire_d2_18),.data_out(wire_d2_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3220(.data_in(wire_d2_19),.data_out(wire_d2_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3221(.data_in(wire_d2_20),.data_out(wire_d2_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3222(.data_in(wire_d2_21),.data_out(wire_d2_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3223(.data_in(wire_d2_22),.data_out(wire_d2_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3224(.data_in(wire_d2_23),.data_out(wire_d2_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3225(.data_in(wire_d2_24),.data_out(wire_d2_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3226(.data_in(wire_d2_25),.data_out(wire_d2_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3227(.data_in(wire_d2_26),.data_out(wire_d2_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3228(.data_in(wire_d2_27),.data_out(wire_d2_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3229(.data_in(wire_d2_28),.data_out(wire_d2_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3230(.data_in(wire_d2_29),.data_out(wire_d2_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3231(.data_in(wire_d2_30),.data_out(wire_d2_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3232(.data_in(wire_d2_31),.data_out(wire_d2_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3233(.data_in(wire_d2_32),.data_out(wire_d2_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3234(.data_in(wire_d2_33),.data_out(wire_d2_34),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3235(.data_in(wire_d2_34),.data_out(wire_d2_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3236(.data_in(wire_d2_35),.data_out(wire_d2_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3237(.data_in(wire_d2_36),.data_out(wire_d2_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3238(.data_in(wire_d2_37),.data_out(wire_d2_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3239(.data_in(wire_d2_38),.data_out(wire_d2_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3240(.data_in(wire_d2_39),.data_out(wire_d2_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3241(.data_in(wire_d2_40),.data_out(wire_d2_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3242(.data_in(wire_d2_41),.data_out(wire_d2_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3243(.data_in(wire_d2_42),.data_out(wire_d2_43),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3244(.data_in(wire_d2_43),.data_out(wire_d2_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3245(.data_in(wire_d2_44),.data_out(wire_d2_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3246(.data_in(wire_d2_45),.data_out(wire_d2_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3247(.data_in(wire_d2_46),.data_out(wire_d2_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3248(.data_in(wire_d2_47),.data_out(wire_d2_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3249(.data_in(wire_d2_48),.data_out(d_out2),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance430(.data_in(d_in3),.data_out(wire_d3_0),.clk(clk),.rst(rst));            //channel 4
	invertion #(.WIDTH(WIDTH)) invertion_instance431(.data_in(wire_d3_0),.data_out(wire_d3_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance432(.data_in(wire_d3_1),.data_out(wire_d3_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance433(.data_in(wire_d3_2),.data_out(wire_d3_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance434(.data_in(wire_d3_3),.data_out(wire_d3_4),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance435(.data_in(wire_d3_4),.data_out(wire_d3_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance436(.data_in(wire_d3_5),.data_out(wire_d3_6),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance437(.data_in(wire_d3_6),.data_out(wire_d3_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance438(.data_in(wire_d3_7),.data_out(wire_d3_8),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance439(.data_in(wire_d3_8),.data_out(wire_d3_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4310(.data_in(wire_d3_9),.data_out(wire_d3_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4311(.data_in(wire_d3_10),.data_out(wire_d3_11),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4312(.data_in(wire_d3_11),.data_out(wire_d3_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4313(.data_in(wire_d3_12),.data_out(wire_d3_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4314(.data_in(wire_d3_13),.data_out(wire_d3_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4315(.data_in(wire_d3_14),.data_out(wire_d3_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4316(.data_in(wire_d3_15),.data_out(wire_d3_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4317(.data_in(wire_d3_16),.data_out(wire_d3_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4318(.data_in(wire_d3_17),.data_out(wire_d3_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4319(.data_in(wire_d3_18),.data_out(wire_d3_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4320(.data_in(wire_d3_19),.data_out(wire_d3_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4321(.data_in(wire_d3_20),.data_out(wire_d3_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4322(.data_in(wire_d3_21),.data_out(wire_d3_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4323(.data_in(wire_d3_22),.data_out(wire_d3_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4324(.data_in(wire_d3_23),.data_out(wire_d3_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4325(.data_in(wire_d3_24),.data_out(wire_d3_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4326(.data_in(wire_d3_25),.data_out(wire_d3_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4327(.data_in(wire_d3_26),.data_out(wire_d3_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4328(.data_in(wire_d3_27),.data_out(wire_d3_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4329(.data_in(wire_d3_28),.data_out(wire_d3_29),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4330(.data_in(wire_d3_29),.data_out(wire_d3_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4331(.data_in(wire_d3_30),.data_out(wire_d3_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4332(.data_in(wire_d3_31),.data_out(wire_d3_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4333(.data_in(wire_d3_32),.data_out(wire_d3_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4334(.data_in(wire_d3_33),.data_out(wire_d3_34),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4335(.data_in(wire_d3_34),.data_out(wire_d3_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4336(.data_in(wire_d3_35),.data_out(wire_d3_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4337(.data_in(wire_d3_36),.data_out(wire_d3_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4338(.data_in(wire_d3_37),.data_out(wire_d3_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4339(.data_in(wire_d3_38),.data_out(wire_d3_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4340(.data_in(wire_d3_39),.data_out(wire_d3_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4341(.data_in(wire_d3_40),.data_out(wire_d3_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4342(.data_in(wire_d3_41),.data_out(wire_d3_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4343(.data_in(wire_d3_42),.data_out(wire_d3_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4344(.data_in(wire_d3_43),.data_out(wire_d3_44),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4345(.data_in(wire_d3_44),.data_out(wire_d3_45),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4346(.data_in(wire_d3_45),.data_out(wire_d3_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4347(.data_in(wire_d3_46),.data_out(wire_d3_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4348(.data_in(wire_d3_47),.data_out(wire_d3_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4349(.data_in(wire_d3_48),.data_out(d_out3),.clk(clk),.rst(rst));

	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance540(.data_in(d_in4),.data_out(wire_d4_0),.clk(clk),.rst(rst));            //channel 5
	large_mux #(.WIDTH(WIDTH)) large_mux_instance541(.data_in(wire_d4_0),.data_out(wire_d4_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance542(.data_in(wire_d4_1),.data_out(wire_d4_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance543(.data_in(wire_d4_2),.data_out(wire_d4_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance544(.data_in(wire_d4_3),.data_out(wire_d4_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance545(.data_in(wire_d4_4),.data_out(wire_d4_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance546(.data_in(wire_d4_5),.data_out(wire_d4_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance547(.data_in(wire_d4_6),.data_out(wire_d4_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance548(.data_in(wire_d4_7),.data_out(wire_d4_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance549(.data_in(wire_d4_8),.data_out(wire_d4_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5410(.data_in(wire_d4_9),.data_out(wire_d4_10),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5411(.data_in(wire_d4_10),.data_out(wire_d4_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5412(.data_in(wire_d4_11),.data_out(wire_d4_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5413(.data_in(wire_d4_12),.data_out(wire_d4_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5414(.data_in(wire_d4_13),.data_out(wire_d4_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5415(.data_in(wire_d4_14),.data_out(wire_d4_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5416(.data_in(wire_d4_15),.data_out(wire_d4_16),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5417(.data_in(wire_d4_16),.data_out(wire_d4_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5418(.data_in(wire_d4_17),.data_out(wire_d4_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5419(.data_in(wire_d4_18),.data_out(wire_d4_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5420(.data_in(wire_d4_19),.data_out(wire_d4_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5421(.data_in(wire_d4_20),.data_out(wire_d4_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5422(.data_in(wire_d4_21),.data_out(wire_d4_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5423(.data_in(wire_d4_22),.data_out(wire_d4_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5424(.data_in(wire_d4_23),.data_out(wire_d4_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5425(.data_in(wire_d4_24),.data_out(wire_d4_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5426(.data_in(wire_d4_25),.data_out(wire_d4_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5427(.data_in(wire_d4_26),.data_out(wire_d4_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5428(.data_in(wire_d4_27),.data_out(wire_d4_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5429(.data_in(wire_d4_28),.data_out(wire_d4_29),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5430(.data_in(wire_d4_29),.data_out(wire_d4_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5431(.data_in(wire_d4_30),.data_out(wire_d4_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5432(.data_in(wire_d4_31),.data_out(wire_d4_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5433(.data_in(wire_d4_32),.data_out(wire_d4_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5434(.data_in(wire_d4_33),.data_out(wire_d4_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5435(.data_in(wire_d4_34),.data_out(wire_d4_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5436(.data_in(wire_d4_35),.data_out(wire_d4_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5437(.data_in(wire_d4_36),.data_out(wire_d4_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5438(.data_in(wire_d4_37),.data_out(wire_d4_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5439(.data_in(wire_d4_38),.data_out(wire_d4_39),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5440(.data_in(wire_d4_39),.data_out(wire_d4_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5441(.data_in(wire_d4_40),.data_out(wire_d4_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5442(.data_in(wire_d4_41),.data_out(wire_d4_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5443(.data_in(wire_d4_42),.data_out(wire_d4_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5444(.data_in(wire_d4_43),.data_out(wire_d4_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5445(.data_in(wire_d4_44),.data_out(wire_d4_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5446(.data_in(wire_d4_45),.data_out(wire_d4_46),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5447(.data_in(wire_d4_46),.data_out(wire_d4_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5448(.data_in(wire_d4_47),.data_out(wire_d4_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5449(.data_in(wire_d4_48),.data_out(d_out4),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance650(.data_in(d_in5),.data_out(wire_d5_0),.clk(clk),.rst(rst));            //channel 6
	invertion #(.WIDTH(WIDTH)) invertion_instance651(.data_in(wire_d5_0),.data_out(wire_d5_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance652(.data_in(wire_d5_1),.data_out(wire_d5_2),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance653(.data_in(wire_d5_2),.data_out(wire_d5_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance654(.data_in(wire_d5_3),.data_out(wire_d5_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance655(.data_in(wire_d5_4),.data_out(wire_d5_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance656(.data_in(wire_d5_5),.data_out(wire_d5_6),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance657(.data_in(wire_d5_6),.data_out(wire_d5_7),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance658(.data_in(wire_d5_7),.data_out(wire_d5_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance659(.data_in(wire_d5_8),.data_out(wire_d5_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6510(.data_in(wire_d5_9),.data_out(wire_d5_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6511(.data_in(wire_d5_10),.data_out(wire_d5_11),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6512(.data_in(wire_d5_11),.data_out(wire_d5_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6513(.data_in(wire_d5_12),.data_out(wire_d5_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6514(.data_in(wire_d5_13),.data_out(wire_d5_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6515(.data_in(wire_d5_14),.data_out(wire_d5_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6516(.data_in(wire_d5_15),.data_out(wire_d5_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6517(.data_in(wire_d5_16),.data_out(wire_d5_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6518(.data_in(wire_d5_17),.data_out(wire_d5_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6519(.data_in(wire_d5_18),.data_out(wire_d5_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6520(.data_in(wire_d5_19),.data_out(wire_d5_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6521(.data_in(wire_d5_20),.data_out(wire_d5_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6522(.data_in(wire_d5_21),.data_out(wire_d5_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6523(.data_in(wire_d5_22),.data_out(wire_d5_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6524(.data_in(wire_d5_23),.data_out(wire_d5_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6525(.data_in(wire_d5_24),.data_out(wire_d5_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6526(.data_in(wire_d5_25),.data_out(wire_d5_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6527(.data_in(wire_d5_26),.data_out(wire_d5_27),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance6528(.data_in(wire_d5_27),.data_out(wire_d5_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6529(.data_in(wire_d5_28),.data_out(wire_d5_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6530(.data_in(wire_d5_29),.data_out(wire_d5_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance6531(.data_in(wire_d5_30),.data_out(wire_d5_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6532(.data_in(wire_d5_31),.data_out(wire_d5_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6533(.data_in(wire_d5_32),.data_out(wire_d5_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance6534(.data_in(wire_d5_33),.data_out(wire_d5_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance6535(.data_in(wire_d5_34),.data_out(wire_d5_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6536(.data_in(wire_d5_35),.data_out(wire_d5_36),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance6537(.data_in(wire_d5_36),.data_out(wire_d5_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance6538(.data_in(wire_d5_37),.data_out(wire_d5_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6539(.data_in(wire_d5_38),.data_out(wire_d5_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance6540(.data_in(wire_d5_39),.data_out(wire_d5_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance6541(.data_in(wire_d5_40),.data_out(wire_d5_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6542(.data_in(wire_d5_41),.data_out(wire_d5_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6543(.data_in(wire_d5_42),.data_out(wire_d5_43),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6544(.data_in(wire_d5_43),.data_out(wire_d5_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6545(.data_in(wire_d5_44),.data_out(wire_d5_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance6546(.data_in(wire_d5_45),.data_out(wire_d5_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance6547(.data_in(wire_d5_46),.data_out(wire_d5_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance6548(.data_in(wire_d5_47),.data_out(wire_d5_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance6549(.data_in(wire_d5_48),.data_out(d_out5),.clk(clk),.rst(rst));

	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance760(.data_in(d_in6),.data_out(wire_d6_0),.clk(clk),.rst(rst));            //channel 7
	decoder_top #(.WIDTH(WIDTH)) decoder_instance761(.data_in(wire_d6_0),.data_out(wire_d6_1),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance762(.data_in(wire_d6_1),.data_out(wire_d6_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance763(.data_in(wire_d6_2),.data_out(wire_d6_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance764(.data_in(wire_d6_3),.data_out(wire_d6_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance765(.data_in(wire_d6_4),.data_out(wire_d6_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance766(.data_in(wire_d6_5),.data_out(wire_d6_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance767(.data_in(wire_d6_6),.data_out(wire_d6_7),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance768(.data_in(wire_d6_7),.data_out(wire_d6_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance769(.data_in(wire_d6_8),.data_out(wire_d6_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7610(.data_in(wire_d6_9),.data_out(wire_d6_10),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7611(.data_in(wire_d6_10),.data_out(wire_d6_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7612(.data_in(wire_d6_11),.data_out(wire_d6_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7613(.data_in(wire_d6_12),.data_out(wire_d6_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7614(.data_in(wire_d6_13),.data_out(wire_d6_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7615(.data_in(wire_d6_14),.data_out(wire_d6_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7616(.data_in(wire_d6_15),.data_out(wire_d6_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7617(.data_in(wire_d6_16),.data_out(wire_d6_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7618(.data_in(wire_d6_17),.data_out(wire_d6_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7619(.data_in(wire_d6_18),.data_out(wire_d6_19),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7620(.data_in(wire_d6_19),.data_out(wire_d6_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance7621(.data_in(wire_d6_20),.data_out(wire_d6_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7622(.data_in(wire_d6_21),.data_out(wire_d6_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7623(.data_in(wire_d6_22),.data_out(wire_d6_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7624(.data_in(wire_d6_23),.data_out(wire_d6_24),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance7625(.data_in(wire_d6_24),.data_out(wire_d6_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7626(.data_in(wire_d6_25),.data_out(wire_d6_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7627(.data_in(wire_d6_26),.data_out(wire_d6_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7628(.data_in(wire_d6_27),.data_out(wire_d6_28),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7629(.data_in(wire_d6_28),.data_out(wire_d6_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7630(.data_in(wire_d6_29),.data_out(wire_d6_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7631(.data_in(wire_d6_30),.data_out(wire_d6_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7632(.data_in(wire_d6_31),.data_out(wire_d6_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance7633(.data_in(wire_d6_32),.data_out(wire_d6_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance7634(.data_in(wire_d6_33),.data_out(wire_d6_34),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance7635(.data_in(wire_d6_34),.data_out(wire_d6_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7636(.data_in(wire_d6_35),.data_out(wire_d6_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance7637(.data_in(wire_d6_36),.data_out(wire_d6_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7638(.data_in(wire_d6_37),.data_out(wire_d6_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7639(.data_in(wire_d6_38),.data_out(wire_d6_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7640(.data_in(wire_d6_39),.data_out(wire_d6_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance7641(.data_in(wire_d6_40),.data_out(wire_d6_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7642(.data_in(wire_d6_41),.data_out(wire_d6_42),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7643(.data_in(wire_d6_42),.data_out(wire_d6_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance7644(.data_in(wire_d6_43),.data_out(wire_d6_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance7645(.data_in(wire_d6_44),.data_out(wire_d6_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7646(.data_in(wire_d6_45),.data_out(wire_d6_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance7647(.data_in(wire_d6_46),.data_out(wire_d6_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance7648(.data_in(wire_d6_47),.data_out(wire_d6_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance7649(.data_in(wire_d6_48),.data_out(d_out6),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance870(.data_in(d_in7),.data_out(wire_d7_0),.clk(clk),.rst(rst));            //channel 8
	encoder #(.WIDTH(WIDTH)) encoder_instance871(.data_in(wire_d7_0),.data_out(wire_d7_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance872(.data_in(wire_d7_1),.data_out(wire_d7_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance873(.data_in(wire_d7_2),.data_out(wire_d7_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance874(.data_in(wire_d7_3),.data_out(wire_d7_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance875(.data_in(wire_d7_4),.data_out(wire_d7_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance876(.data_in(wire_d7_5),.data_out(wire_d7_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance877(.data_in(wire_d7_6),.data_out(wire_d7_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance878(.data_in(wire_d7_7),.data_out(wire_d7_8),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance879(.data_in(wire_d7_8),.data_out(wire_d7_9),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8710(.data_in(wire_d7_9),.data_out(wire_d7_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8711(.data_in(wire_d7_10),.data_out(wire_d7_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8712(.data_in(wire_d7_11),.data_out(wire_d7_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8713(.data_in(wire_d7_12),.data_out(wire_d7_13),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8714(.data_in(wire_d7_13),.data_out(wire_d7_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8715(.data_in(wire_d7_14),.data_out(wire_d7_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8716(.data_in(wire_d7_15),.data_out(wire_d7_16),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8717(.data_in(wire_d7_16),.data_out(wire_d7_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8718(.data_in(wire_d7_17),.data_out(wire_d7_18),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8719(.data_in(wire_d7_18),.data_out(wire_d7_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8720(.data_in(wire_d7_19),.data_out(wire_d7_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance8721(.data_in(wire_d7_20),.data_out(wire_d7_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance8722(.data_in(wire_d7_21),.data_out(wire_d7_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8723(.data_in(wire_d7_22),.data_out(wire_d7_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8724(.data_in(wire_d7_23),.data_out(wire_d7_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8725(.data_in(wire_d7_24),.data_out(wire_d7_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8726(.data_in(wire_d7_25),.data_out(wire_d7_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8727(.data_in(wire_d7_26),.data_out(wire_d7_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8728(.data_in(wire_d7_27),.data_out(wire_d7_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8729(.data_in(wire_d7_28),.data_out(wire_d7_29),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8730(.data_in(wire_d7_29),.data_out(wire_d7_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8731(.data_in(wire_d7_30),.data_out(wire_d7_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance8732(.data_in(wire_d7_31),.data_out(wire_d7_32),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8733(.data_in(wire_d7_32),.data_out(wire_d7_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8734(.data_in(wire_d7_33),.data_out(wire_d7_34),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance8735(.data_in(wire_d7_34),.data_out(wire_d7_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8736(.data_in(wire_d7_35),.data_out(wire_d7_36),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8737(.data_in(wire_d7_36),.data_out(wire_d7_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8738(.data_in(wire_d7_37),.data_out(wire_d7_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8739(.data_in(wire_d7_38),.data_out(wire_d7_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance8740(.data_in(wire_d7_39),.data_out(wire_d7_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8741(.data_in(wire_d7_40),.data_out(wire_d7_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8742(.data_in(wire_d7_41),.data_out(wire_d7_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance8743(.data_in(wire_d7_42),.data_out(wire_d7_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance8744(.data_in(wire_d7_43),.data_out(wire_d7_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance8745(.data_in(wire_d7_44),.data_out(wire_d7_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance8746(.data_in(wire_d7_45),.data_out(wire_d7_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance8747(.data_in(wire_d7_46),.data_out(wire_d7_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance8748(.data_in(wire_d7_47),.data_out(wire_d7_48),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance8749(.data_in(wire_d7_48),.data_out(d_out7),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance980(.data_in(d_in8),.data_out(wire_d8_0),.clk(clk),.rst(rst));            //channel 9
	large_adder #(.WIDTH(WIDTH)) large_adder_instance981(.data_in(wire_d8_0),.data_out(wire_d8_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance982(.data_in(wire_d8_1),.data_out(wire_d8_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance983(.data_in(wire_d8_2),.data_out(wire_d8_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance984(.data_in(wire_d8_3),.data_out(wire_d8_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance985(.data_in(wire_d8_4),.data_out(wire_d8_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance986(.data_in(wire_d8_5),.data_out(wire_d8_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance987(.data_in(wire_d8_6),.data_out(wire_d8_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance988(.data_in(wire_d8_7),.data_out(wire_d8_8),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance989(.data_in(wire_d8_8),.data_out(wire_d8_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9810(.data_in(wire_d8_9),.data_out(wire_d8_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9811(.data_in(wire_d8_10),.data_out(wire_d8_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9812(.data_in(wire_d8_11),.data_out(wire_d8_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9813(.data_in(wire_d8_12),.data_out(wire_d8_13),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9814(.data_in(wire_d8_13),.data_out(wire_d8_14),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9815(.data_in(wire_d8_14),.data_out(wire_d8_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9816(.data_in(wire_d8_15),.data_out(wire_d8_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9817(.data_in(wire_d8_16),.data_out(wire_d8_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9818(.data_in(wire_d8_17),.data_out(wire_d8_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9819(.data_in(wire_d8_18),.data_out(wire_d8_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance9820(.data_in(wire_d8_19),.data_out(wire_d8_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9821(.data_in(wire_d8_20),.data_out(wire_d8_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9822(.data_in(wire_d8_21),.data_out(wire_d8_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9823(.data_in(wire_d8_22),.data_out(wire_d8_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9824(.data_in(wire_d8_23),.data_out(wire_d8_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9825(.data_in(wire_d8_24),.data_out(wire_d8_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9826(.data_in(wire_d8_25),.data_out(wire_d8_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance9827(.data_in(wire_d8_26),.data_out(wire_d8_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9828(.data_in(wire_d8_27),.data_out(wire_d8_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9829(.data_in(wire_d8_28),.data_out(wire_d8_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9830(.data_in(wire_d8_29),.data_out(wire_d8_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9831(.data_in(wire_d8_30),.data_out(wire_d8_31),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9832(.data_in(wire_d8_31),.data_out(wire_d8_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance9833(.data_in(wire_d8_32),.data_out(wire_d8_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance9834(.data_in(wire_d8_33),.data_out(wire_d8_34),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance9835(.data_in(wire_d8_34),.data_out(wire_d8_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9836(.data_in(wire_d8_35),.data_out(wire_d8_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9837(.data_in(wire_d8_36),.data_out(wire_d8_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9838(.data_in(wire_d8_37),.data_out(wire_d8_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance9839(.data_in(wire_d8_38),.data_out(wire_d8_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9840(.data_in(wire_d8_39),.data_out(wire_d8_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9841(.data_in(wire_d8_40),.data_out(wire_d8_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance9842(.data_in(wire_d8_41),.data_out(wire_d8_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance9843(.data_in(wire_d8_42),.data_out(wire_d8_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9844(.data_in(wire_d8_43),.data_out(wire_d8_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance9845(.data_in(wire_d8_44),.data_out(wire_d8_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance9846(.data_in(wire_d8_45),.data_out(wire_d8_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9847(.data_in(wire_d8_46),.data_out(wire_d8_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance9848(.data_in(wire_d8_47),.data_out(wire_d8_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance9849(.data_in(wire_d8_48),.data_out(d_out8),.clk(clk),.rst(rst));

	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance10090(.data_in(d_in9),.data_out(wire_d9_0),.clk(clk),.rst(rst));            //channel 10
	invertion #(.WIDTH(WIDTH)) invertion_instance10091(.data_in(wire_d9_0),.data_out(wire_d9_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10092(.data_in(wire_d9_1),.data_out(wire_d9_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance10093(.data_in(wire_d9_2),.data_out(wire_d9_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance10094(.data_in(wire_d9_3),.data_out(wire_d9_4),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance10095(.data_in(wire_d9_4),.data_out(wire_d9_5),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance10096(.data_in(wire_d9_5),.data_out(wire_d9_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance10097(.data_in(wire_d9_6),.data_out(wire_d9_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance10098(.data_in(wire_d9_7),.data_out(wire_d9_8),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance10099(.data_in(wire_d9_8),.data_out(wire_d9_9),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance100910(.data_in(wire_d9_9),.data_out(wire_d9_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance100911(.data_in(wire_d9_10),.data_out(wire_d9_11),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance100912(.data_in(wire_d9_11),.data_out(wire_d9_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100913(.data_in(wire_d9_12),.data_out(wire_d9_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100914(.data_in(wire_d9_13),.data_out(wire_d9_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100915(.data_in(wire_d9_14),.data_out(wire_d9_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100916(.data_in(wire_d9_15),.data_out(wire_d9_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100917(.data_in(wire_d9_16),.data_out(wire_d9_17),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance100918(.data_in(wire_d9_17),.data_out(wire_d9_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100919(.data_in(wire_d9_18),.data_out(wire_d9_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100920(.data_in(wire_d9_19),.data_out(wire_d9_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100921(.data_in(wire_d9_20),.data_out(wire_d9_21),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance100922(.data_in(wire_d9_21),.data_out(wire_d9_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100923(.data_in(wire_d9_22),.data_out(wire_d9_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100924(.data_in(wire_d9_23),.data_out(wire_d9_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100925(.data_in(wire_d9_24),.data_out(wire_d9_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100926(.data_in(wire_d9_25),.data_out(wire_d9_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100927(.data_in(wire_d9_26),.data_out(wire_d9_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance100928(.data_in(wire_d9_27),.data_out(wire_d9_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100929(.data_in(wire_d9_28),.data_out(wire_d9_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance100930(.data_in(wire_d9_29),.data_out(wire_d9_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100931(.data_in(wire_d9_30),.data_out(wire_d9_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100932(.data_in(wire_d9_31),.data_out(wire_d9_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100933(.data_in(wire_d9_32),.data_out(wire_d9_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance100934(.data_in(wire_d9_33),.data_out(wire_d9_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100935(.data_in(wire_d9_34),.data_out(wire_d9_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100936(.data_in(wire_d9_35),.data_out(wire_d9_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance100937(.data_in(wire_d9_36),.data_out(wire_d9_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100938(.data_in(wire_d9_37),.data_out(wire_d9_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance100939(.data_in(wire_d9_38),.data_out(wire_d9_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance100940(.data_in(wire_d9_39),.data_out(wire_d9_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100941(.data_in(wire_d9_40),.data_out(wire_d9_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance100942(.data_in(wire_d9_41),.data_out(wire_d9_42),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100943(.data_in(wire_d9_42),.data_out(wire_d9_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100944(.data_in(wire_d9_43),.data_out(wire_d9_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance100945(.data_in(wire_d9_44),.data_out(wire_d9_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100946(.data_in(wire_d9_45),.data_out(wire_d9_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance100947(.data_in(wire_d9_46),.data_out(wire_d9_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance100948(.data_in(wire_d9_47),.data_out(wire_d9_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance100949(.data_in(wire_d9_48),.data_out(d_out9),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance110100(.data_in(d_in10),.data_out(wire_d10_0),.clk(clk),.rst(rst));            //channel 11
	large_mux #(.WIDTH(WIDTH)) large_mux_instance110101(.data_in(wire_d10_0),.data_out(wire_d10_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance110102(.data_in(wire_d10_1),.data_out(wire_d10_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance110103(.data_in(wire_d10_2),.data_out(wire_d10_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance110104(.data_in(wire_d10_3),.data_out(wire_d10_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance110105(.data_in(wire_d10_4),.data_out(wire_d10_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance110106(.data_in(wire_d10_5),.data_out(wire_d10_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance110107(.data_in(wire_d10_6),.data_out(wire_d10_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance110108(.data_in(wire_d10_7),.data_out(wire_d10_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance110109(.data_in(wire_d10_8),.data_out(wire_d10_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1101010(.data_in(wire_d10_9),.data_out(wire_d10_10),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1101011(.data_in(wire_d10_10),.data_out(wire_d10_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101012(.data_in(wire_d10_11),.data_out(wire_d10_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101013(.data_in(wire_d10_12),.data_out(wire_d10_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101014(.data_in(wire_d10_13),.data_out(wire_d10_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101015(.data_in(wire_d10_14),.data_out(wire_d10_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1101016(.data_in(wire_d10_15),.data_out(wire_d10_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1101017(.data_in(wire_d10_16),.data_out(wire_d10_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1101018(.data_in(wire_d10_17),.data_out(wire_d10_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101019(.data_in(wire_d10_18),.data_out(wire_d10_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101020(.data_in(wire_d10_19),.data_out(wire_d10_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1101021(.data_in(wire_d10_20),.data_out(wire_d10_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1101022(.data_in(wire_d10_21),.data_out(wire_d10_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1101023(.data_in(wire_d10_22),.data_out(wire_d10_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1101024(.data_in(wire_d10_23),.data_out(wire_d10_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1101025(.data_in(wire_d10_24),.data_out(wire_d10_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101026(.data_in(wire_d10_25),.data_out(wire_d10_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101027(.data_in(wire_d10_26),.data_out(wire_d10_27),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101028(.data_in(wire_d10_27),.data_out(wire_d10_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1101029(.data_in(wire_d10_28),.data_out(wire_d10_29),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1101030(.data_in(wire_d10_29),.data_out(wire_d10_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101031(.data_in(wire_d10_30),.data_out(wire_d10_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101032(.data_in(wire_d10_31),.data_out(wire_d10_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1101033(.data_in(wire_d10_32),.data_out(wire_d10_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101034(.data_in(wire_d10_33),.data_out(wire_d10_34),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1101035(.data_in(wire_d10_34),.data_out(wire_d10_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1101036(.data_in(wire_d10_35),.data_out(wire_d10_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1101037(.data_in(wire_d10_36),.data_out(wire_d10_37),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1101038(.data_in(wire_d10_37),.data_out(wire_d10_38),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101039(.data_in(wire_d10_38),.data_out(wire_d10_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101040(.data_in(wire_d10_39),.data_out(wire_d10_40),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1101041(.data_in(wire_d10_40),.data_out(wire_d10_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1101042(.data_in(wire_d10_41),.data_out(wire_d10_42),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1101043(.data_in(wire_d10_42),.data_out(wire_d10_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1101044(.data_in(wire_d10_43),.data_out(wire_d10_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1101045(.data_in(wire_d10_44),.data_out(wire_d10_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1101046(.data_in(wire_d10_45),.data_out(wire_d10_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1101047(.data_in(wire_d10_46),.data_out(wire_d10_47),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101048(.data_in(wire_d10_47),.data_out(wire_d10_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1101049(.data_in(wire_d10_48),.data_out(d_out10),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance120110(.data_in(d_in11),.data_out(wire_d11_0),.clk(clk),.rst(rst));            //channel 12
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance120111(.data_in(wire_d11_0),.data_out(wire_d11_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance120112(.data_in(wire_d11_1),.data_out(wire_d11_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance120113(.data_in(wire_d11_2),.data_out(wire_d11_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance120114(.data_in(wire_d11_3),.data_out(wire_d11_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance120115(.data_in(wire_d11_4),.data_out(wire_d11_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance120116(.data_in(wire_d11_5),.data_out(wire_d11_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance120117(.data_in(wire_d11_6),.data_out(wire_d11_7),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance120118(.data_in(wire_d11_7),.data_out(wire_d11_8),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance120119(.data_in(wire_d11_8),.data_out(wire_d11_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1201110(.data_in(wire_d11_9),.data_out(wire_d11_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201111(.data_in(wire_d11_10),.data_out(wire_d11_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201112(.data_in(wire_d11_11),.data_out(wire_d11_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201113(.data_in(wire_d11_12),.data_out(wire_d11_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201114(.data_in(wire_d11_13),.data_out(wire_d11_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1201115(.data_in(wire_d11_14),.data_out(wire_d11_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1201116(.data_in(wire_d11_15),.data_out(wire_d11_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201117(.data_in(wire_d11_16),.data_out(wire_d11_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1201118(.data_in(wire_d11_17),.data_out(wire_d11_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201119(.data_in(wire_d11_18),.data_out(wire_d11_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1201120(.data_in(wire_d11_19),.data_out(wire_d11_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201121(.data_in(wire_d11_20),.data_out(wire_d11_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201122(.data_in(wire_d11_21),.data_out(wire_d11_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201123(.data_in(wire_d11_22),.data_out(wire_d11_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201124(.data_in(wire_d11_23),.data_out(wire_d11_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1201125(.data_in(wire_d11_24),.data_out(wire_d11_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201126(.data_in(wire_d11_25),.data_out(wire_d11_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201127(.data_in(wire_d11_26),.data_out(wire_d11_27),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201128(.data_in(wire_d11_27),.data_out(wire_d11_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201129(.data_in(wire_d11_28),.data_out(wire_d11_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201130(.data_in(wire_d11_29),.data_out(wire_d11_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201131(.data_in(wire_d11_30),.data_out(wire_d11_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201132(.data_in(wire_d11_31),.data_out(wire_d11_32),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1201133(.data_in(wire_d11_32),.data_out(wire_d11_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201134(.data_in(wire_d11_33),.data_out(wire_d11_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1201135(.data_in(wire_d11_34),.data_out(wire_d11_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201136(.data_in(wire_d11_35),.data_out(wire_d11_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1201137(.data_in(wire_d11_36),.data_out(wire_d11_37),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1201138(.data_in(wire_d11_37),.data_out(wire_d11_38),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1201139(.data_in(wire_d11_38),.data_out(wire_d11_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1201140(.data_in(wire_d11_39),.data_out(wire_d11_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1201141(.data_in(wire_d11_40),.data_out(wire_d11_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1201142(.data_in(wire_d11_41),.data_out(wire_d11_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1201143(.data_in(wire_d11_42),.data_out(wire_d11_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1201144(.data_in(wire_d11_43),.data_out(wire_d11_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1201145(.data_in(wire_d11_44),.data_out(wire_d11_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1201146(.data_in(wire_d11_45),.data_out(wire_d11_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1201147(.data_in(wire_d11_46),.data_out(wire_d11_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1201148(.data_in(wire_d11_47),.data_out(wire_d11_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1201149(.data_in(wire_d11_48),.data_out(d_out11),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance130120(.data_in(d_in12),.data_out(wire_d12_0),.clk(clk),.rst(rst));            //channel 13
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance130121(.data_in(wire_d12_0),.data_out(wire_d12_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance130122(.data_in(wire_d12_1),.data_out(wire_d12_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance130123(.data_in(wire_d12_2),.data_out(wire_d12_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance130124(.data_in(wire_d12_3),.data_out(wire_d12_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance130125(.data_in(wire_d12_4),.data_out(wire_d12_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance130126(.data_in(wire_d12_5),.data_out(wire_d12_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance130127(.data_in(wire_d12_6),.data_out(wire_d12_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance130128(.data_in(wire_d12_7),.data_out(wire_d12_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance130129(.data_in(wire_d12_8),.data_out(wire_d12_9),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301210(.data_in(wire_d12_9),.data_out(wire_d12_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301211(.data_in(wire_d12_10),.data_out(wire_d12_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301212(.data_in(wire_d12_11),.data_out(wire_d12_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1301213(.data_in(wire_d12_12),.data_out(wire_d12_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1301214(.data_in(wire_d12_13),.data_out(wire_d12_14),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1301215(.data_in(wire_d12_14),.data_out(wire_d12_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301216(.data_in(wire_d12_15),.data_out(wire_d12_16),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301217(.data_in(wire_d12_16),.data_out(wire_d12_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301218(.data_in(wire_d12_17),.data_out(wire_d12_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1301219(.data_in(wire_d12_18),.data_out(wire_d12_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301220(.data_in(wire_d12_19),.data_out(wire_d12_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1301221(.data_in(wire_d12_20),.data_out(wire_d12_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301222(.data_in(wire_d12_21),.data_out(wire_d12_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301223(.data_in(wire_d12_22),.data_out(wire_d12_23),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301224(.data_in(wire_d12_23),.data_out(wire_d12_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1301225(.data_in(wire_d12_24),.data_out(wire_d12_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301226(.data_in(wire_d12_25),.data_out(wire_d12_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1301227(.data_in(wire_d12_26),.data_out(wire_d12_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301228(.data_in(wire_d12_27),.data_out(wire_d12_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1301229(.data_in(wire_d12_28),.data_out(wire_d12_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301230(.data_in(wire_d12_29),.data_out(wire_d12_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301231(.data_in(wire_d12_30),.data_out(wire_d12_31),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1301232(.data_in(wire_d12_31),.data_out(wire_d12_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301233(.data_in(wire_d12_32),.data_out(wire_d12_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301234(.data_in(wire_d12_33),.data_out(wire_d12_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301235(.data_in(wire_d12_34),.data_out(wire_d12_35),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1301236(.data_in(wire_d12_35),.data_out(wire_d12_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301237(.data_in(wire_d12_36),.data_out(wire_d12_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1301238(.data_in(wire_d12_37),.data_out(wire_d12_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1301239(.data_in(wire_d12_38),.data_out(wire_d12_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1301240(.data_in(wire_d12_39),.data_out(wire_d12_40),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1301241(.data_in(wire_d12_40),.data_out(wire_d12_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1301242(.data_in(wire_d12_41),.data_out(wire_d12_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1301243(.data_in(wire_d12_42),.data_out(wire_d12_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1301244(.data_in(wire_d12_43),.data_out(wire_d12_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1301245(.data_in(wire_d12_44),.data_out(wire_d12_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1301246(.data_in(wire_d12_45),.data_out(wire_d12_46),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1301247(.data_in(wire_d12_46),.data_out(wire_d12_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1301248(.data_in(wire_d12_47),.data_out(wire_d12_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1301249(.data_in(wire_d12_48),.data_out(d_out12),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance140130(.data_in(d_in13),.data_out(wire_d13_0),.clk(clk),.rst(rst));            //channel 14
	invertion #(.WIDTH(WIDTH)) invertion_instance140131(.data_in(wire_d13_0),.data_out(wire_d13_1),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance140132(.data_in(wire_d13_1),.data_out(wire_d13_2),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance140133(.data_in(wire_d13_2),.data_out(wire_d13_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance140134(.data_in(wire_d13_3),.data_out(wire_d13_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance140135(.data_in(wire_d13_4),.data_out(wire_d13_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance140136(.data_in(wire_d13_5),.data_out(wire_d13_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance140137(.data_in(wire_d13_6),.data_out(wire_d13_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance140138(.data_in(wire_d13_7),.data_out(wire_d13_8),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance140139(.data_in(wire_d13_8),.data_out(wire_d13_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401310(.data_in(wire_d13_9),.data_out(wire_d13_10),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401311(.data_in(wire_d13_10),.data_out(wire_d13_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401312(.data_in(wire_d13_11),.data_out(wire_d13_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1401313(.data_in(wire_d13_12),.data_out(wire_d13_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1401314(.data_in(wire_d13_13),.data_out(wire_d13_14),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1401315(.data_in(wire_d13_14),.data_out(wire_d13_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401316(.data_in(wire_d13_15),.data_out(wire_d13_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401317(.data_in(wire_d13_16),.data_out(wire_d13_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401318(.data_in(wire_d13_17),.data_out(wire_d13_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401319(.data_in(wire_d13_18),.data_out(wire_d13_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401320(.data_in(wire_d13_19),.data_out(wire_d13_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401321(.data_in(wire_d13_20),.data_out(wire_d13_21),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1401322(.data_in(wire_d13_21),.data_out(wire_d13_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1401323(.data_in(wire_d13_22),.data_out(wire_d13_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1401324(.data_in(wire_d13_23),.data_out(wire_d13_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401325(.data_in(wire_d13_24),.data_out(wire_d13_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401326(.data_in(wire_d13_25),.data_out(wire_d13_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1401327(.data_in(wire_d13_26),.data_out(wire_d13_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401328(.data_in(wire_d13_27),.data_out(wire_d13_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401329(.data_in(wire_d13_28),.data_out(wire_d13_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401330(.data_in(wire_d13_29),.data_out(wire_d13_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401331(.data_in(wire_d13_30),.data_out(wire_d13_31),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1401332(.data_in(wire_d13_31),.data_out(wire_d13_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1401333(.data_in(wire_d13_32),.data_out(wire_d13_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401334(.data_in(wire_d13_33),.data_out(wire_d13_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401335(.data_in(wire_d13_34),.data_out(wire_d13_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1401336(.data_in(wire_d13_35),.data_out(wire_d13_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1401337(.data_in(wire_d13_36),.data_out(wire_d13_37),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1401338(.data_in(wire_d13_37),.data_out(wire_d13_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1401339(.data_in(wire_d13_38),.data_out(wire_d13_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1401340(.data_in(wire_d13_39),.data_out(wire_d13_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1401341(.data_in(wire_d13_40),.data_out(wire_d13_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1401342(.data_in(wire_d13_41),.data_out(wire_d13_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1401343(.data_in(wire_d13_42),.data_out(wire_d13_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1401344(.data_in(wire_d13_43),.data_out(wire_d13_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1401345(.data_in(wire_d13_44),.data_out(wire_d13_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1401346(.data_in(wire_d13_45),.data_out(wire_d13_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1401347(.data_in(wire_d13_46),.data_out(wire_d13_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1401348(.data_in(wire_d13_47),.data_out(wire_d13_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1401349(.data_in(wire_d13_48),.data_out(d_out13),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance150140(.data_in(d_in14),.data_out(wire_d14_0),.clk(clk),.rst(rst));            //channel 15
	decoder_top #(.WIDTH(WIDTH)) decoder_instance150141(.data_in(wire_d14_0),.data_out(wire_d14_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance150142(.data_in(wire_d14_1),.data_out(wire_d14_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance150143(.data_in(wire_d14_2),.data_out(wire_d14_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance150144(.data_in(wire_d14_3),.data_out(wire_d14_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance150145(.data_in(wire_d14_4),.data_out(wire_d14_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance150146(.data_in(wire_d14_5),.data_out(wire_d14_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance150147(.data_in(wire_d14_6),.data_out(wire_d14_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance150148(.data_in(wire_d14_7),.data_out(wire_d14_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance150149(.data_in(wire_d14_8),.data_out(wire_d14_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501410(.data_in(wire_d14_9),.data_out(wire_d14_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1501411(.data_in(wire_d14_10),.data_out(wire_d14_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1501412(.data_in(wire_d14_11),.data_out(wire_d14_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501413(.data_in(wire_d14_12),.data_out(wire_d14_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501414(.data_in(wire_d14_13),.data_out(wire_d14_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501415(.data_in(wire_d14_14),.data_out(wire_d14_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1501416(.data_in(wire_d14_15),.data_out(wire_d14_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501417(.data_in(wire_d14_16),.data_out(wire_d14_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501418(.data_in(wire_d14_17),.data_out(wire_d14_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501419(.data_in(wire_d14_18),.data_out(wire_d14_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501420(.data_in(wire_d14_19),.data_out(wire_d14_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1501421(.data_in(wire_d14_20),.data_out(wire_d14_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1501422(.data_in(wire_d14_21),.data_out(wire_d14_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501423(.data_in(wire_d14_22),.data_out(wire_d14_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501424(.data_in(wire_d14_23),.data_out(wire_d14_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1501425(.data_in(wire_d14_24),.data_out(wire_d14_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501426(.data_in(wire_d14_25),.data_out(wire_d14_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501427(.data_in(wire_d14_26),.data_out(wire_d14_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1501428(.data_in(wire_d14_27),.data_out(wire_d14_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1501429(.data_in(wire_d14_28),.data_out(wire_d14_29),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1501430(.data_in(wire_d14_29),.data_out(wire_d14_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501431(.data_in(wire_d14_30),.data_out(wire_d14_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1501432(.data_in(wire_d14_31),.data_out(wire_d14_32),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1501433(.data_in(wire_d14_32),.data_out(wire_d14_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1501434(.data_in(wire_d14_33),.data_out(wire_d14_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1501435(.data_in(wire_d14_34),.data_out(wire_d14_35),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1501436(.data_in(wire_d14_35),.data_out(wire_d14_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1501437(.data_in(wire_d14_36),.data_out(wire_d14_37),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501438(.data_in(wire_d14_37),.data_out(wire_d14_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1501439(.data_in(wire_d14_38),.data_out(wire_d14_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1501440(.data_in(wire_d14_39),.data_out(wire_d14_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1501441(.data_in(wire_d14_40),.data_out(wire_d14_41),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1501442(.data_in(wire_d14_41),.data_out(wire_d14_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1501443(.data_in(wire_d14_42),.data_out(wire_d14_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1501444(.data_in(wire_d14_43),.data_out(wire_d14_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1501445(.data_in(wire_d14_44),.data_out(wire_d14_45),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1501446(.data_in(wire_d14_45),.data_out(wire_d14_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1501447(.data_in(wire_d14_46),.data_out(wire_d14_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1501448(.data_in(wire_d14_47),.data_out(wire_d14_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1501449(.data_in(wire_d14_48),.data_out(d_out14),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance160150(.data_in(d_in15),.data_out(wire_d15_0),.clk(clk),.rst(rst));            //channel 16
	register #(.WIDTH(WIDTH)) register_instance160151(.data_in(wire_d15_0),.data_out(wire_d15_1),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance160152(.data_in(wire_d15_1),.data_out(wire_d15_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance160153(.data_in(wire_d15_2),.data_out(wire_d15_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance160154(.data_in(wire_d15_3),.data_out(wire_d15_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance160155(.data_in(wire_d15_4),.data_out(wire_d15_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance160156(.data_in(wire_d15_5),.data_out(wire_d15_6),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance160157(.data_in(wire_d15_6),.data_out(wire_d15_7),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance160158(.data_in(wire_d15_7),.data_out(wire_d15_8),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance160159(.data_in(wire_d15_8),.data_out(wire_d15_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1601510(.data_in(wire_d15_9),.data_out(wire_d15_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1601511(.data_in(wire_d15_10),.data_out(wire_d15_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601512(.data_in(wire_d15_11),.data_out(wire_d15_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601513(.data_in(wire_d15_12),.data_out(wire_d15_13),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601514(.data_in(wire_d15_13),.data_out(wire_d15_14),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601515(.data_in(wire_d15_14),.data_out(wire_d15_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601516(.data_in(wire_d15_15),.data_out(wire_d15_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601517(.data_in(wire_d15_16),.data_out(wire_d15_17),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1601518(.data_in(wire_d15_17),.data_out(wire_d15_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601519(.data_in(wire_d15_18),.data_out(wire_d15_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601520(.data_in(wire_d15_19),.data_out(wire_d15_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601521(.data_in(wire_d15_20),.data_out(wire_d15_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1601522(.data_in(wire_d15_21),.data_out(wire_d15_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601523(.data_in(wire_d15_22),.data_out(wire_d15_23),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1601524(.data_in(wire_d15_23),.data_out(wire_d15_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601525(.data_in(wire_d15_24),.data_out(wire_d15_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1601526(.data_in(wire_d15_25),.data_out(wire_d15_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1601527(.data_in(wire_d15_26),.data_out(wire_d15_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601528(.data_in(wire_d15_27),.data_out(wire_d15_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1601529(.data_in(wire_d15_28),.data_out(wire_d15_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1601530(.data_in(wire_d15_29),.data_out(wire_d15_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1601531(.data_in(wire_d15_30),.data_out(wire_d15_31),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1601532(.data_in(wire_d15_31),.data_out(wire_d15_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1601533(.data_in(wire_d15_32),.data_out(wire_d15_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1601534(.data_in(wire_d15_33),.data_out(wire_d15_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1601535(.data_in(wire_d15_34),.data_out(wire_d15_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1601536(.data_in(wire_d15_35),.data_out(wire_d15_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1601537(.data_in(wire_d15_36),.data_out(wire_d15_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601538(.data_in(wire_d15_37),.data_out(wire_d15_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601539(.data_in(wire_d15_38),.data_out(wire_d15_39),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1601540(.data_in(wire_d15_39),.data_out(wire_d15_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601541(.data_in(wire_d15_40),.data_out(wire_d15_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601542(.data_in(wire_d15_41),.data_out(wire_d15_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1601543(.data_in(wire_d15_42),.data_out(wire_d15_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1601544(.data_in(wire_d15_43),.data_out(wire_d15_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1601545(.data_in(wire_d15_44),.data_out(wire_d15_45),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1601546(.data_in(wire_d15_45),.data_out(wire_d15_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1601547(.data_in(wire_d15_46),.data_out(wire_d15_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1601548(.data_in(wire_d15_47),.data_out(wire_d15_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1601549(.data_in(wire_d15_48),.data_out(d_out15),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance170160(.data_in(d_in16),.data_out(wire_d16_0),.clk(clk),.rst(rst));            //channel 17
	large_mux #(.WIDTH(WIDTH)) large_mux_instance170161(.data_in(wire_d16_0),.data_out(wire_d16_1),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance170162(.data_in(wire_d16_1),.data_out(wire_d16_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance170163(.data_in(wire_d16_2),.data_out(wire_d16_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance170164(.data_in(wire_d16_3),.data_out(wire_d16_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance170165(.data_in(wire_d16_4),.data_out(wire_d16_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance170166(.data_in(wire_d16_5),.data_out(wire_d16_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance170167(.data_in(wire_d16_6),.data_out(wire_d16_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance170168(.data_in(wire_d16_7),.data_out(wire_d16_8),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance170169(.data_in(wire_d16_8),.data_out(wire_d16_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701610(.data_in(wire_d16_9),.data_out(wire_d16_10),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1701611(.data_in(wire_d16_10),.data_out(wire_d16_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701612(.data_in(wire_d16_11),.data_out(wire_d16_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701613(.data_in(wire_d16_12),.data_out(wire_d16_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701614(.data_in(wire_d16_13),.data_out(wire_d16_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701615(.data_in(wire_d16_14),.data_out(wire_d16_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701616(.data_in(wire_d16_15),.data_out(wire_d16_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701617(.data_in(wire_d16_16),.data_out(wire_d16_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1701618(.data_in(wire_d16_17),.data_out(wire_d16_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1701619(.data_in(wire_d16_18),.data_out(wire_d16_19),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701620(.data_in(wire_d16_19),.data_out(wire_d16_20),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701621(.data_in(wire_d16_20),.data_out(wire_d16_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701622(.data_in(wire_d16_21),.data_out(wire_d16_22),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701623(.data_in(wire_d16_22),.data_out(wire_d16_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701624(.data_in(wire_d16_23),.data_out(wire_d16_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701625(.data_in(wire_d16_24),.data_out(wire_d16_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1701626(.data_in(wire_d16_25),.data_out(wire_d16_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1701627(.data_in(wire_d16_26),.data_out(wire_d16_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1701628(.data_in(wire_d16_27),.data_out(wire_d16_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701629(.data_in(wire_d16_28),.data_out(wire_d16_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1701630(.data_in(wire_d16_29),.data_out(wire_d16_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1701631(.data_in(wire_d16_30),.data_out(wire_d16_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701632(.data_in(wire_d16_31),.data_out(wire_d16_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701633(.data_in(wire_d16_32),.data_out(wire_d16_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1701634(.data_in(wire_d16_33),.data_out(wire_d16_34),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1701635(.data_in(wire_d16_34),.data_out(wire_d16_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1701636(.data_in(wire_d16_35),.data_out(wire_d16_36),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1701637(.data_in(wire_d16_36),.data_out(wire_d16_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1701638(.data_in(wire_d16_37),.data_out(wire_d16_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1701639(.data_in(wire_d16_38),.data_out(wire_d16_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1701640(.data_in(wire_d16_39),.data_out(wire_d16_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701641(.data_in(wire_d16_40),.data_out(wire_d16_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1701642(.data_in(wire_d16_41),.data_out(wire_d16_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1701643(.data_in(wire_d16_42),.data_out(wire_d16_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701644(.data_in(wire_d16_43),.data_out(wire_d16_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1701645(.data_in(wire_d16_44),.data_out(wire_d16_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1701646(.data_in(wire_d16_45),.data_out(wire_d16_46),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1701647(.data_in(wire_d16_46),.data_out(wire_d16_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1701648(.data_in(wire_d16_47),.data_out(wire_d16_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1701649(.data_in(wire_d16_48),.data_out(d_out16),.clk(clk),.rst(rst));

	large_adder #(.WIDTH(WIDTH)) large_adder_instance180170(.data_in(d_in17),.data_out(wire_d17_0),.clk(clk),.rst(rst));            //channel 18
	large_mux #(.WIDTH(WIDTH)) large_mux_instance180171(.data_in(wire_d17_0),.data_out(wire_d17_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance180172(.data_in(wire_d17_1),.data_out(wire_d17_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance180173(.data_in(wire_d17_2),.data_out(wire_d17_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance180174(.data_in(wire_d17_3),.data_out(wire_d17_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance180175(.data_in(wire_d17_4),.data_out(wire_d17_5),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance180176(.data_in(wire_d17_5),.data_out(wire_d17_6),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance180177(.data_in(wire_d17_6),.data_out(wire_d17_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance180178(.data_in(wire_d17_7),.data_out(wire_d17_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance180179(.data_in(wire_d17_8),.data_out(wire_d17_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801710(.data_in(wire_d17_9),.data_out(wire_d17_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1801711(.data_in(wire_d17_10),.data_out(wire_d17_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801712(.data_in(wire_d17_11),.data_out(wire_d17_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1801713(.data_in(wire_d17_12),.data_out(wire_d17_13),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801714(.data_in(wire_d17_13),.data_out(wire_d17_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801715(.data_in(wire_d17_14),.data_out(wire_d17_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801716(.data_in(wire_d17_15),.data_out(wire_d17_16),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1801717(.data_in(wire_d17_16),.data_out(wire_d17_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1801718(.data_in(wire_d17_17),.data_out(wire_d17_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1801719(.data_in(wire_d17_18),.data_out(wire_d17_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801720(.data_in(wire_d17_19),.data_out(wire_d17_20),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801721(.data_in(wire_d17_20),.data_out(wire_d17_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801722(.data_in(wire_d17_21),.data_out(wire_d17_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1801723(.data_in(wire_d17_22),.data_out(wire_d17_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1801724(.data_in(wire_d17_23),.data_out(wire_d17_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801725(.data_in(wire_d17_24),.data_out(wire_d17_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801726(.data_in(wire_d17_25),.data_out(wire_d17_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1801727(.data_in(wire_d17_26),.data_out(wire_d17_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801728(.data_in(wire_d17_27),.data_out(wire_d17_28),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1801729(.data_in(wire_d17_28),.data_out(wire_d17_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801730(.data_in(wire_d17_29),.data_out(wire_d17_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1801731(.data_in(wire_d17_30),.data_out(wire_d17_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801732(.data_in(wire_d17_31),.data_out(wire_d17_32),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801733(.data_in(wire_d17_32),.data_out(wire_d17_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801734(.data_in(wire_d17_33),.data_out(wire_d17_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1801735(.data_in(wire_d17_34),.data_out(wire_d17_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801736(.data_in(wire_d17_35),.data_out(wire_d17_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801737(.data_in(wire_d17_36),.data_out(wire_d17_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1801738(.data_in(wire_d17_37),.data_out(wire_d17_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1801739(.data_in(wire_d17_38),.data_out(wire_d17_39),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801740(.data_in(wire_d17_39),.data_out(wire_d17_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1801741(.data_in(wire_d17_40),.data_out(wire_d17_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1801742(.data_in(wire_d17_41),.data_out(wire_d17_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801743(.data_in(wire_d17_42),.data_out(wire_d17_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1801744(.data_in(wire_d17_43),.data_out(wire_d17_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1801745(.data_in(wire_d17_44),.data_out(wire_d17_45),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1801746(.data_in(wire_d17_45),.data_out(wire_d17_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1801747(.data_in(wire_d17_46),.data_out(wire_d17_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1801748(.data_in(wire_d17_47),.data_out(wire_d17_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1801749(.data_in(wire_d17_48),.data_out(d_out17),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance190180(.data_in(d_in18),.data_out(wire_d18_0),.clk(clk),.rst(rst));            //channel 19
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance190181(.data_in(wire_d18_0),.data_out(wire_d18_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance190182(.data_in(wire_d18_1),.data_out(wire_d18_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance190183(.data_in(wire_d18_2),.data_out(wire_d18_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance190184(.data_in(wire_d18_3),.data_out(wire_d18_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance190185(.data_in(wire_d18_4),.data_out(wire_d18_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance190186(.data_in(wire_d18_5),.data_out(wire_d18_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance190187(.data_in(wire_d18_6),.data_out(wire_d18_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance190188(.data_in(wire_d18_7),.data_out(wire_d18_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance190189(.data_in(wire_d18_8),.data_out(wire_d18_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1901810(.data_in(wire_d18_9),.data_out(wire_d18_10),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901811(.data_in(wire_d18_10),.data_out(wire_d18_11),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1901812(.data_in(wire_d18_11),.data_out(wire_d18_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1901813(.data_in(wire_d18_12),.data_out(wire_d18_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1901814(.data_in(wire_d18_13),.data_out(wire_d18_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901815(.data_in(wire_d18_14),.data_out(wire_d18_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901816(.data_in(wire_d18_15),.data_out(wire_d18_16),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1901817(.data_in(wire_d18_16),.data_out(wire_d18_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901818(.data_in(wire_d18_17),.data_out(wire_d18_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901819(.data_in(wire_d18_18),.data_out(wire_d18_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901820(.data_in(wire_d18_19),.data_out(wire_d18_20),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1901821(.data_in(wire_d18_20),.data_out(wire_d18_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901822(.data_in(wire_d18_21),.data_out(wire_d18_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901823(.data_in(wire_d18_22),.data_out(wire_d18_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901824(.data_in(wire_d18_23),.data_out(wire_d18_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901825(.data_in(wire_d18_24),.data_out(wire_d18_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance1901826(.data_in(wire_d18_25),.data_out(wire_d18_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901827(.data_in(wire_d18_26),.data_out(wire_d18_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901828(.data_in(wire_d18_27),.data_out(wire_d18_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1901829(.data_in(wire_d18_28),.data_out(wire_d18_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance1901830(.data_in(wire_d18_29),.data_out(wire_d18_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901831(.data_in(wire_d18_30),.data_out(wire_d18_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance1901832(.data_in(wire_d18_31),.data_out(wire_d18_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901833(.data_in(wire_d18_32),.data_out(wire_d18_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901834(.data_in(wire_d18_33),.data_out(wire_d18_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901835(.data_in(wire_d18_34),.data_out(wire_d18_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance1901836(.data_in(wire_d18_35),.data_out(wire_d18_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1901837(.data_in(wire_d18_36),.data_out(wire_d18_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance1901838(.data_in(wire_d18_37),.data_out(wire_d18_38),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901839(.data_in(wire_d18_38),.data_out(wire_d18_39),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1901840(.data_in(wire_d18_39),.data_out(wire_d18_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance1901841(.data_in(wire_d18_40),.data_out(wire_d18_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901842(.data_in(wire_d18_41),.data_out(wire_d18_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1901843(.data_in(wire_d18_42),.data_out(wire_d18_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance1901844(.data_in(wire_d18_43),.data_out(wire_d18_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance1901845(.data_in(wire_d18_44),.data_out(wire_d18_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance1901846(.data_in(wire_d18_45),.data_out(wire_d18_46),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance1901847(.data_in(wire_d18_46),.data_out(wire_d18_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance1901848(.data_in(wire_d18_47),.data_out(wire_d18_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance1901849(.data_in(wire_d18_48),.data_out(d_out18),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance200190(.data_in(d_in19),.data_out(wire_d19_0),.clk(clk),.rst(rst));            //channel 20
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance200191(.data_in(wire_d19_0),.data_out(wire_d19_1),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance200192(.data_in(wire_d19_1),.data_out(wire_d19_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance200193(.data_in(wire_d19_2),.data_out(wire_d19_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance200194(.data_in(wire_d19_3),.data_out(wire_d19_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance200195(.data_in(wire_d19_4),.data_out(wire_d19_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance200196(.data_in(wire_d19_5),.data_out(wire_d19_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance200197(.data_in(wire_d19_6),.data_out(wire_d19_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance200198(.data_in(wire_d19_7),.data_out(wire_d19_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance200199(.data_in(wire_d19_8),.data_out(wire_d19_9),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001910(.data_in(wire_d19_9),.data_out(wire_d19_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2001911(.data_in(wire_d19_10),.data_out(wire_d19_11),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2001912(.data_in(wire_d19_11),.data_out(wire_d19_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2001913(.data_in(wire_d19_12),.data_out(wire_d19_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001914(.data_in(wire_d19_13),.data_out(wire_d19_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001915(.data_in(wire_d19_14),.data_out(wire_d19_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001916(.data_in(wire_d19_15),.data_out(wire_d19_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2001917(.data_in(wire_d19_16),.data_out(wire_d19_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2001918(.data_in(wire_d19_17),.data_out(wire_d19_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001919(.data_in(wire_d19_18),.data_out(wire_d19_19),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2001920(.data_in(wire_d19_19),.data_out(wire_d19_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2001921(.data_in(wire_d19_20),.data_out(wire_d19_21),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001922(.data_in(wire_d19_21),.data_out(wire_d19_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2001923(.data_in(wire_d19_22),.data_out(wire_d19_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2001924(.data_in(wire_d19_23),.data_out(wire_d19_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001925(.data_in(wire_d19_24),.data_out(wire_d19_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001926(.data_in(wire_d19_25),.data_out(wire_d19_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2001927(.data_in(wire_d19_26),.data_out(wire_d19_27),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2001928(.data_in(wire_d19_27),.data_out(wire_d19_28),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2001929(.data_in(wire_d19_28),.data_out(wire_d19_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001930(.data_in(wire_d19_29),.data_out(wire_d19_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2001931(.data_in(wire_d19_30),.data_out(wire_d19_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2001932(.data_in(wire_d19_31),.data_out(wire_d19_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2001933(.data_in(wire_d19_32),.data_out(wire_d19_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2001934(.data_in(wire_d19_33),.data_out(wire_d19_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2001935(.data_in(wire_d19_34),.data_out(wire_d19_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2001936(.data_in(wire_d19_35),.data_out(wire_d19_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001937(.data_in(wire_d19_36),.data_out(wire_d19_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2001938(.data_in(wire_d19_37),.data_out(wire_d19_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001939(.data_in(wire_d19_38),.data_out(wire_d19_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001940(.data_in(wire_d19_39),.data_out(wire_d19_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2001941(.data_in(wire_d19_40),.data_out(wire_d19_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2001942(.data_in(wire_d19_41),.data_out(wire_d19_42),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2001943(.data_in(wire_d19_42),.data_out(wire_d19_43),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2001944(.data_in(wire_d19_43),.data_out(wire_d19_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2001945(.data_in(wire_d19_44),.data_out(wire_d19_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2001946(.data_in(wire_d19_45),.data_out(wire_d19_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2001947(.data_in(wire_d19_46),.data_out(wire_d19_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2001948(.data_in(wire_d19_47),.data_out(wire_d19_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2001949(.data_in(wire_d19_48),.data_out(d_out19),.clk(clk),.rst(rst));

	large_adder #(.WIDTH(WIDTH)) large_adder_instance210200(.data_in(d_in20),.data_out(wire_d20_0),.clk(clk),.rst(rst));            //channel 21
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance210201(.data_in(wire_d20_0),.data_out(wire_d20_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance210202(.data_in(wire_d20_1),.data_out(wire_d20_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance210203(.data_in(wire_d20_2),.data_out(wire_d20_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance210204(.data_in(wire_d20_3),.data_out(wire_d20_4),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance210205(.data_in(wire_d20_4),.data_out(wire_d20_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance210206(.data_in(wire_d20_5),.data_out(wire_d20_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance210207(.data_in(wire_d20_6),.data_out(wire_d20_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance210208(.data_in(wire_d20_7),.data_out(wire_d20_8),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance210209(.data_in(wire_d20_8),.data_out(wire_d20_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102010(.data_in(wire_d20_9),.data_out(wire_d20_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2102011(.data_in(wire_d20_10),.data_out(wire_d20_11),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2102012(.data_in(wire_d20_11),.data_out(wire_d20_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102013(.data_in(wire_d20_12),.data_out(wire_d20_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2102014(.data_in(wire_d20_13),.data_out(wire_d20_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2102015(.data_in(wire_d20_14),.data_out(wire_d20_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102016(.data_in(wire_d20_15),.data_out(wire_d20_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102017(.data_in(wire_d20_16),.data_out(wire_d20_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102018(.data_in(wire_d20_17),.data_out(wire_d20_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2102019(.data_in(wire_d20_18),.data_out(wire_d20_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102020(.data_in(wire_d20_19),.data_out(wire_d20_20),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2102021(.data_in(wire_d20_20),.data_out(wire_d20_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2102022(.data_in(wire_d20_21),.data_out(wire_d20_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102023(.data_in(wire_d20_22),.data_out(wire_d20_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102024(.data_in(wire_d20_23),.data_out(wire_d20_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102025(.data_in(wire_d20_24),.data_out(wire_d20_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102026(.data_in(wire_d20_25),.data_out(wire_d20_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102027(.data_in(wire_d20_26),.data_out(wire_d20_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102028(.data_in(wire_d20_27),.data_out(wire_d20_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2102029(.data_in(wire_d20_28),.data_out(wire_d20_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2102030(.data_in(wire_d20_29),.data_out(wire_d20_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102031(.data_in(wire_d20_30),.data_out(wire_d20_31),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102032(.data_in(wire_d20_31),.data_out(wire_d20_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2102033(.data_in(wire_d20_32),.data_out(wire_d20_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102034(.data_in(wire_d20_33),.data_out(wire_d20_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102035(.data_in(wire_d20_34),.data_out(wire_d20_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102036(.data_in(wire_d20_35),.data_out(wire_d20_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2102037(.data_in(wire_d20_36),.data_out(wire_d20_37),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102038(.data_in(wire_d20_37),.data_out(wire_d20_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102039(.data_in(wire_d20_38),.data_out(wire_d20_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2102040(.data_in(wire_d20_39),.data_out(wire_d20_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2102041(.data_in(wire_d20_40),.data_out(wire_d20_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2102042(.data_in(wire_d20_41),.data_out(wire_d20_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2102043(.data_in(wire_d20_42),.data_out(wire_d20_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2102044(.data_in(wire_d20_43),.data_out(wire_d20_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2102045(.data_in(wire_d20_44),.data_out(wire_d20_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102046(.data_in(wire_d20_45),.data_out(wire_d20_46),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2102047(.data_in(wire_d20_46),.data_out(wire_d20_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2102048(.data_in(wire_d20_47),.data_out(wire_d20_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2102049(.data_in(wire_d20_48),.data_out(d_out20),.clk(clk),.rst(rst));

	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance220210(.data_in(d_in21),.data_out(wire_d21_0),.clk(clk),.rst(rst));            //channel 22
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance220211(.data_in(wire_d21_0),.data_out(wire_d21_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance220212(.data_in(wire_d21_1),.data_out(wire_d21_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance220213(.data_in(wire_d21_2),.data_out(wire_d21_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance220214(.data_in(wire_d21_3),.data_out(wire_d21_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance220215(.data_in(wire_d21_4),.data_out(wire_d21_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance220216(.data_in(wire_d21_5),.data_out(wire_d21_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance220217(.data_in(wire_d21_6),.data_out(wire_d21_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance220218(.data_in(wire_d21_7),.data_out(wire_d21_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance220219(.data_in(wire_d21_8),.data_out(wire_d21_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2202110(.data_in(wire_d21_9),.data_out(wire_d21_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2202111(.data_in(wire_d21_10),.data_out(wire_d21_11),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2202112(.data_in(wire_d21_11),.data_out(wire_d21_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2202113(.data_in(wire_d21_12),.data_out(wire_d21_13),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202114(.data_in(wire_d21_13),.data_out(wire_d21_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2202115(.data_in(wire_d21_14),.data_out(wire_d21_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202116(.data_in(wire_d21_15),.data_out(wire_d21_16),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202117(.data_in(wire_d21_16),.data_out(wire_d21_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202118(.data_in(wire_d21_17),.data_out(wire_d21_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2202119(.data_in(wire_d21_18),.data_out(wire_d21_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202120(.data_in(wire_d21_19),.data_out(wire_d21_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202121(.data_in(wire_d21_20),.data_out(wire_d21_21),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2202122(.data_in(wire_d21_21),.data_out(wire_d21_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202123(.data_in(wire_d21_22),.data_out(wire_d21_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202124(.data_in(wire_d21_23),.data_out(wire_d21_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202125(.data_in(wire_d21_24),.data_out(wire_d21_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202126(.data_in(wire_d21_25),.data_out(wire_d21_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202127(.data_in(wire_d21_26),.data_out(wire_d21_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2202128(.data_in(wire_d21_27),.data_out(wire_d21_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2202129(.data_in(wire_d21_28),.data_out(wire_d21_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202130(.data_in(wire_d21_29),.data_out(wire_d21_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202131(.data_in(wire_d21_30),.data_out(wire_d21_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202132(.data_in(wire_d21_31),.data_out(wire_d21_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2202133(.data_in(wire_d21_32),.data_out(wire_d21_33),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202134(.data_in(wire_d21_33),.data_out(wire_d21_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2202135(.data_in(wire_d21_34),.data_out(wire_d21_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2202136(.data_in(wire_d21_35),.data_out(wire_d21_36),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2202137(.data_in(wire_d21_36),.data_out(wire_d21_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2202138(.data_in(wire_d21_37),.data_out(wire_d21_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2202139(.data_in(wire_d21_38),.data_out(wire_d21_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202140(.data_in(wire_d21_39),.data_out(wire_d21_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2202141(.data_in(wire_d21_40),.data_out(wire_d21_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2202142(.data_in(wire_d21_41),.data_out(wire_d21_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2202143(.data_in(wire_d21_42),.data_out(wire_d21_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2202144(.data_in(wire_d21_43),.data_out(wire_d21_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2202145(.data_in(wire_d21_44),.data_out(wire_d21_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2202146(.data_in(wire_d21_45),.data_out(wire_d21_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2202147(.data_in(wire_d21_46),.data_out(wire_d21_47),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2202148(.data_in(wire_d21_47),.data_out(wire_d21_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2202149(.data_in(wire_d21_48),.data_out(d_out21),.clk(clk),.rst(rst));

	large_adder #(.WIDTH(WIDTH)) large_adder_instance230220(.data_in(d_in22),.data_out(wire_d22_0),.clk(clk),.rst(rst));            //channel 23
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance230221(.data_in(wire_d22_0),.data_out(wire_d22_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance230222(.data_in(wire_d22_1),.data_out(wire_d22_2),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance230223(.data_in(wire_d22_2),.data_out(wire_d22_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance230224(.data_in(wire_d22_3),.data_out(wire_d22_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance230225(.data_in(wire_d22_4),.data_out(wire_d22_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance230226(.data_in(wire_d22_5),.data_out(wire_d22_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance230227(.data_in(wire_d22_6),.data_out(wire_d22_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance230228(.data_in(wire_d22_7),.data_out(wire_d22_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance230229(.data_in(wire_d22_8),.data_out(wire_d22_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302210(.data_in(wire_d22_9),.data_out(wire_d22_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302211(.data_in(wire_d22_10),.data_out(wire_d22_11),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2302212(.data_in(wire_d22_11),.data_out(wire_d22_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302213(.data_in(wire_d22_12),.data_out(wire_d22_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302214(.data_in(wire_d22_13),.data_out(wire_d22_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302215(.data_in(wire_d22_14),.data_out(wire_d22_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302216(.data_in(wire_d22_15),.data_out(wire_d22_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302217(.data_in(wire_d22_16),.data_out(wire_d22_17),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2302218(.data_in(wire_d22_17),.data_out(wire_d22_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302219(.data_in(wire_d22_18),.data_out(wire_d22_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302220(.data_in(wire_d22_19),.data_out(wire_d22_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302221(.data_in(wire_d22_20),.data_out(wire_d22_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2302222(.data_in(wire_d22_21),.data_out(wire_d22_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2302223(.data_in(wire_d22_22),.data_out(wire_d22_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2302224(.data_in(wire_d22_23),.data_out(wire_d22_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302225(.data_in(wire_d22_24),.data_out(wire_d22_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302226(.data_in(wire_d22_25),.data_out(wire_d22_26),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2302227(.data_in(wire_d22_26),.data_out(wire_d22_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2302228(.data_in(wire_d22_27),.data_out(wire_d22_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2302229(.data_in(wire_d22_28),.data_out(wire_d22_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302230(.data_in(wire_d22_29),.data_out(wire_d22_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2302231(.data_in(wire_d22_30),.data_out(wire_d22_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302232(.data_in(wire_d22_31),.data_out(wire_d22_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302233(.data_in(wire_d22_32),.data_out(wire_d22_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302234(.data_in(wire_d22_33),.data_out(wire_d22_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2302235(.data_in(wire_d22_34),.data_out(wire_d22_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302236(.data_in(wire_d22_35),.data_out(wire_d22_36),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302237(.data_in(wire_d22_36),.data_out(wire_d22_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2302238(.data_in(wire_d22_37),.data_out(wire_d22_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2302239(.data_in(wire_d22_38),.data_out(wire_d22_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2302240(.data_in(wire_d22_39),.data_out(wire_d22_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2302241(.data_in(wire_d22_40),.data_out(wire_d22_41),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2302242(.data_in(wire_d22_41),.data_out(wire_d22_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2302243(.data_in(wire_d22_42),.data_out(wire_d22_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2302244(.data_in(wire_d22_43),.data_out(wire_d22_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302245(.data_in(wire_d22_44),.data_out(wire_d22_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302246(.data_in(wire_d22_45),.data_out(wire_d22_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2302247(.data_in(wire_d22_46),.data_out(wire_d22_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2302248(.data_in(wire_d22_47),.data_out(wire_d22_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2302249(.data_in(wire_d22_48),.data_out(d_out22),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance240230(.data_in(d_in23),.data_out(wire_d23_0),.clk(clk),.rst(rst));            //channel 24
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance240231(.data_in(wire_d23_0),.data_out(wire_d23_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance240232(.data_in(wire_d23_1),.data_out(wire_d23_2),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance240233(.data_in(wire_d23_2),.data_out(wire_d23_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance240234(.data_in(wire_d23_3),.data_out(wire_d23_4),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance240235(.data_in(wire_d23_4),.data_out(wire_d23_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance240236(.data_in(wire_d23_5),.data_out(wire_d23_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance240237(.data_in(wire_d23_6),.data_out(wire_d23_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance240238(.data_in(wire_d23_7),.data_out(wire_d23_8),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance240239(.data_in(wire_d23_8),.data_out(wire_d23_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402310(.data_in(wire_d23_9),.data_out(wire_d23_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402311(.data_in(wire_d23_10),.data_out(wire_d23_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402312(.data_in(wire_d23_11),.data_out(wire_d23_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402313(.data_in(wire_d23_12),.data_out(wire_d23_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402314(.data_in(wire_d23_13),.data_out(wire_d23_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2402315(.data_in(wire_d23_14),.data_out(wire_d23_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2402316(.data_in(wire_d23_15),.data_out(wire_d23_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2402317(.data_in(wire_d23_16),.data_out(wire_d23_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2402318(.data_in(wire_d23_17),.data_out(wire_d23_18),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2402319(.data_in(wire_d23_18),.data_out(wire_d23_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402320(.data_in(wire_d23_19),.data_out(wire_d23_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402321(.data_in(wire_d23_20),.data_out(wire_d23_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2402322(.data_in(wire_d23_21),.data_out(wire_d23_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402323(.data_in(wire_d23_22),.data_out(wire_d23_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402324(.data_in(wire_d23_23),.data_out(wire_d23_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2402325(.data_in(wire_d23_24),.data_out(wire_d23_25),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2402326(.data_in(wire_d23_25),.data_out(wire_d23_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402327(.data_in(wire_d23_26),.data_out(wire_d23_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402328(.data_in(wire_d23_27),.data_out(wire_d23_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402329(.data_in(wire_d23_28),.data_out(wire_d23_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2402330(.data_in(wire_d23_29),.data_out(wire_d23_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2402331(.data_in(wire_d23_30),.data_out(wire_d23_31),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2402332(.data_in(wire_d23_31),.data_out(wire_d23_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2402333(.data_in(wire_d23_32),.data_out(wire_d23_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2402334(.data_in(wire_d23_33),.data_out(wire_d23_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2402335(.data_in(wire_d23_34),.data_out(wire_d23_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402336(.data_in(wire_d23_35),.data_out(wire_d23_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402337(.data_in(wire_d23_36),.data_out(wire_d23_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402338(.data_in(wire_d23_37),.data_out(wire_d23_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2402339(.data_in(wire_d23_38),.data_out(wire_d23_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402340(.data_in(wire_d23_39),.data_out(wire_d23_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2402341(.data_in(wire_d23_40),.data_out(wire_d23_41),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2402342(.data_in(wire_d23_41),.data_out(wire_d23_42),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402343(.data_in(wire_d23_42),.data_out(wire_d23_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2402344(.data_in(wire_d23_43),.data_out(wire_d23_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2402345(.data_in(wire_d23_44),.data_out(wire_d23_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2402346(.data_in(wire_d23_45),.data_out(wire_d23_46),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2402347(.data_in(wire_d23_46),.data_out(wire_d23_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2402348(.data_in(wire_d23_47),.data_out(wire_d23_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2402349(.data_in(wire_d23_48),.data_out(d_out23),.clk(clk),.rst(rst));

	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance250240(.data_in(d_in24),.data_out(wire_d24_0),.clk(clk),.rst(rst));            //channel 25
	decoder_top #(.WIDTH(WIDTH)) decoder_instance250241(.data_in(wire_d24_0),.data_out(wire_d24_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance250242(.data_in(wire_d24_1),.data_out(wire_d24_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance250243(.data_in(wire_d24_2),.data_out(wire_d24_3),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance250244(.data_in(wire_d24_3),.data_out(wire_d24_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance250245(.data_in(wire_d24_4),.data_out(wire_d24_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance250246(.data_in(wire_d24_5),.data_out(wire_d24_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance250247(.data_in(wire_d24_6),.data_out(wire_d24_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance250248(.data_in(wire_d24_7),.data_out(wire_d24_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance250249(.data_in(wire_d24_8),.data_out(wire_d24_9),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2502410(.data_in(wire_d24_9),.data_out(wire_d24_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2502411(.data_in(wire_d24_10),.data_out(wire_d24_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502412(.data_in(wire_d24_11),.data_out(wire_d24_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502413(.data_in(wire_d24_12),.data_out(wire_d24_13),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502414(.data_in(wire_d24_13),.data_out(wire_d24_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2502415(.data_in(wire_d24_14),.data_out(wire_d24_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2502416(.data_in(wire_d24_15),.data_out(wire_d24_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2502417(.data_in(wire_d24_16),.data_out(wire_d24_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502418(.data_in(wire_d24_17),.data_out(wire_d24_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502419(.data_in(wire_d24_18),.data_out(wire_d24_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2502420(.data_in(wire_d24_19),.data_out(wire_d24_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2502421(.data_in(wire_d24_20),.data_out(wire_d24_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502422(.data_in(wire_d24_21),.data_out(wire_d24_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502423(.data_in(wire_d24_22),.data_out(wire_d24_23),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2502424(.data_in(wire_d24_23),.data_out(wire_d24_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502425(.data_in(wire_d24_24),.data_out(wire_d24_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2502426(.data_in(wire_d24_25),.data_out(wire_d24_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502427(.data_in(wire_d24_26),.data_out(wire_d24_27),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502428(.data_in(wire_d24_27),.data_out(wire_d24_28),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502429(.data_in(wire_d24_28),.data_out(wire_d24_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2502430(.data_in(wire_d24_29),.data_out(wire_d24_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2502431(.data_in(wire_d24_30),.data_out(wire_d24_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502432(.data_in(wire_d24_31),.data_out(wire_d24_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2502433(.data_in(wire_d24_32),.data_out(wire_d24_33),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502434(.data_in(wire_d24_33),.data_out(wire_d24_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2502435(.data_in(wire_d24_34),.data_out(wire_d24_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502436(.data_in(wire_d24_35),.data_out(wire_d24_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2502437(.data_in(wire_d24_36),.data_out(wire_d24_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2502438(.data_in(wire_d24_37),.data_out(wire_d24_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502439(.data_in(wire_d24_38),.data_out(wire_d24_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2502440(.data_in(wire_d24_39),.data_out(wire_d24_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502441(.data_in(wire_d24_40),.data_out(wire_d24_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2502442(.data_in(wire_d24_41),.data_out(wire_d24_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2502443(.data_in(wire_d24_42),.data_out(wire_d24_43),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2502444(.data_in(wire_d24_43),.data_out(wire_d24_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2502445(.data_in(wire_d24_44),.data_out(wire_d24_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2502446(.data_in(wire_d24_45),.data_out(wire_d24_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2502447(.data_in(wire_d24_46),.data_out(wire_d24_47),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2502448(.data_in(wire_d24_47),.data_out(wire_d24_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2502449(.data_in(wire_d24_48),.data_out(d_out24),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance260250(.data_in(d_in25),.data_out(wire_d25_0),.clk(clk),.rst(rst));            //channel 26
	encoder #(.WIDTH(WIDTH)) encoder_instance260251(.data_in(wire_d25_0),.data_out(wire_d25_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance260252(.data_in(wire_d25_1),.data_out(wire_d25_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance260253(.data_in(wire_d25_2),.data_out(wire_d25_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance260254(.data_in(wire_d25_3),.data_out(wire_d25_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance260255(.data_in(wire_d25_4),.data_out(wire_d25_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance260256(.data_in(wire_d25_5),.data_out(wire_d25_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance260257(.data_in(wire_d25_6),.data_out(wire_d25_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance260258(.data_in(wire_d25_7),.data_out(wire_d25_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance260259(.data_in(wire_d25_8),.data_out(wire_d25_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602510(.data_in(wire_d25_9),.data_out(wire_d25_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602511(.data_in(wire_d25_10),.data_out(wire_d25_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2602512(.data_in(wire_d25_11),.data_out(wire_d25_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2602513(.data_in(wire_d25_12),.data_out(wire_d25_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602514(.data_in(wire_d25_13),.data_out(wire_d25_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602515(.data_in(wire_d25_14),.data_out(wire_d25_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2602516(.data_in(wire_d25_15),.data_out(wire_d25_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602517(.data_in(wire_d25_16),.data_out(wire_d25_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602518(.data_in(wire_d25_17),.data_out(wire_d25_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602519(.data_in(wire_d25_18),.data_out(wire_d25_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2602520(.data_in(wire_d25_19),.data_out(wire_d25_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602521(.data_in(wire_d25_20),.data_out(wire_d25_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602522(.data_in(wire_d25_21),.data_out(wire_d25_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602523(.data_in(wire_d25_22),.data_out(wire_d25_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602524(.data_in(wire_d25_23),.data_out(wire_d25_24),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2602525(.data_in(wire_d25_24),.data_out(wire_d25_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602526(.data_in(wire_d25_25),.data_out(wire_d25_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2602527(.data_in(wire_d25_26),.data_out(wire_d25_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602528(.data_in(wire_d25_27),.data_out(wire_d25_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602529(.data_in(wire_d25_28),.data_out(wire_d25_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2602530(.data_in(wire_d25_29),.data_out(wire_d25_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602531(.data_in(wire_d25_30),.data_out(wire_d25_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602532(.data_in(wire_d25_31),.data_out(wire_d25_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2602533(.data_in(wire_d25_32),.data_out(wire_d25_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2602534(.data_in(wire_d25_33),.data_out(wire_d25_34),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2602535(.data_in(wire_d25_34),.data_out(wire_d25_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2602536(.data_in(wire_d25_35),.data_out(wire_d25_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602537(.data_in(wire_d25_36),.data_out(wire_d25_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2602538(.data_in(wire_d25_37),.data_out(wire_d25_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602539(.data_in(wire_d25_38),.data_out(wire_d25_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2602540(.data_in(wire_d25_39),.data_out(wire_d25_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602541(.data_in(wire_d25_40),.data_out(wire_d25_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602542(.data_in(wire_d25_41),.data_out(wire_d25_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2602543(.data_in(wire_d25_42),.data_out(wire_d25_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2602544(.data_in(wire_d25_43),.data_out(wire_d25_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2602545(.data_in(wire_d25_44),.data_out(wire_d25_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2602546(.data_in(wire_d25_45),.data_out(wire_d25_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2602547(.data_in(wire_d25_46),.data_out(wire_d25_47),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2602548(.data_in(wire_d25_47),.data_out(wire_d25_48),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2602549(.data_in(wire_d25_48),.data_out(d_out25),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance270260(.data_in(d_in26),.data_out(wire_d26_0),.clk(clk),.rst(rst));            //channel 27
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance270261(.data_in(wire_d26_0),.data_out(wire_d26_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance270262(.data_in(wire_d26_1),.data_out(wire_d26_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance270263(.data_in(wire_d26_2),.data_out(wire_d26_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance270264(.data_in(wire_d26_3),.data_out(wire_d26_4),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance270265(.data_in(wire_d26_4),.data_out(wire_d26_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance270266(.data_in(wire_d26_5),.data_out(wire_d26_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance270267(.data_in(wire_d26_6),.data_out(wire_d26_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance270268(.data_in(wire_d26_7),.data_out(wire_d26_8),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance270269(.data_in(wire_d26_8),.data_out(wire_d26_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702610(.data_in(wire_d26_9),.data_out(wire_d26_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2702611(.data_in(wire_d26_10),.data_out(wire_d26_11),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2702612(.data_in(wire_d26_11),.data_out(wire_d26_12),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2702613(.data_in(wire_d26_12),.data_out(wire_d26_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702614(.data_in(wire_d26_13),.data_out(wire_d26_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702615(.data_in(wire_d26_14),.data_out(wire_d26_15),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702616(.data_in(wire_d26_15),.data_out(wire_d26_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702617(.data_in(wire_d26_16),.data_out(wire_d26_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702618(.data_in(wire_d26_17),.data_out(wire_d26_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2702619(.data_in(wire_d26_18),.data_out(wire_d26_19),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702620(.data_in(wire_d26_19),.data_out(wire_d26_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702621(.data_in(wire_d26_20),.data_out(wire_d26_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2702622(.data_in(wire_d26_21),.data_out(wire_d26_22),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702623(.data_in(wire_d26_22),.data_out(wire_d26_23),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2702624(.data_in(wire_d26_23),.data_out(wire_d26_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702625(.data_in(wire_d26_24),.data_out(wire_d26_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2702626(.data_in(wire_d26_25),.data_out(wire_d26_26),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2702627(.data_in(wire_d26_26),.data_out(wire_d26_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2702628(.data_in(wire_d26_27),.data_out(wire_d26_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2702629(.data_in(wire_d26_28),.data_out(wire_d26_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2702630(.data_in(wire_d26_29),.data_out(wire_d26_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702631(.data_in(wire_d26_30),.data_out(wire_d26_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2702632(.data_in(wire_d26_31),.data_out(wire_d26_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2702633(.data_in(wire_d26_32),.data_out(wire_d26_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702634(.data_in(wire_d26_33),.data_out(wire_d26_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702635(.data_in(wire_d26_34),.data_out(wire_d26_35),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702636(.data_in(wire_d26_35),.data_out(wire_d26_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2702637(.data_in(wire_d26_36),.data_out(wire_d26_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2702638(.data_in(wire_d26_37),.data_out(wire_d26_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2702639(.data_in(wire_d26_38),.data_out(wire_d26_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2702640(.data_in(wire_d26_39),.data_out(wire_d26_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2702641(.data_in(wire_d26_40),.data_out(wire_d26_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702642(.data_in(wire_d26_41),.data_out(wire_d26_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2702643(.data_in(wire_d26_42),.data_out(wire_d26_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702644(.data_in(wire_d26_43),.data_out(wire_d26_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702645(.data_in(wire_d26_44),.data_out(wire_d26_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2702646(.data_in(wire_d26_45),.data_out(wire_d26_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2702647(.data_in(wire_d26_46),.data_out(wire_d26_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2702648(.data_in(wire_d26_47),.data_out(wire_d26_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2702649(.data_in(wire_d26_48),.data_out(d_out26),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance280270(.data_in(d_in27),.data_out(wire_d27_0),.clk(clk),.rst(rst));            //channel 28
	large_adder #(.WIDTH(WIDTH)) large_adder_instance280271(.data_in(wire_d27_0),.data_out(wire_d27_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance280272(.data_in(wire_d27_1),.data_out(wire_d27_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance280273(.data_in(wire_d27_2),.data_out(wire_d27_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance280274(.data_in(wire_d27_3),.data_out(wire_d27_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance280275(.data_in(wire_d27_4),.data_out(wire_d27_5),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance280276(.data_in(wire_d27_5),.data_out(wire_d27_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance280277(.data_in(wire_d27_6),.data_out(wire_d27_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance280278(.data_in(wire_d27_7),.data_out(wire_d27_8),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance280279(.data_in(wire_d27_8),.data_out(wire_d27_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802710(.data_in(wire_d27_9),.data_out(wire_d27_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2802711(.data_in(wire_d27_10),.data_out(wire_d27_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802712(.data_in(wire_d27_11),.data_out(wire_d27_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802713(.data_in(wire_d27_12),.data_out(wire_d27_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802714(.data_in(wire_d27_13),.data_out(wire_d27_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802715(.data_in(wire_d27_14),.data_out(wire_d27_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802716(.data_in(wire_d27_15),.data_out(wire_d27_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802717(.data_in(wire_d27_16),.data_out(wire_d27_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802718(.data_in(wire_d27_17),.data_out(wire_d27_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802719(.data_in(wire_d27_18),.data_out(wire_d27_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2802720(.data_in(wire_d27_19),.data_out(wire_d27_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802721(.data_in(wire_d27_20),.data_out(wire_d27_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802722(.data_in(wire_d27_21),.data_out(wire_d27_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802723(.data_in(wire_d27_22),.data_out(wire_d27_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802724(.data_in(wire_d27_23),.data_out(wire_d27_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802725(.data_in(wire_d27_24),.data_out(wire_d27_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802726(.data_in(wire_d27_25),.data_out(wire_d27_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802727(.data_in(wire_d27_26),.data_out(wire_d27_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802728(.data_in(wire_d27_27),.data_out(wire_d27_28),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802729(.data_in(wire_d27_28),.data_out(wire_d27_29),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2802730(.data_in(wire_d27_29),.data_out(wire_d27_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2802731(.data_in(wire_d27_30),.data_out(wire_d27_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2802732(.data_in(wire_d27_31),.data_out(wire_d27_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2802733(.data_in(wire_d27_32),.data_out(wire_d27_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802734(.data_in(wire_d27_33),.data_out(wire_d27_34),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2802735(.data_in(wire_d27_34),.data_out(wire_d27_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2802736(.data_in(wire_d27_35),.data_out(wire_d27_36),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2802737(.data_in(wire_d27_36),.data_out(wire_d27_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2802738(.data_in(wire_d27_37),.data_out(wire_d27_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802739(.data_in(wire_d27_38),.data_out(wire_d27_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2802740(.data_in(wire_d27_39),.data_out(wire_d27_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2802741(.data_in(wire_d27_40),.data_out(wire_d27_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2802742(.data_in(wire_d27_41),.data_out(wire_d27_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802743(.data_in(wire_d27_42),.data_out(wire_d27_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2802744(.data_in(wire_d27_43),.data_out(wire_d27_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2802745(.data_in(wire_d27_44),.data_out(wire_d27_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2802746(.data_in(wire_d27_45),.data_out(wire_d27_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2802747(.data_in(wire_d27_46),.data_out(wire_d27_47),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2802748(.data_in(wire_d27_47),.data_out(wire_d27_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2802749(.data_in(wire_d27_48),.data_out(d_out27),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance290280(.data_in(d_in28),.data_out(wire_d28_0),.clk(clk),.rst(rst));            //channel 29
	encoder #(.WIDTH(WIDTH)) encoder_instance290281(.data_in(wire_d28_0),.data_out(wire_d28_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance290282(.data_in(wire_d28_1),.data_out(wire_d28_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance290283(.data_in(wire_d28_2),.data_out(wire_d28_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance290284(.data_in(wire_d28_3),.data_out(wire_d28_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance290285(.data_in(wire_d28_4),.data_out(wire_d28_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance290286(.data_in(wire_d28_5),.data_out(wire_d28_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance290287(.data_in(wire_d28_6),.data_out(wire_d28_7),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance290288(.data_in(wire_d28_7),.data_out(wire_d28_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance290289(.data_in(wire_d28_8),.data_out(wire_d28_9),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902810(.data_in(wire_d28_9),.data_out(wire_d28_10),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902811(.data_in(wire_d28_10),.data_out(wire_d28_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902812(.data_in(wire_d28_11),.data_out(wire_d28_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902813(.data_in(wire_d28_12),.data_out(wire_d28_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2902814(.data_in(wire_d28_13),.data_out(wire_d28_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902815(.data_in(wire_d28_14),.data_out(wire_d28_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2902816(.data_in(wire_d28_15),.data_out(wire_d28_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902817(.data_in(wire_d28_16),.data_out(wire_d28_17),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902818(.data_in(wire_d28_17),.data_out(wire_d28_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902819(.data_in(wire_d28_18),.data_out(wire_d28_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2902820(.data_in(wire_d28_19),.data_out(wire_d28_20),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance2902821(.data_in(wire_d28_20),.data_out(wire_d28_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902822(.data_in(wire_d28_21),.data_out(wire_d28_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2902823(.data_in(wire_d28_22),.data_out(wire_d28_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance2902824(.data_in(wire_d28_23),.data_out(wire_d28_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902825(.data_in(wire_d28_24),.data_out(wire_d28_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902826(.data_in(wire_d28_25),.data_out(wire_d28_26),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2902827(.data_in(wire_d28_26),.data_out(wire_d28_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902828(.data_in(wire_d28_27),.data_out(wire_d28_28),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902829(.data_in(wire_d28_28),.data_out(wire_d28_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance2902830(.data_in(wire_d28_29),.data_out(wire_d28_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902831(.data_in(wire_d28_30),.data_out(wire_d28_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902832(.data_in(wire_d28_31),.data_out(wire_d28_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902833(.data_in(wire_d28_32),.data_out(wire_d28_33),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2902834(.data_in(wire_d28_33),.data_out(wire_d28_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902835(.data_in(wire_d28_34),.data_out(wire_d28_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902836(.data_in(wire_d28_35),.data_out(wire_d28_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance2902837(.data_in(wire_d28_36),.data_out(wire_d28_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2902838(.data_in(wire_d28_37),.data_out(wire_d28_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902839(.data_in(wire_d28_38),.data_out(wire_d28_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance2902840(.data_in(wire_d28_39),.data_out(wire_d28_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance2902841(.data_in(wire_d28_40),.data_out(wire_d28_41),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance2902842(.data_in(wire_d28_41),.data_out(wire_d28_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance2902843(.data_in(wire_d28_42),.data_out(wire_d28_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902844(.data_in(wire_d28_43),.data_out(wire_d28_44),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance2902845(.data_in(wire_d28_44),.data_out(wire_d28_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance2902846(.data_in(wire_d28_45),.data_out(wire_d28_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance2902847(.data_in(wire_d28_46),.data_out(wire_d28_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902848(.data_in(wire_d28_47),.data_out(wire_d28_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance2902849(.data_in(wire_d28_48),.data_out(d_out28),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance300290(.data_in(d_in29),.data_out(wire_d29_0),.clk(clk),.rst(rst));            //channel 30
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance300291(.data_in(wire_d29_0),.data_out(wire_d29_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance300292(.data_in(wire_d29_1),.data_out(wire_d29_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance300293(.data_in(wire_d29_2),.data_out(wire_d29_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance300294(.data_in(wire_d29_3),.data_out(wire_d29_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance300295(.data_in(wire_d29_4),.data_out(wire_d29_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance300296(.data_in(wire_d29_5),.data_out(wire_d29_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance300297(.data_in(wire_d29_6),.data_out(wire_d29_7),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance300298(.data_in(wire_d29_7),.data_out(wire_d29_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance300299(.data_in(wire_d29_8),.data_out(wire_d29_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002910(.data_in(wire_d29_9),.data_out(wire_d29_10),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3002911(.data_in(wire_d29_10),.data_out(wire_d29_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002912(.data_in(wire_d29_11),.data_out(wire_d29_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3002913(.data_in(wire_d29_12),.data_out(wire_d29_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002914(.data_in(wire_d29_13),.data_out(wire_d29_14),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3002915(.data_in(wire_d29_14),.data_out(wire_d29_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3002916(.data_in(wire_d29_15),.data_out(wire_d29_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002917(.data_in(wire_d29_16),.data_out(wire_d29_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002918(.data_in(wire_d29_17),.data_out(wire_d29_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002919(.data_in(wire_d29_18),.data_out(wire_d29_19),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3002920(.data_in(wire_d29_19),.data_out(wire_d29_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3002921(.data_in(wire_d29_20),.data_out(wire_d29_21),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3002922(.data_in(wire_d29_21),.data_out(wire_d29_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3002923(.data_in(wire_d29_22),.data_out(wire_d29_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002924(.data_in(wire_d29_23),.data_out(wire_d29_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3002925(.data_in(wire_d29_24),.data_out(wire_d29_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002926(.data_in(wire_d29_25),.data_out(wire_d29_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3002927(.data_in(wire_d29_26),.data_out(wire_d29_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002928(.data_in(wire_d29_27),.data_out(wire_d29_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3002929(.data_in(wire_d29_28),.data_out(wire_d29_29),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3002930(.data_in(wire_d29_29),.data_out(wire_d29_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002931(.data_in(wire_d29_30),.data_out(wire_d29_31),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002932(.data_in(wire_d29_31),.data_out(wire_d29_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002933(.data_in(wire_d29_32),.data_out(wire_d29_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002934(.data_in(wire_d29_33),.data_out(wire_d29_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002935(.data_in(wire_d29_34),.data_out(wire_d29_35),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3002936(.data_in(wire_d29_35),.data_out(wire_d29_36),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002937(.data_in(wire_d29_36),.data_out(wire_d29_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3002938(.data_in(wire_d29_37),.data_out(wire_d29_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3002939(.data_in(wire_d29_38),.data_out(wire_d29_39),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002940(.data_in(wire_d29_39),.data_out(wire_d29_40),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3002941(.data_in(wire_d29_40),.data_out(wire_d29_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3002942(.data_in(wire_d29_41),.data_out(wire_d29_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002943(.data_in(wire_d29_42),.data_out(wire_d29_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3002944(.data_in(wire_d29_43),.data_out(wire_d29_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3002945(.data_in(wire_d29_44),.data_out(wire_d29_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3002946(.data_in(wire_d29_45),.data_out(wire_d29_46),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3002947(.data_in(wire_d29_46),.data_out(wire_d29_47),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3002948(.data_in(wire_d29_47),.data_out(wire_d29_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3002949(.data_in(wire_d29_48),.data_out(d_out29),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance310300(.data_in(d_in30),.data_out(wire_d30_0),.clk(clk),.rst(rst));            //channel 31
	large_adder #(.WIDTH(WIDTH)) large_adder_instance310301(.data_in(wire_d30_0),.data_out(wire_d30_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance310302(.data_in(wire_d30_1),.data_out(wire_d30_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance310303(.data_in(wire_d30_2),.data_out(wire_d30_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance310304(.data_in(wire_d30_3),.data_out(wire_d30_4),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance310305(.data_in(wire_d30_4),.data_out(wire_d30_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance310306(.data_in(wire_d30_5),.data_out(wire_d30_6),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance310307(.data_in(wire_d30_6),.data_out(wire_d30_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance310308(.data_in(wire_d30_7),.data_out(wire_d30_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance310309(.data_in(wire_d30_8),.data_out(wire_d30_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103010(.data_in(wire_d30_9),.data_out(wire_d30_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103011(.data_in(wire_d30_10),.data_out(wire_d30_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3103012(.data_in(wire_d30_11),.data_out(wire_d30_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103013(.data_in(wire_d30_12),.data_out(wire_d30_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103014(.data_in(wire_d30_13),.data_out(wire_d30_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103015(.data_in(wire_d30_14),.data_out(wire_d30_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3103016(.data_in(wire_d30_15),.data_out(wire_d30_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3103017(.data_in(wire_d30_16),.data_out(wire_d30_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103018(.data_in(wire_d30_17),.data_out(wire_d30_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3103019(.data_in(wire_d30_18),.data_out(wire_d30_19),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103020(.data_in(wire_d30_19),.data_out(wire_d30_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3103021(.data_in(wire_d30_20),.data_out(wire_d30_21),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3103022(.data_in(wire_d30_21),.data_out(wire_d30_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103023(.data_in(wire_d30_22),.data_out(wire_d30_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103024(.data_in(wire_d30_23),.data_out(wire_d30_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103025(.data_in(wire_d30_24),.data_out(wire_d30_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103026(.data_in(wire_d30_25),.data_out(wire_d30_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103027(.data_in(wire_d30_26),.data_out(wire_d30_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3103028(.data_in(wire_d30_27),.data_out(wire_d30_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3103029(.data_in(wire_d30_28),.data_out(wire_d30_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103030(.data_in(wire_d30_29),.data_out(wire_d30_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103031(.data_in(wire_d30_30),.data_out(wire_d30_31),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3103032(.data_in(wire_d30_31),.data_out(wire_d30_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3103033(.data_in(wire_d30_32),.data_out(wire_d30_33),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3103034(.data_in(wire_d30_33),.data_out(wire_d30_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3103035(.data_in(wire_d30_34),.data_out(wire_d30_35),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103036(.data_in(wire_d30_35),.data_out(wire_d30_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103037(.data_in(wire_d30_36),.data_out(wire_d30_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103038(.data_in(wire_d30_37),.data_out(wire_d30_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3103039(.data_in(wire_d30_38),.data_out(wire_d30_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103040(.data_in(wire_d30_39),.data_out(wire_d30_40),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3103041(.data_in(wire_d30_40),.data_out(wire_d30_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103042(.data_in(wire_d30_41),.data_out(wire_d30_42),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3103043(.data_in(wire_d30_42),.data_out(wire_d30_43),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3103044(.data_in(wire_d30_43),.data_out(wire_d30_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3103045(.data_in(wire_d30_44),.data_out(wire_d30_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3103046(.data_in(wire_d30_45),.data_out(wire_d30_46),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3103047(.data_in(wire_d30_46),.data_out(wire_d30_47),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3103048(.data_in(wire_d30_47),.data_out(wire_d30_48),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3103049(.data_in(wire_d30_48),.data_out(d_out30),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance320310(.data_in(d_in31),.data_out(wire_d31_0),.clk(clk),.rst(rst));            //channel 32
	encoder #(.WIDTH(WIDTH)) encoder_instance320311(.data_in(wire_d31_0),.data_out(wire_d31_1),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance320312(.data_in(wire_d31_1),.data_out(wire_d31_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance320313(.data_in(wire_d31_2),.data_out(wire_d31_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance320314(.data_in(wire_d31_3),.data_out(wire_d31_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance320315(.data_in(wire_d31_4),.data_out(wire_d31_5),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance320316(.data_in(wire_d31_5),.data_out(wire_d31_6),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance320317(.data_in(wire_d31_6),.data_out(wire_d31_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance320318(.data_in(wire_d31_7),.data_out(wire_d31_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance320319(.data_in(wire_d31_8),.data_out(wire_d31_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3203110(.data_in(wire_d31_9),.data_out(wire_d31_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203111(.data_in(wire_d31_10),.data_out(wire_d31_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203112(.data_in(wire_d31_11),.data_out(wire_d31_12),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203113(.data_in(wire_d31_12),.data_out(wire_d31_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3203114(.data_in(wire_d31_13),.data_out(wire_d31_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203115(.data_in(wire_d31_14),.data_out(wire_d31_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3203116(.data_in(wire_d31_15),.data_out(wire_d31_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203117(.data_in(wire_d31_16),.data_out(wire_d31_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203118(.data_in(wire_d31_17),.data_out(wire_d31_18),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203119(.data_in(wire_d31_18),.data_out(wire_d31_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203120(.data_in(wire_d31_19),.data_out(wire_d31_20),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203121(.data_in(wire_d31_20),.data_out(wire_d31_21),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3203122(.data_in(wire_d31_21),.data_out(wire_d31_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203123(.data_in(wire_d31_22),.data_out(wire_d31_23),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203124(.data_in(wire_d31_23),.data_out(wire_d31_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203125(.data_in(wire_d31_24),.data_out(wire_d31_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203126(.data_in(wire_d31_25),.data_out(wire_d31_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203127(.data_in(wire_d31_26),.data_out(wire_d31_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203128(.data_in(wire_d31_27),.data_out(wire_d31_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203129(.data_in(wire_d31_28),.data_out(wire_d31_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3203130(.data_in(wire_d31_29),.data_out(wire_d31_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203131(.data_in(wire_d31_30),.data_out(wire_d31_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203132(.data_in(wire_d31_31),.data_out(wire_d31_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203133(.data_in(wire_d31_32),.data_out(wire_d31_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203134(.data_in(wire_d31_33),.data_out(wire_d31_34),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3203135(.data_in(wire_d31_34),.data_out(wire_d31_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203136(.data_in(wire_d31_35),.data_out(wire_d31_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3203137(.data_in(wire_d31_36),.data_out(wire_d31_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3203138(.data_in(wire_d31_37),.data_out(wire_d31_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203139(.data_in(wire_d31_38),.data_out(wire_d31_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203140(.data_in(wire_d31_39),.data_out(wire_d31_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3203141(.data_in(wire_d31_40),.data_out(wire_d31_41),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3203142(.data_in(wire_d31_41),.data_out(wire_d31_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3203143(.data_in(wire_d31_42),.data_out(wire_d31_43),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203144(.data_in(wire_d31_43),.data_out(wire_d31_44),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3203145(.data_in(wire_d31_44),.data_out(wire_d31_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3203146(.data_in(wire_d31_45),.data_out(wire_d31_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3203147(.data_in(wire_d31_46),.data_out(wire_d31_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3203148(.data_in(wire_d31_47),.data_out(wire_d31_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3203149(.data_in(wire_d31_48),.data_out(d_out31),.clk(clk),.rst(rst));

	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance330320(.data_in(d_in32),.data_out(wire_d32_0),.clk(clk),.rst(rst));            //channel 33
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance330321(.data_in(wire_d32_0),.data_out(wire_d32_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance330322(.data_in(wire_d32_1),.data_out(wire_d32_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance330323(.data_in(wire_d32_2),.data_out(wire_d32_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance330324(.data_in(wire_d32_3),.data_out(wire_d32_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance330325(.data_in(wire_d32_4),.data_out(wire_d32_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance330326(.data_in(wire_d32_5),.data_out(wire_d32_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance330327(.data_in(wire_d32_6),.data_out(wire_d32_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance330328(.data_in(wire_d32_7),.data_out(wire_d32_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance330329(.data_in(wire_d32_8),.data_out(wire_d32_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303210(.data_in(wire_d32_9),.data_out(wire_d32_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303211(.data_in(wire_d32_10),.data_out(wire_d32_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303212(.data_in(wire_d32_11),.data_out(wire_d32_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3303213(.data_in(wire_d32_12),.data_out(wire_d32_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303214(.data_in(wire_d32_13),.data_out(wire_d32_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303215(.data_in(wire_d32_14),.data_out(wire_d32_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303216(.data_in(wire_d32_15),.data_out(wire_d32_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303217(.data_in(wire_d32_16),.data_out(wire_d32_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3303218(.data_in(wire_d32_17),.data_out(wire_d32_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303219(.data_in(wire_d32_18),.data_out(wire_d32_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303220(.data_in(wire_d32_19),.data_out(wire_d32_20),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3303221(.data_in(wire_d32_20),.data_out(wire_d32_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3303222(.data_in(wire_d32_21),.data_out(wire_d32_22),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303223(.data_in(wire_d32_22),.data_out(wire_d32_23),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303224(.data_in(wire_d32_23),.data_out(wire_d32_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3303225(.data_in(wire_d32_24),.data_out(wire_d32_25),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303226(.data_in(wire_d32_25),.data_out(wire_d32_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303227(.data_in(wire_d32_26),.data_out(wire_d32_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3303228(.data_in(wire_d32_27),.data_out(wire_d32_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3303229(.data_in(wire_d32_28),.data_out(wire_d32_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303230(.data_in(wire_d32_29),.data_out(wire_d32_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3303231(.data_in(wire_d32_30),.data_out(wire_d32_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303232(.data_in(wire_d32_31),.data_out(wire_d32_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303233(.data_in(wire_d32_32),.data_out(wire_d32_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3303234(.data_in(wire_d32_33),.data_out(wire_d32_34),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3303235(.data_in(wire_d32_34),.data_out(wire_d32_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3303236(.data_in(wire_d32_35),.data_out(wire_d32_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3303237(.data_in(wire_d32_36),.data_out(wire_d32_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3303238(.data_in(wire_d32_37),.data_out(wire_d32_38),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3303239(.data_in(wire_d32_38),.data_out(wire_d32_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303240(.data_in(wire_d32_39),.data_out(wire_d32_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303241(.data_in(wire_d32_40),.data_out(wire_d32_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303242(.data_in(wire_d32_41),.data_out(wire_d32_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3303243(.data_in(wire_d32_42),.data_out(wire_d32_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3303244(.data_in(wire_d32_43),.data_out(wire_d32_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3303245(.data_in(wire_d32_44),.data_out(wire_d32_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3303246(.data_in(wire_d32_45),.data_out(wire_d32_46),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3303247(.data_in(wire_d32_46),.data_out(wire_d32_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3303248(.data_in(wire_d32_47),.data_out(wire_d32_48),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3303249(.data_in(wire_d32_48),.data_out(d_out32),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance340330(.data_in(d_in33),.data_out(wire_d33_0),.clk(clk),.rst(rst));            //channel 34
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance340331(.data_in(wire_d33_0),.data_out(wire_d33_1),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance340332(.data_in(wire_d33_1),.data_out(wire_d33_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance340333(.data_in(wire_d33_2),.data_out(wire_d33_3),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance340334(.data_in(wire_d33_3),.data_out(wire_d33_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance340335(.data_in(wire_d33_4),.data_out(wire_d33_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance340336(.data_in(wire_d33_5),.data_out(wire_d33_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance340337(.data_in(wire_d33_6),.data_out(wire_d33_7),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance340338(.data_in(wire_d33_7),.data_out(wire_d33_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance340339(.data_in(wire_d33_8),.data_out(wire_d33_9),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3403310(.data_in(wire_d33_9),.data_out(wire_d33_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3403311(.data_in(wire_d33_10),.data_out(wire_d33_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403312(.data_in(wire_d33_11),.data_out(wire_d33_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403313(.data_in(wire_d33_12),.data_out(wire_d33_13),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3403314(.data_in(wire_d33_13),.data_out(wire_d33_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403315(.data_in(wire_d33_14),.data_out(wire_d33_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403316(.data_in(wire_d33_15),.data_out(wire_d33_16),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403317(.data_in(wire_d33_16),.data_out(wire_d33_17),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3403318(.data_in(wire_d33_17),.data_out(wire_d33_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3403319(.data_in(wire_d33_18),.data_out(wire_d33_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403320(.data_in(wire_d33_19),.data_out(wire_d33_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3403321(.data_in(wire_d33_20),.data_out(wire_d33_21),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3403322(.data_in(wire_d33_21),.data_out(wire_d33_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3403323(.data_in(wire_d33_22),.data_out(wire_d33_23),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403324(.data_in(wire_d33_23),.data_out(wire_d33_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403325(.data_in(wire_d33_24),.data_out(wire_d33_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403326(.data_in(wire_d33_25),.data_out(wire_d33_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403327(.data_in(wire_d33_26),.data_out(wire_d33_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3403328(.data_in(wire_d33_27),.data_out(wire_d33_28),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3403329(.data_in(wire_d33_28),.data_out(wire_d33_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3403330(.data_in(wire_d33_29),.data_out(wire_d33_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3403331(.data_in(wire_d33_30),.data_out(wire_d33_31),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3403332(.data_in(wire_d33_31),.data_out(wire_d33_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403333(.data_in(wire_d33_32),.data_out(wire_d33_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3403334(.data_in(wire_d33_33),.data_out(wire_d33_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3403335(.data_in(wire_d33_34),.data_out(wire_d33_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3403336(.data_in(wire_d33_35),.data_out(wire_d33_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403337(.data_in(wire_d33_36),.data_out(wire_d33_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403338(.data_in(wire_d33_37),.data_out(wire_d33_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3403339(.data_in(wire_d33_38),.data_out(wire_d33_39),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3403340(.data_in(wire_d33_39),.data_out(wire_d33_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3403341(.data_in(wire_d33_40),.data_out(wire_d33_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403342(.data_in(wire_d33_41),.data_out(wire_d33_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3403343(.data_in(wire_d33_42),.data_out(wire_d33_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3403344(.data_in(wire_d33_43),.data_out(wire_d33_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3403345(.data_in(wire_d33_44),.data_out(wire_d33_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3403346(.data_in(wire_d33_45),.data_out(wire_d33_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3403347(.data_in(wire_d33_46),.data_out(wire_d33_47),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3403348(.data_in(wire_d33_47),.data_out(wire_d33_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3403349(.data_in(wire_d33_48),.data_out(d_out33),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance350340(.data_in(d_in34),.data_out(wire_d34_0),.clk(clk),.rst(rst));            //channel 35
	decoder_top #(.WIDTH(WIDTH)) decoder_instance350341(.data_in(wire_d34_0),.data_out(wire_d34_1),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance350342(.data_in(wire_d34_1),.data_out(wire_d34_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance350343(.data_in(wire_d34_2),.data_out(wire_d34_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance350344(.data_in(wire_d34_3),.data_out(wire_d34_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance350345(.data_in(wire_d34_4),.data_out(wire_d34_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance350346(.data_in(wire_d34_5),.data_out(wire_d34_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance350347(.data_in(wire_d34_6),.data_out(wire_d34_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance350348(.data_in(wire_d34_7),.data_out(wire_d34_8),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance350349(.data_in(wire_d34_8),.data_out(wire_d34_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3503410(.data_in(wire_d34_9),.data_out(wire_d34_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503411(.data_in(wire_d34_10),.data_out(wire_d34_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503412(.data_in(wire_d34_11),.data_out(wire_d34_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3503413(.data_in(wire_d34_12),.data_out(wire_d34_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503414(.data_in(wire_d34_13),.data_out(wire_d34_14),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3503415(.data_in(wire_d34_14),.data_out(wire_d34_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503416(.data_in(wire_d34_15),.data_out(wire_d34_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3503417(.data_in(wire_d34_16),.data_out(wire_d34_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503418(.data_in(wire_d34_17),.data_out(wire_d34_18),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503419(.data_in(wire_d34_18),.data_out(wire_d34_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503420(.data_in(wire_d34_19),.data_out(wire_d34_20),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3503421(.data_in(wire_d34_20),.data_out(wire_d34_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503422(.data_in(wire_d34_21),.data_out(wire_d34_22),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3503423(.data_in(wire_d34_22),.data_out(wire_d34_23),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503424(.data_in(wire_d34_23),.data_out(wire_d34_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3503425(.data_in(wire_d34_24),.data_out(wire_d34_25),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503426(.data_in(wire_d34_25),.data_out(wire_d34_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503427(.data_in(wire_d34_26),.data_out(wire_d34_27),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503428(.data_in(wire_d34_27),.data_out(wire_d34_28),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503429(.data_in(wire_d34_28),.data_out(wire_d34_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503430(.data_in(wire_d34_29),.data_out(wire_d34_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3503431(.data_in(wire_d34_30),.data_out(wire_d34_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503432(.data_in(wire_d34_31),.data_out(wire_d34_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3503433(.data_in(wire_d34_32),.data_out(wire_d34_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503434(.data_in(wire_d34_33),.data_out(wire_d34_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3503435(.data_in(wire_d34_34),.data_out(wire_d34_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3503436(.data_in(wire_d34_35),.data_out(wire_d34_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503437(.data_in(wire_d34_36),.data_out(wire_d34_37),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3503438(.data_in(wire_d34_37),.data_out(wire_d34_38),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503439(.data_in(wire_d34_38),.data_out(wire_d34_39),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3503440(.data_in(wire_d34_39),.data_out(wire_d34_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3503441(.data_in(wire_d34_40),.data_out(wire_d34_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3503442(.data_in(wire_d34_41),.data_out(wire_d34_42),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3503443(.data_in(wire_d34_42),.data_out(wire_d34_43),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503444(.data_in(wire_d34_43),.data_out(wire_d34_44),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3503445(.data_in(wire_d34_44),.data_out(wire_d34_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3503446(.data_in(wire_d34_45),.data_out(wire_d34_46),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3503447(.data_in(wire_d34_46),.data_out(wire_d34_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3503448(.data_in(wire_d34_47),.data_out(wire_d34_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3503449(.data_in(wire_d34_48),.data_out(d_out34),.clk(clk),.rst(rst));

	large_adder #(.WIDTH(WIDTH)) large_adder_instance360350(.data_in(d_in35),.data_out(wire_d35_0),.clk(clk),.rst(rst));            //channel 36
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance360351(.data_in(wire_d35_0),.data_out(wire_d35_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance360352(.data_in(wire_d35_1),.data_out(wire_d35_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance360353(.data_in(wire_d35_2),.data_out(wire_d35_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance360354(.data_in(wire_d35_3),.data_out(wire_d35_4),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance360355(.data_in(wire_d35_4),.data_out(wire_d35_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance360356(.data_in(wire_d35_5),.data_out(wire_d35_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance360357(.data_in(wire_d35_6),.data_out(wire_d35_7),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance360358(.data_in(wire_d35_7),.data_out(wire_d35_8),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance360359(.data_in(wire_d35_8),.data_out(wire_d35_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603510(.data_in(wire_d35_9),.data_out(wire_d35_10),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603511(.data_in(wire_d35_10),.data_out(wire_d35_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3603512(.data_in(wire_d35_11),.data_out(wire_d35_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603513(.data_in(wire_d35_12),.data_out(wire_d35_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3603514(.data_in(wire_d35_13),.data_out(wire_d35_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603515(.data_in(wire_d35_14),.data_out(wire_d35_15),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603516(.data_in(wire_d35_15),.data_out(wire_d35_16),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3603517(.data_in(wire_d35_16),.data_out(wire_d35_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603518(.data_in(wire_d35_17),.data_out(wire_d35_18),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603519(.data_in(wire_d35_18),.data_out(wire_d35_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603520(.data_in(wire_d35_19),.data_out(wire_d35_20),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3603521(.data_in(wire_d35_20),.data_out(wire_d35_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3603522(.data_in(wire_d35_21),.data_out(wire_d35_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3603523(.data_in(wire_d35_22),.data_out(wire_d35_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603524(.data_in(wire_d35_23),.data_out(wire_d35_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603525(.data_in(wire_d35_24),.data_out(wire_d35_25),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3603526(.data_in(wire_d35_25),.data_out(wire_d35_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603527(.data_in(wire_d35_26),.data_out(wire_d35_27),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3603528(.data_in(wire_d35_27),.data_out(wire_d35_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603529(.data_in(wire_d35_28),.data_out(wire_d35_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603530(.data_in(wire_d35_29),.data_out(wire_d35_30),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603531(.data_in(wire_d35_30),.data_out(wire_d35_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3603532(.data_in(wire_d35_31),.data_out(wire_d35_32),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603533(.data_in(wire_d35_32),.data_out(wire_d35_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603534(.data_in(wire_d35_33),.data_out(wire_d35_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3603535(.data_in(wire_d35_34),.data_out(wire_d35_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3603536(.data_in(wire_d35_35),.data_out(wire_d35_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3603537(.data_in(wire_d35_36),.data_out(wire_d35_37),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3603538(.data_in(wire_d35_37),.data_out(wire_d35_38),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603539(.data_in(wire_d35_38),.data_out(wire_d35_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603540(.data_in(wire_d35_39),.data_out(wire_d35_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603541(.data_in(wire_d35_40),.data_out(wire_d35_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603542(.data_in(wire_d35_41),.data_out(wire_d35_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3603543(.data_in(wire_d35_42),.data_out(wire_d35_43),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603544(.data_in(wire_d35_43),.data_out(wire_d35_44),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3603545(.data_in(wire_d35_44),.data_out(wire_d35_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3603546(.data_in(wire_d35_45),.data_out(wire_d35_46),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3603547(.data_in(wire_d35_46),.data_out(wire_d35_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3603548(.data_in(wire_d35_47),.data_out(wire_d35_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3603549(.data_in(wire_d35_48),.data_out(d_out35),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance370360(.data_in(d_in36),.data_out(wire_d36_0),.clk(clk),.rst(rst));            //channel 37
	register #(.WIDTH(WIDTH)) register_instance370361(.data_in(wire_d36_0),.data_out(wire_d36_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance370362(.data_in(wire_d36_1),.data_out(wire_d36_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance370363(.data_in(wire_d36_2),.data_out(wire_d36_3),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance370364(.data_in(wire_d36_3),.data_out(wire_d36_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance370365(.data_in(wire_d36_4),.data_out(wire_d36_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance370366(.data_in(wire_d36_5),.data_out(wire_d36_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance370367(.data_in(wire_d36_6),.data_out(wire_d36_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance370368(.data_in(wire_d36_7),.data_out(wire_d36_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance370369(.data_in(wire_d36_8),.data_out(wire_d36_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703610(.data_in(wire_d36_9),.data_out(wire_d36_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703611(.data_in(wire_d36_10),.data_out(wire_d36_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3703612(.data_in(wire_d36_11),.data_out(wire_d36_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703613(.data_in(wire_d36_12),.data_out(wire_d36_13),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703614(.data_in(wire_d36_13),.data_out(wire_d36_14),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703615(.data_in(wire_d36_14),.data_out(wire_d36_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703616(.data_in(wire_d36_15),.data_out(wire_d36_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703617(.data_in(wire_d36_16),.data_out(wire_d36_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703618(.data_in(wire_d36_17),.data_out(wire_d36_18),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3703619(.data_in(wire_d36_18),.data_out(wire_d36_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703620(.data_in(wire_d36_19),.data_out(wire_d36_20),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3703621(.data_in(wire_d36_20),.data_out(wire_d36_21),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3703622(.data_in(wire_d36_21),.data_out(wire_d36_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703623(.data_in(wire_d36_22),.data_out(wire_d36_23),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3703624(.data_in(wire_d36_23),.data_out(wire_d36_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3703625(.data_in(wire_d36_24),.data_out(wire_d36_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703626(.data_in(wire_d36_25),.data_out(wire_d36_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703627(.data_in(wire_d36_26),.data_out(wire_d36_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3703628(.data_in(wire_d36_27),.data_out(wire_d36_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3703629(.data_in(wire_d36_28),.data_out(wire_d36_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3703630(.data_in(wire_d36_29),.data_out(wire_d36_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3703631(.data_in(wire_d36_30),.data_out(wire_d36_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3703632(.data_in(wire_d36_31),.data_out(wire_d36_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703633(.data_in(wire_d36_32),.data_out(wire_d36_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3703634(.data_in(wire_d36_33),.data_out(wire_d36_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3703635(.data_in(wire_d36_34),.data_out(wire_d36_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703636(.data_in(wire_d36_35),.data_out(wire_d36_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703637(.data_in(wire_d36_36),.data_out(wire_d36_37),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3703638(.data_in(wire_d36_37),.data_out(wire_d36_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3703639(.data_in(wire_d36_38),.data_out(wire_d36_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3703640(.data_in(wire_d36_39),.data_out(wire_d36_40),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3703641(.data_in(wire_d36_40),.data_out(wire_d36_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703642(.data_in(wire_d36_41),.data_out(wire_d36_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3703643(.data_in(wire_d36_42),.data_out(wire_d36_43),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3703644(.data_in(wire_d36_43),.data_out(wire_d36_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3703645(.data_in(wire_d36_44),.data_out(wire_d36_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3703646(.data_in(wire_d36_45),.data_out(wire_d36_46),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3703647(.data_in(wire_d36_46),.data_out(wire_d36_47),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3703648(.data_in(wire_d36_47),.data_out(wire_d36_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3703649(.data_in(wire_d36_48),.data_out(d_out36),.clk(clk),.rst(rst));

	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance380370(.data_in(d_in37),.data_out(wire_d37_0),.clk(clk),.rst(rst));            //channel 38
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance380371(.data_in(wire_d37_0),.data_out(wire_d37_1),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance380372(.data_in(wire_d37_1),.data_out(wire_d37_2),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance380373(.data_in(wire_d37_2),.data_out(wire_d37_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance380374(.data_in(wire_d37_3),.data_out(wire_d37_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance380375(.data_in(wire_d37_4),.data_out(wire_d37_5),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance380376(.data_in(wire_d37_5),.data_out(wire_d37_6),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance380377(.data_in(wire_d37_6),.data_out(wire_d37_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance380378(.data_in(wire_d37_7),.data_out(wire_d37_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance380379(.data_in(wire_d37_8),.data_out(wire_d37_9),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3803710(.data_in(wire_d37_9),.data_out(wire_d37_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803711(.data_in(wire_d37_10),.data_out(wire_d37_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803712(.data_in(wire_d37_11),.data_out(wire_d37_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3803713(.data_in(wire_d37_12),.data_out(wire_d37_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803714(.data_in(wire_d37_13),.data_out(wire_d37_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803715(.data_in(wire_d37_14),.data_out(wire_d37_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803716(.data_in(wire_d37_15),.data_out(wire_d37_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803717(.data_in(wire_d37_16),.data_out(wire_d37_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803718(.data_in(wire_d37_17),.data_out(wire_d37_18),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803719(.data_in(wire_d37_18),.data_out(wire_d37_19),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3803720(.data_in(wire_d37_19),.data_out(wire_d37_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803721(.data_in(wire_d37_20),.data_out(wire_d37_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803722(.data_in(wire_d37_21),.data_out(wire_d37_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803723(.data_in(wire_d37_22),.data_out(wire_d37_23),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3803724(.data_in(wire_d37_23),.data_out(wire_d37_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803725(.data_in(wire_d37_24),.data_out(wire_d37_25),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3803726(.data_in(wire_d37_25),.data_out(wire_d37_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3803727(.data_in(wire_d37_26),.data_out(wire_d37_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803728(.data_in(wire_d37_27),.data_out(wire_d37_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3803729(.data_in(wire_d37_28),.data_out(wire_d37_29),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3803730(.data_in(wire_d37_29),.data_out(wire_d37_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803731(.data_in(wire_d37_30),.data_out(wire_d37_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803732(.data_in(wire_d37_31),.data_out(wire_d37_32),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3803733(.data_in(wire_d37_32),.data_out(wire_d37_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803734(.data_in(wire_d37_33),.data_out(wire_d37_34),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803735(.data_in(wire_d37_34),.data_out(wire_d37_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803736(.data_in(wire_d37_35),.data_out(wire_d37_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3803737(.data_in(wire_d37_36),.data_out(wire_d37_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3803738(.data_in(wire_d37_37),.data_out(wire_d37_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803739(.data_in(wire_d37_38),.data_out(wire_d37_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3803740(.data_in(wire_d37_39),.data_out(wire_d37_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803741(.data_in(wire_d37_40),.data_out(wire_d37_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3803742(.data_in(wire_d37_41),.data_out(wire_d37_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3803743(.data_in(wire_d37_42),.data_out(wire_d37_43),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3803744(.data_in(wire_d37_43),.data_out(wire_d37_44),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3803745(.data_in(wire_d37_44),.data_out(wire_d37_45),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3803746(.data_in(wire_d37_45),.data_out(wire_d37_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3803747(.data_in(wire_d37_46),.data_out(wire_d37_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3803748(.data_in(wire_d37_47),.data_out(wire_d37_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3803749(.data_in(wire_d37_48),.data_out(d_out37),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance390380(.data_in(d_in38),.data_out(wire_d38_0),.clk(clk),.rst(rst));            //channel 39
	large_mux #(.WIDTH(WIDTH)) large_mux_instance390381(.data_in(wire_d38_0),.data_out(wire_d38_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance390382(.data_in(wire_d38_1),.data_out(wire_d38_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance390383(.data_in(wire_d38_2),.data_out(wire_d38_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance390384(.data_in(wire_d38_3),.data_out(wire_d38_4),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance390385(.data_in(wire_d38_4),.data_out(wire_d38_5),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance390386(.data_in(wire_d38_5),.data_out(wire_d38_6),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance390387(.data_in(wire_d38_6),.data_out(wire_d38_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance390388(.data_in(wire_d38_7),.data_out(wire_d38_8),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance390389(.data_in(wire_d38_8),.data_out(wire_d38_9),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903810(.data_in(wire_d38_9),.data_out(wire_d38_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903811(.data_in(wire_d38_10),.data_out(wire_d38_11),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903812(.data_in(wire_d38_11),.data_out(wire_d38_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3903813(.data_in(wire_d38_12),.data_out(wire_d38_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903814(.data_in(wire_d38_13),.data_out(wire_d38_14),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903815(.data_in(wire_d38_14),.data_out(wire_d38_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903816(.data_in(wire_d38_15),.data_out(wire_d38_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3903817(.data_in(wire_d38_16),.data_out(wire_d38_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903818(.data_in(wire_d38_17),.data_out(wire_d38_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3903819(.data_in(wire_d38_18),.data_out(wire_d38_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903820(.data_in(wire_d38_19),.data_out(wire_d38_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3903821(.data_in(wire_d38_20),.data_out(wire_d38_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903822(.data_in(wire_d38_21),.data_out(wire_d38_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3903823(.data_in(wire_d38_22),.data_out(wire_d38_23),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903824(.data_in(wire_d38_23),.data_out(wire_d38_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3903825(.data_in(wire_d38_24),.data_out(wire_d38_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3903826(.data_in(wire_d38_25),.data_out(wire_d38_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903827(.data_in(wire_d38_26),.data_out(wire_d38_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3903828(.data_in(wire_d38_27),.data_out(wire_d38_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance3903829(.data_in(wire_d38_28),.data_out(wire_d38_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903830(.data_in(wire_d38_29),.data_out(wire_d38_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903831(.data_in(wire_d38_30),.data_out(wire_d38_31),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3903832(.data_in(wire_d38_31),.data_out(wire_d38_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903833(.data_in(wire_d38_32),.data_out(wire_d38_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903834(.data_in(wire_d38_33),.data_out(wire_d38_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance3903835(.data_in(wire_d38_34),.data_out(wire_d38_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance3903836(.data_in(wire_d38_35),.data_out(wire_d38_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3903837(.data_in(wire_d38_36),.data_out(wire_d38_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance3903838(.data_in(wire_d38_37),.data_out(wire_d38_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance3903839(.data_in(wire_d38_38),.data_out(wire_d38_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance3903840(.data_in(wire_d38_39),.data_out(wire_d38_40),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903841(.data_in(wire_d38_40),.data_out(wire_d38_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903842(.data_in(wire_d38_41),.data_out(wire_d38_42),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903843(.data_in(wire_d38_42),.data_out(wire_d38_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance3903844(.data_in(wire_d38_43),.data_out(wire_d38_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance3903845(.data_in(wire_d38_44),.data_out(wire_d38_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance3903846(.data_in(wire_d38_45),.data_out(wire_d38_46),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance3903847(.data_in(wire_d38_46),.data_out(wire_d38_47),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance3903848(.data_in(wire_d38_47),.data_out(wire_d38_48),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance3903849(.data_in(wire_d38_48),.data_out(d_out38),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance400390(.data_in(d_in39),.data_out(wire_d39_0),.clk(clk),.rst(rst));            //channel 40
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance400391(.data_in(wire_d39_0),.data_out(wire_d39_1),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance400392(.data_in(wire_d39_1),.data_out(wire_d39_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance400393(.data_in(wire_d39_2),.data_out(wire_d39_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance400394(.data_in(wire_d39_3),.data_out(wire_d39_4),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance400395(.data_in(wire_d39_4),.data_out(wire_d39_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance400396(.data_in(wire_d39_5),.data_out(wire_d39_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance400397(.data_in(wire_d39_6),.data_out(wire_d39_7),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance400398(.data_in(wire_d39_7),.data_out(wire_d39_8),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance400399(.data_in(wire_d39_8),.data_out(wire_d39_9),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003910(.data_in(wire_d39_9),.data_out(wire_d39_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003911(.data_in(wire_d39_10),.data_out(wire_d39_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003912(.data_in(wire_d39_11),.data_out(wire_d39_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4003913(.data_in(wire_d39_12),.data_out(wire_d39_13),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003914(.data_in(wire_d39_13),.data_out(wire_d39_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4003915(.data_in(wire_d39_14),.data_out(wire_d39_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003916(.data_in(wire_d39_15),.data_out(wire_d39_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003917(.data_in(wire_d39_16),.data_out(wire_d39_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003918(.data_in(wire_d39_17),.data_out(wire_d39_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003919(.data_in(wire_d39_18),.data_out(wire_d39_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003920(.data_in(wire_d39_19),.data_out(wire_d39_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4003921(.data_in(wire_d39_20),.data_out(wire_d39_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003922(.data_in(wire_d39_21),.data_out(wire_d39_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4003923(.data_in(wire_d39_22),.data_out(wire_d39_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4003924(.data_in(wire_d39_23),.data_out(wire_d39_24),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003925(.data_in(wire_d39_24),.data_out(wire_d39_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003926(.data_in(wire_d39_25),.data_out(wire_d39_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003927(.data_in(wire_d39_26),.data_out(wire_d39_27),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4003928(.data_in(wire_d39_27),.data_out(wire_d39_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4003929(.data_in(wire_d39_28),.data_out(wire_d39_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003930(.data_in(wire_d39_29),.data_out(wire_d39_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003931(.data_in(wire_d39_30),.data_out(wire_d39_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003932(.data_in(wire_d39_31),.data_out(wire_d39_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003933(.data_in(wire_d39_32),.data_out(wire_d39_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003934(.data_in(wire_d39_33),.data_out(wire_d39_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4003935(.data_in(wire_d39_34),.data_out(wire_d39_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4003936(.data_in(wire_d39_35),.data_out(wire_d39_36),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003937(.data_in(wire_d39_36),.data_out(wire_d39_37),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4003938(.data_in(wire_d39_37),.data_out(wire_d39_38),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4003939(.data_in(wire_d39_38),.data_out(wire_d39_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4003940(.data_in(wire_d39_39),.data_out(wire_d39_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4003941(.data_in(wire_d39_40),.data_out(wire_d39_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4003942(.data_in(wire_d39_41),.data_out(wire_d39_42),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4003943(.data_in(wire_d39_42),.data_out(wire_d39_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4003944(.data_in(wire_d39_43),.data_out(wire_d39_44),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4003945(.data_in(wire_d39_44),.data_out(wire_d39_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4003946(.data_in(wire_d39_45),.data_out(wire_d39_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4003947(.data_in(wire_d39_46),.data_out(wire_d39_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003948(.data_in(wire_d39_47),.data_out(wire_d39_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4003949(.data_in(wire_d39_48),.data_out(d_out39),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance410400(.data_in(d_in40),.data_out(wire_d40_0),.clk(clk),.rst(rst));            //channel 41
	invertion #(.WIDTH(WIDTH)) invertion_instance410401(.data_in(wire_d40_0),.data_out(wire_d40_1),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance410402(.data_in(wire_d40_1),.data_out(wire_d40_2),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance410403(.data_in(wire_d40_2),.data_out(wire_d40_3),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance410404(.data_in(wire_d40_3),.data_out(wire_d40_4),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance410405(.data_in(wire_d40_4),.data_out(wire_d40_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance410406(.data_in(wire_d40_5),.data_out(wire_d40_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance410407(.data_in(wire_d40_6),.data_out(wire_d40_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance410408(.data_in(wire_d40_7),.data_out(wire_d40_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance410409(.data_in(wire_d40_8),.data_out(wire_d40_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104010(.data_in(wire_d40_9),.data_out(wire_d40_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104011(.data_in(wire_d40_10),.data_out(wire_d40_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4104012(.data_in(wire_d40_11),.data_out(wire_d40_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104013(.data_in(wire_d40_12),.data_out(wire_d40_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4104014(.data_in(wire_d40_13),.data_out(wire_d40_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104015(.data_in(wire_d40_14),.data_out(wire_d40_15),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4104016(.data_in(wire_d40_15),.data_out(wire_d40_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4104017(.data_in(wire_d40_16),.data_out(wire_d40_17),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104018(.data_in(wire_d40_17),.data_out(wire_d40_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4104019(.data_in(wire_d40_18),.data_out(wire_d40_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4104020(.data_in(wire_d40_19),.data_out(wire_d40_20),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4104021(.data_in(wire_d40_20),.data_out(wire_d40_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4104022(.data_in(wire_d40_21),.data_out(wire_d40_22),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4104023(.data_in(wire_d40_22),.data_out(wire_d40_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4104024(.data_in(wire_d40_23),.data_out(wire_d40_24),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104025(.data_in(wire_d40_24),.data_out(wire_d40_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104026(.data_in(wire_d40_25),.data_out(wire_d40_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4104027(.data_in(wire_d40_26),.data_out(wire_d40_27),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4104028(.data_in(wire_d40_27),.data_out(wire_d40_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104029(.data_in(wire_d40_28),.data_out(wire_d40_29),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104030(.data_in(wire_d40_29),.data_out(wire_d40_30),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104031(.data_in(wire_d40_30),.data_out(wire_d40_31),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104032(.data_in(wire_d40_31),.data_out(wire_d40_32),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4104033(.data_in(wire_d40_32),.data_out(wire_d40_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4104034(.data_in(wire_d40_33),.data_out(wire_d40_34),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104035(.data_in(wire_d40_34),.data_out(wire_d40_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4104036(.data_in(wire_d40_35),.data_out(wire_d40_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4104037(.data_in(wire_d40_36),.data_out(wire_d40_37),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4104038(.data_in(wire_d40_37),.data_out(wire_d40_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104039(.data_in(wire_d40_38),.data_out(wire_d40_39),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4104040(.data_in(wire_d40_39),.data_out(wire_d40_40),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4104041(.data_in(wire_d40_40),.data_out(wire_d40_41),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4104042(.data_in(wire_d40_41),.data_out(wire_d40_42),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4104043(.data_in(wire_d40_42),.data_out(wire_d40_43),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4104044(.data_in(wire_d40_43),.data_out(wire_d40_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4104045(.data_in(wire_d40_44),.data_out(wire_d40_45),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104046(.data_in(wire_d40_45),.data_out(wire_d40_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4104047(.data_in(wire_d40_46),.data_out(wire_d40_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4104048(.data_in(wire_d40_47),.data_out(wire_d40_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4104049(.data_in(wire_d40_48),.data_out(d_out40),.clk(clk),.rst(rst));

	large_adder #(.WIDTH(WIDTH)) large_adder_instance420410(.data_in(d_in41),.data_out(wire_d41_0),.clk(clk),.rst(rst));            //channel 42
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance420411(.data_in(wire_d41_0),.data_out(wire_d41_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance420412(.data_in(wire_d41_1),.data_out(wire_d41_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance420413(.data_in(wire_d41_2),.data_out(wire_d41_3),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance420414(.data_in(wire_d41_3),.data_out(wire_d41_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance420415(.data_in(wire_d41_4),.data_out(wire_d41_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance420416(.data_in(wire_d41_5),.data_out(wire_d41_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance420417(.data_in(wire_d41_6),.data_out(wire_d41_7),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance420418(.data_in(wire_d41_7),.data_out(wire_d41_8),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance420419(.data_in(wire_d41_8),.data_out(wire_d41_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204110(.data_in(wire_d41_9),.data_out(wire_d41_10),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204111(.data_in(wire_d41_10),.data_out(wire_d41_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4204112(.data_in(wire_d41_11),.data_out(wire_d41_12),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4204113(.data_in(wire_d41_12),.data_out(wire_d41_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4204114(.data_in(wire_d41_13),.data_out(wire_d41_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204115(.data_in(wire_d41_14),.data_out(wire_d41_15),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4204116(.data_in(wire_d41_15),.data_out(wire_d41_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204117(.data_in(wire_d41_16),.data_out(wire_d41_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4204118(.data_in(wire_d41_17),.data_out(wire_d41_18),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4204119(.data_in(wire_d41_18),.data_out(wire_d41_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4204120(.data_in(wire_d41_19),.data_out(wire_d41_20),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4204121(.data_in(wire_d41_20),.data_out(wire_d41_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204122(.data_in(wire_d41_21),.data_out(wire_d41_22),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4204123(.data_in(wire_d41_22),.data_out(wire_d41_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204124(.data_in(wire_d41_23),.data_out(wire_d41_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204125(.data_in(wire_d41_24),.data_out(wire_d41_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4204126(.data_in(wire_d41_25),.data_out(wire_d41_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4204127(.data_in(wire_d41_26),.data_out(wire_d41_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204128(.data_in(wire_d41_27),.data_out(wire_d41_28),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204129(.data_in(wire_d41_28),.data_out(wire_d41_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204130(.data_in(wire_d41_29),.data_out(wire_d41_30),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204131(.data_in(wire_d41_30),.data_out(wire_d41_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204132(.data_in(wire_d41_31),.data_out(wire_d41_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204133(.data_in(wire_d41_32),.data_out(wire_d41_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204134(.data_in(wire_d41_33),.data_out(wire_d41_34),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4204135(.data_in(wire_d41_34),.data_out(wire_d41_35),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4204136(.data_in(wire_d41_35),.data_out(wire_d41_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204137(.data_in(wire_d41_36),.data_out(wire_d41_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204138(.data_in(wire_d41_37),.data_out(wire_d41_38),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4204139(.data_in(wire_d41_38),.data_out(wire_d41_39),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4204140(.data_in(wire_d41_39),.data_out(wire_d41_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4204141(.data_in(wire_d41_40),.data_out(wire_d41_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4204142(.data_in(wire_d41_41),.data_out(wire_d41_42),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204143(.data_in(wire_d41_42),.data_out(wire_d41_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4204144(.data_in(wire_d41_43),.data_out(wire_d41_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4204145(.data_in(wire_d41_44),.data_out(wire_d41_45),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4204146(.data_in(wire_d41_45),.data_out(wire_d41_46),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4204147(.data_in(wire_d41_46),.data_out(wire_d41_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4204148(.data_in(wire_d41_47),.data_out(wire_d41_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4204149(.data_in(wire_d41_48),.data_out(d_out41),.clk(clk),.rst(rst));

	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance430420(.data_in(d_in42),.data_out(wire_d42_0),.clk(clk),.rst(rst));            //channel 43
	decoder_top #(.WIDTH(WIDTH)) decoder_instance430421(.data_in(wire_d42_0),.data_out(wire_d42_1),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance430422(.data_in(wire_d42_1),.data_out(wire_d42_2),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance430423(.data_in(wire_d42_2),.data_out(wire_d42_3),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance430424(.data_in(wire_d42_3),.data_out(wire_d42_4),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance430425(.data_in(wire_d42_4),.data_out(wire_d42_5),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance430426(.data_in(wire_d42_5),.data_out(wire_d42_6),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance430427(.data_in(wire_d42_6),.data_out(wire_d42_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance430428(.data_in(wire_d42_7),.data_out(wire_d42_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance430429(.data_in(wire_d42_8),.data_out(wire_d42_9),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304210(.data_in(wire_d42_9),.data_out(wire_d42_10),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4304211(.data_in(wire_d42_10),.data_out(wire_d42_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304212(.data_in(wire_d42_11),.data_out(wire_d42_12),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304213(.data_in(wire_d42_12),.data_out(wire_d42_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304214(.data_in(wire_d42_13),.data_out(wire_d42_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304215(.data_in(wire_d42_14),.data_out(wire_d42_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304216(.data_in(wire_d42_15),.data_out(wire_d42_16),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304217(.data_in(wire_d42_16),.data_out(wire_d42_17),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304218(.data_in(wire_d42_17),.data_out(wire_d42_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4304219(.data_in(wire_d42_18),.data_out(wire_d42_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304220(.data_in(wire_d42_19),.data_out(wire_d42_20),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4304221(.data_in(wire_d42_20),.data_out(wire_d42_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304222(.data_in(wire_d42_21),.data_out(wire_d42_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4304223(.data_in(wire_d42_22),.data_out(wire_d42_23),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4304224(.data_in(wire_d42_23),.data_out(wire_d42_24),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4304225(.data_in(wire_d42_24),.data_out(wire_d42_25),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304226(.data_in(wire_d42_25),.data_out(wire_d42_26),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304227(.data_in(wire_d42_26),.data_out(wire_d42_27),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304228(.data_in(wire_d42_27),.data_out(wire_d42_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4304229(.data_in(wire_d42_28),.data_out(wire_d42_29),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4304230(.data_in(wire_d42_29),.data_out(wire_d42_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304231(.data_in(wire_d42_30),.data_out(wire_d42_31),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304232(.data_in(wire_d42_31),.data_out(wire_d42_32),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4304233(.data_in(wire_d42_32),.data_out(wire_d42_33),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4304234(.data_in(wire_d42_33),.data_out(wire_d42_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304235(.data_in(wire_d42_34),.data_out(wire_d42_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304236(.data_in(wire_d42_35),.data_out(wire_d42_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4304237(.data_in(wire_d42_36),.data_out(wire_d42_37),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304238(.data_in(wire_d42_37),.data_out(wire_d42_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304239(.data_in(wire_d42_38),.data_out(wire_d42_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4304240(.data_in(wire_d42_39),.data_out(wire_d42_40),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304241(.data_in(wire_d42_40),.data_out(wire_d42_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4304242(.data_in(wire_d42_41),.data_out(wire_d42_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304243(.data_in(wire_d42_42),.data_out(wire_d42_43),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4304244(.data_in(wire_d42_43),.data_out(wire_d42_44),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4304245(.data_in(wire_d42_44),.data_out(wire_d42_45),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4304246(.data_in(wire_d42_45),.data_out(wire_d42_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4304247(.data_in(wire_d42_46),.data_out(wire_d42_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4304248(.data_in(wire_d42_47),.data_out(wire_d42_48),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4304249(.data_in(wire_d42_48),.data_out(d_out42),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance440430(.data_in(d_in43),.data_out(wire_d43_0),.clk(clk),.rst(rst));            //channel 44
	encoder #(.WIDTH(WIDTH)) encoder_instance440431(.data_in(wire_d43_0),.data_out(wire_d43_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance440432(.data_in(wire_d43_1),.data_out(wire_d43_2),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance440433(.data_in(wire_d43_2),.data_out(wire_d43_3),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance440434(.data_in(wire_d43_3),.data_out(wire_d43_4),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance440435(.data_in(wire_d43_4),.data_out(wire_d43_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance440436(.data_in(wire_d43_5),.data_out(wire_d43_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance440437(.data_in(wire_d43_6),.data_out(wire_d43_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance440438(.data_in(wire_d43_7),.data_out(wire_d43_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance440439(.data_in(wire_d43_8),.data_out(wire_d43_9),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4404310(.data_in(wire_d43_9),.data_out(wire_d43_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404311(.data_in(wire_d43_10),.data_out(wire_d43_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404312(.data_in(wire_d43_11),.data_out(wire_d43_12),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4404313(.data_in(wire_d43_12),.data_out(wire_d43_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404314(.data_in(wire_d43_13),.data_out(wire_d43_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4404315(.data_in(wire_d43_14),.data_out(wire_d43_15),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404316(.data_in(wire_d43_15),.data_out(wire_d43_16),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4404317(.data_in(wire_d43_16),.data_out(wire_d43_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4404318(.data_in(wire_d43_17),.data_out(wire_d43_18),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4404319(.data_in(wire_d43_18),.data_out(wire_d43_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404320(.data_in(wire_d43_19),.data_out(wire_d43_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404321(.data_in(wire_d43_20),.data_out(wire_d43_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404322(.data_in(wire_d43_21),.data_out(wire_d43_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404323(.data_in(wire_d43_22),.data_out(wire_d43_23),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404324(.data_in(wire_d43_23),.data_out(wire_d43_24),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404325(.data_in(wire_d43_24),.data_out(wire_d43_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404326(.data_in(wire_d43_25),.data_out(wire_d43_26),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404327(.data_in(wire_d43_26),.data_out(wire_d43_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4404328(.data_in(wire_d43_27),.data_out(wire_d43_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4404329(.data_in(wire_d43_28),.data_out(wire_d43_29),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404330(.data_in(wire_d43_29),.data_out(wire_d43_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4404331(.data_in(wire_d43_30),.data_out(wire_d43_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4404332(.data_in(wire_d43_31),.data_out(wire_d43_32),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4404333(.data_in(wire_d43_32),.data_out(wire_d43_33),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4404334(.data_in(wire_d43_33),.data_out(wire_d43_34),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404335(.data_in(wire_d43_34),.data_out(wire_d43_35),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404336(.data_in(wire_d43_35),.data_out(wire_d43_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4404337(.data_in(wire_d43_36),.data_out(wire_d43_37),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4404338(.data_in(wire_d43_37),.data_out(wire_d43_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404339(.data_in(wire_d43_38),.data_out(wire_d43_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404340(.data_in(wire_d43_39),.data_out(wire_d43_40),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4404341(.data_in(wire_d43_40),.data_out(wire_d43_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4404342(.data_in(wire_d43_41),.data_out(wire_d43_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4404343(.data_in(wire_d43_42),.data_out(wire_d43_43),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4404344(.data_in(wire_d43_43),.data_out(wire_d43_44),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4404345(.data_in(wire_d43_44),.data_out(wire_d43_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4404346(.data_in(wire_d43_45),.data_out(wire_d43_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4404347(.data_in(wire_d43_46),.data_out(wire_d43_47),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4404348(.data_in(wire_d43_47),.data_out(wire_d43_48),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4404349(.data_in(wire_d43_48),.data_out(d_out43),.clk(clk),.rst(rst));

	decoder_top #(.WIDTH(WIDTH)) decoder_instance450440(.data_in(d_in44),.data_out(wire_d44_0),.clk(clk),.rst(rst));            //channel 45
	large_mux #(.WIDTH(WIDTH)) large_mux_instance450441(.data_in(wire_d44_0),.data_out(wire_d44_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance450442(.data_in(wire_d44_1),.data_out(wire_d44_2),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance450443(.data_in(wire_d44_2),.data_out(wire_d44_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance450444(.data_in(wire_d44_3),.data_out(wire_d44_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance450445(.data_in(wire_d44_4),.data_out(wire_d44_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance450446(.data_in(wire_d44_5),.data_out(wire_d44_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance450447(.data_in(wire_d44_6),.data_out(wire_d44_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance450448(.data_in(wire_d44_7),.data_out(wire_d44_8),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance450449(.data_in(wire_d44_8),.data_out(wire_d44_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504410(.data_in(wire_d44_9),.data_out(wire_d44_10),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504411(.data_in(wire_d44_10),.data_out(wire_d44_11),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504412(.data_in(wire_d44_11),.data_out(wire_d44_12),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4504413(.data_in(wire_d44_12),.data_out(wire_d44_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504414(.data_in(wire_d44_13),.data_out(wire_d44_14),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504415(.data_in(wire_d44_14),.data_out(wire_d44_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4504416(.data_in(wire_d44_15),.data_out(wire_d44_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4504417(.data_in(wire_d44_16),.data_out(wire_d44_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4504418(.data_in(wire_d44_17),.data_out(wire_d44_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4504419(.data_in(wire_d44_18),.data_out(wire_d44_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4504420(.data_in(wire_d44_19),.data_out(wire_d44_20),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4504421(.data_in(wire_d44_20),.data_out(wire_d44_21),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4504422(.data_in(wire_d44_21),.data_out(wire_d44_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504423(.data_in(wire_d44_22),.data_out(wire_d44_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504424(.data_in(wire_d44_23),.data_out(wire_d44_24),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4504425(.data_in(wire_d44_24),.data_out(wire_d44_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4504426(.data_in(wire_d44_25),.data_out(wire_d44_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504427(.data_in(wire_d44_26),.data_out(wire_d44_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504428(.data_in(wire_d44_27),.data_out(wire_d44_28),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4504429(.data_in(wire_d44_28),.data_out(wire_d44_29),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4504430(.data_in(wire_d44_29),.data_out(wire_d44_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4504431(.data_in(wire_d44_30),.data_out(wire_d44_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504432(.data_in(wire_d44_31),.data_out(wire_d44_32),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504433(.data_in(wire_d44_32),.data_out(wire_d44_33),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4504434(.data_in(wire_d44_33),.data_out(wire_d44_34),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504435(.data_in(wire_d44_34),.data_out(wire_d44_35),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4504436(.data_in(wire_d44_35),.data_out(wire_d44_36),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4504437(.data_in(wire_d44_36),.data_out(wire_d44_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504438(.data_in(wire_d44_37),.data_out(wire_d44_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4504439(.data_in(wire_d44_38),.data_out(wire_d44_39),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504440(.data_in(wire_d44_39),.data_out(wire_d44_40),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4504441(.data_in(wire_d44_40),.data_out(wire_d44_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4504442(.data_in(wire_d44_41),.data_out(wire_d44_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4504443(.data_in(wire_d44_42),.data_out(wire_d44_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4504444(.data_in(wire_d44_43),.data_out(wire_d44_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4504445(.data_in(wire_d44_44),.data_out(wire_d44_45),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4504446(.data_in(wire_d44_45),.data_out(wire_d44_46),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4504447(.data_in(wire_d44_46),.data_out(wire_d44_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4504448(.data_in(wire_d44_47),.data_out(wire_d44_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4504449(.data_in(wire_d44_48),.data_out(d_out44),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance460450(.data_in(d_in45),.data_out(wire_d45_0),.clk(clk),.rst(rst));            //channel 46
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance460451(.data_in(wire_d45_0),.data_out(wire_d45_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance460452(.data_in(wire_d45_1),.data_out(wire_d45_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance460453(.data_in(wire_d45_2),.data_out(wire_d45_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance460454(.data_in(wire_d45_3),.data_out(wire_d45_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance460455(.data_in(wire_d45_4),.data_out(wire_d45_5),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance460456(.data_in(wire_d45_5),.data_out(wire_d45_6),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance460457(.data_in(wire_d45_6),.data_out(wire_d45_7),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance460458(.data_in(wire_d45_7),.data_out(wire_d45_8),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance460459(.data_in(wire_d45_8),.data_out(wire_d45_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4604510(.data_in(wire_d45_9),.data_out(wire_d45_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604511(.data_in(wire_d45_10),.data_out(wire_d45_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604512(.data_in(wire_d45_11),.data_out(wire_d45_12),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4604513(.data_in(wire_d45_12),.data_out(wire_d45_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604514(.data_in(wire_d45_13),.data_out(wire_d45_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4604515(.data_in(wire_d45_14),.data_out(wire_d45_15),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4604516(.data_in(wire_d45_15),.data_out(wire_d45_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4604517(.data_in(wire_d45_16),.data_out(wire_d45_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604518(.data_in(wire_d45_17),.data_out(wire_d45_18),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4604519(.data_in(wire_d45_18),.data_out(wire_d45_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604520(.data_in(wire_d45_19),.data_out(wire_d45_20),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4604521(.data_in(wire_d45_20),.data_out(wire_d45_21),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604522(.data_in(wire_d45_21),.data_out(wire_d45_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4604523(.data_in(wire_d45_22),.data_out(wire_d45_23),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604524(.data_in(wire_d45_23),.data_out(wire_d45_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4604525(.data_in(wire_d45_24),.data_out(wire_d45_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4604526(.data_in(wire_d45_25),.data_out(wire_d45_26),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604527(.data_in(wire_d45_26),.data_out(wire_d45_27),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4604528(.data_in(wire_d45_27),.data_out(wire_d45_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604529(.data_in(wire_d45_28),.data_out(wire_d45_29),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604530(.data_in(wire_d45_29),.data_out(wire_d45_30),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604531(.data_in(wire_d45_30),.data_out(wire_d45_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4604532(.data_in(wire_d45_31),.data_out(wire_d45_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4604533(.data_in(wire_d45_32),.data_out(wire_d45_33),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4604534(.data_in(wire_d45_33),.data_out(wire_d45_34),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604535(.data_in(wire_d45_34),.data_out(wire_d45_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4604536(.data_in(wire_d45_35),.data_out(wire_d45_36),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604537(.data_in(wire_d45_36),.data_out(wire_d45_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4604538(.data_in(wire_d45_37),.data_out(wire_d45_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4604539(.data_in(wire_d45_38),.data_out(wire_d45_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4604540(.data_in(wire_d45_39),.data_out(wire_d45_40),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4604541(.data_in(wire_d45_40),.data_out(wire_d45_41),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4604542(.data_in(wire_d45_41),.data_out(wire_d45_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4604543(.data_in(wire_d45_42),.data_out(wire_d45_43),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4604544(.data_in(wire_d45_43),.data_out(wire_d45_44),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4604545(.data_in(wire_d45_44),.data_out(wire_d45_45),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4604546(.data_in(wire_d45_45),.data_out(wire_d45_46),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4604547(.data_in(wire_d45_46),.data_out(wire_d45_47),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4604548(.data_in(wire_d45_47),.data_out(wire_d45_48),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4604549(.data_in(wire_d45_48),.data_out(d_out45),.clk(clk),.rst(rst));

	invertion #(.WIDTH(WIDTH)) invertion_instance470460(.data_in(d_in46),.data_out(wire_d46_0),.clk(clk),.rst(rst));            //channel 47
	large_mux #(.WIDTH(WIDTH)) large_mux_instance470461(.data_in(wire_d46_0),.data_out(wire_d46_1),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance470462(.data_in(wire_d46_1),.data_out(wire_d46_2),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance470463(.data_in(wire_d46_2),.data_out(wire_d46_3),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance470464(.data_in(wire_d46_3),.data_out(wire_d46_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance470465(.data_in(wire_d46_4),.data_out(wire_d46_5),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance470466(.data_in(wire_d46_5),.data_out(wire_d46_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance470467(.data_in(wire_d46_6),.data_out(wire_d46_7),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance470468(.data_in(wire_d46_7),.data_out(wire_d46_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance470469(.data_in(wire_d46_8),.data_out(wire_d46_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704610(.data_in(wire_d46_9),.data_out(wire_d46_10),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4704611(.data_in(wire_d46_10),.data_out(wire_d46_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704612(.data_in(wire_d46_11),.data_out(wire_d46_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704613(.data_in(wire_d46_12),.data_out(wire_d46_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4704614(.data_in(wire_d46_13),.data_out(wire_d46_14),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704615(.data_in(wire_d46_14),.data_out(wire_d46_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704616(.data_in(wire_d46_15),.data_out(wire_d46_16),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4704617(.data_in(wire_d46_16),.data_out(wire_d46_17),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704618(.data_in(wire_d46_17),.data_out(wire_d46_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4704619(.data_in(wire_d46_18),.data_out(wire_d46_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704620(.data_in(wire_d46_19),.data_out(wire_d46_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704621(.data_in(wire_d46_20),.data_out(wire_d46_21),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4704622(.data_in(wire_d46_21),.data_out(wire_d46_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4704623(.data_in(wire_d46_22),.data_out(wire_d46_23),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704624(.data_in(wire_d46_23),.data_out(wire_d46_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4704625(.data_in(wire_d46_24),.data_out(wire_d46_25),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704626(.data_in(wire_d46_25),.data_out(wire_d46_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4704627(.data_in(wire_d46_26),.data_out(wire_d46_27),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4704628(.data_in(wire_d46_27),.data_out(wire_d46_28),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704629(.data_in(wire_d46_28),.data_out(wire_d46_29),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704630(.data_in(wire_d46_29),.data_out(wire_d46_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4704631(.data_in(wire_d46_30),.data_out(wire_d46_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704632(.data_in(wire_d46_31),.data_out(wire_d46_32),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4704633(.data_in(wire_d46_32),.data_out(wire_d46_33),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4704634(.data_in(wire_d46_33),.data_out(wire_d46_34),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4704635(.data_in(wire_d46_34),.data_out(wire_d46_35),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704636(.data_in(wire_d46_35),.data_out(wire_d46_36),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704637(.data_in(wire_d46_36),.data_out(wire_d46_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704638(.data_in(wire_d46_37),.data_out(wire_d46_38),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4704639(.data_in(wire_d46_38),.data_out(wire_d46_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4704640(.data_in(wire_d46_39),.data_out(wire_d46_40),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4704641(.data_in(wire_d46_40),.data_out(wire_d46_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4704642(.data_in(wire_d46_41),.data_out(wire_d46_42),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704643(.data_in(wire_d46_42),.data_out(wire_d46_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704644(.data_in(wire_d46_43),.data_out(wire_d46_44),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4704645(.data_in(wire_d46_44),.data_out(wire_d46_45),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4704646(.data_in(wire_d46_45),.data_out(wire_d46_46),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4704647(.data_in(wire_d46_46),.data_out(wire_d46_47),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704648(.data_in(wire_d46_47),.data_out(wire_d46_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4704649(.data_in(wire_d46_48),.data_out(d_out46),.clk(clk),.rst(rst));

	large_mux #(.WIDTH(WIDTH)) large_mux_instance480470(.data_in(d_in47),.data_out(wire_d47_0),.clk(clk),.rst(rst));            //channel 48
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance480471(.data_in(wire_d47_0),.data_out(wire_d47_1),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance480472(.data_in(wire_d47_1),.data_out(wire_d47_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance480473(.data_in(wire_d47_2),.data_out(wire_d47_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance480474(.data_in(wire_d47_3),.data_out(wire_d47_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance480475(.data_in(wire_d47_4),.data_out(wire_d47_5),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance480476(.data_in(wire_d47_5),.data_out(wire_d47_6),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance480477(.data_in(wire_d47_6),.data_out(wire_d47_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance480478(.data_in(wire_d47_7),.data_out(wire_d47_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance480479(.data_in(wire_d47_8),.data_out(wire_d47_9),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4804710(.data_in(wire_d47_9),.data_out(wire_d47_10),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4804711(.data_in(wire_d47_10),.data_out(wire_d47_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804712(.data_in(wire_d47_11),.data_out(wire_d47_12),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804713(.data_in(wire_d47_12),.data_out(wire_d47_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804714(.data_in(wire_d47_13),.data_out(wire_d47_14),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804715(.data_in(wire_d47_14),.data_out(wire_d47_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4804716(.data_in(wire_d47_15),.data_out(wire_d47_16),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804717(.data_in(wire_d47_16),.data_out(wire_d47_17),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4804718(.data_in(wire_d47_17),.data_out(wire_d47_18),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804719(.data_in(wire_d47_18),.data_out(wire_d47_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4804720(.data_in(wire_d47_19),.data_out(wire_d47_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4804721(.data_in(wire_d47_20),.data_out(wire_d47_21),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4804722(.data_in(wire_d47_21),.data_out(wire_d47_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804723(.data_in(wire_d47_22),.data_out(wire_d47_23),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4804724(.data_in(wire_d47_23),.data_out(wire_d47_24),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804725(.data_in(wire_d47_24),.data_out(wire_d47_25),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804726(.data_in(wire_d47_25),.data_out(wire_d47_26),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4804727(.data_in(wire_d47_26),.data_out(wire_d47_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804728(.data_in(wire_d47_27),.data_out(wire_d47_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4804729(.data_in(wire_d47_28),.data_out(wire_d47_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4804730(.data_in(wire_d47_29),.data_out(wire_d47_30),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804731(.data_in(wire_d47_30),.data_out(wire_d47_31),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4804732(.data_in(wire_d47_31),.data_out(wire_d47_32),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4804733(.data_in(wire_d47_32),.data_out(wire_d47_33),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804734(.data_in(wire_d47_33),.data_out(wire_d47_34),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4804735(.data_in(wire_d47_34),.data_out(wire_d47_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4804736(.data_in(wire_d47_35),.data_out(wire_d47_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4804737(.data_in(wire_d47_36),.data_out(wire_d47_37),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804738(.data_in(wire_d47_37),.data_out(wire_d47_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804739(.data_in(wire_d47_38),.data_out(wire_d47_39),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804740(.data_in(wire_d47_39),.data_out(wire_d47_40),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4804741(.data_in(wire_d47_40),.data_out(wire_d47_41),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804742(.data_in(wire_d47_41),.data_out(wire_d47_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4804743(.data_in(wire_d47_42),.data_out(wire_d47_43),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804744(.data_in(wire_d47_43),.data_out(wire_d47_44),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4804745(.data_in(wire_d47_44),.data_out(wire_d47_45),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4804746(.data_in(wire_d47_45),.data_out(wire_d47_46),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4804747(.data_in(wire_d47_46),.data_out(wire_d47_47),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4804748(.data_in(wire_d47_47),.data_out(wire_d47_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4804749(.data_in(wire_d47_48),.data_out(d_out47),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance490480(.data_in(d_in48),.data_out(wire_d48_0),.clk(clk),.rst(rst));            //channel 49
	large_mux #(.WIDTH(WIDTH)) large_mux_instance490481(.data_in(wire_d48_0),.data_out(wire_d48_1),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance490482(.data_in(wire_d48_1),.data_out(wire_d48_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance490483(.data_in(wire_d48_2),.data_out(wire_d48_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance490484(.data_in(wire_d48_3),.data_out(wire_d48_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance490485(.data_in(wire_d48_4),.data_out(wire_d48_5),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance490486(.data_in(wire_d48_5),.data_out(wire_d48_6),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance490487(.data_in(wire_d48_6),.data_out(wire_d48_7),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance490488(.data_in(wire_d48_7),.data_out(wire_d48_8),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance490489(.data_in(wire_d48_8),.data_out(wire_d48_9),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4904810(.data_in(wire_d48_9),.data_out(wire_d48_10),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904811(.data_in(wire_d48_10),.data_out(wire_d48_11),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4904812(.data_in(wire_d48_11),.data_out(wire_d48_12),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904813(.data_in(wire_d48_12),.data_out(wire_d48_13),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904814(.data_in(wire_d48_13),.data_out(wire_d48_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4904815(.data_in(wire_d48_14),.data_out(wire_d48_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904816(.data_in(wire_d48_15),.data_out(wire_d48_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904817(.data_in(wire_d48_16),.data_out(wire_d48_17),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904818(.data_in(wire_d48_17),.data_out(wire_d48_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904819(.data_in(wire_d48_18),.data_out(wire_d48_19),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4904820(.data_in(wire_d48_19),.data_out(wire_d48_20),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4904821(.data_in(wire_d48_20),.data_out(wire_d48_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904822(.data_in(wire_d48_21),.data_out(wire_d48_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904823(.data_in(wire_d48_22),.data_out(wire_d48_23),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904824(.data_in(wire_d48_23),.data_out(wire_d48_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4904825(.data_in(wire_d48_24),.data_out(wire_d48_25),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4904826(.data_in(wire_d48_25),.data_out(wire_d48_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904827(.data_in(wire_d48_26),.data_out(wire_d48_27),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance4904828(.data_in(wire_d48_27),.data_out(wire_d48_28),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904829(.data_in(wire_d48_28),.data_out(wire_d48_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance4904830(.data_in(wire_d48_29),.data_out(wire_d48_30),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4904831(.data_in(wire_d48_30),.data_out(wire_d48_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904832(.data_in(wire_d48_31),.data_out(wire_d48_32),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904833(.data_in(wire_d48_32),.data_out(wire_d48_33),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance4904834(.data_in(wire_d48_33),.data_out(wire_d48_34),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4904835(.data_in(wire_d48_34),.data_out(wire_d48_35),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4904836(.data_in(wire_d48_35),.data_out(wire_d48_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904837(.data_in(wire_d48_36),.data_out(wire_d48_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance4904838(.data_in(wire_d48_37),.data_out(wire_d48_38),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4904839(.data_in(wire_d48_38),.data_out(wire_d48_39),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance4904840(.data_in(wire_d48_39),.data_out(wire_d48_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance4904841(.data_in(wire_d48_40),.data_out(wire_d48_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance4904842(.data_in(wire_d48_41),.data_out(wire_d48_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance4904843(.data_in(wire_d48_42),.data_out(wire_d48_43),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance4904844(.data_in(wire_d48_43),.data_out(wire_d48_44),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4904845(.data_in(wire_d48_44),.data_out(wire_d48_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4904846(.data_in(wire_d48_45),.data_out(wire_d48_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance4904847(.data_in(wire_d48_46),.data_out(wire_d48_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance4904848(.data_in(wire_d48_47),.data_out(wire_d48_48),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance4904849(.data_in(wire_d48_48),.data_out(d_out48),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance500490(.data_in(d_in49),.data_out(wire_d49_0),.clk(clk),.rst(rst));            //channel 50
	large_adder #(.WIDTH(WIDTH)) large_adder_instance500491(.data_in(wire_d49_0),.data_out(wire_d49_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance500492(.data_in(wire_d49_1),.data_out(wire_d49_2),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance500493(.data_in(wire_d49_2),.data_out(wire_d49_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance500494(.data_in(wire_d49_3),.data_out(wire_d49_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance500495(.data_in(wire_d49_4),.data_out(wire_d49_5),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance500496(.data_in(wire_d49_5),.data_out(wire_d49_6),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance500497(.data_in(wire_d49_6),.data_out(wire_d49_7),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance500498(.data_in(wire_d49_7),.data_out(wire_d49_8),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance500499(.data_in(wire_d49_8),.data_out(wire_d49_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004910(.data_in(wire_d49_9),.data_out(wire_d49_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004911(.data_in(wire_d49_10),.data_out(wire_d49_11),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004912(.data_in(wire_d49_11),.data_out(wire_d49_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004913(.data_in(wire_d49_12),.data_out(wire_d49_13),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004914(.data_in(wire_d49_13),.data_out(wire_d49_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004915(.data_in(wire_d49_14),.data_out(wire_d49_15),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004916(.data_in(wire_d49_15),.data_out(wire_d49_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5004917(.data_in(wire_d49_16),.data_out(wire_d49_17),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5004918(.data_in(wire_d49_17),.data_out(wire_d49_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004919(.data_in(wire_d49_18),.data_out(wire_d49_19),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5004920(.data_in(wire_d49_19),.data_out(wire_d49_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004921(.data_in(wire_d49_20),.data_out(wire_d49_21),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004922(.data_in(wire_d49_21),.data_out(wire_d49_22),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004923(.data_in(wire_d49_22),.data_out(wire_d49_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004924(.data_in(wire_d49_23),.data_out(wire_d49_24),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004925(.data_in(wire_d49_24),.data_out(wire_d49_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5004926(.data_in(wire_d49_25),.data_out(wire_d49_26),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004927(.data_in(wire_d49_26),.data_out(wire_d49_27),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5004928(.data_in(wire_d49_27),.data_out(wire_d49_28),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5004929(.data_in(wire_d49_28),.data_out(wire_d49_29),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5004930(.data_in(wire_d49_29),.data_out(wire_d49_30),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5004931(.data_in(wire_d49_30),.data_out(wire_d49_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004932(.data_in(wire_d49_31),.data_out(wire_d49_32),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004933(.data_in(wire_d49_32),.data_out(wire_d49_33),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004934(.data_in(wire_d49_33),.data_out(wire_d49_34),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004935(.data_in(wire_d49_34),.data_out(wire_d49_35),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5004936(.data_in(wire_d49_35),.data_out(wire_d49_36),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004937(.data_in(wire_d49_36),.data_out(wire_d49_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5004938(.data_in(wire_d49_37),.data_out(wire_d49_38),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004939(.data_in(wire_d49_38),.data_out(wire_d49_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5004940(.data_in(wire_d49_39),.data_out(wire_d49_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5004941(.data_in(wire_d49_40),.data_out(wire_d49_41),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5004942(.data_in(wire_d49_41),.data_out(wire_d49_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5004943(.data_in(wire_d49_42),.data_out(wire_d49_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5004944(.data_in(wire_d49_43),.data_out(wire_d49_44),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5004945(.data_in(wire_d49_44),.data_out(wire_d49_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004946(.data_in(wire_d49_45),.data_out(wire_d49_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5004947(.data_in(wire_d49_46),.data_out(wire_d49_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5004948(.data_in(wire_d49_47),.data_out(wire_d49_48),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5004949(.data_in(wire_d49_48),.data_out(d_out49),.clk(clk),.rst(rst));

	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance510500(.data_in(d_in50),.data_out(wire_d50_0),.clk(clk),.rst(rst));            //channel 51
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance510501(.data_in(wire_d50_0),.data_out(wire_d50_1),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance510502(.data_in(wire_d50_1),.data_out(wire_d50_2),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance510503(.data_in(wire_d50_2),.data_out(wire_d50_3),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance510504(.data_in(wire_d50_3),.data_out(wire_d50_4),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance510505(.data_in(wire_d50_4),.data_out(wire_d50_5),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance510506(.data_in(wire_d50_5),.data_out(wire_d50_6),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance510507(.data_in(wire_d50_6),.data_out(wire_d50_7),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance510508(.data_in(wire_d50_7),.data_out(wire_d50_8),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance510509(.data_in(wire_d50_8),.data_out(wire_d50_9),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5105010(.data_in(wire_d50_9),.data_out(wire_d50_10),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105011(.data_in(wire_d50_10),.data_out(wire_d50_11),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105012(.data_in(wire_d50_11),.data_out(wire_d50_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5105013(.data_in(wire_d50_12),.data_out(wire_d50_13),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5105014(.data_in(wire_d50_13),.data_out(wire_d50_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105015(.data_in(wire_d50_14),.data_out(wire_d50_15),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105016(.data_in(wire_d50_15),.data_out(wire_d50_16),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5105017(.data_in(wire_d50_16),.data_out(wire_d50_17),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105018(.data_in(wire_d50_17),.data_out(wire_d50_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105019(.data_in(wire_d50_18),.data_out(wire_d50_19),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105020(.data_in(wire_d50_19),.data_out(wire_d50_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5105021(.data_in(wire_d50_20),.data_out(wire_d50_21),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5105022(.data_in(wire_d50_21),.data_out(wire_d50_22),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105023(.data_in(wire_d50_22),.data_out(wire_d50_23),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5105024(.data_in(wire_d50_23),.data_out(wire_d50_24),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105025(.data_in(wire_d50_24),.data_out(wire_d50_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5105026(.data_in(wire_d50_25),.data_out(wire_d50_26),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5105027(.data_in(wire_d50_26),.data_out(wire_d50_27),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5105028(.data_in(wire_d50_27),.data_out(wire_d50_28),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105029(.data_in(wire_d50_28),.data_out(wire_d50_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105030(.data_in(wire_d50_29),.data_out(wire_d50_30),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5105031(.data_in(wire_d50_30),.data_out(wire_d50_31),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5105032(.data_in(wire_d50_31),.data_out(wire_d50_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105033(.data_in(wire_d50_32),.data_out(wire_d50_33),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5105034(.data_in(wire_d50_33),.data_out(wire_d50_34),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5105035(.data_in(wire_d50_34),.data_out(wire_d50_35),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5105036(.data_in(wire_d50_35),.data_out(wire_d50_36),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105037(.data_in(wire_d50_36),.data_out(wire_d50_37),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5105038(.data_in(wire_d50_37),.data_out(wire_d50_38),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105039(.data_in(wire_d50_38),.data_out(wire_d50_39),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5105040(.data_in(wire_d50_39),.data_out(wire_d50_40),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5105041(.data_in(wire_d50_40),.data_out(wire_d50_41),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5105042(.data_in(wire_d50_41),.data_out(wire_d50_42),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5105043(.data_in(wire_d50_42),.data_out(wire_d50_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5105044(.data_in(wire_d50_43),.data_out(wire_d50_44),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5105045(.data_in(wire_d50_44),.data_out(wire_d50_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5105046(.data_in(wire_d50_45),.data_out(wire_d50_46),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5105047(.data_in(wire_d50_46),.data_out(wire_d50_47),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5105048(.data_in(wire_d50_47),.data_out(wire_d50_48),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5105049(.data_in(wire_d50_48),.data_out(d_out50),.clk(clk),.rst(rst));

	register #(.WIDTH(WIDTH)) register_instance520510(.data_in(d_in51),.data_out(wire_d51_0),.clk(clk),.rst(rst));            //channel 52
	decoder_top #(.WIDTH(WIDTH)) decoder_instance520511(.data_in(wire_d51_0),.data_out(wire_d51_1),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance520512(.data_in(wire_d51_1),.data_out(wire_d51_2),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance520513(.data_in(wire_d51_2),.data_out(wire_d51_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance520514(.data_in(wire_d51_3),.data_out(wire_d51_4),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance520515(.data_in(wire_d51_4),.data_out(wire_d51_5),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance520516(.data_in(wire_d51_5),.data_out(wire_d51_6),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance520517(.data_in(wire_d51_6),.data_out(wire_d51_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance520518(.data_in(wire_d51_7),.data_out(wire_d51_8),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance520519(.data_in(wire_d51_8),.data_out(wire_d51_9),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205110(.data_in(wire_d51_9),.data_out(wire_d51_10),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5205111(.data_in(wire_d51_10),.data_out(wire_d51_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5205112(.data_in(wire_d51_11),.data_out(wire_d51_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205113(.data_in(wire_d51_12),.data_out(wire_d51_13),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5205114(.data_in(wire_d51_13),.data_out(wire_d51_14),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205115(.data_in(wire_d51_14),.data_out(wire_d51_15),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205116(.data_in(wire_d51_15),.data_out(wire_d51_16),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205117(.data_in(wire_d51_16),.data_out(wire_d51_17),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205118(.data_in(wire_d51_17),.data_out(wire_d51_18),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5205119(.data_in(wire_d51_18),.data_out(wire_d51_19),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205120(.data_in(wire_d51_19),.data_out(wire_d51_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5205121(.data_in(wire_d51_20),.data_out(wire_d51_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5205122(.data_in(wire_d51_21),.data_out(wire_d51_22),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5205123(.data_in(wire_d51_22),.data_out(wire_d51_23),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5205124(.data_in(wire_d51_23),.data_out(wire_d51_24),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5205125(.data_in(wire_d51_24),.data_out(wire_d51_25),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205126(.data_in(wire_d51_25),.data_out(wire_d51_26),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5205127(.data_in(wire_d51_26),.data_out(wire_d51_27),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5205128(.data_in(wire_d51_27),.data_out(wire_d51_28),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5205129(.data_in(wire_d51_28),.data_out(wire_d51_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5205130(.data_in(wire_d51_29),.data_out(wire_d51_30),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205131(.data_in(wire_d51_30),.data_out(wire_d51_31),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5205132(.data_in(wire_d51_31),.data_out(wire_d51_32),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205133(.data_in(wire_d51_32),.data_out(wire_d51_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5205134(.data_in(wire_d51_33),.data_out(wire_d51_34),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5205135(.data_in(wire_d51_34),.data_out(wire_d51_35),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5205136(.data_in(wire_d51_35),.data_out(wire_d51_36),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5205137(.data_in(wire_d51_36),.data_out(wire_d51_37),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205138(.data_in(wire_d51_37),.data_out(wire_d51_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5205139(.data_in(wire_d51_38),.data_out(wire_d51_39),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5205140(.data_in(wire_d51_39),.data_out(wire_d51_40),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5205141(.data_in(wire_d51_40),.data_out(wire_d51_41),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5205142(.data_in(wire_d51_41),.data_out(wire_d51_42),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205143(.data_in(wire_d51_42),.data_out(wire_d51_43),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205144(.data_in(wire_d51_43),.data_out(wire_d51_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205145(.data_in(wire_d51_44),.data_out(wire_d51_45),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5205146(.data_in(wire_d51_45),.data_out(wire_d51_46),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5205147(.data_in(wire_d51_46),.data_out(wire_d51_47),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5205148(.data_in(wire_d51_47),.data_out(wire_d51_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5205149(.data_in(wire_d51_48),.data_out(d_out51),.clk(clk),.rst(rst));

	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance530520(.data_in(d_in52),.data_out(wire_d52_0),.clk(clk),.rst(rst));            //channel 53
	decoder_top #(.WIDTH(WIDTH)) decoder_instance530521(.data_in(wire_d52_0),.data_out(wire_d52_1),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance530522(.data_in(wire_d52_1),.data_out(wire_d52_2),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance530523(.data_in(wire_d52_2),.data_out(wire_d52_3),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance530524(.data_in(wire_d52_3),.data_out(wire_d52_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance530525(.data_in(wire_d52_4),.data_out(wire_d52_5),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance530526(.data_in(wire_d52_5),.data_out(wire_d52_6),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance530527(.data_in(wire_d52_6),.data_out(wire_d52_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance530528(.data_in(wire_d52_7),.data_out(wire_d52_8),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance530529(.data_in(wire_d52_8),.data_out(wire_d52_9),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5305210(.data_in(wire_d52_9),.data_out(wire_d52_10),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305211(.data_in(wire_d52_10),.data_out(wire_d52_11),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5305212(.data_in(wire_d52_11),.data_out(wire_d52_12),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305213(.data_in(wire_d52_12),.data_out(wire_d52_13),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305214(.data_in(wire_d52_13),.data_out(wire_d52_14),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305215(.data_in(wire_d52_14),.data_out(wire_d52_15),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5305216(.data_in(wire_d52_15),.data_out(wire_d52_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305217(.data_in(wire_d52_16),.data_out(wire_d52_17),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305218(.data_in(wire_d52_17),.data_out(wire_d52_18),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5305219(.data_in(wire_d52_18),.data_out(wire_d52_19),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5305220(.data_in(wire_d52_19),.data_out(wire_d52_20),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305221(.data_in(wire_d52_20),.data_out(wire_d52_21),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305222(.data_in(wire_d52_21),.data_out(wire_d52_22),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5305223(.data_in(wire_d52_22),.data_out(wire_d52_23),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305224(.data_in(wire_d52_23),.data_out(wire_d52_24),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5305225(.data_in(wire_d52_24),.data_out(wire_d52_25),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5305226(.data_in(wire_d52_25),.data_out(wire_d52_26),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5305227(.data_in(wire_d52_26),.data_out(wire_d52_27),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5305228(.data_in(wire_d52_27),.data_out(wire_d52_28),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305229(.data_in(wire_d52_28),.data_out(wire_d52_29),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305230(.data_in(wire_d52_29),.data_out(wire_d52_30),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5305231(.data_in(wire_d52_30),.data_out(wire_d52_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305232(.data_in(wire_d52_31),.data_out(wire_d52_32),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5305233(.data_in(wire_d52_32),.data_out(wire_d52_33),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305234(.data_in(wire_d52_33),.data_out(wire_d52_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305235(.data_in(wire_d52_34),.data_out(wire_d52_35),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5305236(.data_in(wire_d52_35),.data_out(wire_d52_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5305237(.data_in(wire_d52_36),.data_out(wire_d52_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305238(.data_in(wire_d52_37),.data_out(wire_d52_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305239(.data_in(wire_d52_38),.data_out(wire_d52_39),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305240(.data_in(wire_d52_39),.data_out(wire_d52_40),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305241(.data_in(wire_d52_40),.data_out(wire_d52_41),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5305242(.data_in(wire_d52_41),.data_out(wire_d52_42),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305243(.data_in(wire_d52_42),.data_out(wire_d52_43),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5305244(.data_in(wire_d52_43),.data_out(wire_d52_44),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5305245(.data_in(wire_d52_44),.data_out(wire_d52_45),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5305246(.data_in(wire_d52_45),.data_out(wire_d52_46),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5305247(.data_in(wire_d52_46),.data_out(wire_d52_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5305248(.data_in(wire_d52_47),.data_out(wire_d52_48),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5305249(.data_in(wire_d52_48),.data_out(d_out52),.clk(clk),.rst(rst));

	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance540530(.data_in(d_in53),.data_out(wire_d53_0),.clk(clk),.rst(rst));            //channel 54
	large_adder #(.WIDTH(WIDTH)) large_adder_instance540531(.data_in(wire_d53_0),.data_out(wire_d53_1),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance540532(.data_in(wire_d53_1),.data_out(wire_d53_2),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance540533(.data_in(wire_d53_2),.data_out(wire_d53_3),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance540534(.data_in(wire_d53_3),.data_out(wire_d53_4),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance540535(.data_in(wire_d53_4),.data_out(wire_d53_5),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance540536(.data_in(wire_d53_5),.data_out(wire_d53_6),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance540537(.data_in(wire_d53_6),.data_out(wire_d53_7),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance540538(.data_in(wire_d53_7),.data_out(wire_d53_8),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance540539(.data_in(wire_d53_8),.data_out(wire_d53_9),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405310(.data_in(wire_d53_9),.data_out(wire_d53_10),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405311(.data_in(wire_d53_10),.data_out(wire_d53_11),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405312(.data_in(wire_d53_11),.data_out(wire_d53_12),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405313(.data_in(wire_d53_12),.data_out(wire_d53_13),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405314(.data_in(wire_d53_13),.data_out(wire_d53_14),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5405315(.data_in(wire_d53_14),.data_out(wire_d53_15),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405316(.data_in(wire_d53_15),.data_out(wire_d53_16),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5405317(.data_in(wire_d53_16),.data_out(wire_d53_17),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5405318(.data_in(wire_d53_17),.data_out(wire_d53_18),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405319(.data_in(wire_d53_18),.data_out(wire_d53_19),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405320(.data_in(wire_d53_19),.data_out(wire_d53_20),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5405321(.data_in(wire_d53_20),.data_out(wire_d53_21),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405322(.data_in(wire_d53_21),.data_out(wire_d53_22),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405323(.data_in(wire_d53_22),.data_out(wire_d53_23),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405324(.data_in(wire_d53_23),.data_out(wire_d53_24),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405325(.data_in(wire_d53_24),.data_out(wire_d53_25),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405326(.data_in(wire_d53_25),.data_out(wire_d53_26),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405327(.data_in(wire_d53_26),.data_out(wire_d53_27),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5405328(.data_in(wire_d53_27),.data_out(wire_d53_28),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5405329(.data_in(wire_d53_28),.data_out(wire_d53_29),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405330(.data_in(wire_d53_29),.data_out(wire_d53_30),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405331(.data_in(wire_d53_30),.data_out(wire_d53_31),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405332(.data_in(wire_d53_31),.data_out(wire_d53_32),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5405333(.data_in(wire_d53_32),.data_out(wire_d53_33),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5405334(.data_in(wire_d53_33),.data_out(wire_d53_34),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5405335(.data_in(wire_d53_34),.data_out(wire_d53_35),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5405336(.data_in(wire_d53_35),.data_out(wire_d53_36),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5405337(.data_in(wire_d53_36),.data_out(wire_d53_37),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5405338(.data_in(wire_d53_37),.data_out(wire_d53_38),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5405339(.data_in(wire_d53_38),.data_out(wire_d53_39),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5405340(.data_in(wire_d53_39),.data_out(wire_d53_40),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5405341(.data_in(wire_d53_40),.data_out(wire_d53_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5405342(.data_in(wire_d53_41),.data_out(wire_d53_42),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5405343(.data_in(wire_d53_42),.data_out(wire_d53_43),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5405344(.data_in(wire_d53_43),.data_out(wire_d53_44),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405345(.data_in(wire_d53_44),.data_out(wire_d53_45),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5405346(.data_in(wire_d53_45),.data_out(wire_d53_46),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5405347(.data_in(wire_d53_46),.data_out(wire_d53_47),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5405348(.data_in(wire_d53_47),.data_out(wire_d53_48),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5405349(.data_in(wire_d53_48),.data_out(d_out53),.clk(clk),.rst(rst));

	encoder #(.WIDTH(WIDTH)) encoder_instance550540(.data_in(d_in54),.data_out(wire_d54_0),.clk(clk),.rst(rst));            //channel 55
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance550541(.data_in(wire_d54_0),.data_out(wire_d54_1),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance550542(.data_in(wire_d54_1),.data_out(wire_d54_2),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance550543(.data_in(wire_d54_2),.data_out(wire_d54_3),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance550544(.data_in(wire_d54_3),.data_out(wire_d54_4),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance550545(.data_in(wire_d54_4),.data_out(wire_d54_5),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance550546(.data_in(wire_d54_5),.data_out(wire_d54_6),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance550547(.data_in(wire_d54_6),.data_out(wire_d54_7),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance550548(.data_in(wire_d54_7),.data_out(wire_d54_8),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance550549(.data_in(wire_d54_8),.data_out(wire_d54_9),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5505410(.data_in(wire_d54_9),.data_out(wire_d54_10),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505411(.data_in(wire_d54_10),.data_out(wire_d54_11),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505412(.data_in(wire_d54_11),.data_out(wire_d54_12),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505413(.data_in(wire_d54_12),.data_out(wire_d54_13),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5505414(.data_in(wire_d54_13),.data_out(wire_d54_14),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505415(.data_in(wire_d54_14),.data_out(wire_d54_15),.clk(clk),.rst(rst));
	full_adder_top #(.WIDTH(WIDTH)) full_adder_instance5505416(.data_in(wire_d54_15),.data_out(wire_d54_16),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5505417(.data_in(wire_d54_16),.data_out(wire_d54_17),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5505418(.data_in(wire_d54_17),.data_out(wire_d54_18),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505419(.data_in(wire_d54_18),.data_out(wire_d54_19),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505420(.data_in(wire_d54_19),.data_out(wire_d54_20),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505421(.data_in(wire_d54_20),.data_out(wire_d54_21),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505422(.data_in(wire_d54_21),.data_out(wire_d54_22),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505423(.data_in(wire_d54_22),.data_out(wire_d54_23),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505424(.data_in(wire_d54_23),.data_out(wire_d54_24),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5505425(.data_in(wire_d54_24),.data_out(wire_d54_25),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505426(.data_in(wire_d54_25),.data_out(wire_d54_26),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505427(.data_in(wire_d54_26),.data_out(wire_d54_27),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5505428(.data_in(wire_d54_27),.data_out(wire_d54_28),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5505429(.data_in(wire_d54_28),.data_out(wire_d54_29),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505430(.data_in(wire_d54_29),.data_out(wire_d54_30),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505431(.data_in(wire_d54_30),.data_out(wire_d54_31),.clk(clk),.rst(rst));
	invertion #(.WIDTH(WIDTH)) invertion_instance5505432(.data_in(wire_d54_31),.data_out(wire_d54_32),.clk(clk),.rst(rst));
	d_latch_top #(.WIDTH(WIDTH)) d_latch_instance5505433(.data_in(wire_d54_32),.data_out(wire_d54_33),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505434(.data_in(wire_d54_33),.data_out(wire_d54_34),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5505435(.data_in(wire_d54_34),.data_out(wire_d54_35),.clk(clk),.rst(rst));
	memory_cntrl #(.WIDTH(WIDTH)) memory_cntrl_instance5505436(.data_in(wire_d54_35),.data_out(wire_d54_36),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505437(.data_in(wire_d54_36),.data_out(wire_d54_37),.clk(clk),.rst(rst));
	shift_reg_top #(.WIDTH(WIDTH)) shift_reg_instance5505438(.data_in(wire_d54_37),.data_out(wire_d54_38),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505439(.data_in(wire_d54_38),.data_out(wire_d54_39),.clk(clk),.rst(rst));
	large_adder #(.WIDTH(WIDTH)) large_adder_instance5505440(.data_in(wire_d54_39),.data_out(wire_d54_40),.clk(clk),.rst(rst));
	register #(.WIDTH(WIDTH)) register_instance5505441(.data_in(wire_d54_40),.data_out(wire_d54_41),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505442(.data_in(wire_d54_41),.data_out(wire_d54_42),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5505443(.data_in(wire_d54_42),.data_out(wire_d54_43),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505444(.data_in(wire_d54_43),.data_out(wire_d54_44),.clk(clk),.rst(rst));
	decoder_top #(.WIDTH(WIDTH)) decoder_instance5505445(.data_in(wire_d54_44),.data_out(wire_d54_45),.clk(clk),.rst(rst));
	encoder #(.WIDTH(WIDTH)) encoder_instance5505446(.data_in(wire_d54_45),.data_out(wire_d54_46),.clk(clk),.rst(rst));
	paritygenerator_top #(.WIDTH(WIDTH)) parity_generator_instance5505447(.data_in(wire_d54_46),.data_out(wire_d54_47),.clk(clk),.rst(rst));
	mod_n_counter #(.WIDTH(WIDTH)) mod_n_counter_instance5505448(.data_in(wire_d54_47),.data_out(wire_d54_48),.clk(clk),.rst(rst));
	large_mux #(.WIDTH(WIDTH)) large_mux_instance5505449(.data_in(wire_d54_48),.data_out(d_out54),.clk(clk),.rst(rst));


endmodule