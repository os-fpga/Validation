
module SOC_FPGA_INTF_AXI_M0 (
    // AXI master 0
    input  logic [        31:0] M0_ARADDR   ,
    input  logic [         1:0] M0_ARBURST  ,
    input  logic [         3:0] M0_ARCACHE  ,
    input  logic [         3:0] M0_ARID     ,
    input  logic [         2:0] M0_ARLEN    ,
    input  logic                M0_ARLOCK   ,
    input  logic [         2:0] M0_ARPROT   ,
    output logic                M0_ARREADY  ,
    input  logic [         2:0] M0_ARSIZE   ,
    input  logic                M0_ARVALID  ,
    input  logic [        31:0] M0_AWADDR   ,
    input  logic [         1:0] M0_AWBURST  ,
    input  logic [         3:0] M0_AWCACHE  ,
    input  logic [         3:0] M0_AWID     ,
    input  logic [         2:0] M0_AWLEN    ,
    input  logic                M0_AWLOCK   ,
    input  logic [         2:0] M0_AWPROT   ,
    output logic                M0_AWREADY  ,
    input  logic [         2:0] M0_AWSIZE   ,
    input  logic                M0_AWVALID  ,
    output logic [         3:0] M0_BID      ,
    input  logic                M0_BREADY   ,
    output logic [         1:0] M0_BRESP    ,
    output logic                M0_BVALID   ,
    output logic [        63:0] M0_RDATA    ,
    output logic [         3:0] M0_RID      ,
    output logic                M0_RLAST    ,
    input  logic                M0_RREADY   ,
    output logic [         1:0] M0_RRESP    ,
    output logic                M0_RVALID   ,
    input  logic [        63:0] M0_WDATA    ,
    input  logic                M0_WLAST    ,
    output logic                M0_WREADY   ,
    input  logic [         7:0] M0_WSTRB    ,
    input  logic                M0_WVALID   ,
    input                  	M0_ACLK     ,
    output                  	M0_ARESETN_I 
);
/*
module top(
input reset_n,
input reset_rtl_0_1,
input clk,
input [31:0]C_M_TARGET_SLAVE_BASE_ADDR_0_1,
input m00_axi_init_axi_txn_0_1


);

wire [31:0]C_M_TARGET_SLAVE_BASE_ADDR_0_1;
  wire [31:0]axi_interconnect_wra_0_m00_axi_ARADDR;
  wire [1:0]axi_interconnect_wra_0_m00_axi_ARBURST;
  wire [3:0]axi_interconnect_wra_0_m00_axi_ARCACHE;
  wire [7:0]axi_interconnect_wra_0_m00_axi_ARID;
  wire [7:0]axi_interconnect_wra_0_m00_axi_ARLEN;
  wire axi_interconnect_wra_0_m00_axi_ARLOCK;
  wire [2:0]axi_interconnect_wra_0_m00_axi_ARPROT;
  wire [3:0]axi_interconnect_wra_0_m00_axi_ARQOS;
  wire axi_interconnect_wra_0_m00_axi_ARREADY;
  wire [3:0]axi_interconnect_wra_0_m00_axi_ARREGION;
  wire [2:0]axi_interconnect_wra_0_m00_axi_ARSIZE;
  wire axi_interconnect_wra_0_m00_axi_ARUSER;
  wire axi_interconnect_wra_0_m00_axi_ARVALID;
  wire [31:0]axi_interconnect_wra_0_m00_axi_AWADDR;
  wire [1:0]axi_interconnect_wra_0_m00_axi_AWBURST;
  wire [3:0]axi_interconnect_wra_0_m00_axi_AWCACHE;
  wire [7:0]axi_interconnect_wra_0_m00_axi_AWID;
  wire [7:0]axi_interconnect_wra_0_m00_axi_AWLEN;
  wire axi_interconnect_wra_0_m00_axi_AWLOCK;
  wire [2:0]axi_interconnect_wra_0_m00_axi_AWPROT;
  wire [3:0]axi_interconnect_wra_0_m00_axi_AWQOS;
  wire axi_interconnect_wra_0_m00_axi_AWREADY;
  wire [3:0]axi_interconnect_wra_0_m00_axi_AWREGION;
  wire [2:0]axi_interconnect_wra_0_m00_axi_AWSIZE;
  wire axi_interconnect_wra_0_m00_axi_AWUSER;
  wire axi_interconnect_wra_0_m00_axi_AWVALID;
  wire [7:0]axi_interconnect_wra_0_m00_axi_BID;
  wire axi_interconnect_wra_0_m00_axi_BREADY;
  wire [1:0]axi_interconnect_wra_0_m00_axi_BRESP;
  wire axi_interconnect_wra_0_m00_axi_BUSER;
  wire axi_interconnect_wra_0_m00_axi_BVALID;
  wire [31:0]axi_interconnect_wra_0_m00_axi_RDATA;
  wire [7:0]axi_interconnect_wra_0_m00_axi_RID;
  wire axi_interconnect_wra_0_m00_axi_RLAST;
  wire axi_interconnect_wra_0_m00_axi_RREADY;
  wire [1:0]axi_interconnect_wra_0_m00_axi_RRESP;
  wire axi_interconnect_wra_0_m00_axi_RUSER;
  wire axi_interconnect_wra_0_m00_axi_RVALID;
  wire [31:0]axi_interconnect_wra_0_m00_axi_WDATA;
  wire axi_interconnect_wra_0_m00_axi_WLAST;
  wire axi_interconnect_wra_0_m00_axi_WREADY;
  wire [3:0]axi_interconnect_wra_0_m00_axi_WSTRB;
  wire axi_interconnect_wra_0_m00_axi_WUSER;
  wire axi_interconnect_wra_0_m00_axi_WVALID;
  wire [31:0]axi_interconnect_wra_0_m01_axi_ARADDR;
  wire [1:0]axi_interconnect_wra_0_m01_axi_ARBURST;
  wire [3:0]axi_interconnect_wra_0_m01_axi_ARCACHE;
  wire [7:0]axi_interconnect_wra_0_m01_axi_ARID;
  wire [7:0]axi_interconnect_wra_0_m01_axi_ARLEN;
  wire axi_interconnect_wra_0_m01_axi_ARLOCK;
  wire [2:0]axi_interconnect_wra_0_m01_axi_ARPROT;
  wire [3:0]axi_interconnect_wra_0_m01_axi_ARQOS;
  wire axi_interconnect_wra_0_m01_axi_ARREADY;
  wire [3:0]axi_interconnect_wra_0_m01_axi_ARREGION;
  wire [2:0]axi_interconnect_wra_0_m01_axi_ARSIZE;
  wire axi_interconnect_wra_0_m01_axi_ARUSER;
  wire axi_interconnect_wra_0_m01_axi_ARVALID;
  wire [31:0]axi_interconnect_wra_0_m01_axi_AWADDR;
  wire [1:0]axi_interconnect_wra_0_m01_axi_AWBURST;
  wire [3:0]axi_interconnect_wra_0_m01_axi_AWCACHE;
  wire [7:0]axi_interconnect_wra_0_m01_axi_AWID;
  wire [7:0]axi_interconnect_wra_0_m01_axi_AWLEN;
  wire axi_interconnect_wra_0_m01_axi_AWLOCK;
  wire [2:0]axi_interconnect_wra_0_m01_axi_AWPROT;
  wire [3:0]axi_interconnect_wra_0_m01_axi_AWQOS;
  wire axi_interconnect_wra_0_m01_axi_AWREADY;
  wire [3:0]axi_interconnect_wra_0_m01_axi_AWREGION;
  wire [2:0]axi_interconnect_wra_0_m01_axi_AWSIZE;
  wire axi_interconnect_wra_0_m01_axi_AWUSER;
  wire axi_interconnect_wra_0_m01_axi_AWVALID;
  wire [7:0]axi_interconnect_wra_0_m01_axi_BID;
  wire axi_interconnect_wra_0_m01_axi_BREADY;
  wire [1:0]axi_interconnect_wra_0_m01_axi_BRESP;
  wire axi_interconnect_wra_0_m01_axi_BUSER;
  wire axi_interconnect_wra_0_m01_axi_BVALID;
  wire [31:0]axi_interconnect_wra_0_m01_axi_RDATA;
  wire [7:0]axi_interconnect_wra_0_m01_axi_RID;
  wire axi_interconnect_wra_0_m01_axi_RLAST;
  wire axi_interconnect_wra_0_m01_axi_RREADY;
  wire [1:0]axi_interconnect_wra_0_m01_axi_RRESP;
  wire axi_interconnect_wra_0_m01_axi_RUSER;
  wire axi_interconnect_wra_0_m01_axi_RVALID;
  wire [31:0]axi_interconnect_wra_0_m01_axi_WDATA;
  wire axi_interconnect_wra_0_m01_axi_WLAST;
  wire axi_interconnect_wra_0_m01_axi_WREADY;
  wire [3:0]axi_interconnect_wra_0_m01_axi_WSTRB;
  wire axi_interconnect_wra_0_m01_axi_WUSER;
  wire axi_interconnect_wra_0_m01_axi_WVALID;
  wire clk_100MHz_1;
  wire clk_wiz_clk_out1;
  wire clk_wiz_locked;
  wire m00_axi_init_axi_txn_0_1;
  wire [31:0]myip_0_M00_AXI_ARADDR;
  wire [1:0]myip_0_M00_AXI_ARBURST;
  wire [3:0]myip_0_M00_AXI_ARCACHE;
  wire [0:0]myip_0_M00_AXI_ARID;
  wire [7:0]myip_0_M00_AXI_ARLEN;
  wire myip_0_M00_AXI_ARLOCK;
  wire [2:0]myip_0_M00_AXI_ARPROT;
  wire [3:0]myip_0_M00_AXI_ARQOS;
  wire myip_0_M00_AXI_ARREADY;
  wire [2:0]myip_0_M00_AXI_ARSIZE;
  wire [0:0]myip_0_M00_AXI_ARUSER;
  wire myip_0_M00_AXI_ARVALID;
  wire [31:0]myip_0_M00_AXI_AWADDR;
  wire [1:0]myip_0_M00_AXI_AWBURST;
  wire [3:0]myip_0_M00_AXI_AWCACHE;
  wire [0:0]myip_0_M00_AXI_AWID;
  wire [7:0]myip_0_M00_AXI_AWLEN;
  wire myip_0_M00_AXI_AWLOCK;
  wire [2:0]myip_0_M00_AXI_AWPROT;
  wire [3:0]myip_0_M00_AXI_AWQOS;
  wire myip_0_M00_AXI_AWREADY;
  wire [2:0]myip_0_M00_AXI_AWSIZE;
  wire [0:0]myip_0_M00_AXI_AWUSER;
  wire myip_0_M00_AXI_AWVALID;
  wire [7:0]myip_0_M00_AXI_BID;
  wire myip_0_M00_AXI_BREADY;
  wire [1:0]myip_0_M00_AXI_BRESP;
  wire myip_0_M00_AXI_BUSER;
  wire myip_0_M00_AXI_BVALID;
  wire [31:0]myip_0_M00_AXI_RDATA;
  wire [7:0]myip_0_M00_AXI_RID;
  wire myip_0_M00_AXI_RLAST;
  wire myip_0_M00_AXI_RREADY;
  wire [1:0]myip_0_M00_AXI_RRESP;
  wire myip_0_M00_AXI_RUSER;
  wire myip_0_M00_AXI_RVALID;
  wire [31:0]myip_0_M00_AXI_WDATA;
  wire myip_0_M00_AXI_WLAST;
  wire myip_0_M00_AXI_WREADY;
  wire [3:0]myip_0_M00_AXI_WSTRB;
  wire [0:0]myip_0_M00_AXI_WUSER;
  wire myip_0_M00_AXI_WVALID;
  wire reset_rtl_0_1;
  wire [0:0]rst_clk_wiz_100M_peripheral_aresetn;










design_1_myip_0_0 myip_0
       (.C_M_TARGET_SLAVE_BASE_ADDR_0(C_M_TARGET_SLAVE_BASE_ADDR_0_1),
        .m00_axi_aclk(M0_ACLK),
        .m00_axi_araddr(M0_ARADDR),
        .m00_axi_arburst(M0_ARBURST),
        .m00_axi_arcache(M0_ARCACHE),
        .m00_axi_aresetn(M0_ARESETN_I ),
        .m00_axi_arid(M0_ARID),
        .m00_axi_arlen(M0_ARLEN),
        .m00_axi_arlock(M0_ARLOCK),
        .m00_axi_arprot(M0_ARPROT),
        .m00_axi_arqos(myip_0_M00_AXI_ARQOS),
        .m00_axi_arready(M0_ARREADY),
        .m00_axi_arsize(M0_ARSIZE),
        .m00_axi_aruser(myip_0_M00_AXI_ARUSER),
        .m00_axi_arvalid(M0_ARVALID),
        .m00_axi_awaddr(M0_AWADDR),
        .m00_axi_awburst(M0_AWBURST),
        .m00_axi_awcache(M0_AWCACHE),
        .m00_axi_awid(M0_AWID),
        .m00_axi_awlen(M0_AWLEN),
        .m00_axi_awlock(M0_AWLOCK),
        .m00_axi_awprot(M0_AWPROT),
        .m00_axi_awqos(myip_0_M00_AXI_AWQOS),
        .m00_axi_awready(M0_AWREADY),
        .m00_axi_awsize(M0_AWSIZE),
        .m00_axi_awuser(myip_0_M00_AXI_AWUSER),
        .m00_axi_awvalid(M0_AWVALID),
        .m00_axi_bid(myip_0_M00_AXI_BID[0]),
        .m00_axi_bready(M0_BREADY),
        .m00_axi_bresp(M0_BRESP),
        .m00_axi_buser(myip_0_M00_AXI_BUSER),
        .m00_axi_bvalid(M0_BVALID),
        .m00_axi_init_axi_txn(m00_axi_init_axi_txn_0_1),
        .m00_axi_rdata(M0_RDATA),
        .m00_axi_rid(M0_RID),
        .m00_axi_rlast(M0_RLAST),
        .m00_axi_rready(M0_RREADY),
        .m00_axi_rresp(M0_RRESP),
        .m00_axi_ruser(myip_0_M00_AXI_RUSER),
        .m00_axi_rvalid(M0_RVALID),
        .m00_axi_wdata(M0_WDATA),
        .m00_axi_wlast(M0_WLAST),
        .m00_axi_wready(M0_WREADY),
        .m00_axi_wstrb(M0_WSTRB),
        .m00_axi_wuser(myip_0_M00_AXI_WUSER),
        .m00_axi_wvalid(M0_WVALID));   */

design_1_axi_interconnect_wra_0_0 axi_interconnect_wra_0
       (.clk(clk),
        .m00_axi_araddr(axi_interconnect_wra_0_m00_axi_ARADDR),
        .m00_axi_arburst(axi_interconnect_wra_0_m00_axi_ARBURST),
        .m00_axi_arcache(axi_interconnect_wra_0_m00_axi_ARCACHE),
        .m00_axi_arid(axi_interconnect_wra_0_m00_axi_ARID),
        .m00_axi_arlen(axi_interconnect_wra_0_m00_axi_ARLEN),
        .m00_axi_arlock(axi_interconnect_wra_0_m00_axi_ARLOCK),
        .m00_axi_arprot(axi_interconnect_wra_0_m00_axi_ARPROT),
        .m00_axi_arqos(axi_interconnect_wra_0_m00_axi_ARQOS),
        .m00_axi_arready(axi_interconnect_wra_0_m00_axi_ARREADY),
        .m00_axi_arregion(axi_interconnect_wra_0_m00_axi_ARREGION),
        .m00_axi_arsize(axi_interconnect_wra_0_m00_axi_ARSIZE),
        .m00_axi_aruser(axi_interconnect_wra_0_m00_axi_ARUSER),
        .m00_axi_arvalid(axi_interconnect_wra_0_m00_axi_ARVALID),
        .m00_axi_awaddr(axi_interconnect_wra_0_m00_axi_AWADDR),
        .m00_axi_awburst(axi_interconnect_wra_0_m00_axi_AWBURST),
        .m00_axi_awcache(axi_interconnect_wra_0_m00_axi_AWCACHE),
        .m00_axi_awid(axi_interconnect_wra_0_m00_axi_AWID),
        .m00_axi_awlen(axi_interconnect_wra_0_m00_axi_AWLEN),
        .m00_axi_awlock(axi_interconnect_wra_0_m00_axi_AWLOCK),
        .m00_axi_awprot(axi_interconnect_wra_0_m00_axi_AWPROT),
        .m00_axi_awqos(axi_interconnect_wra_0_m00_axi_AWQOS),
        .m00_axi_awready(axi_interconnect_wra_0_m00_axi_AWREADY),
        .m00_axi_awregion(axi_interconnect_wra_0_m00_axi_AWREGION),
        .m00_axi_awsize(axi_interconnect_wra_0_m00_axi_AWSIZE),
        .m00_axi_awuser(axi_interconnect_wra_0_m00_axi_AWUSER),
        .m00_axi_awvalid(axi_interconnect_wra_0_m00_axi_AWVALID),
        .m00_axi_bid(axi_interconnect_wra_0_m00_axi_BID),
        .m00_axi_bready(axi_interconnect_wra_0_m00_axi_BREADY),
        .m00_axi_bresp(axi_interconnect_wra_0_m00_axi_BRESP),
        .m00_axi_buser(axi_interconnect_wra_0_m00_axi_BUSER),
        .m00_axi_bvalid(axi_interconnect_wra_0_m00_axi_BVALID),
        .m00_axi_rdata(axi_interconnect_wra_0_m00_axi_RDATA),
        .m00_axi_rid(axi_interconnect_wra_0_m00_axi_RID),
        .m00_axi_rlast(axi_interconnect_wra_0_m00_axi_RLAST),
        .m00_axi_rready(axi_interconnect_wra_0_m00_axi_RREADY),
        .m00_axi_rresp(axi_interconnect_wra_0_m00_axi_RRESP),
        .m00_axi_ruser(axi_interconnect_wra_0_m00_axi_RUSER),
        .m00_axi_rvalid(axi_interconnect_wra_0_m00_axi_RVALID),
        .m00_axi_wdata(axi_interconnect_wra_0_m00_axi_WDATA),
        .m00_axi_wlast(axi_interconnect_wra_0_m00_axi_WLAST),
        .m00_axi_wready(axi_interconnect_wra_0_m00_axi_WREADY),
        .m00_axi_wstrb(axi_interconnect_wra_0_m00_axi_WSTRB),
        .m00_axi_wuser(axi_interconnect_wra_0_m00_axi_WUSER),
        .m00_axi_wvalid(axi_interconnect_wra_0_m00_axi_WVALID),
        .m01_axi_araddr(axi_interconnect_wra_0_m01_axi_ARADDR),
        .m01_axi_arburst(axi_interconnect_wra_0_m01_axi_ARBURST),
        .m01_axi_arcache(axi_interconnect_wra_0_m01_axi_ARCACHE),
        .m01_axi_arid(axi_interconnect_wra_0_m01_axi_ARID),
        .m01_axi_arlen(axi_interconnect_wra_0_m01_axi_ARLEN),
        .m01_axi_arlock(axi_interconnect_wra_0_m01_axi_ARLOCK),
        .m01_axi_arprot(axi_interconnect_wra_0_m01_axi_ARPROT),
        .m01_axi_arqos(axi_interconnect_wra_0_m01_axi_ARQOS),
        .m01_axi_arready(axi_interconnect_wra_0_m01_axi_ARREADY),
        .m01_axi_arregion(axi_interconnect_wra_0_m01_axi_ARREGION),
        .m01_axi_arsize(axi_interconnect_wra_0_m01_axi_ARSIZE),
        .m01_axi_aruser(axi_interconnect_wra_0_m01_axi_ARUSER),
        .m01_axi_arvalid(axi_interconnect_wra_0_m01_axi_ARVALID),
        .m01_axi_awaddr(axi_interconnect_wra_0_m01_axi_AWADDR),
        .m01_axi_awburst(axi_interconnect_wra_0_m01_axi_AWBURST),
        .m01_axi_awcache(axi_interconnect_wra_0_m01_axi_AWCACHE),
        .m01_axi_awid(axi_interconnect_wra_0_m01_axi_AWID),
        .m01_axi_awlen(axi_interconnect_wra_0_m01_axi_AWLEN),
        .m01_axi_awlock(axi_interconnect_wra_0_m01_axi_AWLOCK),
        .m01_axi_awprot(axi_interconnect_wra_0_m01_axi_AWPROT),
        .m01_axi_awqos(axi_interconnect_wra_0_m01_axi_AWQOS),
        .m01_axi_awready(axi_interconnect_wra_0_m01_axi_AWREADY),
        .m01_axi_awregion(axi_interconnect_wra_0_m01_axi_AWREGION),
        .m01_axi_awsize(axi_interconnect_wra_0_m01_axi_AWSIZE),
        .m01_axi_awuser(axi_interconnect_wra_0_m01_axi_AWUSER),
        .m01_axi_awvalid(axi_interconnect_wra_0_m01_axi_AWVALID),
        .m01_axi_bid(axi_interconnect_wra_0_m01_axi_BID),
        .m01_axi_bready(axi_interconnect_wra_0_m01_axi_BREADY),
        .m01_axi_bresp(axi_interconnect_wra_0_m01_axi_BRESP),
        .m01_axi_buser(axi_interconnect_wra_0_m01_axi_BUSER),
        .m01_axi_bvalid(axi_interconnect_wra_0_m01_axi_BVALID),
        .m01_axi_rdata(axi_interconnect_wra_0_m01_axi_RDATA),
        .m01_axi_rid(axi_interconnect_wra_0_m01_axi_RID),
        .m01_axi_rlast(axi_interconnect_wra_0_m01_axi_RLAST),
        .m01_axi_rready(axi_interconnect_wra_0_m01_axi_RREADY),
        .m01_axi_rresp(axi_interconnect_wra_0_m01_axi_RRESP),
        .m01_axi_ruser(axi_interconnect_wra_0_m01_axi_RUSER),
        .m01_axi_rvalid(axi_interconnect_wra_0_m01_axi_RVALID),
        .m01_axi_wdata(axi_interconnect_wra_0_m01_axi_WDATA),
        .m01_axi_wlast(axi_interconnect_wra_0_m01_axi_WLAST),
        .m01_axi_wready(axi_interconnect_wra_0_m01_axi_WREADY),
        .m01_axi_wstrb(axi_interconnect_wra_0_m01_axi_WSTRB),
        .m01_axi_wuser(axi_interconnect_wra_0_m01_axi_WUSER),
        .m01_axi_wvalid(axi_interconnect_wra_0_m01_axi_WVALID),
        .m02_axi_arready(1'b0),
        .m02_axi_awready(1'b0),
        .m02_axi_bid({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .m02_axi_bresp({1'b0,1'b0}),
        .m02_axi_buser(1'b0),
        .m02_axi_bvalid(1'b0),
        .m02_axi_rdata({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .m02_axi_rid({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .m02_axi_rlast(1'b0),
        .m02_axi_rresp({1'b0,1'b0}),
        .m02_axi_ruser(1'b0),
        .m02_axi_rvalid(1'b0),
        .m02_axi_wready(1'b0),
        .m03_axi_arready(1'b0),
        .m03_axi_awready(1'b0),
        .m03_axi_bid({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .m03_axi_bresp({1'b0,1'b0}),
        .m03_axi_buser(1'b0),
        .m03_axi_bvalid(1'b0),
        .m03_axi_rdata({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .m03_axi_rid({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .m03_axi_rlast(1'b0),
        .m03_axi_rresp({1'b0,1'b0}),
        .m03_axi_ruser(1'b0),
        .m03_axi_rvalid(1'b0),
        .m03_axi_wready(1'b0),
        .rst(reset_rtl_0_1),
        .s00_axi_araddr(myip_0_M00_AXI_ARADDR),
        .s00_axi_arburst(myip_0_M00_AXI_ARBURST),
        .s00_axi_arcache(myip_0_M00_AXI_ARCACHE),
        .s00_axi_arid({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,myip_0_M00_AXI_ARID}),
        .s00_axi_arlen(myip_0_M00_AXI_ARLEN),
        .s00_axi_arlock(myip_0_M00_AXI_ARLOCK),
        .s00_axi_arprot(myip_0_M00_AXI_ARPROT),
        .s00_axi_arqos(myip_0_M00_AXI_ARQOS),
        .s00_axi_arready(myip_0_M00_AXI_ARREADY),
        .s00_axi_arregion({1'b0,1'b0,1'b0,1'b0}),
        .s00_axi_arsize(myip_0_M00_AXI_ARSIZE),
        .s00_axi_aruser(myip_0_M00_AXI_ARUSER),
        .s00_axi_arvalid(myip_0_M00_AXI_ARVALID),
        .s00_axi_awaddr(myip_0_M00_AXI_AWADDR),
        .s00_axi_awburst(myip_0_M00_AXI_AWBURST),
        .s00_axi_awcache(myip_0_M00_AXI_AWCACHE),
        .s00_axi_awid({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,myip_0_M00_AXI_AWID}),
        .s00_axi_awlen(myip_0_M00_AXI_AWLEN),
        .s00_axi_awlock(myip_0_M00_AXI_AWLOCK),
        .s00_axi_awprot(myip_0_M00_AXI_AWPROT),
        .s00_axi_awqos(myip_0_M00_AXI_AWQOS),
        .s00_axi_awready(myip_0_M00_AXI_AWREADY),
        .s00_axi_awregion({1'b0,1'b0,1'b0,1'b0}),
        .s00_axi_awsize(myip_0_M00_AXI_AWSIZE),
        .s00_axi_awuser(myip_0_M00_AXI_AWUSER),
        .s00_axi_awvalid(myip_0_M00_AXI_AWVALID),
        .s00_axi_bid(myip_0_M00_AXI_BID),
        .s00_axi_bready(myip_0_M00_AXI_BREADY),
        .s00_axi_bresp(myip_0_M00_AXI_BRESP),
        .s00_axi_buser(myip_0_M00_AXI_BUSER),
        .s00_axi_bvalid(myip_0_M00_AXI_BVALID),
        .s00_axi_rdata(myip_0_M00_AXI_RDATA),
        .s00_axi_rid(myip_0_M00_AXI_RID),
        .s00_axi_rlast(myip_0_M00_AXI_RLAST),
        .s00_axi_rready(myip_0_M00_AXI_RREADY),
        .s00_axi_rresp(myip_0_M00_AXI_RRESP),
        .s00_axi_ruser(myip_0_M00_AXI_RUSER),
        .s00_axi_rvalid(myip_0_M00_AXI_RVALID),
        .s00_axi_wdata(myip_0_M00_AXI_WDATA),
        .s00_axi_wlast(myip_0_M00_AXI_WLAST),
        .s00_axi_wready(myip_0_M00_AXI_WREADY),
        .s00_axi_wstrb(myip_0_M00_AXI_WSTRB),
        .s00_axi_wuser(myip_0_M00_AXI_WUSER),
        .s00_axi_wvalid(myip_0_M00_AXI_WVALID),
        .s01_axi_araddr({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .s01_axi_arburst({1'b0,1'b1}),
        .s01_axi_arcache({1'b0,1'b0,1'b1,1'b1}),
        .s01_axi_arid({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .s01_axi_arlen({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .s01_axi_arlock(1'b0),
        .s01_axi_arprot({1'b0,1'b0,1'b0}),
        .s01_axi_arqos({1'b0,1'b0,1'b0,1'b0}),
        .s01_axi_arregion({1'b0,1'b0,1'b0,1'b0}),
        .s01_axi_arsize({1'b0,1'b1,1'b0}),
        .s01_axi_aruser(1'b0),
        .s01_axi_arvalid(1'b0),
        .s01_axi_awaddr({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .s01_axi_awburst({1'b0,1'b1}),
        .s01_axi_awcache({1'b0,1'b0,1'b1,1'b1}),
        .s01_axi_awid({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .s01_axi_awlen({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .s01_axi_awlock(1'b0),
        .s01_axi_awprot({1'b0,1'b0,1'b0}),
        .s01_axi_awqos({1'b0,1'b0,1'b0,1'b0}),
        .s01_axi_awregion({1'b0,1'b0,1'b0,1'b0}),
        .s01_axi_awsize({1'b0,1'b1,1'b0}),
        .s01_axi_awuser(1'b0),
        .s01_axi_awvalid(1'b0),
        .s01_axi_bready(1'b0),
        .s01_axi_rready(1'b0),
        .s01_axi_wdata({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .s01_axi_wlast(1'b0),
        .s01_axi_wstrb({1'b1,1'b1,1'b1,1'b1}),
        .s01_axi_wuser(1'b0),
        .s01_axi_wvalid(1'b0),
        .s02_axi_araddr({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .s02_axi_arburst({1'b0,1'b1}),
        .s02_axi_arcache({1'b0,1'b0,1'b1,1'b1}),
        .s02_axi_arid({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .s02_axi_arlen({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .s02_axi_arlock(1'b0),
        .s02_axi_arprot({1'b0,1'b0,1'b0}),
        .s02_axi_arqos({1'b0,1'b0,1'b0,1'b0}),
        .s02_axi_arregion({1'b0,1'b0,1'b0,1'b0}),
        .s02_axi_arsize({1'b0,1'b1,1'b0}),
        .s02_axi_aruser(1'b0),
        .s02_axi_arvalid(1'b0),
        .s02_axi_awaddr({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .s02_axi_awburst({1'b0,1'b1}),
        .s02_axi_awcache({1'b0,1'b0,1'b1,1'b1}),
        .s02_axi_awid({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .s02_axi_awlen({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .s02_axi_awlock(1'b0),
        .s02_axi_awprot({1'b0,1'b0,1'b0}),
        .s02_axi_awqos({1'b0,1'b0,1'b0,1'b0}),
        .s02_axi_awregion({1'b0,1'b0,1'b0,1'b0}),
        .s02_axi_awsize({1'b0,1'b1,1'b0}),
        .s02_axi_awuser(1'b0),
        .s02_axi_awvalid(1'b0),
        .s02_axi_bready(1'b0),
        .s02_axi_rready(1'b0),
        .s02_axi_wdata({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .s02_axi_wlast(1'b0),
        .s02_axi_wstrb({1'b1,1'b1,1'b1,1'b1}),
        .s02_axi_wuser(1'b0),
        .s02_axi_wvalid(1'b0),
        .s03_axi_araddr({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .s03_axi_arburst({1'b0,1'b1}),
        .s03_axi_arcache({1'b0,1'b0,1'b1,1'b1}),
        .s03_axi_arid({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .s03_axi_arlen({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .s03_axi_arlock(1'b0),
        .s03_axi_arprot({1'b0,1'b0,1'b0}),
        .s03_axi_arqos({1'b0,1'b0,1'b0,1'b0}),
        .s03_axi_arregion({1'b0,1'b0,1'b0,1'b0}),
        .s03_axi_arsize({1'b0,1'b1,1'b0}),
        .s03_axi_aruser(1'b0),
        .s03_axi_arvalid(1'b0),
        .s03_axi_awaddr({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .s03_axi_awburst({1'b0,1'b1}),
        .s03_axi_awcache({1'b0,1'b0,1'b1,1'b1}),
        .s03_axi_awid({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .s03_axi_awlen({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .s03_axi_awlock(1'b0),
        .s03_axi_awprot({1'b0,1'b0,1'b0}),
        .s03_axi_awqos({1'b0,1'b0,1'b0,1'b0}),
        .s03_axi_awregion({1'b0,1'b0,1'b0,1'b0}),
        .s03_axi_awsize({1'b0,1'b1,1'b0}),
        .s03_axi_awuser(1'b0),
        .s03_axi_awvalid(1'b0),
        .s03_axi_bready(1'b0),
        .s03_axi_rready(1'b0),
        .s03_axi_wdata({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),
        .s03_axi_wlast(1'b0),
        .s03_axi_wstrb({1'b1,1'b1,1'b1,1'b1}),
        .s03_axi_wuser(1'b0),
        .s03_axi_wvalid(1'b0));
  design_1_axi_ram_wrapper_0_1 axi_ram_wrapper_0
       (.clk(clk),
        .rst(reset_rtl_0_1),
        .s_axi_araddr(axi_interconnect_wra_0_m00_axi_ARADDR),
        .s_axi_arburst(axi_interconnect_wra_0_m00_axi_ARBURST),
        .s_axi_arcache(axi_interconnect_wra_0_m00_axi_ARCACHE),
        .s_axi_arid(axi_interconnect_wra_0_m00_axi_ARID),
        .s_axi_arlen(axi_interconnect_wra_0_m00_axi_ARLEN),
        .s_axi_arlock(axi_interconnect_wra_0_m00_axi_ARLOCK),
        .s_axi_arprot(axi_interconnect_wra_0_m00_axi_ARPROT),
        .s_axi_arqos(axi_interconnect_wra_0_m00_axi_ARQOS),
        .s_axi_arready(axi_interconnect_wra_0_m00_axi_ARREADY),
        .s_axi_arregion(axi_interconnect_wra_0_m00_axi_ARREGION),
        .s_axi_arsize(axi_interconnect_wra_0_m00_axi_ARSIZE),
        .s_axi_aruser(axi_interconnect_wra_0_m00_axi_ARUSER),
        .s_axi_arvalid(axi_interconnect_wra_0_m00_axi_ARVALID),
        .s_axi_awaddr(axi_interconnect_wra_0_m00_axi_AWADDR),
        .s_axi_awburst(axi_interconnect_wra_0_m00_axi_AWBURST),
        .s_axi_awcache(axi_interconnect_wra_0_m00_axi_AWCACHE),
        .s_axi_awid(axi_interconnect_wra_0_m00_axi_AWID),
        .s_axi_awlen(axi_interconnect_wra_0_m00_axi_AWLEN),
        .s_axi_awlock(axi_interconnect_wra_0_m00_axi_AWLOCK),
        .s_axi_awprot(axi_interconnect_wra_0_m00_axi_AWPROT),
        .s_axi_awqos(axi_interconnect_wra_0_m00_axi_AWQOS),
        .s_axi_awready(axi_interconnect_wra_0_m00_axi_AWREADY),
        .s_axi_awregion(axi_interconnect_wra_0_m00_axi_AWREGION),
        .s_axi_awsize(axi_interconnect_wra_0_m00_axi_AWSIZE),
        .s_axi_awuser(axi_interconnect_wra_0_m00_axi_AWUSER),
        .s_axi_awvalid(axi_interconnect_wra_0_m00_axi_AWVALID),
        .s_axi_bid(axi_interconnect_wra_0_m00_axi_BID),
        .s_axi_bready(axi_interconnect_wra_0_m00_axi_BREADY),
        .s_axi_bresp(axi_interconnect_wra_0_m00_axi_BRESP),
        .s_axi_buser(axi_interconnect_wra_0_m00_axi_BUSER),
        .s_axi_bvalid(axi_interconnect_wra_0_m00_axi_BVALID),
        .s_axi_rdata(axi_interconnect_wra_0_m00_axi_RDATA),
        .s_axi_rid(axi_interconnect_wra_0_m00_axi_RID),
        .s_axi_rlast(axi_interconnect_wra_0_m00_axi_RLAST),
        .s_axi_rready(axi_interconnect_wra_0_m00_axi_RREADY),
        .s_axi_rresp(axi_interconnect_wra_0_m00_axi_RRESP),
        .s_axi_ruser(axi_interconnect_wra_0_m00_axi_RUSER),
        .s_axi_rvalid(axi_interconnect_wra_0_m00_axi_RVALID),
        .s_axi_wdata(axi_interconnect_wra_0_m00_axi_WDATA),
        .s_axi_wlast(axi_interconnect_wra_0_m00_axi_WLAST),
        .s_axi_wready(axi_interconnect_wra_0_m00_axi_WREADY),
        .s_axi_wstrb(axi_interconnect_wra_0_m00_axi_WSTRB),
        .s_axi_wuser(axi_interconnect_wra_0_m00_axi_WUSER),
        .s_axi_wvalid(axi_interconnect_wra_0_m00_axi_WVALID));
  design_1_axi_ram_wrapper_1_0 axi_ram_wrapper_1
       (.clk(clk),
        .rst(reset_rtl_0_1),
        .s_axi_araddr(axi_interconnect_wra_0_m01_axi_ARADDR),
        .s_axi_arburst(axi_interconnect_wra_0_m01_axi_ARBURST),
        .s_axi_arcache(axi_interconnect_wra_0_m01_axi_ARCACHE),
        .s_axi_arid(axi_interconnect_wra_0_m01_axi_ARID),
        .s_axi_arlen(axi_interconnect_wra_0_m01_axi_ARLEN),
        .s_axi_arlock(axi_interconnect_wra_0_m01_axi_ARLOCK),
        .s_axi_arprot(axi_interconnect_wra_0_m01_axi_ARPROT),
        .s_axi_arqos(axi_interconnect_wra_0_m01_axi_ARQOS),
        .s_axi_arready(axi_interconnect_wra_0_m01_axi_ARREADY),
        .s_axi_arregion(axi_interconnect_wra_0_m01_axi_ARREGION),
        .s_axi_arsize(axi_interconnect_wra_0_m01_axi_ARSIZE),
        .s_axi_aruser(axi_interconnect_wra_0_m01_axi_ARUSER),
        .s_axi_arvalid(axi_interconnect_wra_0_m01_axi_ARVALID),
        .s_axi_awaddr(axi_interconnect_wra_0_m01_axi_AWADDR),
        .s_axi_awburst(axi_interconnect_wra_0_m01_axi_AWBURST),
        .s_axi_awcache(axi_interconnect_wra_0_m01_axi_AWCACHE),
        .s_axi_awid(axi_interconnect_wra_0_m01_axi_AWID),
        .s_axi_awlen(axi_interconnect_wra_0_m01_axi_AWLEN),
        .s_axi_awlock(axi_interconnect_wra_0_m01_axi_AWLOCK),
        .s_axi_awprot(axi_interconnect_wra_0_m01_axi_AWPROT),
        .s_axi_awqos(axi_interconnect_wra_0_m01_axi_AWQOS),
        .s_axi_awready(axi_interconnect_wra_0_m01_axi_AWREADY),
        .s_axi_awregion(axi_interconnect_wra_0_m01_axi_AWREGION),
        .s_axi_awsize(axi_interconnect_wra_0_m01_axi_AWSIZE),
        .s_axi_awuser(axi_interconnect_wra_0_m01_axi_AWUSER),
        .s_axi_awvalid(axi_interconnect_wra_0_m01_axi_AWVALID),
        .s_axi_bid(axi_interconnect_wra_0_m01_axi_BID),
        .s_axi_bready(axi_interconnect_wra_0_m01_axi_BREADY),
        .s_axi_bresp(axi_interconnect_wra_0_m01_axi_BRESP),
        .s_axi_buser(axi_interconnect_wra_0_m01_axi_BUSER),
        .s_axi_bvalid(axi_interconnect_wra_0_m01_axi_BVALID),
        .s_axi_rdata(axi_interconnect_wra_0_m01_axi_RDATA),
        .s_axi_rid(axi_interconnect_wra_0_m01_axi_RID),
        .s_axi_rlast(axi_interconnect_wra_0_m01_axi_RLAST),
        .s_axi_rready(axi_interconnect_wra_0_m01_axi_RREADY),
        .s_axi_rresp(axi_interconnect_wra_0_m01_axi_RRESP),
        .s_axi_ruser(axi_interconnect_wra_0_m01_axi_RUSER),
        .s_axi_rvalid(axi_interconnect_wra_0_m01_axi_RVALID),
        .s_axi_wdata(axi_interconnect_wra_0_m01_axi_WDATA),
        .s_axi_wlast(axi_interconnect_wra_0_m01_axi_WLAST),
        .s_axi_wready(axi_interconnect_wra_0_m01_axi_WREADY),
        .s_axi_wstrb(axi_interconnect_wra_0_m01_axi_WSTRB),
        .s_axi_wuser(axi_interconnect_wra_0_m01_axi_WUSER),
        .s_axi_wvalid(axi_interconnect_wra_0_m01_axi_WVALID));

endmodule 