module soc_fpga_intf_inst (
    
    input         clk_fpga_fabric_irq       ,
    input         clk_fpga_fabric_dma       ,
    input         clk_fpga_fabric_gpio       ,
    input         rst_n_fpga_fabric_irq     ,
    input         rst_n_fpga_fabric_dma     ,
    input         rst_n_fpga_fabric_gpio    ,
    output        rst_n_fpga0             ,
    output        rst_n_fpga1             ,
    output        rst_n_fpga_s             ,
    input         clk_fpga_fabric_m0,
    input         clk_fpga_fabric_m1,
    input         clk_fpga_fabric_s0,
    output [31:0] fpga_clk_ahb_s0_haddr     ,
    output [ 2:0] fpga_clk_ahb_s0_hburst    ,
    output        fpga_clk_ahb_s0_hmastlock ,
    input         fpga_clk_ahb_s0_hready    ,
    output [ 3:0] fpga_clk_ahb_s0_hprot     ,
    input  [31:0] fpga_clk_ahb_s0_hrdata    ,
    input         fpga_clk_ahb_s0_hresp     ,
    output        fpga_clk_ahb_s0_hsel      ,
    output [ 2:0] fpga_clk_ahb_s0_hsize     ,
    output [ 1:0] fpga_clk_ahb_s0_htrans    ,
    output [ 3:0] fpga_clk_ahb_s0_hwbe      ,
    output [31:0] fpga_clk_ahb_s0_hwdata    ,
    output        fpga_clk_ahb_s0_hwrite    ,
    input  [31:0] fpga_clk_axi_m0_ar_addr   ,
    input  [ 1:0] fpga_clk_axi_m0_ar_burst  ,
    input  [ 3:0] fpga_clk_axi_m0_ar_cache  ,
    input  [ 3:0] fpga_clk_axi_m0_ar_id     ,
    input  [ 2:0] fpga_clk_axi_m0_ar_len    ,
    input         fpga_clk_axi_m0_ar_lock   ,
    input  [ 2:0] fpga_clk_axi_m0_ar_prot   ,
    output        fpga_clk_axi_m0_ar_ready  ,
    input  [ 2:0] fpga_clk_axi_m0_ar_size   ,
    input         fpga_clk_axi_m0_ar_valid  ,
    input  [31:0] fpga_clk_axi_m0_aw_addr   ,
    input  [ 1:0] fpga_clk_axi_m0_aw_burst  ,
    input  [ 3:0] fpga_clk_axi_m0_aw_cache  ,
    input  [ 3:0] fpga_clk_axi_m0_aw_id     ,
    input  [ 2:0] fpga_clk_axi_m0_aw_len    ,
    input         fpga_clk_axi_m0_aw_lock   ,
    input  [ 2:0] fpga_clk_axi_m0_aw_prot   ,
    output        fpga_clk_axi_m0_aw_ready  ,
    input  [ 2:0] fpga_clk_axi_m0_aw_size   ,
    input         fpga_clk_axi_m0_aw_valid  ,
    output [ 3:0] fpga_clk_axi_m0_b_id      ,
    input         fpga_clk_axi_m0_b_ready   ,
    output [ 1:0] fpga_clk_axi_m0_b_resp    ,
    output        fpga_clk_axi_m0_b_valid   ,
    output [63:0] fpga_clk_axi_m0_r_data    ,
    output [ 3:0] fpga_clk_axi_m0_r_id      ,
    output        fpga_clk_axi_m0_r_last    ,
    input         fpga_clk_axi_m0_r_ready   ,
    output [ 1:0] fpga_clk_axi_m0_r_resp    ,
    output        fpga_clk_axi_m0_r_valid   ,
    input  [63:0] fpga_clk_axi_m0_w_data    ,
    input         fpga_clk_axi_m0_w_last    ,
    output        fpga_clk_axi_m0_w_ready   ,
    input  [ 7:0] fpga_clk_axi_m0_w_strb    ,
    input         fpga_clk_axi_m0_w_valid   ,
    input  [31:0] fpga_clk_axi_m1_ar_addr   ,
    input  [ 1:0] fpga_clk_axi_m1_ar_burst  ,
    input  [ 3:0] fpga_clk_axi_m1_ar_cache  ,
    input  [ 3:0] fpga_clk_axi_m1_ar_id     ,
    input  [ 3:0] fpga_clk_axi_m1_ar_len    ,
    input         fpga_clk_axi_m1_ar_lock   ,
    input  [ 2:0] fpga_clk_axi_m1_ar_prot   ,
    output        fpga_clk_axi_m1_ar_ready  ,
    input  [ 2:0] fpga_clk_axi_m1_ar_size   ,
    input         fpga_clk_axi_m1_ar_valid  ,
    input  [31:0] fpga_clk_axi_m1_aw_addr   ,
    input  [ 1:0] fpga_clk_axi_m1_aw_burst  ,
    input  [ 3:0] fpga_clk_axi_m1_aw_cache  ,
    input  [ 3:0] fpga_clk_axi_m1_aw_id     ,
    input  [ 3:0] fpga_clk_axi_m1_aw_len    ,
    input         fpga_clk_axi_m1_aw_lock   ,
    input  [ 2:0] fpga_clk_axi_m1_aw_prot   ,
    output        fpga_clk_axi_m1_aw_ready  ,
    input  [ 2:0] fpga_clk_axi_m1_aw_size   ,
    input         fpga_clk_axi_m1_aw_valid  ,
    output [ 3:0] fpga_clk_axi_m1_b_id      ,
    input         fpga_clk_axi_m1_b_ready   ,
    output [ 1:0] fpga_clk_axi_m1_b_resp    ,
    output        fpga_clk_axi_m1_b_valid   ,
    output [31:0] fpga_clk_axi_m1_r_data    ,
    output [ 3:0] fpga_clk_axi_m1_r_id      ,
    output        fpga_clk_axi_m1_r_last    ,
    input         fpga_clk_axi_m1_r_ready   ,
    output [ 1:0] fpga_clk_axi_m1_r_resp    ,
    output        fpga_clk_axi_m1_r_valid   ,
    input  [31:0] fpga_clk_axi_m1_w_data    ,
    input         fpga_clk_axi_m1_w_last    ,
    output        fpga_clk_axi_m1_w_ready   ,
    input  [ 3:0] fpga_clk_axi_m1_w_strb    ,
    input         fpga_clk_axi_m1_w_valid   ,
    input  [15:0] fpga_clk_irq_src          ,
    output [15:0] fpga_clk_irq_set          ,
    input  [ 3:0] fpga_clk_dma_req          ,
    output [ 3:0] fpga_clk_dma_ack          ,
    input         fpga_jtag_tck                ,
    output        fpga_jtag_tdi                ,
    input         fpga_jtag_tdo                ,
    output        fpga_jtag_tms                ,
    output        fpga_jtag_trstn              ,
    input         fpga_jtag_en                 ,
    input         soc_fpga_jtag_tdi                ,
    output        soc_fpga_jtag_tdo                ,
    input         soc_fpga_jtag_tms                ,
    input         soc_fpga_jtag_trstn              ,
    output [39:0] fpga_pad_c       ,
    input  [39:0] fpga_pad_i       ,
    input  [39:0] fpga_pad_oen     

);

soc_fpga_intf inst (
    .clk_fpga_fabric_irq(clk_fpga_fabric_irq),
    .clk_fpga_fabric_dma(clk_fpga_fabric_dma),
    .clk_fpga_fabric_gpio(clk_fpga_fabric_gpio),
    .rst_n_fpga_fabric_irq(rst_n_fpga_fabric_irq),
    .rst_n_fpga_fabric_dma(rst_n_fpga_fabric_dma),
    .rst_n_fpga_fabric_gpio(rst_n_fpga_fabric_gpio),
    .rst_n_fpga0(rst_n_fpga0),
    .rst_n_fpga1(rst_n_fpga1),
    .rst_n_fpga_s(rst_n_fpga_s),
    .clk_fpga_fabric_m0(clk_fpga_fabric_m0),
    .clk_fpga_fabric_m1(clk_fpga_fabric_m1),
    .clk_fpga_fabric_s0(clk_fpga_fabric_s0),
    .fpga_clk_ahb_s0_haddr(fpga_clk_ahb_s0_haddr),
    .fpga_clk_ahb_s0_hburst(fpga_clk_ahb_s0_hburst),
    .fpga_clk_ahb_s0_hmastlock(fpga_clk_ahb_s0_hmastlock),
    .fpga_clk_ahb_s0_hready(fpga_clk_ahb_s0_hready),
    .fpga_clk_ahb_s0_hprot(fpga_clk_ahb_s0_hprot),
    .fpga_clk_ahb_s0_hrdata(fpga_clk_ahb_s0_hrdata),
    .fpga_clk_ahb_s0_hresp(fpga_clk_ahb_s0_hresp),
    .fpga_clk_ahb_s0_hsel(fpga_clk_ahb_s0_hsel),
    .fpga_clk_ahb_s0_hsize(fpga_clk_ahb_s0_hsize),
    .fpga_clk_ahb_s0_htrans(fpga_clk_ahb_s0_htrans),
    .fpga_clk_ahb_s0_hwbe(fpga_clk_ahb_s0_hwbe),
    .fpga_clk_ahb_s0_hwdata(fpga_clk_ahb_s0_hwdata),
    .fpga_clk_ahb_s0_hwrite(fpga_clk_ahb_s0_hwrite),
    .fpga_clk_axi_m0_ar_addr(fpga_clk_axi_m0_ar_addr),
    .fpga_clk_axi_m0_ar_burst(fpga_clk_axi_m0_ar_burst),
    .fpga_clk_axi_m0_ar_cache(fpga_clk_axi_m0_ar_cache),
    .fpga_clk_axi_m0_ar_id(fpga_clk_axi_m0_ar_id),
    .fpga_clk_axi_m0_ar_len(fpga_clk_axi_m0_ar_len),
    .fpga_clk_axi_m0_ar_lock(fpga_clk_axi_m0_ar_lock),
    .fpga_clk_axi_m0_ar_prot(fpga_clk_axi_m0_ar_prot),
    .fpga_clk_axi_m0_ar_ready(fpga_clk_axi_m0_ar_ready),
    .fpga_clk_axi_m0_ar_size(fpga_clk_axi_m0_ar_size),
    .fpga_clk_axi_m0_ar_valid(fpga_clk_axi_m0_ar_valid),
    .fpga_clk_axi_m0_aw_addr(fpga_clk_axi_m0_aw_addr),
    .fpga_clk_axi_m0_aw_burst(fpga_clk_axi_m0_aw_burst),
    .fpga_clk_axi_m0_aw_cache(fpga_clk_axi_m0_aw_cache),
    .fpga_clk_axi_m0_aw_id(fpga_clk_axi_m0_aw_id),
    .fpga_clk_axi_m0_aw_len(fpga_clk_axi_m0_aw_len),
    .fpga_clk_axi_m0_aw_lock(fpga_clk_axi_m0_aw_lock),
    .fpga_clk_axi_m0_aw_prot(fpga_clk_axi_m0_aw_prot),
    .fpga_clk_axi_m0_aw_ready(fpga_clk_axi_m0_aw_ready),
    .fpga_clk_axi_m0_aw_size(fpga_clk_axi_m0_aw_size),
    .fpga_clk_axi_m0_aw_valid(fpga_clk_axi_m0_aw_valid),
    .fpga_clk_axi_m0_b_id(fpga_clk_axi_m0_b_id),
    .fpga_clk_axi_m0_b_ready(fpga_clk_axi_m0_b_ready),
    .fpga_clk_axi_m0_b_resp(fpga_clk_axi_m0_b_resp),
    .fpga_clk_axi_m0_b_valid(fpga_clk_axi_m0_b_valid),
    .fpga_clk_axi_m0_r_data(fpga_clk_axi_m0_r_data),
    .fpga_clk_axi_m0_r_id(fpga_clk_axi_m0_r_id),
    .fpga_clk_axi_m0_r_last(fpga_clk_axi_m0_r_last),
    .fpga_clk_axi_m0_r_ready(fpga_clk_axi_m0_r_ready),
    .fpga_clk_axi_m0_r_resp(fpga_clk_axi_m0_r_resp),
    .fpga_clk_axi_m0_r_valid(fpga_clk_axi_m0_r_valid),
    .fpga_clk_axi_m0_w_data(fpga_clk_axi_m0_w_data),
    .fpga_clk_axi_m0_w_last(fpga_clk_axi_m0_w_last),
    .fpga_clk_axi_m0_w_ready(fpga_clk_axi_m0_w_ready),
    .fpga_clk_axi_m0_w_strb(fpga_clk_axi_m0_w_strb),
    .fpga_clk_axi_m0_w_valid(fpga_clk_axi_m0_w_valid),
    .fpga_clk_axi_m1_ar_addr(fpga_clk_axi_m1_ar_addr),
    .fpga_clk_axi_m1_ar_burst(fpga_clk_axi_m1_ar_burst),
    .fpga_clk_axi_m1_ar_cache(fpga_clk_axi_m1_ar_cache),
    .fpga_clk_axi_m1_ar_id(fpga_clk_axi_m1_ar_id),
    .fpga_clk_axi_m1_ar_len(fpga_clk_axi_m1_ar_len),
    .fpga_clk_axi_m1_ar_lock(fpga_clk_axi_m1_ar_lock),
    .fpga_clk_axi_m1_ar_prot(fpga_clk_axi_m1_ar_prot),
    .fpga_clk_axi_m1_ar_ready(fpga_clk_axi_m1_ar_ready),
    .fpga_clk_axi_m1_ar_size(fpga_clk_axi_m1_ar_size),
    .fpga_clk_axi_m1_ar_valid(fpga_clk_axi_m1_ar_valid),
    .fpga_clk_axi_m1_aw_addr(fpga_clk_axi_m1_aw_addr),
    .fpga_clk_axi_m1_aw_burst(fpga_clk_axi_m1_aw_burst),
    .fpga_clk_axi_m1_aw_cache(fpga_clk_axi_m1_aw_cache),
    .fpga_clk_axi_m1_aw_id(fpga_clk_axi_m1_aw_id),
    .fpga_clk_axi_m1_aw_len(fpga_clk_axi_m1_aw_len),
    .fpga_clk_axi_m1_aw_lock(fpga_clk_axi_m1_aw_lock),
    .fpga_clk_axi_m1_aw_prot(fpga_clk_axi_m1_aw_prot),
    .fpga_clk_axi_m1_aw_ready(fpga_clk_axi_m1_aw_ready),
    .fpga_clk_axi_m1_aw_size(fpga_clk_axi_m1_aw_size),
    .fpga_clk_axi_m1_aw_valid(fpga_clk_axi_m1_aw_valid),
    .fpga_clk_axi_m1_b_id(fpga_clk_axi_m1_b_id),
    .fpga_clk_axi_m1_b_ready(fpga_clk_axi_m1_b_ready),
    .fpga_clk_axi_m1_b_resp(fpga_clk_axi_m1_b_resp),
    .fpga_clk_axi_m1_b_valid(fpga_clk_axi_m1_b_valid),
    .fpga_clk_axi_m1_r_data(fpga_clk_axi_m1_r_data),
    .fpga_clk_axi_m1_r_id(fpga_clk_axi_m1_r_id),
    .fpga_clk_axi_m1_r_last(fpga_clk_axi_m1_r_last),
    .fpga_clk_axi_m1_r_ready(fpga_clk_axi_m1_r_ready),
    .fpga_clk_axi_m1_r_resp(fpga_clk_axi_m1_r_resp),
    .fpga_clk_axi_m1_r_valid(fpga_clk_axi_m1_r_valid),
    .fpga_clk_axi_m1_w_data(fpga_clk_axi_m1_w_data),
    .fpga_clk_axi_m1_w_last(fpga_clk_axi_m1_w_last),
    .fpga_clk_axi_m1_w_ready(fpga_clk_axi_m1_w_ready),
    .fpga_clk_axi_m1_w_strb(fpga_clk_axi_m1_w_strb),
    .fpga_clk_axi_m1_w_valid(fpga_clk_axi_m1_w_valid),
    .fpga_clk_irq_src(fpga_clk_irq_src),
    .fpga_clk_irq_set(fpga_clk_irq_set),
    .fpga_clk_dma_req(fpga_clk_dma_req),
    .fpga_clk_dma_ack(fpga_clk_dma_ack),
    .fpga_jtag_tck(fpga_jtag_tck),
    .fpga_jtag_tdi(fpga_jtag_tdi),
    .fpga_jtag_tdo(fpga_jtag_tdo),
    .fpga_jtag_tms(fpga_jtag_tms),
    .fpga_jtag_trstn(fpga_jtag_trstn),
    .fpga_jtag_en(fpga_jtag_en),
    .soc_fpga_jtag_tdi(soc_fpga_jtag_tdi),
    .soc_fpga_jtag_tdo(soc_fpga_jtag_tdo),
    .soc_fpga_jtag_tms(soc_fpga_jtag_tms),
    .soc_fpga_jtag_trstn(soc_fpga_jtag_trstn),
    .fpga_pad_c(fpga_pad_c),
    .fpga_pad_i(fpga_pad_i),
    .fpga_pad_oen(fpga_pad_oen)
);

endmodule 
