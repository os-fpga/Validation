/////////////////////////////////////////
//  Functionality: feedthrough path
//  Author:        George Chen
////////////////////////////////////////
// `timescale 1ns / 1ps


module GJC9( din, dout);

  input din;
  output dout;

  assign dout = din ;
   
endmodule
