-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb6",
     9 => x"9c080b0b",
    10 => x"0bb6a008",
    11 => x"0b0b0bb6",
    12 => x"a4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b6a40c0b",
    16 => x"0b0bb6a0",
    17 => x"0c0b0b0b",
    18 => x"b69c0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bafc4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b69c7080",
    57 => x"c0cc278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"5188b004",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bb6ac0c",
    65 => x"9f0bb6b0",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"b6b008ff",
    69 => x"05b6b00c",
    70 => x"b6b00880",
    71 => x"25eb38b6",
    72 => x"ac08ff05",
    73 => x"b6ac0cb6",
    74 => x"ac088025",
    75 => x"d738800b",
    76 => x"b6b00c80",
    77 => x"0bb6ac0c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bb6ac08",
    97 => x"258f3882",
    98 => x"bd2db6ac",
    99 => x"08ff05b6",
   100 => x"ac0c82ff",
   101 => x"04b6ac08",
   102 => x"b6b00853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"b6ac08a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134b6b0",
   111 => x"088105b6",
   112 => x"b00cb6b0",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bb6b00c",
   116 => x"b6ac0881",
   117 => x"05b6ac0c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134b6",
   122 => x"b0088105",
   123 => x"b6b00cb6",
   124 => x"b008a02e",
   125 => x"0981068e",
   126 => x"38800bb6",
   127 => x"b00cb6ac",
   128 => x"088105b6",
   129 => x"ac0c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bb6b4",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bb6b40c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872b6",
   169 => x"b4088407",
   170 => x"b6b40c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb2f0",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfdfc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"b6b40852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"b69c0c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"81808051",
   203 => x"c0115170",
   204 => x"fb380284",
   205 => x"050d0402",
   206 => x"fc050d84",
   207 => x"bf5186a4",
   208 => x"2dff1151",
   209 => x"708025f6",
   210 => x"38028405",
   211 => x"0d0402fc",
   212 => x"050dec51",
   213 => x"83710c86",
   214 => x"a42d8271",
   215 => x"0c028405",
   216 => x"0d0402fc",
   217 => x"050dec51",
   218 => x"a2710c86",
   219 => x"a42d8271",
   220 => x"0c028405",
   221 => x"0d0402dc",
   222 => x"050d8059",
   223 => x"840bec0c",
   224 => x"a00bec0c",
   225 => x"7a52b6b8",
   226 => x"51a7812d",
   227 => x"b69c0879",
   228 => x"2e80eb38",
   229 => x"b6bc0879",
   230 => x"ff125659",
   231 => x"5673792e",
   232 => x"8b388118",
   233 => x"74812a55",
   234 => x"5873f738",
   235 => x"f7185881",
   236 => x"59807625",
   237 => x"80c83877",
   238 => x"52735184",
   239 => x"8b2db784",
   240 => x"52b6b851",
   241 => x"a9b72db6",
   242 => x"9c08802e",
   243 => x"9a38b784",
   244 => x"5783fc55",
   245 => x"76708405",
   246 => x"5808e80c",
   247 => x"fc155574",
   248 => x"8025f138",
   249 => x"87ee04b6",
   250 => x"9c085984",
   251 => x"8056b6b8",
   252 => x"51a98a2d",
   253 => x"fc801681",
   254 => x"15555687",
   255 => x"b104b6bc",
   256 => x"08f80c86",
   257 => x"b72d8051",
   258 => x"86e22d80",
   259 => x"5186ce2d",
   260 => x"78802e8d",
   261 => x"38b2f451",
   262 => x"8fdf2d8d",
   263 => x"e32d88a7",
   264 => x"04b3ec51",
   265 => x"8fdf2d78",
   266 => x"b69c0c02",
   267 => x"a4050d04",
   268 => x"02f0050d",
   269 => x"840bec0c",
   270 => x"8dc42d8a",
   271 => x"932d81f8",
   272 => x"2d83528d",
   273 => x"a92d8151",
   274 => x"84f02dff",
   275 => x"12527180",
   276 => x"25f13884",
   277 => x"0bec0cb0",
   278 => x"ec5185fe",
   279 => x"2d9e9e2d",
   280 => x"b69c0880",
   281 => x"2e819738",
   282 => x"810bfc0c",
   283 => x"b0fc5185",
   284 => x"fe2db194",
   285 => x"5186f62d",
   286 => x"86b72d86",
   287 => x"f651afbe",
   288 => x"2db2f451",
   289 => x"8fdf2d8d",
   290 => x"e32d8a9f",
   291 => x"2d8fef2d",
   292 => x"b3880b80",
   293 => x"f52db4d8",
   294 => x"08708106",
   295 => x"54555371",
   296 => x"802e8538",
   297 => x"72810753",
   298 => x"73812a70",
   299 => x"81065152",
   300 => x"71802e85",
   301 => x"38728207",
   302 => x"5373822a",
   303 => x"70810651",
   304 => x"5271802e",
   305 => x"85387284",
   306 => x"07537383",
   307 => x"2a708106",
   308 => x"51527180",
   309 => x"2e853872",
   310 => x"88075373",
   311 => x"842a7081",
   312 => x"06515271",
   313 => x"802e8538",
   314 => x"72900753",
   315 => x"72fc0c86",
   316 => x"52b69c08",
   317 => x"83388452",
   318 => x"71ec0c89",
   319 => x"8a04800b",
   320 => x"b69c0c02",
   321 => x"90050d04",
   322 => x"71980c04",
   323 => x"ffb008b6",
   324 => x"9c0c0481",
   325 => x"0bffb00c",
   326 => x"04800bff",
   327 => x"b00c0402",
   328 => x"f4050d8b",
   329 => x"a104b69c",
   330 => x"0881f02e",
   331 => x"09810689",
   332 => x"38810bb4",
   333 => x"d00c8ba1",
   334 => x"04b69c08",
   335 => x"81e02e09",
   336 => x"81068938",
   337 => x"810bb4d4",
   338 => x"0c8ba104",
   339 => x"b69c0852",
   340 => x"b4d40880",
   341 => x"2e8838b6",
   342 => x"9c088180",
   343 => x"05527184",
   344 => x"2c728f06",
   345 => x"5353b4d0",
   346 => x"08802e99",
   347 => x"38728429",
   348 => x"b4900572",
   349 => x"1381712b",
   350 => x"70097308",
   351 => x"06730c51",
   352 => x"53538b97",
   353 => x"04728429",
   354 => x"b4900572",
   355 => x"1383712b",
   356 => x"72080772",
   357 => x"0c535380",
   358 => x"0bb4d40c",
   359 => x"800bb4d0",
   360 => x"0cb6c451",
   361 => x"8ca22db6",
   362 => x"9c08ff24",
   363 => x"fef83880",
   364 => x"0bb69c0c",
   365 => x"028c050d",
   366 => x"0402f805",
   367 => x"0db49052",
   368 => x"8f518072",
   369 => x"70840554",
   370 => x"0cff1151",
   371 => x"708025f2",
   372 => x"38028805",
   373 => x"0d0402f0",
   374 => x"050d7551",
   375 => x"8a992d70",
   376 => x"822cfc06",
   377 => x"b4901172",
   378 => x"109e0671",
   379 => x"0870722a",
   380 => x"70830682",
   381 => x"742b7009",
   382 => x"7406760c",
   383 => x"54515657",
   384 => x"5351538a",
   385 => x"932d71b6",
   386 => x"9c0c0290",
   387 => x"050d0402",
   388 => x"fc050d72",
   389 => x"5180710c",
   390 => x"800b8412",
   391 => x"0c028405",
   392 => x"0d0402f0",
   393 => x"050d7570",
   394 => x"08841208",
   395 => x"535353ff",
   396 => x"5471712e",
   397 => x"a8388a99",
   398 => x"2d841308",
   399 => x"70842914",
   400 => x"88117008",
   401 => x"7081ff06",
   402 => x"84180881",
   403 => x"11870684",
   404 => x"1a0c5351",
   405 => x"55515151",
   406 => x"8a932d71",
   407 => x"5473b69c",
   408 => x"0c029005",
   409 => x"0d0402f8",
   410 => x"050d8a99",
   411 => x"2de00870",
   412 => x"8b2a7081",
   413 => x"06515252",
   414 => x"70802e9d",
   415 => x"38b6c408",
   416 => x"708429b6",
   417 => x"cc057381",
   418 => x"ff06710c",
   419 => x"5151b6c4",
   420 => x"08811187",
   421 => x"06b6c40c",
   422 => x"51800bb6",
   423 => x"ec0c8a8c",
   424 => x"2d8a932d",
   425 => x"0288050d",
   426 => x"0402fc05",
   427 => x"0d8a992d",
   428 => x"810bb6ec",
   429 => x"0c8a932d",
   430 => x"b6ec0851",
   431 => x"70fa3802",
   432 => x"84050d04",
   433 => x"02fc050d",
   434 => x"b6c4518c",
   435 => x"8f2d8bb9",
   436 => x"2d8ce651",
   437 => x"8a882d02",
   438 => x"84050d04",
   439 => x"b6f008b6",
   440 => x"9c0c0402",
   441 => x"fc050d8d",
   442 => x"ed048a9f",
   443 => x"2d87518b",
   444 => x"d62db69c",
   445 => x"08f43880",
   446 => x"da518bd6",
   447 => x"2db69c08",
   448 => x"e938b69c",
   449 => x"08b4dc0c",
   450 => x"b69c0851",
   451 => x"84f02d02",
   452 => x"84050d04",
   453 => x"02ec050d",
   454 => x"76548052",
   455 => x"870b8815",
   456 => x"80f52d56",
   457 => x"53747224",
   458 => x"8338a053",
   459 => x"725182f9",
   460 => x"2d81128b",
   461 => x"1580f52d",
   462 => x"54527272",
   463 => x"25de3802",
   464 => x"94050d04",
   465 => x"02f0050d",
   466 => x"b6f00854",
   467 => x"81f82d80",
   468 => x"0bb6f40c",
   469 => x"7308802e",
   470 => x"81803882",
   471 => x"0bb6b00c",
   472 => x"b6f4088f",
   473 => x"06b6ac0c",
   474 => x"73085271",
   475 => x"832e9638",
   476 => x"71832689",
   477 => x"3871812e",
   478 => x"af388fc5",
   479 => x"0471852e",
   480 => x"9f388fc5",
   481 => x"04881480",
   482 => x"f52d8415",
   483 => x"08b1a053",
   484 => x"545285fe",
   485 => x"2d718429",
   486 => x"13700852",
   487 => x"528fc904",
   488 => x"73518e94",
   489 => x"2d8fc504",
   490 => x"b4d80888",
   491 => x"15082c70",
   492 => x"81065152",
   493 => x"71802e87",
   494 => x"38b1a451",
   495 => x"8fc204b1",
   496 => x"a85185fe",
   497 => x"2d841408",
   498 => x"5185fe2d",
   499 => x"b6f40881",
   500 => x"05b6f40c",
   501 => x"8c14548e",
   502 => x"d4040290",
   503 => x"050d0471",
   504 => x"b6f00c8e",
   505 => x"c42db6f4",
   506 => x"08ff05b6",
   507 => x"f80c0402",
   508 => x"e8050db6",
   509 => x"f008b6fc",
   510 => x"08575587",
   511 => x"518bd62d",
   512 => x"b69c0881",
   513 => x"2a708106",
   514 => x"51527180",
   515 => x"2ea03890",
   516 => x"95048a9f",
   517 => x"2d87518b",
   518 => x"d62db69c",
   519 => x"08f438b4",
   520 => x"dc088132",
   521 => x"70b4dc0c",
   522 => x"70525284",
   523 => x"f02db4dc",
   524 => x"08903881",
   525 => x"fd518bd6",
   526 => x"2d81fa51",
   527 => x"8bd62d96",
   528 => x"a50480fe",
   529 => x"518bd62d",
   530 => x"b69c0880",
   531 => x"2ea63880",
   532 => x"0bb4dc0c",
   533 => x"805184f0",
   534 => x"2d90df04",
   535 => x"8a9f2d80",
   536 => x"fe518bd6",
   537 => x"2db69c08",
   538 => x"f338810b",
   539 => x"b4dc0c81",
   540 => x"5184f02d",
   541 => x"81f5518b",
   542 => x"d62db69c",
   543 => x"08812a70",
   544 => x"81065152",
   545 => x"71802eaf",
   546 => x"38b6f808",
   547 => x"5271802e",
   548 => x"8938ff12",
   549 => x"b6f80c91",
   550 => x"b704b6f4",
   551 => x"0810b6f4",
   552 => x"08057084",
   553 => x"29165152",
   554 => x"88120880",
   555 => x"2e8938ff",
   556 => x"51881208",
   557 => x"52712d81",
   558 => x"f2518bd6",
   559 => x"2db69c08",
   560 => x"812a7081",
   561 => x"06515271",
   562 => x"802eb138",
   563 => x"b6f408ff",
   564 => x"11b6f808",
   565 => x"56535373",
   566 => x"72258938",
   567 => x"8114b6f8",
   568 => x"0c91fc04",
   569 => x"72101370",
   570 => x"84291651",
   571 => x"52881208",
   572 => x"802e8938",
   573 => x"fe518812",
   574 => x"0852712d",
   575 => x"81fd518b",
   576 => x"d62db69c",
   577 => x"08812a70",
   578 => x"81065152",
   579 => x"71802ead",
   580 => x"38b6f808",
   581 => x"802e8938",
   582 => x"800bb6f8",
   583 => x"0c92bd04",
   584 => x"b6f40810",
   585 => x"b6f40805",
   586 => x"70842916",
   587 => x"51528812",
   588 => x"08802e89",
   589 => x"38fd5188",
   590 => x"12085271",
   591 => x"2d81fa51",
   592 => x"8bd62db6",
   593 => x"9c08812a",
   594 => x"70810651",
   595 => x"5271802e",
   596 => x"ae38b6f4",
   597 => x"08ff1154",
   598 => x"52b6f808",
   599 => x"73258838",
   600 => x"72b6f80c",
   601 => x"92ff0471",
   602 => x"10127084",
   603 => x"29165152",
   604 => x"88120880",
   605 => x"2e8938fc",
   606 => x"51881208",
   607 => x"52712db6",
   608 => x"f8087053",
   609 => x"5473802e",
   610 => x"8a388c15",
   611 => x"ff155555",
   612 => x"93850482",
   613 => x"0bb6b00c",
   614 => x"718f06b6",
   615 => x"ac0c81eb",
   616 => x"518bd62d",
   617 => x"b69c0881",
   618 => x"2a708106",
   619 => x"51527180",
   620 => x"2ead3874",
   621 => x"08852e09",
   622 => x"8106a438",
   623 => x"881580f5",
   624 => x"2dff0552",
   625 => x"71881681",
   626 => x"b72d7198",
   627 => x"2b527180",
   628 => x"25883880",
   629 => x"0b881681",
   630 => x"b72d7451",
   631 => x"8e942d81",
   632 => x"f4518bd6",
   633 => x"2db69c08",
   634 => x"812a7081",
   635 => x"06515271",
   636 => x"802eb338",
   637 => x"7408852e",
   638 => x"098106aa",
   639 => x"38881580",
   640 => x"f52d8105",
   641 => x"52718816",
   642 => x"81b72d71",
   643 => x"81ff068b",
   644 => x"1680f52d",
   645 => x"54527272",
   646 => x"27873872",
   647 => x"881681b7",
   648 => x"2d74518e",
   649 => x"942d80da",
   650 => x"518bd62d",
   651 => x"b69c0881",
   652 => x"2a708106",
   653 => x"51527180",
   654 => x"2e81a638",
   655 => x"b6f008b6",
   656 => x"f8085553",
   657 => x"73802e8a",
   658 => x"388c13ff",
   659 => x"15555394",
   660 => x"c4047208",
   661 => x"5271822e",
   662 => x"a6387182",
   663 => x"26893871",
   664 => x"812ea938",
   665 => x"95e10471",
   666 => x"832eb138",
   667 => x"71842e09",
   668 => x"810680ed",
   669 => x"38881308",
   670 => x"518fdf2d",
   671 => x"95e104b6",
   672 => x"f8085188",
   673 => x"13085271",
   674 => x"2d95e104",
   675 => x"810b8814",
   676 => x"082bb4d8",
   677 => x"0832b4d8",
   678 => x"0c95b704",
   679 => x"881380f5",
   680 => x"2d81058b",
   681 => x"1480f52d",
   682 => x"53547174",
   683 => x"24833880",
   684 => x"54738814",
   685 => x"81b72d8e",
   686 => x"c42d95e1",
   687 => x"04750880",
   688 => x"2ea23875",
   689 => x"08518bd6",
   690 => x"2db69c08",
   691 => x"81065271",
   692 => x"802e8b38",
   693 => x"b6f80851",
   694 => x"84160852",
   695 => x"712d8816",
   696 => x"5675da38",
   697 => x"8054800b",
   698 => x"b6b00c73",
   699 => x"8f06b6ac",
   700 => x"0ca05273",
   701 => x"b6f8082e",
   702 => x"09810698",
   703 => x"38b6f408",
   704 => x"ff057432",
   705 => x"70098105",
   706 => x"7072079f",
   707 => x"2a917131",
   708 => x"51515353",
   709 => x"715182f9",
   710 => x"2d811454",
   711 => x"8e7425c6",
   712 => x"38b4dc08",
   713 => x"5271b69c",
   714 => x"0c029805",
   715 => x"0d0402f4",
   716 => x"050dd452",
   717 => x"81ff720c",
   718 => x"71085381",
   719 => x"ff720c72",
   720 => x"882b83fe",
   721 => x"80067208",
   722 => x"7081ff06",
   723 => x"51525381",
   724 => x"ff720c72",
   725 => x"7107882b",
   726 => x"72087081",
   727 => x"ff065152",
   728 => x"5381ff72",
   729 => x"0c727107",
   730 => x"882b7208",
   731 => x"7081ff06",
   732 => x"7207b69c",
   733 => x"0c525302",
   734 => x"8c050d04",
   735 => x"02f4050d",
   736 => x"74767181",
   737 => x"ff06d40c",
   738 => x"5353b780",
   739 => x"08853871",
   740 => x"892b5271",
   741 => x"982ad40c",
   742 => x"71902a70",
   743 => x"81ff06d4",
   744 => x"0c517188",
   745 => x"2a7081ff",
   746 => x"06d40c51",
   747 => x"7181ff06",
   748 => x"d40c7290",
   749 => x"2a7081ff",
   750 => x"06d40c51",
   751 => x"d4087081",
   752 => x"ff065151",
   753 => x"82b8bf52",
   754 => x"7081ff2e",
   755 => x"09810694",
   756 => x"3881ff0b",
   757 => x"d40cd408",
   758 => x"7081ff06",
   759 => x"ff145451",
   760 => x"5171e538",
   761 => x"70b69c0c",
   762 => x"028c050d",
   763 => x"0402fc05",
   764 => x"0d81c751",
   765 => x"81ff0bd4",
   766 => x"0cff1151",
   767 => x"708025f4",
   768 => x"38028405",
   769 => x"0d0402f4",
   770 => x"050d81ff",
   771 => x"0bd40c93",
   772 => x"53805287",
   773 => x"fc80c151",
   774 => x"96fc2db6",
   775 => x"9c088b38",
   776 => x"81ff0bd4",
   777 => x"0c815398",
   778 => x"b30497ed",
   779 => x"2dff1353",
   780 => x"72df3872",
   781 => x"b69c0c02",
   782 => x"8c050d04",
   783 => x"02ec050d",
   784 => x"810bb780",
   785 => x"0c8454d0",
   786 => x"08708f2a",
   787 => x"70810651",
   788 => x"515372f3",
   789 => x"3872d00c",
   790 => x"97ed2db1",
   791 => x"ac5185fe",
   792 => x"2dd00870",
   793 => x"8f2a7081",
   794 => x"06515153",
   795 => x"72f33881",
   796 => x"0bd00cb1",
   797 => x"53805284",
   798 => x"d480c051",
   799 => x"96fc2db6",
   800 => x"9c08812e",
   801 => x"93387282",
   802 => x"2ebd38ff",
   803 => x"135372e5",
   804 => x"38ff1454",
   805 => x"73ffb038",
   806 => x"97ed2d83",
   807 => x"aa52849c",
   808 => x"80c85196",
   809 => x"fc2db69c",
   810 => x"08812e09",
   811 => x"81069238",
   812 => x"96ae2db6",
   813 => x"9c0883ff",
   814 => x"ff065372",
   815 => x"83aa2e9d",
   816 => x"3898862d",
   817 => x"99d804b1",
   818 => x"c05185fe",
   819 => x"2d80539b",
   820 => x"a604b1d8",
   821 => x"5185fe2d",
   822 => x"80549af8",
   823 => x"0481ff0b",
   824 => x"d40cb154",
   825 => x"97ed2d8f",
   826 => x"cf538052",
   827 => x"87fc80f7",
   828 => x"5196fc2d",
   829 => x"b69c0855",
   830 => x"b69c0881",
   831 => x"2e098106",
   832 => x"9b3881ff",
   833 => x"0bd40c82",
   834 => x"0a52849c",
   835 => x"80e95196",
   836 => x"fc2db69c",
   837 => x"08802e8d",
   838 => x"3897ed2d",
   839 => x"ff135372",
   840 => x"c9389aeb",
   841 => x"0481ff0b",
   842 => x"d40cb69c",
   843 => x"085287fc",
   844 => x"80fa5196",
   845 => x"fc2db69c",
   846 => x"08b13881",
   847 => x"ff0bd40c",
   848 => x"d4085381",
   849 => x"ff0bd40c",
   850 => x"81ff0bd4",
   851 => x"0c81ff0b",
   852 => x"d40c81ff",
   853 => x"0bd40c72",
   854 => x"862a7081",
   855 => x"06765651",
   856 => x"53729538",
   857 => x"b69c0854",
   858 => x"9af80473",
   859 => x"822efee2",
   860 => x"38ff1454",
   861 => x"73feed38",
   862 => x"73b7800c",
   863 => x"738b3881",
   864 => x"5287fc80",
   865 => x"d05196fc",
   866 => x"2d81ff0b",
   867 => x"d40cd008",
   868 => x"708f2a70",
   869 => x"81065151",
   870 => x"5372f338",
   871 => x"72d00c81",
   872 => x"ff0bd40c",
   873 => x"815372b6",
   874 => x"9c0c0294",
   875 => x"050d0402",
   876 => x"e8050d78",
   877 => x"55805681",
   878 => x"ff0bd40c",
   879 => x"d008708f",
   880 => x"2a708106",
   881 => x"51515372",
   882 => x"f3388281",
   883 => x"0bd00c81",
   884 => x"ff0bd40c",
   885 => x"775287fc",
   886 => x"80d15196",
   887 => x"fc2d80db",
   888 => x"c6df54b6",
   889 => x"9c08802e",
   890 => x"8a38b1fc",
   891 => x"5185fe2d",
   892 => x"9cc60481",
   893 => x"ff0bd40c",
   894 => x"d4087081",
   895 => x"ff065153",
   896 => x"7281fe2e",
   897 => x"0981069d",
   898 => x"3880ff53",
   899 => x"96ae2db6",
   900 => x"9c087570",
   901 => x"8405570c",
   902 => x"ff135372",
   903 => x"8025ed38",
   904 => x"81569cab",
   905 => x"04ff1454",
   906 => x"73c93881",
   907 => x"ff0bd40c",
   908 => x"81ff0bd4",
   909 => x"0cd00870",
   910 => x"8f2a7081",
   911 => x"06515153",
   912 => x"72f33872",
   913 => x"d00c75b6",
   914 => x"9c0c0298",
   915 => x"050d0402",
   916 => x"e8050d77",
   917 => x"797b5855",
   918 => x"55805372",
   919 => x"7625a338",
   920 => x"74708105",
   921 => x"5680f52d",
   922 => x"74708105",
   923 => x"5680f52d",
   924 => x"52527171",
   925 => x"2e863881",
   926 => x"519d8404",
   927 => x"8113539c",
   928 => x"db048051",
   929 => x"70b69c0c",
   930 => x"0298050d",
   931 => x"0402ec05",
   932 => x"0d765574",
   933 => x"802ebb38",
   934 => x"9a1580e0",
   935 => x"2d51aa8d",
   936 => x"2db69c08",
   937 => x"b69c08bd",
   938 => x"b40cb69c",
   939 => x"085454bd",
   940 => x"9008802e",
   941 => x"99389415",
   942 => x"80e02d51",
   943 => x"aa8d2db6",
   944 => x"9c08902b",
   945 => x"83fff00a",
   946 => x"06707507",
   947 => x"515372bd",
   948 => x"b40cbdb4",
   949 => x"08537280",
   950 => x"2e9938bd",
   951 => x"8808fe14",
   952 => x"7129bd9c",
   953 => x"0805bdb8",
   954 => x"0c70842b",
   955 => x"bd940c54",
   956 => x"9e9904bd",
   957 => x"a008bdb4",
   958 => x"0cbda408",
   959 => x"bdb80cbd",
   960 => x"9008802e",
   961 => x"8a38bd88",
   962 => x"08842b53",
   963 => x"9e9504bd",
   964 => x"a808842b",
   965 => x"5372bd94",
   966 => x"0c029405",
   967 => x"0d0402d8",
   968 => x"050d800b",
   969 => x"bd900c84",
   970 => x"5498bc2d",
   971 => x"b69c0880",
   972 => x"2e9538b7",
   973 => x"84528051",
   974 => x"9baf2db6",
   975 => x"9c08802e",
   976 => x"8638fe54",
   977 => x"9ecf04ff",
   978 => x"14547380",
   979 => x"24db3873",
   980 => x"8c38b290",
   981 => x"5185fe2d",
   982 => x"7355a3d8",
   983 => x"04805681",
   984 => x"0bbdbc0c",
   985 => x"8853b2a0",
   986 => x"52b7ba51",
   987 => x"9ccf2db6",
   988 => x"9c08762e",
   989 => x"09810687",
   990 => x"38b69c08",
   991 => x"bdbc0c88",
   992 => x"53b2ac52",
   993 => x"b7d6519c",
   994 => x"cf2db69c",
   995 => x"088738b6",
   996 => x"9c08bdbc",
   997 => x"0cbdbc08",
   998 => x"802e80f6",
   999 => x"38baca0b",
  1000 => x"80f52dba",
  1001 => x"cb0b80f5",
  1002 => x"2d71982b",
  1003 => x"71902b07",
  1004 => x"bacc0b80",
  1005 => x"f52d7088",
  1006 => x"2b7207ba",
  1007 => x"cd0b80f5",
  1008 => x"2d7107bb",
  1009 => x"820b80f5",
  1010 => x"2dbb830b",
  1011 => x"80f52d71",
  1012 => x"882b0753",
  1013 => x"5f54525a",
  1014 => x"56575573",
  1015 => x"81abaa2e",
  1016 => x"0981068d",
  1017 => x"387551a9",
  1018 => x"dd2db69c",
  1019 => x"08569ffe",
  1020 => x"047382d4",
  1021 => x"d52e8738",
  1022 => x"b2b851a0",
  1023 => x"bf04b784",
  1024 => x"5275519b",
  1025 => x"af2db69c",
  1026 => x"0855b69c",
  1027 => x"08802e83",
  1028 => x"c7388853",
  1029 => x"b2ac52b7",
  1030 => x"d6519ccf",
  1031 => x"2db69c08",
  1032 => x"8938810b",
  1033 => x"bd900ca0",
  1034 => x"c5048853",
  1035 => x"b2a052b7",
  1036 => x"ba519ccf",
  1037 => x"2db69c08",
  1038 => x"802e8a38",
  1039 => x"b2d05185",
  1040 => x"fe2da19f",
  1041 => x"04bb820b",
  1042 => x"80f52d54",
  1043 => x"7380d52e",
  1044 => x"09810680",
  1045 => x"ca38bb83",
  1046 => x"0b80f52d",
  1047 => x"547381aa",
  1048 => x"2e098106",
  1049 => x"ba38800b",
  1050 => x"b7840b80",
  1051 => x"f52d5654",
  1052 => x"7481e92e",
  1053 => x"83388154",
  1054 => x"7481eb2e",
  1055 => x"8c388055",
  1056 => x"73752e09",
  1057 => x"810682d0",
  1058 => x"38b78f0b",
  1059 => x"80f52d55",
  1060 => x"748d38b7",
  1061 => x"900b80f5",
  1062 => x"2d547382",
  1063 => x"2e863880",
  1064 => x"55a3d804",
  1065 => x"b7910b80",
  1066 => x"f52d70bd",
  1067 => x"880cff05",
  1068 => x"bd8c0cb7",
  1069 => x"920b80f5",
  1070 => x"2db7930b",
  1071 => x"80f52d58",
  1072 => x"76057782",
  1073 => x"80290570",
  1074 => x"bd980cb7",
  1075 => x"940b80f5",
  1076 => x"2d70bdac",
  1077 => x"0cbd9008",
  1078 => x"59575876",
  1079 => x"802e81a3",
  1080 => x"388853b2",
  1081 => x"ac52b7d6",
  1082 => x"519ccf2d",
  1083 => x"b69c0881",
  1084 => x"e738bd88",
  1085 => x"0870842b",
  1086 => x"bd940c70",
  1087 => x"bda80cb7",
  1088 => x"a90b80f5",
  1089 => x"2db7a80b",
  1090 => x"80f52d71",
  1091 => x"82802905",
  1092 => x"b7aa0b80",
  1093 => x"f52d7084",
  1094 => x"80802912",
  1095 => x"b7ab0b80",
  1096 => x"f52d7081",
  1097 => x"800a2912",
  1098 => x"70bdb00c",
  1099 => x"bdac0871",
  1100 => x"29bd9808",
  1101 => x"0570bd9c",
  1102 => x"0cb7b10b",
  1103 => x"80f52db7",
  1104 => x"b00b80f5",
  1105 => x"2d718280",
  1106 => x"2905b7b2",
  1107 => x"0b80f52d",
  1108 => x"70848080",
  1109 => x"2912b7b3",
  1110 => x"0b80f52d",
  1111 => x"70982b81",
  1112 => x"f00a0672",
  1113 => x"0570bda0",
  1114 => x"0cfe117e",
  1115 => x"297705bd",
  1116 => x"a40c5259",
  1117 => x"5243545e",
  1118 => x"51525952",
  1119 => x"5d575957",
  1120 => x"a3d104b7",
  1121 => x"960b80f5",
  1122 => x"2db7950b",
  1123 => x"80f52d71",
  1124 => x"82802905",
  1125 => x"70bd940c",
  1126 => x"70a02983",
  1127 => x"ff057089",
  1128 => x"2a70bda8",
  1129 => x"0cb79b0b",
  1130 => x"80f52db7",
  1131 => x"9a0b80f5",
  1132 => x"2d718280",
  1133 => x"290570bd",
  1134 => x"b00c7b71",
  1135 => x"291e70bd",
  1136 => x"a40c7dbd",
  1137 => x"a00c7305",
  1138 => x"bd9c0c55",
  1139 => x"5e515155",
  1140 => x"5580519d",
  1141 => x"8d2d8155",
  1142 => x"74b69c0c",
  1143 => x"02a8050d",
  1144 => x"0402ec05",
  1145 => x"0d767087",
  1146 => x"2c7180ff",
  1147 => x"06555654",
  1148 => x"bd90088a",
  1149 => x"3873882c",
  1150 => x"7481ff06",
  1151 => x"5455b784",
  1152 => x"52bd9808",
  1153 => x"15519baf",
  1154 => x"2db69c08",
  1155 => x"54b69c08",
  1156 => x"802eb338",
  1157 => x"bd900880",
  1158 => x"2e983872",
  1159 => x"8429b784",
  1160 => x"05700852",
  1161 => x"53a9dd2d",
  1162 => x"b69c08f0",
  1163 => x"0a0653a4",
  1164 => x"c4047210",
  1165 => x"b7840570",
  1166 => x"80e02d52",
  1167 => x"53aa8d2d",
  1168 => x"b69c0853",
  1169 => x"725473b6",
  1170 => x"9c0c0294",
  1171 => x"050d0402",
  1172 => x"e0050d79",
  1173 => x"70842cbd",
  1174 => x"b8080571",
  1175 => x"8f065255",
  1176 => x"53728938",
  1177 => x"b7845273",
  1178 => x"519baf2d",
  1179 => x"72a029b7",
  1180 => x"84055480",
  1181 => x"7480f52d",
  1182 => x"56537473",
  1183 => x"2e833881",
  1184 => x"537481e5",
  1185 => x"2e81ef38",
  1186 => x"81707406",
  1187 => x"54587280",
  1188 => x"2e81e338",
  1189 => x"8b1480f5",
  1190 => x"2d70832a",
  1191 => x"79065856",
  1192 => x"769838b4",
  1193 => x"e0085372",
  1194 => x"883872bb",
  1195 => x"840b81b7",
  1196 => x"2d76b4e0",
  1197 => x"0c7353a6",
  1198 => x"f804758f",
  1199 => x"2e098106",
  1200 => x"81b43874",
  1201 => x"9f068d29",
  1202 => x"baf71151",
  1203 => x"53811480",
  1204 => x"f52d7370",
  1205 => x"81055581",
  1206 => x"b72d8314",
  1207 => x"80f52d73",
  1208 => x"70810555",
  1209 => x"81b72d85",
  1210 => x"1480f52d",
  1211 => x"73708105",
  1212 => x"5581b72d",
  1213 => x"871480f5",
  1214 => x"2d737081",
  1215 => x"055581b7",
  1216 => x"2d891480",
  1217 => x"f52d7370",
  1218 => x"81055581",
  1219 => x"b72d8e14",
  1220 => x"80f52d73",
  1221 => x"70810555",
  1222 => x"81b72d90",
  1223 => x"1480f52d",
  1224 => x"73708105",
  1225 => x"5581b72d",
  1226 => x"921480f5",
  1227 => x"2d737081",
  1228 => x"055581b7",
  1229 => x"2d941480",
  1230 => x"f52d7370",
  1231 => x"81055581",
  1232 => x"b72d9614",
  1233 => x"80f52d73",
  1234 => x"70810555",
  1235 => x"81b72d98",
  1236 => x"1480f52d",
  1237 => x"73708105",
  1238 => x"5581b72d",
  1239 => x"9c1480f5",
  1240 => x"2d737081",
  1241 => x"055581b7",
  1242 => x"2d9e1480",
  1243 => x"f52d7381",
  1244 => x"b72d77b4",
  1245 => x"e00c8053",
  1246 => x"72b69c0c",
  1247 => x"02a0050d",
  1248 => x"0402cc05",
  1249 => x"0d7e605e",
  1250 => x"5a800bbd",
  1251 => x"b408bdb8",
  1252 => x"08595c56",
  1253 => x"8058bd94",
  1254 => x"08782e81",
  1255 => x"ae38778f",
  1256 => x"06a01757",
  1257 => x"54738f38",
  1258 => x"b7845276",
  1259 => x"51811757",
  1260 => x"9baf2db7",
  1261 => x"84568076",
  1262 => x"80f52d56",
  1263 => x"5474742e",
  1264 => x"83388154",
  1265 => x"7481e52e",
  1266 => x"80f63881",
  1267 => x"70750655",
  1268 => x"5c73802e",
  1269 => x"80ea388b",
  1270 => x"1680f52d",
  1271 => x"98065978",
  1272 => x"80de388b",
  1273 => x"537c5275",
  1274 => x"519ccf2d",
  1275 => x"b69c0880",
  1276 => x"cf389c16",
  1277 => x"0851a9dd",
  1278 => x"2db69c08",
  1279 => x"841b0c9a",
  1280 => x"1680e02d",
  1281 => x"51aa8d2d",
  1282 => x"b69c08b6",
  1283 => x"9c08881c",
  1284 => x"0cb69c08",
  1285 => x"5555bd90",
  1286 => x"08802e98",
  1287 => x"38941680",
  1288 => x"e02d51aa",
  1289 => x"8d2db69c",
  1290 => x"08902b83",
  1291 => x"fff00a06",
  1292 => x"70165154",
  1293 => x"73881b0c",
  1294 => x"787a0c7b",
  1295 => x"54a98104",
  1296 => x"811858bd",
  1297 => x"94087826",
  1298 => x"fed438bd",
  1299 => x"9008802e",
  1300 => x"ae387a51",
  1301 => x"a3e12db6",
  1302 => x"9c08b69c",
  1303 => x"0880ffff",
  1304 => x"fff80655",
  1305 => x"5b7380ff",
  1306 => x"fffff82e",
  1307 => x"9238b69c",
  1308 => x"08fe05bd",
  1309 => x"880829bd",
  1310 => x"9c080557",
  1311 => x"a7940480",
  1312 => x"5473b69c",
  1313 => x"0c02b405",
  1314 => x"0d0402f4",
  1315 => x"050d7470",
  1316 => x"08810571",
  1317 => x"0c7008bd",
  1318 => x"8c080653",
  1319 => x"53718e38",
  1320 => x"88130851",
  1321 => x"a3e12db6",
  1322 => x"9c088814",
  1323 => x"0c810bb6",
  1324 => x"9c0c028c",
  1325 => x"050d0402",
  1326 => x"f0050d75",
  1327 => x"881108fe",
  1328 => x"05bd8808",
  1329 => x"29bd9c08",
  1330 => x"117208bd",
  1331 => x"8c080605",
  1332 => x"79555354",
  1333 => x"549baf2d",
  1334 => x"0290050d",
  1335 => x"0402f405",
  1336 => x"0d747088",
  1337 => x"2a83fe80",
  1338 => x"06707298",
  1339 => x"2a077288",
  1340 => x"2b87fc80",
  1341 => x"80067398",
  1342 => x"2b81f00a",
  1343 => x"06717307",
  1344 => x"07b69c0c",
  1345 => x"56515351",
  1346 => x"028c050d",
  1347 => x"0402f805",
  1348 => x"0d028e05",
  1349 => x"80f52d74",
  1350 => x"882b0770",
  1351 => x"83ffff06",
  1352 => x"b69c0c51",
  1353 => x"0288050d",
  1354 => x"0402f405",
  1355 => x"0d747678",
  1356 => x"53545280",
  1357 => x"71259738",
  1358 => x"72708105",
  1359 => x"5480f52d",
  1360 => x"72708105",
  1361 => x"5481b72d",
  1362 => x"ff115170",
  1363 => x"eb388072",
  1364 => x"81b72d02",
  1365 => x"8c050d04",
  1366 => x"02e8050d",
  1367 => x"77568070",
  1368 => x"56547376",
  1369 => x"24b138bd",
  1370 => x"9408742e",
  1371 => x"aa387351",
  1372 => x"a4cf2db6",
  1373 => x"9c08b69c",
  1374 => x"08098105",
  1375 => x"70b69c08",
  1376 => x"079f2a77",
  1377 => x"05811757",
  1378 => x"57535374",
  1379 => x"76248838",
  1380 => x"bd940874",
  1381 => x"26d83872",
  1382 => x"b69c0c02",
  1383 => x"98050d04",
  1384 => x"02f0050d",
  1385 => x"b6980816",
  1386 => x"51aad82d",
  1387 => x"b69c0880",
  1388 => x"2e9b388b",
  1389 => x"53b69c08",
  1390 => x"52bb8451",
  1391 => x"aaa92dbd",
  1392 => x"c0085473",
  1393 => x"802e8638",
  1394 => x"bb845173",
  1395 => x"2d029005",
  1396 => x"0d0402dc",
  1397 => x"050d8070",
  1398 => x"5a5574b6",
  1399 => x"980825af",
  1400 => x"38bd9408",
  1401 => x"752ea838",
  1402 => x"7851a4cf",
  1403 => x"2db69c08",
  1404 => x"09810570",
  1405 => x"b69c0807",
  1406 => x"9f2a7605",
  1407 => x"811b5b56",
  1408 => x"5474b698",
  1409 => x"08258838",
  1410 => x"bd940879",
  1411 => x"26da3880",
  1412 => x"5578bd94",
  1413 => x"082781cd",
  1414 => x"387851a4",
  1415 => x"cf2db69c",
  1416 => x"08802e81",
  1417 => x"a238b69c",
  1418 => x"088b0580",
  1419 => x"f52d7084",
  1420 => x"2a708106",
  1421 => x"77107884",
  1422 => x"2bbb840b",
  1423 => x"80f52d5c",
  1424 => x"5c535155",
  1425 => x"5673802e",
  1426 => x"80c63874",
  1427 => x"16822bae",
  1428 => x"880bb4ec",
  1429 => x"120c5477",
  1430 => x"753110bd",
  1431 => x"c4115556",
  1432 => x"90747081",
  1433 => x"055681b7",
  1434 => x"2da07481",
  1435 => x"b72d7681",
  1436 => x"ff068116",
  1437 => x"58547380",
  1438 => x"2e89389c",
  1439 => x"53bb8452",
  1440 => x"ad89048b",
  1441 => x"53b69c08",
  1442 => x"52bdc616",
  1443 => x"51adbf04",
  1444 => x"7416822b",
  1445 => x"aba00bb4",
  1446 => x"ec120c54",
  1447 => x"7681ff06",
  1448 => x"81165854",
  1449 => x"73802e89",
  1450 => x"389c53bb",
  1451 => x"8452adb7",
  1452 => x"048b53b6",
  1453 => x"9c085277",
  1454 => x"753110bd",
  1455 => x"c4055176",
  1456 => x"55aaa92d",
  1457 => x"adda0474",
  1458 => x"90297531",
  1459 => x"7010bdc4",
  1460 => x"055154b6",
  1461 => x"9c087481",
  1462 => x"b72d8119",
  1463 => x"59748b24",
  1464 => x"a238ac91",
  1465 => x"04749029",
  1466 => x"75317010",
  1467 => x"bdc4058c",
  1468 => x"77315751",
  1469 => x"54807481",
  1470 => x"b72d9e14",
  1471 => x"ff165654",
  1472 => x"74f33802",
  1473 => x"a4050d04",
  1474 => x"02fc050d",
  1475 => x"b6980813",
  1476 => x"51aad82d",
  1477 => x"b69c0880",
  1478 => x"2e8838b6",
  1479 => x"9c08519d",
  1480 => x"8d2d800b",
  1481 => x"b6980cab",
  1482 => x"d22d8ec4",
  1483 => x"2d028405",
  1484 => x"0d0402fc",
  1485 => x"050d7251",
  1486 => x"70fd2ead",
  1487 => x"3870fd24",
  1488 => x"8a3870fc",
  1489 => x"2e80c438",
  1490 => x"af930470",
  1491 => x"fe2eb138",
  1492 => x"70ff2e09",
  1493 => x"8106bc38",
  1494 => x"b6980851",
  1495 => x"70802eb3",
  1496 => x"38ff11b6",
  1497 => x"980caf93",
  1498 => x"04b69808",
  1499 => x"f00570b6",
  1500 => x"980c5170",
  1501 => x"80259c38",
  1502 => x"800bb698",
  1503 => x"0caf9304",
  1504 => x"b6980881",
  1505 => x"05b6980c",
  1506 => x"af9304b6",
  1507 => x"98089005",
  1508 => x"b6980cab",
  1509 => x"d22d8ec4",
  1510 => x"2d028405",
  1511 => x"0d0402fc",
  1512 => x"050d800b",
  1513 => x"b6980cab",
  1514 => x"d22d8ddc",
  1515 => x"2db69c08",
  1516 => x"b6880cb4",
  1517 => x"e4518fdf",
  1518 => x"2d028405",
  1519 => x"0d0471bd",
  1520 => x"c00c0400",
  1521 => x"00ffffff",
  1522 => x"ff00ffff",
  1523 => x"ffff00ff",
  1524 => x"ffffff00",
  1525 => x"2020202a",
  1526 => x"556e416d",
  1527 => x"6967612a",
  1528 => x"20202000",
  1529 => x"20202020",
  1530 => x"20202020",
  1531 => x"20202020",
  1532 => x"20202000",
  1533 => x"5265696e",
  1534 => x"6963696f",
  1535 => x"00000000",
  1536 => x"45666563",
  1537 => x"746f2054",
  1538 => x"56000000",
  1539 => x"45666563",
  1540 => x"746f2043",
  1541 => x"6f6c6f72",
  1542 => x"00000000",
  1543 => x"496e6963",
  1544 => x"696f2052",
  1545 => x"61706964",
  1546 => x"6f000000",
  1547 => x"466f727a",
  1548 => x"6172204d",
  1549 => x"42433100",
  1550 => x"43617267",
  1551 => x"61722052",
  1552 => x"4f4d2047",
  1553 => x"42201000",
  1554 => x"53616c69",
  1555 => x"72000000",
  1556 => x"46616c6c",
  1557 => x"6f20656e",
  1558 => x"20524f4d",
  1559 => x"20696e69",
  1560 => x"6369616c",
  1561 => x"00000000",
  1562 => x"4f4b0000",
  1563 => x"44657465",
  1564 => x"6374616e",
  1565 => x"646f2053",
  1566 => x"440a0000",
  1567 => x"43617267",
  1568 => x"616e646f",
  1569 => x"20524f4d",
  1570 => x"20707269",
  1571 => x"6e636970",
  1572 => x"616c0a00",
  1573 => x"524f4d20",
  1574 => x"20202020",
  1575 => x"20474200",
  1576 => x"16200000",
  1577 => x"14200000",
  1578 => x"15200000",
  1579 => x"496e6963",
  1580 => x"69616e64",
  1581 => x"6f205344",
  1582 => x"2e2e2e0a",
  1583 => x"00000000",
  1584 => x"4572726f",
  1585 => x"7220616c",
  1586 => x"20696e69",
  1587 => x"63696172",
  1588 => x"20534421",
  1589 => x"0a000000",
  1590 => x"53444843",
  1591 => x"20657272",
  1592 => x"6f72210a",
  1593 => x"00000000",
  1594 => x"4572726f",
  1595 => x"72206465",
  1596 => x"20657363",
  1597 => x"72697475",
  1598 => x"72610a00",
  1599 => x"4572726f",
  1600 => x"72206465",
  1601 => x"206c6563",
  1602 => x"74757261",
  1603 => x"0a000000",
  1604 => x"4572726f",
  1605 => x"7220656e",
  1606 => x"2053440a",
  1607 => x"00000000",
  1608 => x"46415431",
  1609 => x"36202020",
  1610 => x"00000000",
  1611 => x"46415433",
  1612 => x"32202020",
  1613 => x"00000000",
  1614 => x"4e6f2068",
  1615 => x"61792070",
  1616 => x"61727469",
  1617 => x"63696f6e",
  1618 => x"2053440a",
  1619 => x"00000000",
  1620 => x"466f726d",
  1621 => x"61746f20",
  1622 => x"5344204d",
  1623 => x"616c6f0a",
  1624 => x"00000000",
  1625 => x"416e7465",
  1626 => x"72696f72",
  1627 => x"00000000",
  1628 => x"00000002",
  1629 => x"00000002",
  1630 => x"000017d4",
  1631 => x"00000000",
  1632 => x"00000002",
  1633 => x"000017e4",
  1634 => x"00000000",
  1635 => x"00000002",
  1636 => x"000017f4",
  1637 => x"0000034e",
  1638 => x"00000001",
  1639 => x"00001800",
  1640 => x"00000001",
  1641 => x"00000001",
  1642 => x"0000180c",
  1643 => x"00000002",
  1644 => x"00000001",
  1645 => x"0000181c",
  1646 => x"00000003",
  1647 => x"00000001",
  1648 => x"0000182c",
  1649 => x"00000004",
  1650 => x"00000002",
  1651 => x"00001838",
  1652 => x"0000179e",
  1653 => x"00000002",
  1654 => x"00001848",
  1655 => x"000006e3",
  1656 => x"00000000",
  1657 => x"00000000",
  1658 => x"00000000",
  1659 => x"00000004",
  1660 => x"00001850",
  1661 => x"000019ec",
  1662 => x"00000004",
  1663 => x"00001868",
  1664 => x"00001974",
  1665 => x"00000000",
  1666 => x"00000000",
  1667 => x"00000000",
  1668 => x"00000000",
  1669 => x"00000000",
  1670 => x"00000000",
  1671 => x"00000000",
  1672 => x"00000000",
  1673 => x"00000000",
  1674 => x"00000000",
  1675 => x"00000000",
  1676 => x"00000000",
  1677 => x"00000000",
  1678 => x"00000000",
  1679 => x"00000000",
  1680 => x"00000000",
  1681 => x"00000000",
  1682 => x"00000000",
  1683 => x"00000000",
  1684 => x"00000000",
  1685 => x"00000000",
  1686 => x"00000000",
  1687 => x"00000000",
  1688 => x"00000000",
  1689 => x"00000002",
  1690 => x"00001ec4",
  1691 => x"000015a0",
  1692 => x"00000002",
  1693 => x"00001ee2",
  1694 => x"000015a0",
  1695 => x"00000002",
  1696 => x"00001f00",
  1697 => x"000015a0",
  1698 => x"00000002",
  1699 => x"00001f1e",
  1700 => x"000015a0",
  1701 => x"00000002",
  1702 => x"00001f3c",
  1703 => x"000015a0",
  1704 => x"00000002",
  1705 => x"00001f5a",
  1706 => x"000015a0",
  1707 => x"00000002",
  1708 => x"00001f78",
  1709 => x"000015a0",
  1710 => x"00000002",
  1711 => x"00001f96",
  1712 => x"000015a0",
  1713 => x"00000002",
  1714 => x"00001fb4",
  1715 => x"000015a0",
  1716 => x"00000002",
  1717 => x"00001fd2",
  1718 => x"000015a0",
  1719 => x"00000002",
  1720 => x"00001ff0",
  1721 => x"000015a0",
  1722 => x"00000002",
  1723 => x"0000200e",
  1724 => x"000015a0",
  1725 => x"00000002",
  1726 => x"0000202c",
  1727 => x"000015a0",
  1728 => x"00000004",
  1729 => x"00001964",
  1730 => x"00000000",
  1731 => x"00000000",
  1732 => x"00000000",
  1733 => x"00001732",
  1734 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;