module LATCHS_primitive_inst_old(D, G, R, Q);
  input D;
  input G;
  output Q;
  input R;

LATCHS inst (.*);

endmodule
