module ram_simple_dp_synch_wf_readmem_1024x32 (clk, we,re, read_addr, write_addr, din, dout);
    input clk, we, re;
    input [9:0] read_addr, write_addr;
    input [31:0] din;
    `ifdef IVERILOG
         output reg [31:0] dout=0;
    `else
        output reg [31:0] dout;
    `endif
    
    reg [31:0] ram [1023:0];

    initial begin
         $readmemh("mem.init", ram);
    end
    
    always @(posedge clk)
    begin
        if (we)
            ram[write_addr] <= din;
        if (re) begin
            dout <= ram[read_addr];
            if (we && read_addr == write_addr)
                dout <= din;
        end
    end

endmodule