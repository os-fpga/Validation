module puz_bank3 (clk,index,masked,to_check,match);
input clk;
input [7:0] index;
output [323:0] masked;
wire [323:0] masked;
input tri [323:0] to_check;
output match;

reg[15:0] soln_sig;
reg[15:0] soln_sig_r;
reg[15:0] check_sig;
reg[323:0] clue;

assign masked = clue;
function [15:0] signature;
  input [323:0] puz;
  reg [15:0] tmp;
  begin
    tmp[0] = puz[279]^puz[179]^puz[61]^puz[42]^puz[161]^puz[167]^puz[291]^puz[122]^puz[280]^puz[271]^puz[24]^puz[176]^puz[266]^puz[65]^puz[186]^puz[4];
    tmp[1] = puz[166]^puz[240]^puz[104]^puz[68]^puz[1]^puz[210]^puz[318]^puz[80]^puz[303]^puz[279]^puz[87]^puz[169]^puz[301]^puz[123]^puz[214]^puz[243];
    tmp[2] = puz[10]^puz[83]^puz[114]^puz[178]^puz[295]^puz[70]^puz[205]^puz[271]^puz[15]^puz[81]^puz[311]^puz[72]^puz[115]^puz[175]^puz[162]^puz[16];
    tmp[3] = puz[278]^puz[11]^puz[232]^puz[232]^puz[49]^puz[59]^puz[124]^puz[15]^puz[253]^puz[230]^puz[122]^puz[246]^puz[145]^puz[127]^puz[306]^puz[255];
    tmp[4] = puz[142]^puz[160]^puz[163]^puz[234]^puz[163]^puz[162]^puz[141]^puz[38]^puz[282]^puz[58]^puz[299]^puz[131]^puz[96]^puz[312]^puz[184]^puz[269];
    tmp[5] = puz[312]^puz[202]^puz[180]^puz[212]^puz[79]^puz[208]^puz[243]^puz[19]^puz[138]^puz[163]^puz[198]^puz[321]^puz[77]^puz[131]^puz[9]^puz[34];
    tmp[6] = puz[295]^puz[64]^puz[124]^puz[188]^puz[210]^puz[306]^puz[81]^puz[122]^puz[280]^puz[57]^puz[145]^puz[213]^puz[161]^puz[197]^puz[38]^puz[72];
    tmp[7] = puz[23]^puz[314]^puz[68]^puz[212]^puz[248]^puz[178]^puz[159]^puz[289]^puz[215]^puz[5]^puz[301]^puz[211]^puz[226]^puz[150]^puz[279]^puz[237];
    tmp[8] = puz[258]^puz[157]^puz[217]^puz[294]^puz[215]^puz[240]^puz[130]^puz[24]^puz[113]^puz[122]^puz[309]^puz[45]^puz[203]^puz[200]^puz[274]^puz[44];
    tmp[9] = puz[203]^puz[270]^puz[84]^puz[129]^puz[239]^puz[290]^puz[315]^puz[232]^puz[303]^puz[154]^puz[25]^puz[160]^puz[247]^puz[264]^puz[12]^puz[187];
    tmp[10] = puz[29]^puz[57]^puz[142]^puz[28]^puz[266]^puz[27]^puz[187]^puz[179]^puz[290]^puz[28]^puz[171]^puz[240]^puz[97]^puz[95]^puz[270]^puz[291];
    tmp[11] = puz[17]^puz[269]^puz[264]^puz[227]^puz[264]^puz[70]^puz[304]^puz[150]^puz[22]^puz[89]^puz[198]^puz[131]^puz[0]^puz[129]^puz[272]^puz[321];
    tmp[12] = puz[295]^puz[46]^puz[34]^puz[267]^puz[155]^puz[59]^puz[142]^puz[280]^puz[189]^puz[301]^puz[63]^puz[306]^puz[115]^puz[172]^puz[124]^puz[281];
    tmp[13] = puz[224]^puz[201]^puz[19]^puz[225]^puz[64]^puz[127]^puz[118]^puz[200]^puz[177]^puz[170]^puz[202]^puz[193]^puz[125]^puz[113]^puz[194]^puz[154];
    tmp[14] = puz[181]^puz[267]^puz[71]^puz[267]^puz[27]^puz[40]^puz[89]^puz[219]^puz[9]^puz[120]^puz[164]^puz[310]^puz[190]^puz[317]^puz[292]^puz[139];
    tmp[15] = puz[0]^puz[97]^puz[142]^puz[168]^puz[98]^puz[146]^puz[149]^puz[140]^puz[118]^puz[165]^puz[175]^puz[1]^puz[127]^puz[28]^puz[67]^puz[227];
    signature = tmp;
  end
endfunction

// Match comparator - latency one
//  so the signatures can go in ROM
always @(posedge clk) begin
  soln_sig_r <= soln_sig;
  check_sig <= signature (to_check);
end
assign match = (check_sig == soln_sig_r);

always @(index) begin
	case (index)
      0 : begin
         soln_sig = signature(324'h897561423_436297851_251843769_342175698_769384215_518926347_975632184_683419572_124758936);
         // Rules : HARD derived
         clue = 324'h000000000_000007851_050040000_042100090_009080005_010906300_070630000_600009000_120700000;
          // 25 clues
       end
      1 : begin
         soln_sig = signature(324'h417926538_325478961_698135742_762593184_539841627_184267359_951382476_873614295_246759813);
         // Rules : HARD
         clue = 324'h000000000_000078060_000105700_700000004_030040000_180260059_000000000_873004095_200000803;
          // 25 clues
       end
      2 : begin
         soln_sig = signature(324'h478532619_695781423_123694857_857469132_234157968_961823574_782915346_549376281_316248795);
         // Rules : HARD derived
         clue = 324'h000000000_000080423_020600000_007400002_030057900_061003070_080905000_500070000_310008000;
          // 25 clues
       end
      3 : begin
         soln_sig = signature(324'h274568139_381924657_569173428_792485316_458316792_136792584_617839245_943257861_825641973);
         // Rules : HARD derived
         clue = 324'h000000000_000904050_000170400_790085016_400000002_030002000_000000000_943200061_800000903;
          // 25 clues
       end
      4 : begin
         soln_sig = signature(324'h256798431_971463825_384152796_627945183_819376542_435281967_548627319_192534678_763819254);
         // Rules : HARD derived
         clue = 324'h000000000_001403805_000000096_000900180_800000000_035001900_040027000_000030600_700800050;
          // 23 clues
       end
      5 : begin
         soln_sig = signature(324'h687539241_134287956_259614783_765391824_398742615_412856379_926175438_573468192_841923567);
         // Rules : MEDIUM derived
         clue = 324'h000000000_004280006_009610000_000300020_300040005_002006079_000005038_070000190_001000000;
          // 23 clues
       end
      6 : begin
         soln_sig = signature(324'h265941387_718536942_349827561_873264159_524719638_196358274_932475816_451682793_687193425);
         // Rules : MEDIUM derived
         clue = 324'h000000000_008036002_009027000_003200059_000010030_100008004_000400016_050000790_007000000;
          // 23 clues
       end
      7 : begin
         soln_sig = signature(324'h291364578_348175629_765928431_683417952_579682314_124593867_956241783_832759146_417836295);
         // Rules : HARD derived
         clue = 324'h000000000_008075609_000000031_600000000_079080300_000003860_050240000_000700100_400006090;
          // 23 clues
       end
      8 : begin
         soln_sig = signature(324'h613892457_827354961_549167238_931275684_268413795_754689123_176528349_482931576_395746812);
         // Rules : HARD derived
         clue = 324'h000000000_020000961_509007000_901000004_008003000_000600023_100008000_082000506_000740800;
          // 24 clues
       end
      9 : begin
         soln_sig = signature(324'h631492875_429578316_758361249_582916734_197243658_346785192_265139487_973824561_814657923);
         // Rules : MEDIUM derived
         clue = 324'h000000000_020570000_000001009_500000034_007200000_040080190_005130080_903004060_004000000;
          // 23 clues
       end
      10 : begin
         soln_sig = signature(324'h735462918_429871653_618593472_543287169_291634785_876159324_362745891_184926537_957318246);
         // Rules : EASY derived
         clue = 324'h000000000_029070600_600093000_503007060_200030005_800109024_300000001_080020007_050000040;
          // 26 clues
       end
      11 : begin
         soln_sig = signature(324'h628917453_359426781_417385296_763159824_541278369_982634517_296843175_135792648_874561932);
         // Rules : EASY derived
         clue = 324'h000000000_050400000_000005296_060000000_001070369_002004007_200000170_030700000_000560002;
          // 23 clues
       end
      12 : begin
         soln_sig = signature(324'h357862149_261349875_849157236_614528397_938714562_725936481_586273914_492681753_173495628);
         // Rules : EASY derived
         clue = 324'h000000000_061300800_800150000_600500007_900014062_705030080_500000004_090600003_070000020;
          // 26 clues
       end
      13 : begin
         soln_sig = signature(324'h613897452_982435761_547216839_254769183_731582694_869341275_126958347_498173526_375624918);
         // Rules : HARD derived
         clue = 324'h000000000_080000761_507200000_000060083_701000004_009300000_100900000_098000506_000024900;
          // 24 clues
       end
      14 : begin
         soln_sig = signature(324'h186547392_294138567_375926841_468312975_512479683_937685214_841263759_729854136_653791428);
         // Rules : EASY derived
         clue = 324'h000000000_090030000_000900841_008300005_010000000_007005214_800000750_020050000_000091008;
          // 23 clues
       end
      15 : begin
         soln_sig = signature(324'h548197326_791236485_263584971_812749563_475362819_639851247_956418732_124973658_387625194);
         // Rules : MEDIUM derived
         clue = 324'h000000000_090206000_000080001_002009000_070300810_600000047_006408030_104070050_007000000;
          // 23 clues
       end
      16 : begin
         soln_sig = signature(324'h972485631_165372894_348691725_697528413_283147956_514963287_756219348_839754162_421836579);
         // Rules : HARD derived
         clue = 324'h000000000_105070090_008600005_000500413_003007050_004900200_006019040_830000002_000030009;
          // 26 clues
       end
      17 : begin
         soln_sig = signature(324'h754832691_168495273_932167548_813976425_675284319_429513786_586741932_297358164_341629857);
         // Rules : HARD derived
         clue = 324'h000000000_108005070_002060008_003070400_000080319_009500080_006701030_290000004_000009007;
          // 26 clues
       end
      18 : begin
         soln_sig = signature(324'h186954372_257163948_943287165_534618729_791325684_628479531_475831296_812796453_369542817);
         // Rules : HARD derived
         clue = 324'h000000000_250000900_040207000_000600000_701300080_020470031_005000000_010796003_360002800;
          // 26 clues
       end
      19 : begin
         soln_sig = signature(324'h618735429_534289176_792614358_329871645_465392781_187456293_876943512_953127864_241568937);
         // Rules : HARD derived
         clue = 324'h000000000_530000070_092600358_029071045_060000080_000006003_800940000_000000000_001508000;
          // 25 clues
       end
      20 : begin
         soln_sig = signature(324'h612439785_548276931_937185624_896547213_251893476_473612859_384761592_165928347_729354168);
         // Rules : HARD derived
         clue = 324'h000000000_540000900_030085000_806007010_050803076_000002000_004000000_060928007_720050100;
          // 26 clues
       end
      21 : begin
         soln_sig = signature(324'h874659321_563412798_912738654_385126947_749583216_621974835_498361572_156297483_237845169);
         // Rules : HARD derived
         clue = 324'h000000000_560000090_012008654_080000040_000080006_021970035_400301000_000000000_007045000;
          // 25 clues
       end
      22 : begin
         soln_sig = signature(324'h876459321_312867549_459231687_963174258_728395416_145628973_281943765_594786132_637512894);
         // Rules : EASY derived
         clue = 324'h000000001_000060040_450000007_903004000_008090010_000600003_201000060_000086030_007500800;
          // 23 clues
       end
      23 : begin
         soln_sig = signature(324'h653819472_714362598_982745361_147528639_829637145_536194827_391256784_268471953_475983216);
         // Rules : EASY derived
         clue = 324'h000000002_704060000_080700360_000008030_000030005_030100020_000206704_008001900_005000000;
          // 23 clues
       end
      24 : begin
         soln_sig = signature(324'h498562173_631789245_527413698_869174352_273695814_154238967_945321786_782946531_316857429);
         // Rules : MEDIUM derived
         clue = 324'h000000003_000709000_507000600_060004050_003090000_004208900_900000080_780046001_010800020;
          // 25 clues
       end
      25 : begin
         soln_sig = signature(324'h973621854_126548379_548397621_354962718_812475936_697183245_465239187_731856492_289714563);
         // Rules : HARD derived
         clue = 324'h000000004_006008070_000397000_000000000_012000930_690000000_005239180_700056002_000010000;
          // 24 clues
       end
      26 : begin
         soln_sig = signature(324'h281743695_659182734_374659128_892476351_537921486_416835972_925364817_743218569_168597243);
         // Rules : EASY derived
         clue = 324'h000000005_000100030_370000008_002400050_000001006_406030000_905000010_000210060_008007200;
          // 23 clues
       end
      27 : begin
         soln_sig = signature(324'h947813265_831265749_652479138_194782356_765391482_283654971_516937824_478126593_329548617);
         // Rules : HARD derived
         clue = 324'h000000005_001200040_000479000_190000000_000000000_083000970_006937820_400106003_000008000;
          // 24 clues
       end
      28 : begin
         soln_sig = signature(324'h938627145_471589362_625341897_389176254_714235986_256498713_867953421_592714638_143862579);
         // Rules : EASY derived
         clue = 324'h000000005_401009000_020040890_080070050_000200080_000008003_000950401_002700600_003000000;
          // 23 clues
       end
      29 : begin
         soln_sig = signature(324'h318742956_769815432_245963718_456127893_923684175_871539624_132496587_584371269_697258341);
         // Rules : MEDIUM derived
         clue = 324'h000000006_000015000_205000700_006100000_003084100_070030020_100000080_580370009_090008040;
          // 25 clues
       end
      30 : begin
         soln_sig = signature(324'h745368912_126954837_938712465_397846251_462195783_581273694_259637148_814529376_673481529);
         // Rules : HARD derived
         clue = 324'h000000010_000950007_900002005_300840001_060000700_080203090_050600108_004000070_070000020;
          // 25 clues
       end
      31 : begin
         soln_sig = signature(324'h258469317_764123985_391587642_973651428_546872139_182934576_627315894_819746253_435298761);
         // Rules : MEDIUM derived
         clue = 324'h000000010_060003000_390500002_003001420_046072100_000930000_007310804_800006000_000000701;
          // 27 clues
       end
      32 : begin
         soln_sig = signature(324'h968752413_372941586_451836729_627398145_189425637_534617298_793164852_815273964_246589371);
         // Rules : MEDIUM derived
         clue = 324'h000000010_070040000_450006009_027390100_000405000_004010290_003104802_800070000_000000301;
          // 27 clues
       end
      33 : begin
         soln_sig = signature(324'h569738214_742915683_183462759_851293476_637854921_294176538_928541367_416327895_375689142);
         // Rules : MEDIUM derived
         clue = 324'h000000014_000900000_183000000_000203000_600850000_290000030_000500307_416020805_000600100;
          // 25 clues
       end
      34 : begin
         soln_sig = signature(324'h926483715_357196284_184275396_243958671_765321948_891647532_678519423_512734869_439862157);
         // Rules : MEDIUM derived
         clue = 324'h000000015_000006000_184000000_200908000_760000040_000047000_000009403_512700809_000002100;
          // 25 clues
       end
      35 : begin
         soln_sig = signature(324'h278641539_341597628_596238174_163759842_785324961_924186357_857962413_432815796_619473285);
         // Rules : MEDIUM derived
         clue = 324'h000000030_040097600_000208170_063050000_000004900_024100000_057002003_000010000_000000080;
          // 23 clues
       end
      36 : begin
         soln_sig = signature(324'h821694537_356271498_749385261_138726954_564139782_297458613_415867329_982543176_673912845);
         // Rules : MEDIUM derived
         clue = 324'h000000030_350070000_009000201_038000054_000009700_000050000_005800020_900003070_600912000;
          // 24 clues
       end
      37 : begin
         soln_sig = signature(324'h274859631_386127945_519346827_145962783_837415296_692783514_961538472_753294168_428671359);
         // Rules : MEDIUM derived
         clue = 324'h000000031_000020005_009300800_100960000_807005200_090080014_060008402_700000060_008001000;
          // 26 clues
       end
      38 : begin
         soln_sig = signature(324'h328956741_419827563_765413298_291784356_854361972_673295184_187639425_542178639_936542817);
         // Rules : HARD derived
         clue = 324'h000000040_000807003_700010008_090000300_050061070_600205004_080009405_002000030_030000010;
          // 25 clues
       end
      39 : begin
         soln_sig = signature(324'h896317542_375642918_421895367_548729136_937561284_162438795_659174823_284953671_713286459);
         // Rules : HARD derived
         clue = 324'h000000042_005600000_020800307_000700100_900060000_002038005_000000803_204050601_003200000;
          // 25 clues
       end
      40 : begin
         soln_sig = signature(324'h869372451_274519638_513648297_627934185_391285764_458167329_946753812_185426973_732891546);
         // Rules : HARD derived
         clue = 324'h000000051_004009000_010008207_600900000_001280004_000007300_000000802_105400903_002001000;
          // 25 clues
       end
      41 : begin
         soln_sig = signature(324'h356891472_794523861_128476935_483759126_261384597_975162384_842917653_517638249_639245718);
         // Rules : MEDIUM derived
         clue = 324'h000000072_000003001_008070900_080009026_200084000_905100300_040900603_500000040_009200000;
          // 26 clues
       end
      42 : begin
         soln_sig = signature(324'h481692573_325178649_697534821_569417382_174823956_238956417_752349168_946781235_813265794);
         // Rules : EASY derived
         clue = 324'h000000073_020000640_690530000_560000082_004000950_008000007_700300068_000781000_000005000;
          // 26 clues
       end
      43 : begin
         soln_sig = signature(324'h182654379_953782416_467913852_271598634_598346127_346271985_735169248_614827593_829435761);
         // Rules : EASY derived
         clue = 324'h000000079_050000410_460903000_001000630_008000007_340000085_700009048_000827000_000030000;
          // 26 clues
       end
      44 : begin
         soln_sig = signature(324'h459613287_836527149_271948653_743169825_618752934_592384716_925471368_384296571_167835492);
         // Rules : MEDIUM derived
         clue = 324'h000000080_030507100_000940650_043060000_018002000_000300700_025400008_000006000_000000090;
          // 23 clues
       end
      45 : begin
         soln_sig = signature(324'h197653284_385742961_264819735_721368459_439125876_856974123_548296317_613487592_972531648);
         // Rules : HARD derived
         clue = 324'h000000080_305002000_004810700_001008409_030000876_006004020_000090000_600400000_900031000;
          // 25 clues
       end
      46 : begin
         soln_sig = signature(324'h782356491_593142867_461789253_158437926_936218745_247695138_319864572_675921384_824573619);
         // Rules : HARD derived
         clue = 324'h000000090_503040000_001709200_050000926_006010040_007090108_000800000_600001000_800570000;
          // 25 clues
       end
      47 : begin
         soln_sig = signature(324'h453128796_972356184_618794523_586417239_394265871_721839645_137642958_845971362_269583417);
         // Rules : MEDIUM derived
         clue = 324'h000000090_970006000_008000503_000007000_094000071_000800600_007040050_800900060_200583000;
          // 24 clues
       end
      48 : begin
         soln_sig = signature(324'h825694137_397152684_614387925_461239578_259478361_783561249_572943816_146825793_938716452);
         // Rules : HARD derived
         clue = 324'h000000100_300002080_014000000_400030070_209070000_080061240_070040016_000800000_900700002;
          // 25 clues
       end
      49 : begin
         soln_sig = signature(324'h968345127_123769845_574182693_759421368_416837259_382956471_847693512_695218734_231574986);
         // Rules : EASY derived
         clue = 324'h000000120_000060800_504000000_059001000_400000200_002006471_007000000_090200730_200504080;
          // 25 clues
       end
      50 : begin
         soln_sig = signature(324'h376519248_542386971_819427635_498231756_257648319_163975824_925163487_731894562_684752193);
         // Rules : HARD derived
         clue = 324'h000000208_500306071_000000000_000200750_007000000_160005020_000060080_030094000_004700100;
          // 23 clues
       end
      51 : begin
         soln_sig = signature(324'h147563298_692718543_835492716_371654829_958321467_264879135_526137984_413985672_789246351);
         // Rules : HARD derived
         clue = 324'h000000208_600710043_000000000_370600020_000020460_004000000_000007080_010905000_009040300;
          // 23 clues
       end
      52 : begin
         soln_sig = signature(324'h946138275_821574639_573926418_739842561_618759324_254361897_192685743_365497182_487213956);
         // Rules : MEDIUM derived
         clue = 324'h000000275_800000630_500020000_000002000_010709304_000300090_002000040_005490080_007010050;
          // 25 clues
       end
      53 : begin
         soln_sig = signature(324'h157486293_962573841_834219576_428951367_793862154_516734982_689127435_275348619_341695728);
         // Rules : HARD derived
         clue = 324'h000000290_000503000_830009000_000901007_003000050_010704080_600020030_205008000_000600008;
          // 24 clues
       end
      54 : begin
         soln_sig = signature(324'h751824396_268391475_493675812_987436251_514287639_632519784_349168527_126753948_875942163);
         // Rules : MEDIUM derived
         clue = 324'h000000300_200090005_490075000_900006200_510200009_000000080_000008020_006003000_805040060;
          // 24 clues
       end
      55 : begin
         soln_sig = signature(324'h873961452_216754389_594823167_935176824_187542693_462398571_659437218_321689745_748215936);
         // Rules : HARD derived
         clue = 324'h000000400_010750000_090803060_000076000_100002090_000008500_600030008_300000705_008010006;
          // 24 clues
       end
      56 : begin
         soln_sig = signature(324'h936725481_127843695_854169273_293418756_471596832_568372914_785634129_612957348_349281567);
         // Rules : HARD derived
         clue = 324'h000000400_020803000_050069070_200010050_000090800_000370000_700600009_600000308_009200007;
          // 24 clues
       end
      57 : begin
         soln_sig = signature(324'h183529476_457816329_692743518_861392745_924657183_375481962_718235694_546978231_239164857);
         // Rules : MEDIUM derived
         clue = 324'h000000400_050016320_090000508_001002005_000000000_005400902_718035000_000900030_039060000;
          // 26 clues
       end
      58 : begin
         soln_sig = signature(324'h756913428_438562197_129748356_812496573_543871962_967235841_685124739_294387615_371659284);
         // Rules : EASY derived
         clue = 324'h000000420_030000007_000040000_002000073_000071060_900005001_005024700_090007010_301050200;
          // 25 clues
       end
      59 : begin
         soln_sig = signature(324'h796153482_245986173_318427695_483572961_562819347_179364528_924735816_837641259_651298734);
         // Rules : MEDIUM
         clue = 324'h000000480_200006000_010007005_000500900_000010000_079300020_004705006_800041009_050208030;
          // 26 clues
       end
      60 : begin
         soln_sig = signature(324'h917638524_362954718_548172963_826417359_139285647_475396182_683721495_751849236_294563871);
         // Rules : EASY derived
         clue = 324'h000000500_002904010_508100003_000007309_100000040_475006100_000000490_701000000_200060000;
          // 25 clues
       end
      61 : begin
         soln_sig = signature(324'h687231594_394756182_125498763_876129435_549367218_231845976_762984351_418573629_953612847);
         // Rules : MEDIUM derived
         clue = 324'h000000504_090050080_020400003_870009000_000360200_001000000_000904000_008070600_000012007;
          // 23 clues
       end
      62 : begin
         soln_sig = signature(324'h917346528_245781369_386925174_728453916_194867235_653192847_432579681_571638492_869214753);
         // Rules : HARD derived
         clue = 324'h000000520_000081000_380020000_008000010_090067030_000092007_400500080_501030000_000004003;
          // 24 clues
       end
      63 : begin
         soln_sig = signature(324'h948723561_562914837_713658492_286497315_179536248_354182679_831249756_497865123_625371984);
         // Rules : EASY derived
         clue = 324'h000000560_000004800_703000000_006400315_079500000_300000600_001000000_090060120_600370080;
          // 25 clues
       end
      64 : begin
         soln_sig = signature(324'h725394681_984126375_163758249_246831957_579462813_831579426_312647598_697285134_458913762);
         // Rules : HARD derived
         clue = 324'h000000600_000120370_100708049_000000000_000060010_030509000_000000508_007280000_400003060;
          // 23 clues
       end
      65 : begin
         soln_sig = signature(324'h572384619_341695278_698217543_735861492_926543781_814729365_483172956_267958134_159436827);
         // Rules : EASY derived
         clue = 324'h000000600_001095070_608007003_700000090_926040700_000020305_000000950_207000000_100400000;
          // 25 clues
       end
      66 : begin
         soln_sig = signature(324'h482519637_175463298_396872415_659237184_724185369_831694572_568741923_947326851_213958746);
         // Rules : HARD
         clue = 324'h000000600_100400098_090872005_059037004_000080000_001090570_000740003_000000000_200000046;
          // 26 clues
       end
      67 : begin
         soln_sig = signature(324'h351428697_497651382_862973154_734296518_685314729_129587436_213749865_946835271_578162943);
         // Rules : MEDIUM derived
         clue = 324'h000000607_000600080_000003150_700206000_600314020_109080000_003740005_040000070_008102000;
          // 27 clues
       end
      68 : begin
         soln_sig = signature(324'h723518649_549673128_186429375_694735812_851962437_237841956_378294561_912356784_465187293);
         // Rules : MEDIUM derived
         clue = 324'h000000609_040600020_080009005_000705800_001000000_230040000_000094000_002300700_000180003;
          // 23 clues
       end
      69 : begin
         soln_sig = signature(324'h791823645_862954137_543176928_659231874_437689512_128745369_276518493_315497286_984362751);
         // Rules : MEDIUM derived
         clue = 324'h000000645_800000130_500006000_000030070_000600000_020740309_006000090_005097080_004002050;
          // 25 clues
       end
      70 : begin
         soln_sig = signature(324'h251489736_438576921_679132584_124758369_396241857_587963412_965827143_742315698_813694275);
         // Rules : HARD derived
         clue = 324'h000000700_000506920_600032084_000700060_090041000_000000000_000000103_002305000_800090070;
          // 23 clues
       end
      71 : begin
         soln_sig = signature(324'h534169728_218437956_976582134_341856297_852974361_697213485_483621579_769345812_125798643);
         // Rules : HARD derived
         clue = 324'h000000700_200030050_076000000_301800000_050970360_600200080_080600079_000005000_100008003;
          // 25 clues
       end
      72 : begin
         soln_sig = signature(324'h549618732_628397154_137542896_491856273_276934581_385721649_713289465_962475318_854163927);
         // Rules : MEDIUM derived
         clue = 324'h000000700_600300004_130540000_490006003_000000080_300020600_000080060_002070000_804100020;
          // 24 clues
       end
      73 : begin
         soln_sig = signature(324'h473265819_596148327_128379456_715482693_862931574_934657182_687594231_249813765_351726948);
         // Rules : HARD derived
         clue = 324'h000000800_500040027_020379006_005002690_062901004_000007000_000094001_000000000_300000048;
          // 26 clues
       end
      74 : begin
         soln_sig = signature(324'h672159843_914238657_538764192_749826315_283517469_165943728_327691584_856472931_491385276);
         // Rules : HARD derived
         clue = 324'h000000803_010200000_500004100_000820000_083500069_160000020_007090080_050000001_400080070;
          // 25 clues
       end
      75 : begin
         soln_sig = signature(324'h976351824_124768953_583492671_857619432_632547198_491283765_369124587_218975346_745836219);
         // Rules : MEDIUM derived
         clue = 324'h000000804_000008050_000090670_800619030_602500000_400083000_009104007_010000040_005036000;
          // 27 clues
       end
      76 : begin
         soln_sig = signature(324'h296415837_817639452_435872196_981247563_562193784_743568921_679384215_358721649_124956378);
         // Rules : EASY derived
         clue = 324'h000000830_010000002_000800000_000240060_500090004_003000021_009380200_050020040_104900300;
          // 25 clues
       end
      77 : begin
         soln_sig = signature(324'h413287965_976451328_582936741_829765413_367149852_154823697_641372589_795618234_238594176);
         // Rules : MEDIUM derived
         clue = 324'h000000900_070450320_080000701_000000000_007009802_004020007_641370000_000008030_038500000;
          // 26 clues
       end
      78 : begin
         soln_sig = signature(324'h271346958_896175423_345298176_427931685_953862714_618754392_789623541_532419867_164587239);
         // Rules : MEDIUM derived
         clue = 324'h000000950_800100000_040200006_027030080_000060700_000004000_009620001_500409007_060580030;
          // 26 clues
       end
      79 : begin
         soln_sig = signature(324'h857341629_321569874_964287513_498652137_573918462_216734985_185423796_639175248_742896351);
         // Rules : EASY derived
         clue = 324'h000001000_020000004_000000510_008600007_500000402_000704900_080400700_600105040_702006050;
          // 25 clues
       end
      80 : begin
         soln_sig = signature(324'h592781634_183426759_764953821_621847395_479235186_358619247_815364972_247198563_936572418);
         // Rules : HARD derived
         clue = 324'h000001030_100420000_760000801_020000390_000005100_058600000_000004970_000000000_936000008;
          // 24 clues
       end
      81 : begin
         soln_sig = signature(324'h265371948_941285367_387964152_523819674_896547213_714632895_479128536_652793481_138456729);
         // Rules : MEDIUM derived
         clue = 324'h000001040_040085300_300904000_503800070_000007010_000600090_470020500_002003000_008400000;
          // 25 clues
       end
      82 : begin
         soln_sig = signature(324'h435681279_721549368_896723514_689215743_214376985_573498621_967134852_342857196_158962437);
         // Rules : HARD derived
         clue = 324'h000001200_000540360_890000000_080010043_004070005_070008600_000000050_040850000_100902000;
          // 25 clues
       end
      83 : begin
         soln_sig = signature(324'h254391867_963874521_817652934_592763148_431285679_786149352_648517293_375928416_129436785);
         // Rules : MEDIUM derived
         clue = 324'h000001800_900000000_017652000_000000040_031080600_000000052_600500090_000008010_009406700;
          // 24 clues
       end
      84 : begin
         soln_sig = signature(324'h498732516_536914287_217856493_761493852_924587361_853621974_649278135_175349628_382165749);
         // Rules : EASY derived
         clue = 324'h000002000_000904007_010800403_061000800_000000060_800020000_009070100_005300008_002060049;
          // 24 clues
       end
      85 : begin
         soln_sig = signature(324'h539672481_871459623_624381579_167245398_952738146_483196257_215967834_746823915_398514762);
         // Rules : MEDIUM derived
         clue = 324'h000002000_001400000_000301570_060005300_002000040_080090200_000060834_000800010_090004000;
          // 23 clues
       end
      86 : begin
         soln_sig = signature(324'h941672358_853419267_267385194_594827613_182536479_736194825_618953742_475268931_329741586);
         // Rules : MEDIUM derived
         clue = 324'h000002008_050410000_000000000_004000603_100500000_030090820_608003700_400260900_300000000;
          // 23 clues
       end
      87 : begin
         soln_sig = signature(324'h196352478_357846129_842917635_761284593_528139764_934765812_689573241_413628957_275491386);
         // Rules : EASY derived
         clue = 324'h000002008_050800100_040010000_001200590_008030060_000705002_680070040_400000907_005000006;
          // 26 clues
       end
      88 : begin
         soln_sig = signature(324'h513862479_872394165_496157283_365729814_124586397_987413652_231978546_748635921_659241738);
         // Rules : HARD derived
         clue = 324'h000002009_070090060_006050000_300000800_004500000_900013000_201008500_008000020_050040708;
          // 24 clues
       end
      89 : begin
         soln_sig = signature(324'h968142735_213587649_745369821_489253176_156478293_327691458_631924587_574836912_892715364);
         // Rules : MEDIUM
         clue = 324'h000002030_000500000_705060000_080000006_100070200_027000400_630900087_000000010_892000060;
          // 24 clues
       end
      90 : begin
         soln_sig = signature(324'h493672581_825931674_716845239_541289763_932716458_687453912_279168345_368594127_154327896);
         // Rules : MEDIUM derived
         clue = 324'h000002081_005000600_700040000_040089700_030010008_000400900_200000340_300590000_000007806;
          // 25 clues
       end
      91 : begin
         soln_sig = signature(324'h785942316_923716854_146583279_862391547_531674928_497258163_354169782_278435691_619827435);
         // Rules : HARD derived
         clue = 324'h000002310_900000000_006580009_802001500_500600900_400000000_050000780_078030000_000020030;
          // 24 clues
       end
      92 : begin
         soln_sig = signature(324'h149532687_275986314_836471259_963217845_487659123_521843796_754328961_392165478_618794532);
         // Rules : MEDIUM derived
         clue = 324'h000002600_075000000_036470050_903007040_007059023_000840000_700000000_090100408_000004002;
          // 27 clues
       end
      93 : begin
         soln_sig = signature(324'h863142957_592837416_714956238_279483561_436571829_185269374_651394782_928715643_347628195);
         // Rules : HARD derived
         clue = 324'h000002900_000800406_000950008_200400061_030070020_005209004_000000000_000010003_347008000;
          // 25 clues
       end
      94 : begin
         soln_sig = signature(324'h417562938_859173642_326894715_281349576_964758123_573621894_632987451_198435267_745216389);
         // Rules : HARD derived
         clue = 324'h000002900_800100600_020094005_081000000_900758000_000600004_600980001_000400060_740000000;
          // 25 clues
       end
      95 : begin
         soln_sig = signature(324'h498753126_532619487_617842395_865437219_721986534_943125768_284561973_376294851_159378642);
         // Rules : MEDIUM derived
         clue = 324'h000003000_002010087_610840090_860000200_000900000_040005000_200061000_070004000_009300000;
          // 23 clues
       end
      96 : begin
         soln_sig = signature(324'h491873265_386251974_527469831_978325146_234716598_615984723_869542317_742138659_153697482);
         // Rules : MEDIUM derived
         clue = 324'h000003005_000200070_000069800_008000106_000700000_000004003_000002000_700130609_150090080;
          // 23 clues
       end
      97 : begin
         soln_sig = signature(324'h745213968_612589473_398467512_259741836_436852791_187936254_571324689_864195327_923678145);
         // Rules : MEDIUM derived
         clue = 324'h000003060_000500070_008060502_200700830_400002000_100900000_500004000_000105300_003078005;
          // 25 clues
       end
      98 : begin
         soln_sig = signature(324'h827953614_451862739_936471258_674135982_518249376_392687145_145796823_263518497_789324561);
         // Rules : HARD derived
         clue = 324'h000003604_000002000_930000058_604000000_010000070_002080005_100706020_000000097_000304000;
          // 23 clues
       end
      99 : begin
         soln_sig = signature(324'h589463712_137259648_264178539_928731456_413596827_756842391_895614273_372985164_641327985);
         // Rules : HARD derived
         clue = 324'h000003700_100000040_060008500_008000400_003000827_056000390_090004200_000900060_000307000;
          // 24 clues
       end
      100 : begin
         soln_sig = signature(324'h826514397_971326584_435978261_793482615_514639728_682157439_148763952_359241876_267895143);
         // Rules : EASY derived
         clue = 324'h000004007_070326084_400900200_000000010_000009700_080057000_008703900_050000800_200090003;
          // 26 clues
       end
      101 : begin
         soln_sig = signature(324'h132694758_564872391_879135426_316489572_925713864_487256139_798361245_643528917_251947683);
         // Rules : EASY
         clue = 324'h000004008_560000301_800030020_310000500_000700064_087000000_000300000_000020917_200040000;
          // 24 clues
       end
      102 : begin
         soln_sig = signature(324'h359264871_428137695_176859324_697542138_584391267_213786549_941628753_832975416_765413982);
         // Rules : EASY derived
         clue = 324'h000004800_400100605_070859000_007002030_080000000_000000500_901600700_000070410_000010082;
          // 25 clues
       end
      103 : begin
         soln_sig = signature(324'h164935278_928471356_735682194_413856927_857219463_296743581_671524839_382197645_549368712);
         // Rules : HARD derived
         clue = 324'h000005000_000401050_000080090_003800900_850200400_296000001_600024800_002000000_000300710;
          // 25 clues
       end
      104 : begin
         soln_sig = signature(324'h293875641_456913872_178624593_349281756_562497318_817356924_925168437_784532169_631749285);
         // Rules : EASY derived
         clue = 324'h000005000_400910000_000600093_000201700_060090000_800000004_025060437_004030060_001000000;
          // 24 clues
       end
      105 : begin
         soln_sig = signature(324'h849765231_352981467_176234598_621853974_593147682_487629315_935418726_214376859_768592143);
         // Rules : MEDIUM derived
         clue = 324'h000005030_300080460_100004000_001003900_090100602_400000000_005000000_000076809_060090100;
          // 24 clues
       end
      106 : begin
         soln_sig = signature(324'h497285361_625137948_138964725_762813594_841596237_953742816_319678452_574321689_286459173);
         // Rules : HARD derived
         clue = 324'h000005360_600007908_108000000_000003500_840000030_900040000_000600002_000301080_006059000;
          // 24 clues
       end
      107 : begin
         soln_sig = signature(324'h178965423_453872916_926143875_839721654_261584397_547396281_794658132_382417569_615239748);
         // Rules : HARD derived
         clue = 324'h000005420_050800000_900040800_030701000_200000090_500306001_704000000_000007509_000209000;
          // 24 clues
       end
      108 : begin
         soln_sig = signature(324'h581376942_967428513_324195687_459817236_638542791_172963854_743259168_215684379_896731425);
         // Rules : MEDIUM derived
         clue = 324'h000006000_000020500_004005007_400800006_630002000_000900050_700000160_005084079_800700400;
          // 25 clues
       end
      109 : begin
         soln_sig = signature(324'h319846257_452719863_678325419_524971638_167483592_983652741_796234185_235168974_841597326);
         // Rules : EASY derived
         clue = 324'h000006007_052000003_600325400_000071600_000080000_003600701_090034000_000000004_801590000;
          // 26 clues
       end
      110 : begin
         soln_sig = signature(324'h846357219_512649378_739812564_465238197_928761435_173495682_257183946_394576821_681924753);
         // Rules : EASY derived
         clue = 324'h000007209_010000008_039010560_405008000_920000030_100000602_050000040_000006020_600900000;
          // 25 clues
       end
      111 : begin
         soln_sig = signature(324'h134257896_795468312_682391574_279835461_341976285_856142937_513629748_928714653_467583129);
         // Rules : EASY derived
         clue = 324'h000007806_005408000_000090000_070800000_001000005_000042030_500600700_920700653_400000000;
          // 24 clues
       end
      112 : begin
         soln_sig = signature(324'h231978546_794651328_865423719_916387254_547219863_382564197_629835471_158746932_473192685);
         // Rules : MEDIUM derived
         clue = 324'h000008000_700000000_060400019_000080054_000009063_002500000_600000000_108740000_003102005;
          // 23 clues
       end
      113 : begin
         soln_sig = signature(324'h576428913_143569872_892137645_761285439_459376281_328914756_917643528_285791364_634852197);
         // Rules : MEDIUM derived
         clue = 324'h000008013_040060000_002100000_760000009_400300280_000010000_910640008_000000304_600050000;
          // 24 clues
       end
      114 : begin
         soln_sig = signature(324'h954638172_716295348_832471659_167589423_295314786_348726591_421853967_689147235_573962814);
         // Rules : EASY derived
         clue = 324'h000008100_700200040_832400000_167009000_000300000_000720090_020800007_609040000_000000800;
          // 24 clues
       end
      115 : begin
         soln_sig = signature(324'h267539814_419876523_853412769_321957648_598264371_674381952_936125487_185743296_742698135);
         // Rules : MEDIUM derived
         clue = 324'h000009000_010000500_050402069_000900600_000000071_004380050_006100407_005000200_700098100;
          // 26 clues
       end
      116 : begin
         soln_sig = signature(324'h215469783_394178256_768352149_953724861_486531927_127986534_842617395_579843612_631295478);
         // Rules : MEDIUM derived
         clue = 324'h000009000_300070256_000350000_050004061_080000920_107006000_000010300_500000010_600005008;
          // 25 clues
       end
      117 : begin
         soln_sig = signature(324'h851649723_943287156_627351948_362794581_715862439_489513672_596428317_274136895_138975264);
         // Rules : HARD
         clue = 324'h000009000_900087150_600050000_360700000_005000409_009000002_000400300_004030005_100070060;
          // 24 clues
       end
      118 : begin
         soln_sig = signature(324'h537289641_684317259_912645738_891734562_463528197_275961384_749156823_358472916_126893475);
         // Rules : HARD derived
         clue = 324'h000009001_000010009_002000038_000000500_060008000_005900300_700006020_300402900_100000075;
          // 23 clues
       end
      119 : begin
         soln_sig = signature(324'h185469237_697532814_243178965_368245179_519387642_724916583_456721398_832694751_971853426);
         // Rules : EASY derived
         clue = 324'h000009230_007000000_040070005_300045000_000300642_000010000_006700000_000090751_900050400;
          // 24 clues
       end
      120 : begin
         soln_sig = signature(324'h823514796_476983512_951672843_619847325_742359168_385126479_298731654_567498231_134265987);
         // Rules : HARD derived
         clue = 324'h000010000_000083010_000600040_610007300_742000008_005006400_200730600_007000000_000005980;
          // 25 clues
       end
      121 : begin
         soln_sig = signature(324'h739516428_845723619_612849573_563978142_971462385_284135796_158394267_496257831_327681954);
         // Rules : HARD derived
         clue = 324'h000010020_045703000_600000000_003970002_000060005_000100090_008004000_490200800_007080054;
          // 25 clues
       end
      122 : begin
         soln_sig = signature(324'h273419568_649853721_158627349_716398254_482165937_935742816_324971685_867534192_591286473);
         // Rules : MEDIUM
         clue = 324'h000010060_000003020_008600309_700090000_400005000_900002810_300070000_000034100_001280003;
          // 25 clues
       end
      123 : begin
         soln_sig = signature(324'h462518793_185973246_973624158_538146972_794235861_216789534_621457389_347891625_859362417);
         // Rules : HARD derived
         clue = 324'h000010093_100070000_903000008_008006970_004200800_000000500_601007000_040890020_000000400;
          // 24 clues
       end
      124 : begin
         soln_sig = signature(324'h984712635_625843791_317695284_193526478_842179356_756438912_271384569_468957123_539261847);
         // Rules : MEDIUM derived
         clue = 324'h000010630_600003700_010000084_103500400_000079006_050000900_000304069_400000100_000200000;
          // 25 clues
       end
      125 : begin
         soln_sig = signature(324'h654812937_321947568_798365421_867531294_519624873_432798156_975483612_146279385_283156749);
         // Rules : HARD derived
         clue = 324'h000010930_300040508_708000000_860000090_500600000_000090100_000003002_000079080_003150000;
          // 24 clues
       end
      126 : begin
         soln_sig = signature(324'h562813947_814279536_397465218_243596871_159738624_678142359_435681792_981327465_726954183);
         // Rules : EASY derived
         clue = 324'h000013000_000009030_097000008_200000000_050730600_008100000_400000090_081027000_006050083;
          // 24 clues
       end
      127 : begin
         soln_sig = signature(324'h845913672_971462835_236785914_694278351_327159468_158634297_782391546_513846729_469527183);
         // Rules : MEDIUM derived
         clue = 324'h000013000_070460000_200700900_600208000_000000400_000030097_080001006_510000000_009500003;
          // 23 clues
       end
      128 : begin
         soln_sig = signature(324'h534218697_296473158_781965324_948627531_315894276_627351849_473182965_859736412_162549783);
         // Rules : HARD derived
         clue = 324'h000018090_296000008_001000304_900600530_000090070_020000000_003080000_000000412_000500000;
          // 23 clues
       end
      129 : begin
         soln_sig = signature(324'h542718693_719365824_638492715_457986132_981234567_263157489_396541278_175829346_824673951);
         // Rules : HARD derived
         clue = 324'h000018093_000060000_030000010_050006000_980200507_203000000_000500208_100020300_004000001;
          // 24 clues
       end
      130 : begin
         soln_sig = signature(324'h413725986_982164753_765938124_598647312_234891567_671352498_857213649_126479835_349586271);
         // Rules : HARD derived
         clue = 324'h000020000_002104700_060000100_008640002_030001060_071000008_800200009_000009035_000580000;
          // 25 clues
       end
      131 : begin
         soln_sig = signature(324'h485927163_327168459_196543872_769385241_841692537_253471698_674819325_512736984_938254716);
         // Rules : MEDIUM derived
         clue = 324'h000020000_300100459_000503000_060000240_801090000_050070098_000800300_500000080_900050006;
          // 25 clues
       end
      132 : begin
         soln_sig = signature(324'h146728359_785391624_923546718_294853167_678219543_531467982_862975431_359184276_417632895);
         // Rules : MEDIUM derived
         clue = 324'h000020350_705000024_900006000_000800107_600009000_000000980_002900400_050000070_400600800;
          // 24 clues
       end
      133 : begin
         soln_sig = signature(324'h846123795_253976184_917584236_495367821_328419567_671852943_534291678_162738459_789645312);
         // Rules : MEDIUM derived
         clue = 324'h000020700_053000000_017504030_005360021_000409000_601050040_500000000_060008409_000040002;
          // 27 clues
       end
      134 : begin
         soln_sig = signature(324'h695721843_743856291_128493576_812369754_376548912_459172638_281935467_534687129_967214385);
         // Rules : MEDIUM derived
         clue = 324'h000021040_000006200_008000500_010060000_070500000_009000008_000905460_034000009_900210085;
          // 25 clues
       end
      135 : begin
         soln_sig = signature(324'h491623785_752481369_386579412_168954237_235716948_947832651_513247896_674198523_829365174);
         // Rules : MEDIUM derived
         clue = 324'h000023000_002001369_000500000_108900000_030700908_040000650_003000800_000008020_009300004;
          // 25 clues
       end
      136 : begin
         soln_sig = signature(324'h567923481_819647352_243185976_724319568_136258794_958764123_391872645_472536819_685491237);
         // Rules : MEDIUM derived
         clue = 324'h000023480_010640050_000000900_000010060_130008000_950700000_000800000_470030009_000000200;
          // 23 clues
       end
      137 : begin
         soln_sig = signature(324'h973528614_681479532_425163789_892315467_734692851_516847293_359284176_268731945_147956328);
         // Rules : HARD derived
         clue = 324'h000028014_000000032_005100000_090000007_004600850_510000000_300000006_200030940_107006020;
          // 26 clues
       end
      138 : begin
         soln_sig = signature(324'h573429816_461875329_298361475_917543268_382617954_645298731_736954182_854132697_129786543);
         // Rules : HARD derived
         clue = 324'h000029800_000800000_000301070_000040260_300600900_040000030_736004000_000000090_120000503;
          // 24 clues
       end
      139 : begin
         soln_sig = signature(324'h491736258_578412639_632589471_143957826_259168347_867243915_384671592_726395184_915824763);
         // Rules : MEDIUM derived
         clue = 324'h000030000_008002000_000089470_003000020_050100300_060040900_000600592_000005080_010020000;
          // 23 clues
       end
      140 : begin
         soln_sig = signature(324'h842635917_916742835_357891426_569173284_183426759_274589361_735918642_421367598_698254173);
         // Rules : HARD derived
         clue = 324'h000030007_900040000_050800000_500070004_080006009_204000000_030008600_001067008_000000103;
          // 23 clues
       end
      141 : begin
         soln_sig = signature(324'h125837469_374956128_986421573_269318745_513764892_847592316_732645981_658179234_491283657);
         // Rules : HARD derived
         clue = 324'h000030400_000906100_000001000_200300040_013700090_847000006_700000000_008079030_000200650;
          // 25 clues
       end
      142 : begin
         soln_sig = signature(324'h485231679_629748531_173956428_758394162_962175843_314862795_247583916_591627384_836419257);
         // Rules : HARD derived
         clue = 324'h000031009_000740500_100000000_008300002_960005003_010002090_007500000_000000304_806019000;
          // 25 clues
       end
      143 : begin
         soln_sig = signature(324'h126438597_743592861_589167432_271856943_495713286_638924715_852641379_314279658_967385124);
         // Rules : EASY derived
         clue = 324'h000038500_000092001_500100430_200800003_405700006_030004000_002000009_010079000_007000100;
          // 26 clues
       end
      144 : begin
         soln_sig = signature(324'h581642397_724359681_369781452_492867513_653914278_817235964_148526739_276193845_935478126);
         // Rules : MEDIUM derived
         clue = 324'h000040000_000309000_069080002_090067010_000000200_800000904_008506009_200100005_030008006;
          // 25 clues
       end
      145 : begin
         soln_sig = signature(324'h329647185_648125397_517389426_781952643_234861759_956473812_893516274_475238961_162794538);
         // Rules : MEDIUM
         clue = 324'h000040000_008100097_510309020_000002000_030060000_950000800_800510000_070030000_002004000;
          // 23 clues
       end
      146 : begin
         soln_sig = signature(324'h851746239_634921578_297835461_542678193_963512784_178493652_415369827_326187945_789254316);
         // Rules : HARD
         clue = 324'h000040009_030900070_007800000_002008000_900510000_100000600_405060800_006000040_080200306;
          // 24 clues
       end
      147 : begin
         soln_sig = signature(324'h795248613_281563794_634791528_857612439_413985267_926374851_369827145_172459386_548136972);
         // Rules : HARD derived
         clue = 324'h000040010_280500700_630090028_800000030_400000007_006070000_009020005_000009386_000106000;
          // 26 clues
       end
      148 : begin
         soln_sig = signature(324'h217943568_345682179_698157423_756298341_932714685_184365792_579836214_421579836_863421957);
         // Rules : HARD derived
         clue = 324'h000040560_300000000_008107003_700008300_900000000_104060700_070000210_021500000_000400050;
          // 24 clues
       end
      149 : begin
         soln_sig = signature(324'h857341962_942567183_163928754_638794215_495132678_721685349_519473826_276859431_384216597);
         // Rules : HARD derived
         clue = 324'h000040960_040007000_100900700_600000010_400032008_020085000_509000000_000050401_000016000;
          // 24 clues
       end
      150 : begin
         soln_sig = signature(324'h617243589_325918746_984675123_532186974_876459312_149327865_451832697_263791458_798564231);
         // Rules : HARD
         clue = 324'h000043000_000900700_900005100_530000074_870000000_000020000_401800600_000000050_008060230;
          // 23 clues
       end
      151 : begin
         soln_sig = signature(324'h821645379_473219856_956783421_785321694_632894517_194576283_268937145_547162938_319458762);
         // Rules : MEDIUM derived
         clue = 324'h000045070_000200800_000003001_700000094_000800000_000006003_008930045_000002000_019050700;
          // 23 clues
       end
      152 : begin
         soln_sig = signature(324'h216354978_834791625_579826341_387219456_421567893_695438217_753642189_148973562_962185734);
         // Rules : MEDIUM derived
         clue = 324'h000050000_030000000_079000000_007009006_021000800_600400210_050000009_008070500_002180030;
          // 23 clues
       end
      153 : begin
         soln_sig = signature(324'h492658713_368712945_517394628_751423869_649871532_283965174_134587296_826139457_975246381);
         // Rules : EASY derived
         clue = 324'h000050003_060012000_507000600_050400060_000000002_283005070_000000000_826100000_000040001;
          // 23 clues
       end
      154 : begin
         soln_sig = signature(324'h162459783_785321964_934687521_376842159_458916372_219573648_847135296_621794835_593268417);
         // Rules : MEDIUM derived
         clue = 324'h000050080_080320900_900087000_000040050_000006070_209003040_840100200_001090000_003008000;
          // 25 clues
       end
      155 : begin
         soln_sig = signature(324'h426859713_759136842_813247569_265481397_187963254_934572186_592714638_371698425_648325971);
         // Rules : EASY derived
         clue = 324'h000050713_050006000_000000000_200400397_100060004_030000000_090004000_001000420_000305001;
          // 23 clues
       end
      156 : begin
         soln_sig = signature(324'h913752468_652384197_478619253_281567349_536498721_749123685_865231974_127945836_394876512);
         // Rules : HARD derived
         clue = 324'h000052008_000080097_000600050_200560009_006090701_040003600_000001004_000000000_394800000;
          // 25 clues
       end
      157 : begin
         soln_sig = signature(324'h978653214_342791685_651284973_527368491_819542367_436179852_795436128_183927546_264815739);
         // Rules : HARD derived
         clue = 324'h000053014_002090600_601000000_000300091_800000000_030170000_700006008_000020040_060015700;
          // 25 clues
       end
      158 : begin
         soln_sig = signature(324'h416357928_253918476_798462531_821796345_649523187_537841692_362179854_974685213_185234769);
         // Rules : HARD derived
         clue = 324'h000057000_250910400_098000000_820790000_600003100_007800002_000070004_000600003_000004009;
          // 25 clues
       end
      159 : begin
         soln_sig = signature(324'h638457912_794132865_152869734_379516248_826394157_541278396_213745689_467983521_985621473);
         // Rules : MEDIUM derived
         clue = 324'h000057910_000030000_002800004_309000208_800000057_500200000_010000080_400900001_900600000;
          // 24 clues
       end
      160 : begin
         soln_sig = signature(324'h149765283_687329415_325814769_491638527_273951846_568472931_714583692_852196374_936247158);
         // Rules : EASY
         clue = 324'h000060203_007029000_000800000_001000007_000950040_060002000_700003600_850006374_900000000;
          // 24 clues
       end
      161 : begin
         soln_sig = signature(324'h842167395_937845126_615932748_584321967_126579483_379684251_253416879_768293514_491758632);
         // Rules : EASY derived
         clue = 324'h000060300_900005020_615002000_000001000_000509080_379080000_050006009_708200000_000000600;
          // 24 clues
       end
      162 : begin
         soln_sig = signature(324'h279865413_135427689_468391527_782534196_613978254_954216738_527683941_341759862_896142375);
         // Rules : EASY derived
         clue = 324'h000060400_005400600_008000520_082030000_010008250_900010000_000000941_040700000_000002300;
          // 24 clues
       end
      163 : begin
         soln_sig = signature(324'h453768912_726391845_918254637_867419523_142835796_539627184_671942358_394586271_285173469);
         // Rules : HARD derived
         clue = 324'h000060912_720000045_008000000_800009020_002000006_509600000_001042000_300580000_000003000;
          // 24 clues
       end
      164 : begin
         soln_sig = signature(324'h835762491_461389572_279145638_618537249_794218356_523496187_187654923_352971864_946823715);
         // Rules : EASY derived
         clue = 324'h000062090_001300502_070040600_010530000_700008050_003400000_000000920_000071004_940000010;
          // 26 clues
       end
      165 : begin
         soln_sig = signature(324'h387564129_915382647_426179835_839715264_564928713_271643598_158436972_693257481_742891356);
         // Rules : EASY derived
         clue = 324'h000064000_005300007_400000000_030010000_000008700_071000008_100030900_600050400_040091300;
          // 23 clues
       end
      166 : begin
         soln_sig = signature(324'h294675831_876132495_351849276_187253649_529764183_643981752_438526917_965417328_712398564);
         // Rules : EASY derived
         clue = 324'h000070000_006000005_050000206_100050049_520000080_000081000_008006017_000400300_002090060;
          // 24 clues
       end
      167 : begin
         soln_sig = signature(324'h512876439_869324571_437159862_956483217_278561943_341792658_124935786_685217394_793648125);
         // Rules : HARD derived
         clue = 324'h000070000_060020500_430009002_906403007_200001900_000002650_004000000_000000094_700600100;
          // 25 clues
       end
      168 : begin
         soln_sig = signature(324'h318675942_964281537_725439816_491563278_583927164_672148395_847392651_136854729_259716483);
         // Rules : HARD derived
         clue = 324'h000070002_000200007_005000016_090060000_003007100_000000300_800090050_100054700_200000083;
          // 23 clues
       end
      169 : begin
         soln_sig = signature(324'h984371256_627859134_513624978_832416795_146795823_795283641_251948367_469137582_378562419);
         // Rules : HARD derived
         clue = 324'h000070200_000800000_513000000_802400090_006090000_000000001_250000300_009037000_070000419;
          // 23 clues
       end
      170 : begin
         soln_sig = signature(324'h634879521_259461837_187532649_793615284_825347196_461928753_948156372_576293418_312784965);
         // Rules : HARD derived
         clue = 324'h000070501_200000007_080000040_000005000_025300006_400900700_008006370_000290400_010000005;
          // 24 clues
       end
      171 : begin
         soln_sig = signature(324'h635279841_478651293_129834675_947526318_862913754_513748962_356492187_781365429_294187536);
         // Rules : HARD derived
         clue = 324'h000070800_400000090_020030600_007000318_062000750_003000900_050090100_000005020_000087000;
          // 24 clues
       end
      172 : begin
         soln_sig = signature(324'h598473162_146529783_327816495_754982316_283761549_961345827_415297638_672138954_839654271);
         // Rules : EASY derived
         clue = 324'h000073060_100500000_027006000_000082010_200000509_900300807_010000630_000000050_009054001;
          // 26 clues
       end
      173 : begin
         soln_sig = signature(324'h528479361_916235847_473681592_859347126_132956784_764128953_687512439_395764218_241893675);
         // Rules : MEDIUM derived
         clue = 324'h000079300_016200000_403000500_009040000_002906004_060008003_680500000_000004200_001000070;
          // 25 clues
       end
      174 : begin
         soln_sig = signature(324'h732185649_586492173_941637852_198573426_374926581_625841397_257318964_463259718_819764235);
         // Rules : EASY derived
         clue = 324'h000080000_000002070_941007000_000000406_300000081_025040000_007008060_060200000_810000035;
          // 24 clues
       end
      175 : begin
         soln_sig = signature(324'h592784316_143625879_867139245_439816752_218573694_675492183_386957421_754261938_921348567);
         // Rules : MEDIUM derived
         clue = 324'h000080000_000020079_800100000_009006050_210003004_075090000_300007400_000000008_020000560;
          // 23 clues
       end
      176 : begin
         soln_sig = signature(324'h513784269_287916534_496253817_841695723_379842156_652371948_764529381_935168472_128437695);
         // Rules : MEDIUM derived
         clue = 324'h000080000_000900500_006050007_840090000_000002050_600001008_700000380_005160072_100007600;
          // 25 clues
       end
      177 : begin
         soln_sig = signature(324'h327689154_965174382_418352796_684923571_291765438_573418629_742596813_139847265_856231947);
         // Rules : EASY derived
         clue = 324'h000080004_060004300_010300000_004900070_000065008_003008620_740500010_100000205_006000007;
          // 26 clues
       end
      178 : begin
         soln_sig = signature(324'h916482537_385976142_724315869_863127495_192564378_457839621_638791254_571243986_249658713);
         // Rules : MEDIUM derived
         clue = 324'h000080030_300900140_700010000_060007405_100000000_007030600_008000000_000240906_040600700;
          // 24 clues
       end
      179 : begin
         soln_sig = signature(324'h421783569_867915234_359264781_216458397_798326145_543197628_932541876_675839412_184672953);
         // Rules : MEDIUM derived
         clue = 324'h000080069_007905000_350000700_006400007_000320005_540000020_030001006_600000012_004000000;
          // 25 clues
       end
      180 : begin
         soln_sig = signature(324'h391487265_485261973_267593184_752138649_914756832_638924751_579842316_823615497_146379528);
         // Rules : HARD derived
         clue = 324'h000080200_085200900_200003084_050100000_004006000_030904700_000000010_003600000_000079508;
          // 25 clues
       end
      181 : begin
         soln_sig = signature(324'h419785362_256931487_387264591_921456738_538179624_764823915_195348276_673512849_842697153);
         // Rules : MEDIUM derived
         clue = 324'h000080300_050930080_080000000_020450000_000009004_700000910_100008270_003000800_000697000;
          // 24 clues
       end
      182 : begin
         soln_sig = signature(324'h241583769_678192534_935647812_514936287_326478195_897215643_463751928_782369451_159824376);
         // Rules : HARD
         clue = 324'h000080700_000002504_000607002_010900080_006078005_800005043_000000000_000300001_159020000;
          // 25 clues
       end
      183 : begin
         soln_sig = signature(324'h159682347_764359218_382174956_247531869_891267435_536498172_923746581_478915623_615823794);
         // Rules : EASY derived
         clue = 324'h000082047_760050010_300000900_000000800_001260005_000400070_000046000_070000023_600003000;
          // 24 clues
       end
      184 : begin
         soln_sig = signature(324'h392185647_861974325_754362918_628743591_917528436_435691872_573819264_149256783_286437159);
         // Rules : EASY derived
         clue = 324'h000085007_000970320_050000000_600043000_000020000_430600800_500819060_040006000_080000109;
          // 26 clues
       end
      185 : begin
         soln_sig = signature(324'h241786935_983251467_567394281_894573612_735162894_126849753_619425378_458637129_372918546);
         // Rules : HARD derived
         clue = 324'h000086030_900200400_067000000_000570002_000000000_100009000_009000000_450630100_302018000;
          // 23 clues
       end
      186 : begin
         soln_sig = signature(324'h361587924_845239167_279416583_658973412_937124856_412658379_523791648_786345291_194862735);
         // Rules : HARD derived
         clue = 324'h000087020_000230100_000000000_050900000_037104806_002000009_523090608_000000000_004000035;
          // 25 clues
       end
      187 : begin
         soln_sig = signature(324'h352691487_189475326_746328591_521937648_894162735_673584912_935816274_417259863_268743159);
         // Rules : EASY derived
         clue = 324'h000090000_080000006_000000590_500000608_000062700_003004002_030006200_400059060_208040050;
          // 25 clues
       end
      188 : begin
         soln_sig = signature(324'h538296174_961374852_472158693_189537246_257461938_643829517_714685329_396712485_825943761);
         // Rules : EASY derived
         clue = 324'h000090004_001300000_472000000_000007200_000001038_603800007_004005000_306000080_005040060;
          // 24 clues
       end
      189 : begin
         soln_sig = signature(324'h568497321_293816745_417532986_689174532_724385619_351269478_946721853_872653194_135948267);
         // Rules : MEDIUM derived
         clue = 324'h000090021_003000700_400500000_080100002_000005600_050260400_900000850_800603000_000040207;
          // 25 clues
       end
      190 : begin
         soln_sig = signature(324'h478192635_913865247_265437189_527348916_341976852_689521374_194653728_852719463_736284591);
         // Rules : HARD
         clue = 324'h000090030_900805000_260000109_000040900_041006000_080000370_000050720_000000000_736000001;
          // 24 clues
       end
      191 : begin
         soln_sig = signature(324'h162598347_587346291_439127865_326479158_814253976_795861432_678932514_941785623_253614789);
         // Rules : MEDIUM derived
         clue = 324'h000090340_000006200_000000065_006479100_804200000_005061000_070000500_900705003_200014000;
          // 27 clues
       end
      192 : begin
         soln_sig = signature(324'h548791362_792638451_316245978_859426713_231579846_674183529_187352694_463917285_925864137);
         // Rules : EASY derived
         clue = 324'h000090360_002000000_010200008_000006713_000500000_600180000_007002000_000900285_900800100;
          // 24 clues
       end
      193 : begin
         soln_sig = signature(324'h584129763_367584129_129673458_972845316_658931247_431267895_243756981_896312574_715498632);
         // Rules : MEDIUM derived
         clue = 324'h000100003_060084000_000000000_070005310_008000207_400060000_203700900_800012500_700000000;
          // 23 clues
       end
      194 : begin
         soln_sig = signature(324'h253168749_847395612_196427853_362714985_478539126_519286437_931872564_724651398_685943271);
         // Rules : EASY derived
         clue = 324'h000100009_047000002_100427800_002010905_000509100_000006000_030802000_000000008_605043000;
          // 26 clues
       end
      195 : begin
         soln_sig = signature(324'h327185649_658942137_941673285_894231756_536798412_712456398_489367521_173529864_265814973);
         // Rules : HARD derived
         clue = 324'h000105000_000900100_040000005_800231700_000700400_700000308_080007001_000009060_260800903;
          // 26 clues
       end
      196 : begin
         soln_sig = signature(324'h532176948_874293156_961458237_397642581_148539672_625817493_219784365_486325719_753961824);
         // Rules : EASY derived
         clue = 324'h000106048_870003050_900000200_000040080_000000600_005017003_000704000_080000019_700900000;
          // 24 clues
       end
      197 : begin
         soln_sig = signature(324'h342156798_597428631_816397452_758643129_921875346_463219587_284561973_139784265_675932814);
         // Rules : HARD derived
         clue = 324'h000106090_597000001_006000402_050000000_900070340_000009080_004001000_000000265_000030000;
          // 23 clues
       end
      198 : begin
         soln_sig = signature(324'h358129746_761845239_429367185_283691574_547283961_916754823_135478692_892536417_674912358);
         // Rules : EASY derived
         clue = 324'h000129000_000005000_420300100_280000504_507000060_010000020_130000000_000530407_604000008;
          // 26 clues
       end
      199 : begin
         soln_sig = signature(324'h697145328_582963714_143827596_731298465_856431972_429576183_978654231_365712849_214389657);
         // Rules : HARD derived
         clue = 324'h000140300_000003000_000027090_700008400_050000070_000500180_978050000_000000040_210000607;
          // 24 clues
       end
      200 : begin
         soln_sig = signature(324'h273156894_619483257_584729316_128564739_746931528_395872641_952617483_861345972_437298165);
         // Rules : EASY derived
         clue = 324'h000150000_000080050_084000006_020504700_006001000_300000000_900000080_061340000_007200065;
          // 24 clues
       end
      201 : begin
         soln_sig = signature(324'h592164378_478253196_613987245_845732961_729416583_361598427_136829754_287345619_954671832);
         // Rules : MEDIUM derived
         clue = 324'h000160070_000050100_003000200_040002000_009000003_060500000_000029750_087000009_900601032;
          // 25 clues
       end
      202 : begin
         soln_sig = signature(324'h259184673_381967542_476235198_718596324_643721985_592843761_927358416_834619257_165472839);
         // Rules : MEDIUM derived
         clue = 324'h000184000_300000000_076200000_018096004_003701000_090043060_000000410_800009057_005000800;
          // 27 clues
       end
      203 : begin
         soln_sig = signature(324'h876192543_549873621_231456897_315948762_628537914_497621358_953714286_784269135_162385479);
         // Rules : MEDIUM derived
         clue = 324'h000190543_000800601_001006000_000000000_620007900_090020300_950000006_700000000_102380009;
          // 26 clues
       end
      204 : begin
         soln_sig = signature(324'h416239758_537648291_289715634_652974813_894163527_371582946_728491365_943856172_165327489);
         // Rules : MEDIUM derived
         clue = 324'h000200000_000600091_200005000_650070003_094100000_001080040_700090300_000000002_060000480;
          // 23 clues
       end
      205 : begin
         soln_sig = signature(324'h783254961_924671385_651389724_578432196_436918257_192567438_369745812_845123679_217896543);
         // Rules : EASY derived
         clue = 324'h000200000_004000005_050000704_570000090_000910000_100500038_009040012_000003600_007800040;
          // 24 clues
       end
      206 : begin
         soln_sig = signature(324'h513278694_874369521_692541873_328715469_961432758_457896312_136954287_785123946_249687135);
         // Rules : HARD derived
         clue = 324'h000200000_070300500_690040003_300010400_000030750_407096002_006000000_000000046_200007100;
          // 25 clues
       end
      207 : begin
         soln_sig = signature(324'h713264895_928315647_546987213_654832179_391576428_287491356_172658934_469723581_835149762);
         // Rules : EASY derived
         clue = 324'h000200000_900015000_000080013_600000009_000570400_080001000_072008934_009003080_005000000;
          // 24 clues
       end
      208 : begin
         soln_sig = signature(324'h564289173_281473569_397651482_452718936_918364257_673592814_826147395_749835621_135926748);
         // Rules : HARD derived
         clue = 324'h000200100_000073500_000050000_052008030_918000007_600002010_800000000_009830020_000006740;
          // 25 clues
       end
      209 : begin
         soln_sig = signature(324'h789231456_136584927_542967381_375149268_621873549_498625713_863492175_257316894_914758632);
         // Rules : MEDIUM derived
         clue = 324'h000200450_000080900_000000081_305009000_001870000_008625700_060000100_200016004_900750000;
          // 27 clues
       end
      210 : begin
         soln_sig = signature(324'h197236854_834759612_526148397_973612548_648597123_215384769_362975481_789461235_451823976);
         // Rules : MEDIUM derived
         clue = 324'h000200850_800050600_020000097_000610008_040000100_205004700_000075081_700000200_000003000;
          // 25 clues
       end
      211 : begin
         soln_sig = signature(324'h653281947_942537186_781496523_836154279_124679835_579328614_298745361_317962458_465813792);
         // Rules : HARD derived
         clue = 324'h000201907_000030000_081000003_830000200_020609005_009000600_000045060_000960400_000810000;
          // 25 clues
       end
      212 : begin
         soln_sig = signature(324'h871265493_469783512_235914678_794826135_586371249_312459867_648537921_953142786_127698354);
         // Rules : EASY derived
         clue = 324'h000205090_400080000_035900000_700020105_000301040_300000807_040000920_000000080_007608004;
          // 26 clues
       end
      213 : begin
         soln_sig = signature(324'h869245137_172398456_435167892_247951683_681423579_953786241_794812365_518639724_326574918);
         // Rules : MEDIUM derived
         clue = 324'h000240000_002090456_000007000_040001603_080000570_903006000_004000300_000030020_006004008;
          // 25 clues
       end
      214 : begin
         soln_sig = signature(324'h793261548_546938217_281745693_379856124_658412739_124397865_915684372_832179456_467523981);
         // Rules : HARD derived
         clue = 324'h000261008_506000000_200700090_370000020_000400700_000090060_005680300_032000400_000000080;
          // 24 clues
       end
      215 : begin
         soln_sig = signature(324'h945273186_816549327_237816594_452781639_169435278_378692415_623958741_584127963_791364852);
         // Rules : HARD derived
         clue = 324'h000273000_800009300_000000004_000000000_160000270_078000000_003058001_500127960_000060000;
          // 24 clues
       end
      216 : begin
         soln_sig = signature(324'h375291864_896734152_421856793_754328916_168479235_932615487_513942678_289567341_647183529);
         // Rules : HARD derived
         clue = 324'h000290064_000000052_001006000_004008910_160000000_030000007_500000008_200500340_607080020;
          // 26 clues
       end
      217 : begin
         soln_sig = signature(324'h126394758_853276914_794185623_268547391_415639287_937812465_342951876_579468132_681723549);
         // Rules : MEDIUM derived
         clue = 324'h000300000_050000900_090180023_008047090_000030200_000000065_002050806_009000100_600703500;
          // 26 clues
       end
      218 : begin
         soln_sig = signature(324'h497318256_312564879_658729413_164852937_875193642_923647185_736281594_241975368_589436721);
         // Rules : EASY derived
         clue = 324'h000300200_300060809_050729000_000000900_005100040_020000000_706080500_000005360_000006021;
          // 25 clues
       end
      219 : begin
         soln_sig = signature(324'h486391572_217845639_935726814_398654721_562173948_174982365_721569483_853417296_649238157);
         // Rules : HARD derived
         clue = 324'h000300502_000800000_930000014_008004001_502000000_070000060_700560080_000000096_000230000;
          // 23 clues
       end
      220 : begin
         soln_sig = signature(324'h451387629_697251348_238964715_526143897_879526134_314879562_745612983_183495276_962738451);
         // Rules : EASY
         clue = 324'h000387000_000050000_230004700_506000090_070000030_310000502_740000000_000405206_902000001;
          // 26 clues
       end
      221 : begin
         soln_sig = signature(324'h581392476_276854931_394761825_812643759_653279184_749518263_935487612_427136598_168925347);
         // Rules : EASY derived
         clue = 324'h000390006_006000030_090000020_010003750_000070004_040008200_005480000_407006500_060920000;
          // 26 clues
       end
      222 : begin
         soln_sig = signature(324'h597412638_428635791_136789425_254897163_813264957_679351284_941523876_362178549_785946312);
         // Rules : HARD derived
         clue = 324'h000400000_400605790_100009000_004000003_810060000_009000204_000020800_002008009_700006010;
          // 24 clues
       end
      223 : begin
         soln_sig = signature(324'h512479836_938621745_476853921_347916258_129587364_685342179_894735612_761294583_253168497);
         // Rules : EASY derived
         clue = 324'h000400806_030000005_076003920_300000208_109500000_680000070_090000010_000200080_200060000;
          // 25 clues
       end
      224 : begin
         soln_sig = signature(324'h592431768_183765294_647982315_826193547_931574826_754826139_365247981_419358672_278619453);
         // Rules : HARD derived
         clue = 324'h000401060_000065200_000000000_006000007_030070000_054820109_365007901_000000000_008000053;
          // 25 clues
       end
      225 : begin
         soln_sig = signature(324'h765483921_489216537_123975684_631548279_948762153_257139468_396824715_874651392_512397846);
         // Rules : HARD derived
         clue = 324'h000403000_000010500_100900600_000008000_940000053_250000000_306020700_000000090_002007840;
          // 23 clues
       end
      226 : begin
         soln_sig = signature(324'h925463718_861257394_473981265_298134657_346725981_517896432_734519826_189642573_652378149);
         // Rules : MEDIUM derived
         clue = 324'h000403708_001000304_400001000_090104050_006020900_000890400_000509800_009000070_052300000;
          // 27 clues
       end
      227 : begin
         soln_sig = signature(324'h879465231_563821947_421397586_257134698_984652173_136978425_318549762_642713859_795286314);
         // Rules : HARD
         clue = 324'h000405200_000800000_000097080_000030690_004600070_030000400_000000700_642003000_095000014;
          // 24 clues
       end
      228 : begin
         soln_sig = signature(324'h625419873_713586249_894273165_186937452_259641738_347825916_432158697_978364521_561792384);
         // Rules : HARD derived
         clue = 324'h000410000_003080049_090073100_006930000_050000708_000005900_032108600_070000020_000000080;
          // 26 clues
       end
      229 : begin
         soln_sig = signature(324'h378462591_419875362_256319487_941623758_762584913_835197624_627948135_183756249_594231876);
         // Rules : HARD derived
         clue = 324'h000460001_009005060_200300000_000000050_700080903_805007000_027000000_000000000_590031800;
          // 23 clues
       end
      230 : begin
         soln_sig = signature(324'h261489753_479356218_385712694_693148527_528697431_714523869_832964175_956871342_147235986);
         // Rules : EASY derived
         clue = 324'h000480003_000306210_080000000_000100000_520007400_700520000_800964070_050070000_040000906;
          // 26 clues
       end
      231 : begin
         soln_sig = signature(324'h632549178_451827963_879361542_367218459_124795386_985634721_246953817_713482695_598176234);
         // Rules : EASY derived
         clue = 324'h000500000_000020060_879060000_300000059_024700000_000000701_006050010_010002000_590000034;
          // 24 clues
       end
      232 : begin
         soln_sig = signature(324'h213564879_849217536_576938214_384795162_697421385_152683497_921356748_768142953_435879621);
         // Rules : EASY derived
         clue = 324'h000500000_000210006_070030204_300005000_097000300_000000090_001006700_008040003_005009021;
          // 24 clues
       end
      233 : begin
         soln_sig = signature(324'h973561284_168342795_542789136_759824361_634175928_281693547_496257813_325418679_817936452);
         // Rules : MEDIUM derived
         clue = 324'h000500000_100000000_040080036_009020000_000005028_000600047_400000000_305018000_007930002;
          // 23 clues
       end
      234 : begin
         soln_sig = signature(324'h281576934_375149862_496328517_549713286_827654391_613892475_964287153_758431629_132965748);
         // Rules : EASY derived
         clue = 324'h000500004_370000802_400008010_049000000_820000300_000090075_000080000_000001629_100005000;
          // 24 clues
       end
      235 : begin
         soln_sig = signature(324'h216593874_785462193_349178652_671324985_934685721_852917436_497251368_128736549_563849217);
         // Rules : HARD derived
         clue = 324'h000500800_000062190_340000000_070300900_030005021_002007006_000000060_020036000_500840000;
          // 25 clues
       end
      236 : begin
         soln_sig = signature(324'h378591642_241786953_659324817_736915284_185243796_924867135_897452361_463179528_512638479);
         // Rules : EASY derived
         clue = 324'h000501000_000080903_600020800_706000200_005000700_024000000_800052061_000009008_500630070;
          // 26 clues
       end
      237 : begin
         soln_sig = signature(324'h793512648_421869753_568473219_215987364_849356172_376124985_134695827_657238491_982741536);
         // Rules : HARD derived
         clue = 324'h000502000_420069700_068000000_005080004_840056000_300100900_000005007_000030001_000700006;
          // 25 clues
       end
      238 : begin
         soln_sig = signature(324'h193542687_647981325_582673149_251496873_839127564_764358912_418239756_375864291_926715438);
         // Rules : HARD derived
         clue = 324'h000502007_000081300_500000000_050400070_009020004_760300002_008030000_000000201_906705000;
          // 25 clues
       end
      239 : begin
         soln_sig = signature(324'h947538216_185276493_236914587_329745168_564381729_871629354_618457932_453892671_792163845);
         // Rules : HARD derived
         clue = 324'h000508006_000006093_000010080_020700100_500081009_001009304_000400002_000000000_792060000;
          // 25 clues
       end
      240 : begin
         soln_sig = signature(324'h387514962_952368741_146972583_469231875_718659234_523847196_234795618_871426359_695183427);
         // Rules : EASY
         clue = 324'h000510060_002008701_040900500_400030070_008009000_020807000_000000610_000420009_690000020;
          // 26 clues
       end
      241 : begin
         soln_sig = signature(324'h379528614_516947328_428361579_867453291_945182736_132796845_783614952_251879463_694235187);
         // Rules : MEDIUM derived
         clue = 324'h000520010_000007300_000060009_000003000_000080006_100000045_003604052_000070000_094200100;
          // 23 clues
       end
      242 : begin
         soln_sig = signature(324'h796528431_158436927_234197865_421783659_967215348_385649172_673951284_512864793_849372516);
         // Rules : MEDIUM derived
         clue = 324'h000528000_100000000_034007000_001083000_060210040_085640002_000000280_500060093_009000500;
          // 27 clues
       end
      243 : begin
         soln_sig = signature(324'h372586941_956714832_148392765_287945316_614873259_539621487_461239578_823157694_795468123);
         // Rules : HARD derived
         clue = 324'h000580000_000010800_040000005_200000306_600873200_000020400_060200008_000100090_790060103;
          // 26 clues
       end
      244 : begin
         soln_sig = signature(324'h627594831_543168792_981237564_134672985_852913476_769845123_316759248_498321657_275486319);
         // Rules : HARD derived
         clue = 324'h000590800_000060000_000207060_030000900_000003470_009040020_000000200_498300000_075000019;
          // 24 clues
       end
      245 : begin
         soln_sig = signature(324'h143597682_862413975_795628314_621934758_958172463_437865291_279381546_384756129_516249837);
         // Rules : HARD derived
         clue = 324'h000597000_800010900_000000004_620000750_058000000_000000000_009380006_300756120_000200000;
          // 24 clues
       end
      246 : begin
         soln_sig = signature(324'h584619327_613278459_729543168_952137684_178964532_346825971_237451896_861392745_495786213);
         // Rules : EASY derived
         clue = 324'h000600007_003008000_729000000_000030084_108004002_000020900_007050000_801000040_005700010;
          // 24 clues
       end
      247 : begin
         soln_sig = signature(324'h145679382_978325146_326481597_682754931_493162758_751893624_234917865_819546273_567238419);
         // Rules : HARD derived
         clue = 324'h000600080_970005100_320400097_600000001_003100000_700000020_004900005_000040273_000038000;
          // 26 clues
       end
      248 : begin
         soln_sig = signature(324'h219673485_875429613_643185972_536748129_198236754_724951368_481597236_362814597_957362841);
         // Rules : MEDIUM derived
         clue = 324'h000600085_070009000_003080000_000008000_190000004_700050360_480097006_000000507_900002000;
          // 24 clues
       end
      249 : begin
         soln_sig = signature(324'h314682597_692457183_857931264_276198435_538724916_149563872_781345629_925876341_463219758);
         // Rules : MEDIUM
         clue = 324'h000600097_002057000_850000200_000108005_530000010_009003002_080040009_900000041_003000000;
          // 25 clues
       end
      250 : begin
         soln_sig = signature(324'h537629184_812547936_496381572_981763425_754892613_623415897_279154368_165238749_348976251);
         // Rules : HARD derived
         clue = 324'h000600104_800000006_090000070_081003005_700002600_000010000_009050360_000208700_040000001;
          // 24 clues
       end
      251 : begin
         soln_sig = signature(324'h738691542_295438176_461725839_984316257_623547981_517289364_146852793_352974618_879163425);
         // Rules : HARD derived
         clue = 324'h000600500_200030100_060705009_000010007_023000000_500289000_100052003_000070010_870000000;
          // 25 clues
       end
      252 : begin
         soln_sig = signature(324'h431682597_598137426_762549183_857326914_613954278_249871635_175493862_924768351_386215749);
         // Rules : MEDIUM derived
         clue = 324'h000602000_000030400_700000183_050000900_003004000_200000000_005400002_004008301_000210709;
          // 24 clues
       end
      253 : begin
         soln_sig = signature(324'h834679215_165284397_279153684_347968152_591342768_628517943_953426871_712895436_486731529);
         // Rules : HARD derived
         clue = 324'h000609000_005200097_070150600_040000102_000040700_008507000_053026800_010000030_000000020;
          // 26 clues
       end
      254 : begin
         soln_sig = signature(324'h528674139_793152846_461893572_912537684_634289751_857461923_386925417_175346298_249718365);
         // Rules : MEDIUM derived
         clue = 324'h000670100_093002000_401000500_002037004_030080001_007400000_380005000_000040200_009000060;
          // 25 clues
       end
      255 : begin
         soln_sig = signature(324'h134685297_596273184_782149563_879456321_641832759_253917846_917568432_468321975_325794618);
         // Rules : MEDIUM derived
         clue = 324'h000680000_090203000_700009500_000000300_000800059_200017000_010060002_460000000_005004008;
          // 23 clues
       end
   endcase
end
endmodule
